magic
tech sky130A
magscale 1 2
timestamp 1680903108
<< viali >>
rect 14105 24361 14139 24395
rect 18153 24361 18187 24395
rect 3985 24293 4019 24327
rect 6561 24293 6595 24327
rect 11713 24293 11747 24327
rect 15577 24293 15611 24327
rect 3249 24225 3283 24259
rect 8217 24225 8251 24259
rect 10977 24225 11011 24259
rect 12817 24225 12851 24259
rect 16037 24225 16071 24259
rect 16129 24225 16163 24259
rect 17601 24225 17635 24259
rect 18797 24225 18831 24259
rect 21281 24225 21315 24259
rect 25053 24225 25087 24259
rect 25145 24225 25179 24259
rect 1777 24157 1811 24191
rect 2237 24157 2271 24191
rect 4169 24157 4203 24191
rect 4813 24157 4847 24191
rect 6745 24157 6779 24191
rect 7205 24157 7239 24191
rect 9321 24157 9355 24191
rect 9781 24157 9815 24191
rect 11897 24157 11931 24191
rect 12357 24157 12391 24191
rect 14473 24157 14507 24191
rect 15945 24157 15979 24191
rect 17325 24157 17359 24191
rect 20177 24157 20211 24191
rect 22293 24157 22327 24191
rect 5825 24089 5859 24123
rect 15117 24089 15151 24123
rect 20545 24089 20579 24123
rect 22569 24089 22603 24123
rect 9137 24021 9171 24055
rect 16957 24021 16991 24055
rect 17417 24021 17451 24055
rect 17969 24021 18003 24055
rect 18521 24021 18555 24055
rect 18613 24021 18647 24055
rect 19441 24021 19475 24055
rect 21097 24021 21131 24055
rect 21465 24021 21499 24055
rect 21925 24021 21959 24055
rect 24041 24021 24075 24055
rect 24593 24021 24627 24055
rect 24961 24021 24995 24055
rect 11529 23817 11563 23851
rect 13737 23817 13771 23851
rect 14105 23817 14139 23851
rect 14473 23817 14507 23851
rect 16037 23817 16071 23851
rect 20867 23817 20901 23851
rect 3985 23749 4019 23783
rect 5825 23749 5859 23783
rect 9137 23749 9171 23783
rect 10885 23749 10919 23783
rect 11713 23749 11747 23783
rect 24317 23749 24351 23783
rect 24685 23749 24719 23783
rect 24961 23749 24995 23783
rect 25145 23749 25179 23783
rect 1685 23681 1719 23715
rect 2973 23681 3007 23715
rect 4813 23681 4847 23715
rect 7941 23681 7975 23715
rect 9781 23681 9815 23715
rect 12081 23681 12115 23715
rect 14565 23681 14599 23715
rect 15945 23681 15979 23715
rect 17233 23681 17267 23715
rect 22293 23681 22327 23715
rect 6561 23613 6595 23647
rect 6837 23613 6871 23647
rect 12541 23613 12575 23647
rect 14749 23613 14783 23647
rect 16221 23613 16255 23647
rect 17325 23613 17359 23647
rect 17509 23613 17543 23647
rect 18061 23613 18095 23647
rect 18337 23613 18371 23647
rect 20637 23613 20671 23647
rect 22569 23613 22603 23647
rect 24501 23613 24535 23647
rect 1869 23545 1903 23579
rect 15301 23545 15335 23579
rect 24041 23545 24075 23579
rect 2329 23477 2363 23511
rect 2421 23477 2455 23511
rect 15577 23477 15611 23511
rect 16865 23477 16899 23511
rect 19809 23477 19843 23511
rect 20085 23477 20119 23511
rect 20269 23477 20303 23511
rect 21833 23477 21867 23511
rect 25237 23477 25271 23511
rect 1501 23273 1535 23307
rect 1777 23273 1811 23307
rect 16773 23273 16807 23307
rect 21189 23273 21223 23307
rect 23397 23273 23431 23307
rect 13553 23205 13587 23239
rect 3249 23137 3283 23171
rect 6561 23137 6595 23171
rect 8309 23137 8343 23171
rect 10517 23137 10551 23171
rect 12173 23137 12207 23171
rect 15301 23137 15335 23171
rect 17785 23137 17819 23171
rect 18705 23137 18739 23171
rect 19717 23137 19751 23171
rect 21649 23137 21683 23171
rect 25145 23137 25179 23171
rect 2237 23069 2271 23103
rect 4077 23069 4111 23103
rect 5457 23069 5491 23103
rect 7205 23069 7239 23103
rect 9413 23069 9447 23103
rect 9873 23069 9907 23103
rect 11713 23069 11747 23103
rect 13737 23069 13771 23103
rect 15025 23069 15059 23103
rect 17601 23069 17635 23103
rect 19441 23069 19475 23103
rect 4261 23001 4295 23035
rect 14381 23001 14415 23035
rect 17693 23001 17727 23035
rect 18485 23001 18519 23035
rect 21925 23001 21959 23035
rect 25053 23001 25087 23035
rect 4721 22933 4755 22967
rect 9229 22933 9263 22967
rect 14473 22933 14507 22967
rect 17233 22933 17267 22967
rect 19073 22933 19107 22967
rect 23857 22933 23891 22967
rect 24593 22933 24627 22967
rect 24961 22933 24995 22967
rect 12081 22729 12115 22763
rect 13093 22729 13127 22763
rect 15393 22729 15427 22763
rect 16405 22729 16439 22763
rect 18613 22729 18647 22763
rect 2329 22661 2363 22695
rect 3985 22661 4019 22695
rect 5733 22661 5767 22695
rect 7297 22661 7331 22695
rect 8769 22661 8803 22695
rect 1685 22593 1719 22627
rect 2973 22593 3007 22627
rect 4813 22593 4847 22627
rect 6653 22593 6687 22627
rect 7573 22593 7607 22627
rect 12173 22593 12207 22627
rect 13001 22593 13035 22627
rect 13645 22593 13679 22627
rect 15945 22593 15979 22627
rect 16865 22593 16899 22627
rect 19165 22593 19199 22627
rect 19625 22593 19659 22627
rect 20269 22593 20303 22627
rect 22017 22593 22051 22627
rect 2513 22525 2547 22559
rect 9413 22525 9447 22559
rect 9689 22525 9723 22559
rect 12265 22525 12299 22559
rect 13921 22525 13955 22559
rect 17141 22525 17175 22559
rect 20545 22525 20579 22559
rect 22293 22525 22327 22559
rect 23305 22525 23339 22559
rect 23581 22525 23615 22559
rect 19349 22457 19383 22491
rect 1777 22389 1811 22423
rect 6745 22389 6779 22423
rect 11161 22389 11195 22423
rect 11713 22389 11747 22423
rect 16037 22389 16071 22423
rect 25053 22389 25087 22423
rect 25421 22389 25455 22423
rect 1685 22185 1719 22219
rect 10964 22185 10998 22219
rect 14552 22185 14586 22219
rect 18889 22185 18923 22219
rect 16497 22117 16531 22151
rect 2881 22049 2915 22083
rect 6101 22049 6135 22083
rect 8309 22049 8343 22083
rect 10701 22049 10735 22083
rect 12449 22049 12483 22083
rect 14289 22049 14323 22083
rect 17049 22049 17083 22083
rect 18153 22049 18187 22083
rect 18245 22049 18279 22083
rect 19993 22049 20027 22083
rect 25237 22049 25271 22083
rect 2237 21981 2271 22015
rect 3985 21981 4019 22015
rect 4261 21981 4295 22015
rect 5457 21981 5491 22015
rect 7389 21981 7423 22015
rect 8953 21981 8987 22015
rect 9505 21981 9539 22015
rect 13001 21981 13035 22015
rect 20361 21981 20395 22015
rect 22753 21981 22787 22015
rect 23213 21981 23247 22015
rect 23489 21981 23523 22015
rect 13553 21913 13587 21947
rect 16865 21913 16899 21947
rect 19533 21913 19567 21947
rect 20637 21913 20671 21947
rect 24961 21913 24995 21947
rect 9321 21845 9355 21879
rect 10057 21845 10091 21879
rect 12909 21845 12943 21879
rect 13645 21845 13679 21879
rect 16037 21845 16071 21879
rect 16957 21845 16991 21879
rect 17693 21845 17727 21879
rect 18061 21845 18095 21879
rect 18705 21845 18739 21879
rect 19625 21845 19659 21879
rect 22109 21845 22143 21879
rect 22569 21845 22603 21879
rect 24593 21845 24627 21879
rect 25053 21845 25087 21879
rect 2145 21641 2179 21675
rect 12633 21641 12667 21675
rect 13461 21641 13495 21675
rect 20453 21641 20487 21675
rect 22017 21641 22051 21675
rect 1685 21573 1719 21607
rect 11805 21573 11839 21607
rect 14289 21573 14323 21607
rect 18245 21573 18279 21607
rect 23673 21573 23707 21607
rect 2973 21505 3007 21539
rect 4813 21505 4847 21539
rect 6745 21505 6779 21539
rect 7389 21505 7423 21539
rect 9045 21505 9079 21539
rect 13369 21505 13403 21539
rect 14197 21505 14231 21539
rect 15393 21505 15427 21539
rect 15485 21505 15519 21539
rect 16221 21505 16255 21539
rect 17417 21505 17451 21539
rect 20821 21505 20855 21539
rect 21465 21505 21499 21539
rect 22385 21505 22419 21539
rect 23397 21505 23431 21539
rect 3525 21437 3559 21471
rect 5089 21437 5123 21471
rect 7665 21437 7699 21471
rect 9321 21437 9355 21471
rect 12725 21437 12759 21471
rect 12909 21437 12943 21471
rect 14381 21437 14415 21471
rect 15669 21437 15703 21471
rect 17509 21437 17543 21471
rect 17693 21437 17727 21471
rect 20913 21437 20947 21471
rect 21097 21437 21131 21471
rect 22477 21437 22511 21471
rect 22661 21437 22695 21471
rect 23029 21437 23063 21471
rect 25421 21369 25455 21403
rect 1777 21301 1811 21335
rect 6561 21301 6595 21335
rect 10793 21301 10827 21335
rect 11161 21301 11195 21335
rect 11253 21301 11287 21335
rect 11529 21301 11563 21335
rect 11897 21301 11931 21335
rect 12265 21301 12299 21335
rect 13829 21301 13863 21335
rect 15025 21301 15059 21335
rect 16037 21301 16071 21335
rect 16405 21301 16439 21335
rect 16681 21301 16715 21335
rect 17049 21301 17083 21335
rect 19533 21301 19567 21335
rect 25145 21301 25179 21335
rect 12909 21097 12943 21131
rect 16681 21097 16715 21131
rect 24593 21097 24627 21131
rect 6377 21029 6411 21063
rect 9965 21029 9999 21063
rect 15485 21029 15519 21063
rect 18889 21029 18923 21063
rect 21189 21029 21223 21063
rect 21649 21029 21683 21063
rect 23949 21029 23983 21063
rect 24133 21029 24167 21063
rect 2789 20961 2823 20995
rect 4445 20961 4479 20995
rect 7389 20961 7423 20995
rect 8677 20961 8711 20995
rect 10425 20961 10459 20995
rect 10517 20961 10551 20995
rect 11161 20961 11195 20995
rect 11437 20961 11471 20995
rect 15945 20961 15979 20995
rect 16037 20961 16071 20995
rect 17141 20961 17175 20995
rect 17233 20961 17267 20995
rect 18337 20961 18371 20995
rect 18521 20961 18555 20995
rect 19717 20961 19751 20995
rect 22201 20961 22235 20995
rect 23305 20961 23339 20995
rect 23397 20961 23431 20995
rect 25145 20961 25179 20995
rect 2237 20893 2271 20927
rect 4077 20893 4111 20927
rect 6009 20893 6043 20927
rect 7113 20893 7147 20927
rect 10333 20893 10367 20927
rect 14381 20893 14415 20927
rect 19441 20893 19475 20927
rect 23213 20893 23247 20927
rect 9321 20825 9355 20859
rect 13553 20825 13587 20859
rect 18245 20825 18279 20859
rect 25053 20825 25087 20859
rect 5825 20757 5859 20791
rect 6653 20757 6687 20791
rect 8953 20757 8987 20791
rect 13645 20757 13679 20791
rect 14473 20757 14507 20791
rect 14841 20757 14875 20791
rect 15025 20757 15059 20791
rect 15853 20757 15887 20791
rect 17049 20757 17083 20791
rect 17877 20757 17911 20791
rect 22017 20757 22051 20791
rect 22109 20757 22143 20791
rect 22845 20757 22879 20791
rect 24961 20757 24995 20791
rect 2237 20553 2271 20587
rect 4813 20553 4847 20587
rect 5181 20553 5215 20587
rect 6561 20553 6595 20587
rect 6837 20553 6871 20587
rect 7757 20553 7791 20587
rect 12449 20553 12483 20587
rect 18705 20553 18739 20587
rect 21005 20553 21039 20587
rect 11161 20485 11195 20519
rect 11345 20485 11379 20519
rect 11621 20485 11655 20519
rect 13829 20485 13863 20519
rect 16313 20485 16347 20519
rect 22477 20485 22511 20519
rect 23213 20485 23247 20519
rect 23765 20485 23799 20519
rect 1777 20417 1811 20451
rect 2421 20417 2455 20451
rect 3065 20417 3099 20451
rect 6009 20417 6043 20451
rect 7297 20417 7331 20451
rect 8585 20417 8619 20451
rect 9045 20417 9079 20451
rect 13185 20417 13219 20451
rect 13553 20417 13587 20451
rect 15853 20417 15887 20451
rect 22569 20417 22603 20451
rect 23489 20417 23523 20451
rect 3341 20349 3375 20383
rect 9321 20349 9355 20383
rect 11805 20349 11839 20383
rect 12541 20349 12575 20383
rect 12725 20349 12759 20383
rect 16957 20349 16991 20383
rect 17233 20349 17267 20383
rect 19257 20349 19291 20383
rect 19533 20349 19567 20383
rect 22661 20349 22695 20383
rect 21465 20281 21499 20315
rect 1593 20213 1627 20247
rect 5825 20213 5859 20247
rect 7113 20213 7147 20247
rect 8401 20213 8435 20247
rect 10793 20213 10827 20247
rect 12081 20213 12115 20247
rect 15301 20213 15335 20247
rect 15945 20213 15979 20247
rect 21281 20213 21315 20247
rect 22109 20213 22143 20247
rect 25237 20213 25271 20247
rect 10425 20009 10459 20043
rect 14933 20009 14967 20043
rect 17141 20009 17175 20043
rect 20729 20009 20763 20043
rect 4537 19941 4571 19975
rect 13369 19941 13403 19975
rect 17693 19941 17727 19975
rect 2513 19873 2547 19907
rect 5457 19873 5491 19907
rect 7113 19873 7147 19907
rect 7389 19873 7423 19907
rect 10885 19873 10919 19907
rect 10977 19873 11011 19907
rect 11621 19873 11655 19907
rect 15485 19873 15519 19907
rect 18245 19873 18279 19907
rect 20085 19873 20119 19907
rect 21097 19873 21131 19907
rect 23949 19873 23983 19907
rect 25053 19873 25087 19907
rect 25237 19873 25271 19907
rect 2237 19805 2271 19839
rect 4721 19805 4755 19839
rect 5181 19805 5215 19839
rect 6653 19805 6687 19839
rect 13921 19805 13955 19839
rect 14289 19805 14323 19839
rect 18889 19805 18923 19839
rect 20453 19805 20487 19839
rect 23673 19805 23707 19839
rect 8401 19737 8435 19771
rect 10793 19737 10827 19771
rect 11904 19737 11938 19771
rect 13645 19737 13679 19771
rect 15393 19737 15427 19771
rect 16221 19737 16255 19771
rect 17049 19737 17083 19771
rect 18153 19737 18187 19771
rect 19809 19737 19843 19771
rect 21373 19737 21407 19771
rect 23765 19737 23799 19771
rect 6469 19669 6503 19703
rect 9137 19669 9171 19703
rect 9781 19669 9815 19703
rect 15301 19669 15335 19703
rect 16313 19669 16347 19703
rect 18061 19669 18095 19703
rect 18705 19669 18739 19703
rect 19441 19669 19475 19703
rect 19901 19669 19935 19703
rect 22845 19669 22879 19703
rect 23305 19669 23339 19703
rect 24593 19669 24627 19703
rect 24961 19669 24995 19703
rect 3893 19465 3927 19499
rect 5825 19465 5859 19499
rect 8401 19465 8435 19499
rect 14473 19465 14507 19499
rect 14933 19465 14967 19499
rect 15301 19465 15335 19499
rect 18797 19465 18831 19499
rect 19257 19465 19291 19499
rect 19625 19465 19659 19499
rect 20453 19465 20487 19499
rect 20821 19465 20855 19499
rect 22017 19465 22051 19499
rect 22385 19465 22419 19499
rect 25053 19465 25087 19499
rect 15393 19397 15427 19431
rect 1961 19329 1995 19363
rect 4077 19329 4111 19363
rect 4813 19329 4847 19363
rect 6009 19329 6043 19363
rect 7297 19329 7331 19363
rect 7941 19329 7975 19363
rect 8585 19329 8619 19363
rect 9045 19329 9079 19363
rect 12725 19329 12759 19363
rect 16313 19329 16347 19363
rect 17049 19329 17083 19363
rect 19717 19329 19751 19363
rect 20913 19329 20947 19363
rect 23305 19329 23339 19363
rect 2237 19261 2271 19295
rect 4537 19261 4571 19295
rect 6469 19261 6503 19295
rect 6653 19261 6687 19295
rect 6837 19261 6871 19295
rect 9321 19261 9355 19295
rect 12081 19261 12115 19295
rect 13001 19261 13035 19295
rect 15577 19261 15611 19295
rect 17325 19261 17359 19295
rect 19901 19261 19935 19295
rect 21005 19261 21039 19295
rect 21557 19261 21591 19295
rect 22477 19261 22511 19295
rect 22569 19261 22603 19295
rect 23581 19261 23615 19295
rect 7757 19193 7791 19227
rect 11069 19193 11103 19227
rect 11529 19193 11563 19227
rect 16681 19193 16715 19227
rect 7113 19125 7147 19159
rect 10793 19125 10827 19159
rect 11253 19125 11287 19159
rect 11805 19125 11839 19159
rect 16129 19125 16163 19159
rect 21925 19125 21959 19159
rect 25329 19125 25363 19159
rect 1961 18921 1995 18955
rect 5825 18921 5859 18955
rect 6469 18921 6503 18955
rect 8401 18921 8435 18955
rect 9229 18921 9263 18955
rect 13001 18921 13035 18955
rect 14289 18921 14323 18955
rect 24409 18921 24443 18955
rect 2605 18853 2639 18887
rect 3249 18853 3283 18887
rect 5181 18853 5215 18887
rect 17233 18853 17267 18887
rect 7389 18785 7423 18819
rect 9873 18785 9907 18819
rect 13645 18785 13679 18819
rect 14749 18785 14783 18819
rect 14841 18785 14875 18819
rect 18613 18785 18647 18819
rect 23121 18785 23155 18819
rect 25053 18785 25087 18819
rect 25237 18785 25271 18819
rect 1685 18717 1719 18751
rect 2145 18717 2179 18751
rect 2789 18717 2823 18751
rect 3433 18717 3467 18751
rect 4261 18717 4295 18751
rect 4721 18717 4755 18751
rect 5365 18717 5399 18751
rect 6009 18717 6043 18751
rect 6653 18717 6687 18751
rect 7113 18717 7147 18751
rect 8593 18717 8627 18751
rect 9597 18717 9631 18751
rect 10425 18717 10459 18751
rect 15485 18717 15519 18751
rect 17509 18717 17543 18751
rect 18429 18717 18463 18751
rect 19625 18717 19659 18751
rect 20361 18717 20395 18751
rect 24133 18717 24167 18751
rect 24961 18717 24995 18751
rect 3893 18649 3927 18683
rect 4077 18649 4111 18683
rect 9689 18649 9723 18683
rect 13369 18649 13403 18683
rect 15761 18649 15795 18683
rect 20637 18649 20671 18683
rect 23029 18649 23063 18683
rect 23857 18649 23891 18683
rect 24041 18649 24075 18683
rect 4537 18581 4571 18615
rect 11713 18581 11747 18615
rect 12541 18581 12575 18615
rect 12725 18581 12759 18615
rect 13461 18581 13495 18615
rect 14657 18581 14691 18615
rect 17693 18581 17727 18615
rect 18061 18581 18095 18615
rect 18521 18581 18555 18615
rect 19441 18581 19475 18615
rect 19901 18581 19935 18615
rect 22109 18581 22143 18615
rect 22569 18581 22603 18615
rect 22937 18581 22971 18615
rect 24593 18581 24627 18615
rect 1593 18377 1627 18411
rect 3893 18377 3927 18411
rect 5181 18377 5215 18411
rect 5825 18377 5859 18411
rect 8309 18377 8343 18411
rect 12173 18377 12207 18411
rect 14289 18377 14323 18411
rect 15209 18377 15243 18411
rect 15669 18377 15703 18411
rect 16313 18377 16347 18411
rect 19717 18377 19751 18411
rect 21557 18377 21591 18411
rect 23305 18377 23339 18411
rect 24317 18377 24351 18411
rect 25053 18377 25087 18411
rect 2237 18309 2271 18343
rect 2789 18309 2823 18343
rect 9229 18309 9263 18343
rect 11069 18309 11103 18343
rect 13001 18309 13035 18343
rect 16497 18309 16531 18343
rect 20913 18309 20947 18343
rect 22017 18309 22051 18343
rect 24041 18309 24075 18343
rect 24961 18309 24995 18343
rect 1777 18241 1811 18275
rect 2973 18241 3007 18275
rect 3433 18241 3467 18275
rect 4721 18241 4755 18275
rect 5365 18241 5399 18275
rect 6009 18241 6043 18275
rect 7205 18241 7239 18275
rect 7849 18241 7883 18275
rect 8493 18241 8527 18275
rect 8953 18241 8987 18275
rect 15577 18241 15611 18275
rect 17233 18241 17267 18275
rect 18429 18241 18463 18275
rect 19625 18241 19659 18275
rect 20821 18241 20855 18275
rect 6745 18173 6779 18207
rect 12265 18173 12299 18207
rect 12357 18173 12391 18207
rect 15761 18173 15795 18207
rect 17325 18173 17359 18207
rect 17417 18173 17451 18207
rect 18521 18173 18555 18207
rect 18705 18173 18739 18207
rect 19855 18173 19889 18207
rect 21005 18173 21039 18207
rect 25237 18173 25271 18207
rect 4537 18105 4571 18139
rect 7021 18105 7055 18139
rect 11805 18105 11839 18139
rect 16865 18105 16899 18139
rect 24593 18105 24627 18139
rect 3249 18037 3283 18071
rect 6561 18037 6595 18071
rect 7665 18037 7699 18071
rect 10701 18037 10735 18071
rect 11253 18037 11287 18071
rect 18061 18037 18095 18071
rect 19257 18037 19291 18071
rect 20453 18037 20487 18071
rect 3249 17833 3283 17867
rect 6469 17833 6503 17867
rect 7757 17833 7791 17867
rect 17141 17833 17175 17867
rect 20992 17833 21026 17867
rect 22477 17833 22511 17867
rect 24593 17833 24627 17867
rect 18153 17765 18187 17799
rect 5181 17697 5215 17731
rect 9781 17697 9815 17731
rect 11989 17697 12023 17731
rect 12265 17697 12299 17731
rect 14289 17697 14323 17731
rect 14933 17697 14967 17731
rect 16681 17697 16715 17731
rect 17693 17697 17727 17731
rect 19993 17697 20027 17731
rect 20729 17697 20763 17731
rect 23765 17697 23799 17731
rect 23857 17697 23891 17731
rect 25053 17697 25087 17731
rect 25237 17697 25271 17731
rect 3433 17629 3467 17663
rect 4077 17629 4111 17663
rect 4721 17629 4755 17663
rect 5457 17629 5491 17663
rect 6653 17629 6687 17663
rect 7297 17629 7331 17663
rect 7941 17629 7975 17663
rect 8585 17629 8619 17663
rect 9321 17629 9355 17663
rect 17509 17629 17543 17663
rect 18797 17629 18831 17663
rect 19901 17629 19935 17663
rect 23673 17629 23707 17663
rect 10057 17561 10091 17595
rect 15209 17561 15243 17595
rect 22845 17561 22879 17595
rect 23029 17561 23063 17595
rect 4261 17493 4295 17527
rect 4537 17493 4571 17527
rect 7113 17493 7147 17527
rect 8401 17493 8435 17527
rect 9137 17493 9171 17527
rect 11529 17493 11563 17527
rect 13737 17493 13771 17527
rect 17601 17493 17635 17527
rect 18613 17493 18647 17527
rect 19441 17493 19475 17527
rect 19809 17493 19843 17527
rect 23305 17493 23339 17527
rect 24409 17493 24443 17527
rect 24961 17493 24995 17527
rect 3893 17289 3927 17323
rect 7205 17289 7239 17323
rect 7849 17289 7883 17323
rect 15853 17289 15887 17323
rect 20085 17289 20119 17323
rect 20545 17289 20579 17323
rect 9505 17221 9539 17255
rect 11989 17221 12023 17255
rect 17325 17221 17359 17255
rect 21189 17221 21223 17255
rect 21925 17221 21959 17255
rect 22109 17221 22143 17255
rect 22293 17221 22327 17255
rect 4077 17153 4111 17187
rect 6745 17153 6779 17187
rect 7389 17153 7423 17187
rect 8033 17153 8067 17187
rect 8769 17153 8803 17187
rect 9229 17153 9263 17187
rect 11253 17153 11287 17187
rect 11713 17153 11747 17187
rect 14473 17153 14507 17187
rect 15025 17153 15059 17187
rect 17233 17153 17267 17187
rect 18337 17153 18371 17187
rect 22569 17153 22603 17187
rect 24869 17153 24903 17187
rect 25329 17153 25363 17187
rect 4537 17085 4571 17119
rect 4813 17085 4847 17119
rect 10977 17085 11011 17119
rect 13461 17085 13495 17119
rect 13921 17085 13955 17119
rect 15945 17085 15979 17119
rect 16037 17085 16071 17119
rect 17417 17085 17451 17119
rect 17877 17085 17911 17119
rect 18613 17085 18647 17119
rect 25053 17085 25087 17119
rect 16865 17017 16899 17051
rect 24317 17017 24351 17051
rect 6561 16949 6595 16983
rect 8585 16949 8619 16983
rect 14841 16949 14875 16983
rect 15485 16949 15519 16983
rect 22832 16949 22866 16983
rect 7297 16745 7331 16779
rect 8401 16745 8435 16779
rect 9045 16745 9079 16779
rect 16037 16745 16071 16779
rect 19704 16745 19738 16779
rect 21189 16745 21223 16779
rect 22556 16745 22590 16779
rect 6929 16609 6963 16643
rect 9229 16609 9263 16643
rect 11253 16609 11287 16643
rect 11437 16609 11471 16643
rect 12265 16609 12299 16643
rect 14289 16609 14323 16643
rect 17141 16609 17175 16643
rect 17417 16609 17451 16643
rect 19441 16609 19475 16643
rect 22293 16609 22327 16643
rect 4169 16541 4203 16575
rect 4721 16541 4755 16575
rect 7481 16541 7515 16575
rect 7941 16541 7975 16575
rect 8585 16541 8619 16575
rect 9689 16541 9723 16575
rect 11161 16541 11195 16575
rect 11989 16541 12023 16575
rect 16681 16541 16715 16575
rect 21649 16541 21683 16575
rect 24593 16541 24627 16575
rect 25237 16541 25271 16575
rect 14565 16473 14599 16507
rect 3985 16405 4019 16439
rect 7757 16405 7791 16439
rect 9505 16405 9539 16439
rect 10149 16405 10183 16439
rect 10793 16405 10827 16439
rect 13737 16405 13771 16439
rect 16497 16405 16531 16439
rect 18889 16405 18923 16439
rect 24041 16405 24075 16439
rect 4261 16201 4295 16235
rect 8033 16201 8067 16235
rect 10793 16201 10827 16235
rect 10885 16201 10919 16235
rect 15485 16201 15519 16235
rect 15853 16201 15887 16235
rect 16681 16201 16715 16235
rect 18429 16201 18463 16235
rect 19809 16201 19843 16235
rect 20913 16201 20947 16235
rect 22477 16201 22511 16235
rect 25329 16201 25363 16235
rect 15117 16133 15151 16167
rect 23765 16133 23799 16167
rect 8677 16065 8711 16099
rect 9321 16065 9355 16099
rect 9965 16065 9999 16099
rect 14289 16065 14323 16099
rect 17141 16065 17175 16099
rect 19717 16065 19751 16099
rect 21557 16065 21591 16099
rect 22385 16065 22419 16099
rect 24685 16065 24719 16099
rect 25145 16065 25179 16099
rect 8217 15997 8251 16031
rect 11069 15997 11103 16031
rect 11713 15997 11747 16031
rect 11989 15997 12023 16031
rect 13461 15997 13495 16031
rect 14381 15997 14415 16031
rect 14565 15997 14599 16031
rect 15945 15997 15979 16031
rect 16037 15997 16071 16031
rect 19901 15997 19935 16031
rect 21005 15997 21039 16031
rect 21097 15997 21131 16031
rect 22661 15997 22695 16031
rect 23857 15997 23891 16031
rect 23949 15997 23983 16031
rect 9137 15929 9171 15963
rect 9781 15929 9815 15963
rect 19349 15929 19383 15963
rect 23029 15929 23063 15963
rect 24869 15929 24903 15963
rect 8493 15861 8527 15895
rect 10425 15861 10459 15895
rect 13921 15861 13955 15895
rect 14933 15861 14967 15895
rect 20545 15861 20579 15895
rect 22017 15861 22051 15895
rect 23397 15861 23431 15895
rect 9873 15657 9907 15691
rect 12725 15657 12759 15691
rect 13829 15657 13863 15691
rect 16037 15657 16071 15691
rect 16681 15657 16715 15691
rect 18705 15657 18739 15691
rect 23397 15657 23431 15691
rect 24501 15657 24535 15691
rect 9229 15589 9263 15623
rect 12265 15589 12299 15623
rect 16405 15589 16439 15623
rect 20729 15589 20763 15623
rect 24041 15589 24075 15623
rect 10793 15521 10827 15555
rect 13185 15521 13219 15555
rect 13369 15521 13403 15555
rect 14289 15521 14323 15555
rect 17233 15521 17267 15555
rect 20085 15521 20119 15555
rect 21373 15521 21407 15555
rect 8769 15453 8803 15487
rect 9413 15453 9447 15487
rect 10057 15453 10091 15487
rect 10517 15453 10551 15487
rect 13093 15453 13127 15487
rect 16957 15453 16991 15487
rect 19993 15453 20027 15487
rect 21097 15453 21131 15487
rect 22019 15453 22053 15487
rect 22753 15453 22787 15487
rect 23581 15453 23615 15487
rect 14565 15385 14599 15419
rect 19901 15385 19935 15419
rect 22201 15385 22235 15419
rect 23857 15385 23891 15419
rect 24869 15385 24903 15419
rect 25053 15385 25087 15419
rect 18981 15317 19015 15351
rect 19533 15317 19567 15351
rect 21189 15317 21223 15351
rect 22845 15317 22879 15351
rect 25329 15317 25363 15351
rect 9413 15113 9447 15147
rect 9689 15113 9723 15147
rect 10977 15113 11011 15147
rect 13461 15113 13495 15147
rect 13921 15113 13955 15147
rect 15301 15113 15335 15147
rect 15485 15113 15519 15147
rect 18981 15113 19015 15147
rect 21097 15113 21131 15147
rect 21465 15113 21499 15147
rect 21649 15113 21683 15147
rect 24593 15113 24627 15147
rect 9873 15045 9907 15079
rect 17141 15045 17175 15079
rect 23121 15045 23155 15079
rect 10517 14977 10551 15011
rect 11161 14977 11195 15011
rect 14565 14977 14599 15011
rect 15025 14977 15059 15011
rect 16865 14977 16899 15011
rect 22109 14977 22143 15011
rect 11713 14909 11747 14943
rect 11989 14909 12023 14943
rect 16129 14909 16163 14943
rect 19349 14909 19383 14943
rect 19625 14909 19659 14943
rect 22845 14909 22879 14943
rect 25053 14909 25087 14943
rect 10333 14841 10367 14875
rect 14841 14841 14875 14875
rect 22293 14841 22327 14875
rect 10057 14773 10091 14807
rect 18613 14773 18647 14807
rect 10425 14569 10459 14603
rect 12449 14569 12483 14603
rect 12909 14569 12943 14603
rect 13461 14569 13495 14603
rect 19441 14569 19475 14603
rect 20453 14569 20487 14603
rect 22937 14569 22971 14603
rect 25237 14569 25271 14603
rect 16037 14501 16071 14535
rect 18245 14501 18279 14535
rect 25421 14501 25455 14535
rect 10977 14433 11011 14467
rect 13553 14433 13587 14467
rect 14289 14433 14323 14467
rect 14565 14433 14599 14467
rect 16773 14433 16807 14467
rect 19993 14433 20027 14467
rect 23765 14433 23799 14467
rect 23949 14433 23983 14467
rect 10701 14365 10735 14399
rect 13093 14365 13127 14399
rect 16497 14365 16531 14399
rect 19901 14365 19935 14399
rect 20821 14365 20855 14399
rect 24685 14365 24719 14399
rect 18705 14297 18739 14331
rect 19809 14297 19843 14331
rect 22569 14297 22603 14331
rect 23305 14229 23339 14263
rect 23673 14229 23707 14263
rect 24777 14229 24811 14263
rect 11805 14025 11839 14059
rect 12449 14025 12483 14059
rect 13093 14025 13127 14059
rect 15485 14025 15519 14059
rect 16129 14025 16163 14059
rect 17509 14025 17543 14059
rect 19533 14025 19567 14059
rect 20269 14025 20303 14059
rect 21189 14025 21223 14059
rect 11345 13957 11379 13991
rect 18245 13957 18279 13991
rect 21097 13957 21131 13991
rect 25145 13957 25179 13991
rect 11161 13889 11195 13923
rect 11989 13889 12023 13923
rect 12633 13889 12667 13923
rect 13277 13889 13311 13923
rect 13737 13889 13771 13923
rect 15761 13889 15795 13923
rect 16313 13889 16347 13923
rect 17417 13889 17451 13923
rect 22109 13889 22143 13923
rect 22845 13889 22879 13923
rect 16681 13821 16715 13855
rect 17601 13821 17635 13855
rect 21281 13821 21315 13855
rect 22293 13821 22327 13855
rect 23121 13821 23155 13855
rect 24593 13821 24627 13855
rect 25329 13821 25363 13855
rect 14000 13685 14034 13719
rect 17049 13685 17083 13719
rect 20729 13685 20763 13719
rect 13829 13481 13863 13515
rect 16037 13481 16071 13515
rect 18705 13481 18739 13515
rect 21465 13481 21499 13515
rect 22188 13481 22222 13515
rect 23949 13481 23983 13515
rect 13553 13413 13587 13447
rect 24133 13413 24167 13447
rect 12081 13345 12115 13379
rect 14289 13345 14323 13379
rect 16497 13345 16531 13379
rect 16773 13345 16807 13379
rect 21925 13345 21959 13379
rect 25145 13345 25179 13379
rect 11805 13277 11839 13311
rect 18889 13277 18923 13311
rect 19717 13277 19751 13311
rect 25053 13277 25087 13311
rect 9597 13209 9631 13243
rect 14565 13209 14599 13243
rect 19349 13209 19383 13243
rect 19993 13209 20027 13243
rect 24409 13209 24443 13243
rect 24961 13209 24995 13243
rect 10885 13141 10919 13175
rect 18245 13141 18279 13175
rect 23673 13141 23707 13175
rect 24593 13141 24627 13175
rect 11529 12937 11563 12971
rect 12633 12937 12667 12971
rect 14289 12937 14323 12971
rect 16313 12937 16347 12971
rect 20729 12937 20763 12971
rect 21373 12937 21407 12971
rect 23765 12937 23799 12971
rect 25513 12937 25547 12971
rect 13001 12869 13035 12903
rect 17141 12869 17175 12903
rect 25053 12869 25087 12903
rect 25329 12869 25363 12903
rect 16865 12801 16899 12835
rect 19441 12801 19475 12835
rect 20637 12801 20671 12835
rect 21465 12801 21499 12835
rect 22017 12801 22051 12835
rect 24041 12801 24075 12835
rect 24225 12801 24259 12835
rect 24777 12801 24811 12835
rect 15209 12733 15243 12767
rect 15485 12733 15519 12767
rect 19533 12733 19567 12767
rect 19625 12733 19659 12767
rect 20821 12733 20855 12767
rect 22293 12733 22327 12767
rect 18613 12665 18647 12699
rect 24593 12665 24627 12699
rect 19073 12597 19107 12631
rect 20269 12597 20303 12631
rect 13461 12393 13495 12427
rect 13737 12393 13771 12427
rect 13921 12393 13955 12427
rect 15485 12393 15519 12427
rect 17509 12393 17543 12427
rect 24409 12325 24443 12359
rect 24685 12325 24719 12359
rect 14289 12257 14323 12291
rect 15761 12257 15795 12291
rect 17969 12257 18003 12291
rect 21189 12257 21223 12291
rect 22293 12257 22327 12291
rect 22569 12257 22603 12291
rect 25053 12257 25087 12291
rect 14565 12189 14599 12223
rect 19441 12189 19475 12223
rect 16037 12121 16071 12155
rect 18705 12121 18739 12155
rect 19717 12121 19751 12155
rect 21649 12121 21683 12155
rect 18797 12053 18831 12087
rect 24041 12053 24075 12087
rect 14565 11849 14599 11883
rect 15117 11849 15151 11883
rect 15669 11849 15703 11883
rect 21465 11849 21499 11883
rect 13093 11781 13127 11815
rect 19717 11781 19751 11815
rect 23305 11781 23339 11815
rect 25145 11781 25179 11815
rect 12817 11713 12851 11747
rect 15301 11713 15335 11747
rect 16313 11713 16347 11747
rect 19441 11713 19475 11747
rect 22201 11713 22235 11747
rect 23949 11713 23983 11747
rect 17141 11645 17175 11679
rect 17417 11645 17451 11679
rect 16129 11577 16163 11611
rect 21189 11577 21223 11611
rect 15761 11509 15795 11543
rect 16773 11509 16807 11543
rect 18889 11509 18923 11543
rect 14657 11305 14691 11339
rect 15485 11305 15519 11339
rect 16129 11305 16163 11339
rect 16773 11305 16807 11339
rect 17417 11305 17451 11339
rect 19257 11305 19291 11339
rect 19533 11305 19567 11339
rect 20453 11305 20487 11339
rect 20821 11305 20855 11339
rect 21189 11305 21223 11339
rect 24593 11305 24627 11339
rect 25237 11305 25271 11339
rect 25513 11305 25547 11339
rect 18705 11237 18739 11271
rect 22017 11237 22051 11271
rect 25145 11237 25179 11271
rect 18061 11169 18095 11203
rect 23857 11169 23891 11203
rect 15669 11101 15703 11135
rect 16313 11101 16347 11135
rect 16957 11101 16991 11135
rect 17601 11101 17635 11135
rect 18889 11101 18923 11135
rect 19993 11101 20027 11135
rect 21373 11101 21407 11135
rect 22201 11101 22235 11135
rect 22661 11101 22695 11135
rect 24777 11101 24811 11135
rect 20085 10965 20119 10999
rect 20637 10965 20671 10999
rect 21649 10965 21683 10999
rect 15761 10761 15795 10795
rect 16405 10761 16439 10795
rect 17141 10761 17175 10795
rect 17325 10761 17359 10795
rect 17417 10761 17451 10795
rect 18061 10761 18095 10795
rect 19349 10761 19383 10795
rect 23305 10693 23339 10727
rect 16957 10625 16991 10659
rect 18245 10625 18279 10659
rect 18889 10625 18923 10659
rect 19533 10625 19567 10659
rect 20177 10625 20211 10659
rect 20821 10625 20855 10659
rect 21465 10625 21499 10659
rect 22109 10625 22143 10659
rect 23949 10625 23983 10659
rect 24685 10557 24719 10591
rect 18705 10489 18739 10523
rect 19993 10489 20027 10523
rect 20637 10421 20671 10455
rect 21281 10421 21315 10455
rect 17417 10217 17451 10251
rect 20729 10217 20763 10251
rect 24593 10217 24627 10251
rect 19441 10149 19475 10183
rect 18061 10081 18095 10115
rect 21373 10081 21407 10115
rect 21649 10081 21683 10115
rect 23857 10081 23891 10115
rect 25145 10081 25179 10115
rect 17601 10013 17635 10047
rect 18337 10013 18371 10047
rect 19625 10013 19659 10047
rect 20913 10013 20947 10047
rect 20085 9945 20119 9979
rect 24961 9945 24995 9979
rect 25053 9945 25087 9979
rect 23121 9877 23155 9911
rect 23305 9605 23339 9639
rect 18245 9537 18279 9571
rect 18889 9537 18923 9571
rect 19533 9537 19567 9571
rect 20177 9537 20211 9571
rect 20913 9537 20947 9571
rect 21281 9537 21315 9571
rect 21465 9537 21499 9571
rect 21557 9537 21591 9571
rect 22109 9537 22143 9571
rect 23949 9537 23983 9571
rect 24777 9469 24811 9503
rect 18061 9401 18095 9435
rect 19349 9401 19383 9435
rect 18705 9333 18739 9367
rect 19993 9333 20027 9367
rect 20729 9333 20763 9367
rect 11805 9129 11839 9163
rect 19073 9129 19107 9163
rect 21005 9129 21039 9163
rect 25421 9129 25455 9163
rect 21281 9061 21315 9095
rect 10057 8993 10091 9027
rect 19441 8993 19475 9027
rect 19717 8993 19751 9027
rect 23857 8993 23891 9027
rect 21465 8925 21499 8959
rect 22661 8925 22695 8959
rect 10333 8857 10367 8891
rect 12081 8857 12115 8891
rect 24685 8857 24719 8891
rect 22017 8789 22051 8823
rect 24777 8789 24811 8823
rect 19441 8585 19475 8619
rect 23305 8517 23339 8551
rect 19625 8449 19659 8483
rect 20269 8449 20303 8483
rect 20913 8449 20947 8483
rect 21281 8449 21315 8483
rect 22109 8449 22143 8483
rect 23949 8449 23983 8483
rect 21465 8381 21499 8415
rect 24593 8381 24627 8415
rect 20085 8313 20119 8347
rect 20729 8313 20763 8347
rect 21373 8041 21407 8075
rect 22017 8041 22051 8075
rect 19993 7905 20027 7939
rect 20085 7905 20119 7939
rect 23857 7905 23891 7939
rect 20913 7837 20947 7871
rect 21557 7837 21591 7871
rect 22201 7837 22235 7871
rect 22845 7837 22879 7871
rect 24869 7837 24903 7871
rect 20729 7701 20763 7735
rect 24685 7701 24719 7735
rect 21281 7497 21315 7531
rect 23305 7429 23339 7463
rect 20821 7361 20855 7395
rect 21465 7361 21499 7395
rect 22293 7361 22327 7395
rect 23949 7361 23983 7395
rect 24685 7293 24719 7327
rect 20637 7225 20671 7259
rect 20637 6885 20671 6919
rect 23857 6817 23891 6851
rect 20821 6749 20855 6783
rect 21465 6749 21499 6783
rect 22201 6749 22235 6783
rect 22661 6749 22695 6783
rect 24685 6681 24719 6715
rect 24869 6681 24903 6715
rect 21281 6613 21315 6647
rect 22017 6613 22051 6647
rect 9321 6409 9355 6443
rect 21649 6409 21683 6443
rect 23305 6341 23339 6375
rect 8677 6273 8711 6307
rect 22293 6273 22327 6307
rect 23949 6273 23983 6307
rect 24777 6205 24811 6239
rect 22017 5865 22051 5899
rect 21373 5797 21407 5831
rect 21557 5661 21591 5695
rect 22201 5661 22235 5695
rect 22845 5661 22879 5695
rect 24869 5661 24903 5695
rect 23857 5593 23891 5627
rect 24685 5525 24719 5559
rect 23305 5253 23339 5287
rect 22293 5185 22327 5219
rect 23949 5185 23983 5219
rect 24685 5117 24719 5151
rect 22385 4777 22419 4811
rect 22661 4573 22695 4607
rect 24869 4573 24903 4607
rect 23857 4505 23891 4539
rect 24685 4437 24719 4471
rect 20269 4097 20303 4131
rect 22293 4097 22327 4131
rect 24133 4097 24167 4131
rect 21281 4029 21315 4063
rect 23305 4029 23339 4063
rect 24777 4029 24811 4063
rect 20821 3485 20855 3519
rect 22845 3485 22879 3519
rect 24777 3485 24811 3519
rect 22017 3417 22051 3451
rect 23857 3417 23891 3451
rect 24593 3349 24627 3383
rect 6837 3145 6871 3179
rect 23305 3077 23339 3111
rect 25145 3077 25179 3111
rect 7021 3009 7055 3043
rect 18429 3009 18463 3043
rect 20085 3009 20119 3043
rect 22293 3009 22327 3043
rect 24133 3009 24167 3043
rect 19349 2941 19383 2975
rect 21281 2941 21315 2975
rect 7481 2601 7515 2635
rect 19809 2533 19843 2567
rect 6837 2397 6871 2431
rect 20269 2397 20303 2431
rect 22845 2397 22879 2431
rect 21281 2329 21315 2363
rect 23857 2329 23891 2363
rect 6561 2261 6595 2295
<< metal1 >>
rect 3050 26392 3056 26444
rect 3108 26432 3114 26444
rect 3326 26432 3332 26444
rect 3108 26404 3332 26432
rect 3108 26392 3114 26404
rect 3326 26392 3332 26404
rect 3384 26392 3390 26444
rect 2130 26324 2136 26376
rect 2188 26364 2194 26376
rect 22186 26364 22192 26376
rect 2188 26336 22192 26364
rect 2188 26324 2194 26336
rect 22186 26324 22192 26336
rect 22244 26324 22250 26376
rect 9582 26256 9588 26308
rect 9640 26296 9646 26308
rect 21818 26296 21824 26308
rect 9640 26268 21824 26296
rect 9640 26256 9646 26268
rect 21818 26256 21824 26268
rect 21876 26256 21882 26308
rect 7558 25236 7564 25288
rect 7616 25276 7622 25288
rect 26142 25276 26148 25288
rect 7616 25248 26148 25276
rect 7616 25236 7622 25248
rect 26142 25236 26148 25248
rect 26200 25236 26206 25288
rect 3602 25168 3608 25220
rect 3660 25208 3666 25220
rect 25590 25208 25596 25220
rect 3660 25180 25596 25208
rect 3660 25168 3666 25180
rect 25590 25168 25596 25180
rect 25648 25168 25654 25220
rect 5166 25100 5172 25152
rect 5224 25140 5230 25152
rect 15838 25140 15844 25152
rect 5224 25112 15844 25140
rect 5224 25100 5230 25112
rect 15838 25100 15844 25112
rect 15896 25100 15902 25152
rect 1946 25032 1952 25084
rect 2004 25072 2010 25084
rect 13998 25072 14004 25084
rect 2004 25044 14004 25072
rect 2004 25032 2010 25044
rect 13998 25032 14004 25044
rect 14056 25032 14062 25084
rect 6638 24964 6644 25016
rect 6696 25004 6702 25016
rect 6696 24976 23428 25004
rect 6696 24964 6702 24976
rect 9858 24896 9864 24948
rect 9916 24936 9922 24948
rect 17310 24936 17316 24948
rect 9916 24908 17316 24936
rect 9916 24896 9922 24908
rect 17310 24896 17316 24908
rect 17368 24896 17374 24948
rect 8478 24828 8484 24880
rect 8536 24868 8542 24880
rect 18138 24868 18144 24880
rect 8536 24840 18144 24868
rect 8536 24828 8542 24840
rect 18138 24828 18144 24840
rect 18196 24828 18202 24880
rect 20622 24828 20628 24880
rect 20680 24868 20686 24880
rect 23198 24868 23204 24880
rect 20680 24840 23204 24868
rect 20680 24828 20686 24840
rect 23198 24828 23204 24840
rect 23256 24828 23262 24880
rect 5810 24760 5816 24812
rect 5868 24800 5874 24812
rect 8386 24800 8392 24812
rect 5868 24772 8392 24800
rect 5868 24760 5874 24772
rect 8386 24760 8392 24772
rect 8444 24760 8450 24812
rect 9766 24760 9772 24812
rect 9824 24800 9830 24812
rect 16022 24800 16028 24812
rect 9824 24772 16028 24800
rect 9824 24760 9830 24772
rect 16022 24760 16028 24772
rect 16080 24760 16086 24812
rect 23400 24800 23428 24976
rect 25130 24800 25136 24812
rect 23400 24772 25136 24800
rect 25130 24760 25136 24772
rect 25188 24760 25194 24812
rect 5994 24692 6000 24744
rect 6052 24732 6058 24744
rect 14090 24732 14096 24744
rect 6052 24704 14096 24732
rect 6052 24692 6058 24704
rect 14090 24692 14096 24704
rect 14148 24692 14154 24744
rect 7742 24624 7748 24676
rect 7800 24664 7806 24676
rect 7800 24636 12434 24664
rect 7800 24624 7806 24636
rect 5258 24556 5264 24608
rect 5316 24596 5322 24608
rect 8570 24596 8576 24608
rect 5316 24568 8576 24596
rect 5316 24556 5322 24568
rect 8570 24556 8576 24568
rect 8628 24556 8634 24608
rect 12406 24596 12434 24636
rect 16850 24624 16856 24676
rect 16908 24664 16914 24676
rect 20622 24664 20628 24676
rect 16908 24636 20628 24664
rect 16908 24624 16914 24636
rect 20622 24624 20628 24636
rect 20680 24624 20686 24676
rect 19702 24596 19708 24608
rect 12406 24568 19708 24596
rect 19702 24556 19708 24568
rect 19760 24556 19766 24608
rect 1104 24506 25852 24528
rect 1104 24454 2950 24506
rect 3002 24454 3014 24506
rect 3066 24454 3078 24506
rect 3130 24454 3142 24506
rect 3194 24454 3206 24506
rect 3258 24454 12950 24506
rect 13002 24454 13014 24506
rect 13066 24454 13078 24506
rect 13130 24454 13142 24506
rect 13194 24454 13206 24506
rect 13258 24454 22950 24506
rect 23002 24454 23014 24506
rect 23066 24454 23078 24506
rect 23130 24454 23142 24506
rect 23194 24454 23206 24506
rect 23258 24454 25852 24506
rect 1104 24432 25852 24454
rect 13998 24352 14004 24404
rect 14056 24392 14062 24404
rect 14093 24395 14151 24401
rect 14093 24392 14105 24395
rect 14056 24364 14105 24392
rect 14056 24352 14062 24364
rect 14093 24361 14105 24364
rect 14139 24361 14151 24395
rect 14093 24355 14151 24361
rect 3973 24327 4031 24333
rect 3973 24293 3985 24327
rect 4019 24324 4031 24327
rect 6362 24324 6368 24336
rect 4019 24296 6368 24324
rect 4019 24293 4031 24296
rect 3973 24287 4031 24293
rect 6362 24284 6368 24296
rect 6420 24284 6426 24336
rect 6546 24284 6552 24336
rect 6604 24284 6610 24336
rect 8478 24324 8484 24336
rect 8128 24296 8484 24324
rect 3237 24259 3295 24265
rect 3237 24225 3249 24259
rect 3283 24256 3295 24259
rect 6454 24256 6460 24268
rect 3283 24228 6460 24256
rect 3283 24225 3295 24228
rect 3237 24219 3295 24225
rect 6454 24216 6460 24228
rect 6512 24216 6518 24268
rect 8128 24256 8156 24296
rect 8478 24284 8484 24296
rect 8536 24284 8542 24336
rect 8846 24284 8852 24336
rect 8904 24324 8910 24336
rect 11701 24327 11759 24333
rect 11701 24324 11713 24327
rect 8904 24296 11713 24324
rect 8904 24284 8910 24296
rect 11701 24293 11713 24296
rect 11747 24293 11759 24327
rect 11701 24287 11759 24293
rect 12342 24284 12348 24336
rect 12400 24324 12406 24336
rect 12400 24296 12848 24324
rect 12400 24284 12406 24296
rect 6656 24228 8156 24256
rect 8205 24259 8263 24265
rect 1762 24148 1768 24200
rect 1820 24148 1826 24200
rect 2225 24191 2283 24197
rect 2225 24157 2237 24191
rect 2271 24188 2283 24191
rect 3878 24188 3884 24200
rect 2271 24160 3884 24188
rect 2271 24157 2283 24160
rect 2225 24151 2283 24157
rect 3878 24148 3884 24160
rect 3936 24148 3942 24200
rect 4157 24191 4215 24197
rect 4157 24157 4169 24191
rect 4203 24157 4215 24191
rect 4157 24151 4215 24157
rect 4172 24120 4200 24151
rect 4798 24148 4804 24200
rect 4856 24148 4862 24200
rect 6656 24188 6684 24228
rect 8205 24225 8217 24259
rect 8251 24256 8263 24259
rect 9674 24256 9680 24268
rect 8251 24228 9680 24256
rect 8251 24225 8263 24228
rect 8205 24219 8263 24225
rect 9674 24216 9680 24228
rect 9732 24216 9738 24268
rect 10962 24216 10968 24268
rect 11020 24216 11026 24268
rect 11790 24216 11796 24268
rect 11848 24256 11854 24268
rect 12820 24265 12848 24296
rect 12805 24259 12863 24265
rect 11848 24228 12388 24256
rect 11848 24216 11854 24228
rect 5736 24160 6684 24188
rect 5736 24120 5764 24160
rect 6730 24148 6736 24200
rect 6788 24148 6794 24200
rect 7193 24191 7251 24197
rect 7193 24188 7205 24191
rect 6840 24160 7205 24188
rect 4172 24092 5764 24120
rect 5810 24080 5816 24132
rect 5868 24080 5874 24132
rect 3970 24012 3976 24064
rect 4028 24052 4034 24064
rect 6840 24052 6868 24160
rect 7193 24157 7205 24160
rect 7239 24157 7251 24191
rect 7193 24151 7251 24157
rect 9306 24148 9312 24200
rect 9364 24148 9370 24200
rect 12360 24197 12388 24228
rect 12805 24225 12817 24259
rect 12851 24225 12863 24259
rect 14108 24256 14136 24355
rect 18138 24352 18144 24404
rect 18196 24352 18202 24404
rect 18248 24364 18736 24392
rect 15565 24327 15623 24333
rect 15565 24293 15577 24327
rect 15611 24324 15623 24327
rect 16390 24324 16396 24336
rect 15611 24296 16396 24324
rect 15611 24293 15623 24296
rect 15565 24287 15623 24293
rect 16390 24284 16396 24296
rect 16448 24284 16454 24336
rect 18248 24324 18276 24364
rect 17604 24296 18276 24324
rect 18708 24324 18736 24364
rect 18782 24352 18788 24404
rect 18840 24392 18846 24404
rect 19978 24392 19984 24404
rect 18840 24364 19984 24392
rect 18840 24352 18846 24364
rect 19978 24352 19984 24364
rect 20036 24352 20042 24404
rect 20070 24352 20076 24404
rect 20128 24392 20134 24404
rect 22370 24392 22376 24404
rect 20128 24364 22376 24392
rect 20128 24352 20134 24364
rect 22370 24352 22376 24364
rect 22428 24392 22434 24404
rect 22428 24364 25268 24392
rect 22428 24352 22434 24364
rect 18708 24296 22094 24324
rect 16025 24259 16083 24265
rect 16025 24256 16037 24259
rect 14108 24228 16037 24256
rect 12805 24219 12863 24225
rect 16025 24225 16037 24228
rect 16071 24225 16083 24259
rect 16025 24219 16083 24225
rect 16114 24216 16120 24268
rect 16172 24216 16178 24268
rect 17604 24265 17632 24296
rect 17589 24259 17647 24265
rect 16868 24228 17540 24256
rect 9769 24191 9827 24197
rect 9769 24157 9781 24191
rect 9815 24157 9827 24191
rect 9769 24151 9827 24157
rect 11885 24191 11943 24197
rect 11885 24157 11897 24191
rect 11931 24157 11943 24191
rect 11885 24151 11943 24157
rect 12345 24191 12403 24197
rect 12345 24157 12357 24191
rect 12391 24157 12403 24191
rect 12345 24151 12403 24157
rect 14461 24191 14519 24197
rect 14461 24157 14473 24191
rect 14507 24188 14519 24191
rect 15654 24188 15660 24200
rect 14507 24160 15660 24188
rect 14507 24157 14519 24160
rect 14461 24151 14519 24157
rect 9784 24120 9812 24151
rect 8496 24092 9812 24120
rect 11900 24120 11928 24151
rect 15654 24148 15660 24160
rect 15712 24148 15718 24200
rect 15933 24191 15991 24197
rect 15933 24157 15945 24191
rect 15979 24188 15991 24191
rect 16868 24188 16896 24228
rect 15979 24160 16896 24188
rect 15979 24157 15991 24160
rect 15933 24151 15991 24157
rect 16942 24148 16948 24200
rect 17000 24188 17006 24200
rect 17313 24191 17371 24197
rect 17313 24188 17325 24191
rect 17000 24160 17325 24188
rect 17000 24148 17006 24160
rect 17313 24157 17325 24160
rect 17359 24157 17371 24191
rect 17512 24188 17540 24228
rect 17589 24225 17601 24259
rect 17635 24225 17647 24259
rect 17589 24219 17647 24225
rect 17770 24216 17776 24268
rect 17828 24256 17834 24268
rect 18690 24256 18696 24268
rect 17828 24228 18696 24256
rect 17828 24216 17834 24228
rect 18690 24216 18696 24228
rect 18748 24216 18754 24268
rect 18782 24216 18788 24268
rect 18840 24216 18846 24268
rect 19978 24216 19984 24268
rect 20036 24256 20042 24268
rect 21269 24259 21327 24265
rect 21269 24256 21281 24259
rect 20036 24228 21281 24256
rect 20036 24216 20042 24228
rect 21269 24225 21281 24228
rect 21315 24225 21327 24259
rect 22066 24256 22094 24296
rect 22554 24256 22560 24268
rect 22066 24228 22560 24256
rect 21269 24219 21327 24225
rect 22554 24216 22560 24228
rect 22612 24216 22618 24268
rect 25038 24216 25044 24268
rect 25096 24216 25102 24268
rect 25133 24259 25191 24265
rect 25133 24225 25145 24259
rect 25179 24225 25191 24259
rect 25133 24219 25191 24225
rect 20070 24188 20076 24200
rect 17512 24160 20076 24188
rect 17313 24151 17371 24157
rect 20070 24148 20076 24160
rect 20128 24148 20134 24200
rect 20165 24191 20223 24197
rect 20165 24157 20177 24191
rect 20211 24157 20223 24191
rect 20165 24151 20223 24157
rect 14642 24120 14648 24132
rect 11900 24092 14648 24120
rect 4028 24024 6868 24052
rect 4028 24012 4034 24024
rect 7466 24012 7472 24064
rect 7524 24052 7530 24064
rect 8496 24052 8524 24092
rect 14642 24080 14648 24092
rect 14700 24080 14706 24132
rect 15105 24123 15163 24129
rect 15105 24089 15117 24123
rect 15151 24120 15163 24123
rect 20180 24120 20208 24151
rect 22278 24148 22284 24200
rect 22336 24148 22342 24200
rect 23842 24148 23848 24200
rect 23900 24188 23906 24200
rect 25148 24188 25176 24219
rect 23900 24160 25176 24188
rect 23900 24148 23906 24160
rect 15151 24092 20208 24120
rect 15151 24089 15163 24092
rect 15105 24083 15163 24089
rect 20254 24080 20260 24132
rect 20312 24120 20318 24132
rect 20533 24123 20591 24129
rect 20533 24120 20545 24123
rect 20312 24092 20545 24120
rect 20312 24080 20318 24092
rect 20533 24089 20545 24092
rect 20579 24089 20591 24123
rect 20533 24083 20591 24089
rect 22557 24123 22615 24129
rect 22557 24089 22569 24123
rect 22603 24089 22615 24123
rect 25038 24120 25044 24132
rect 23782 24092 23980 24120
rect 22557 24083 22615 24089
rect 7524 24024 8524 24052
rect 7524 24012 7530 24024
rect 9122 24012 9128 24064
rect 9180 24012 9186 24064
rect 11330 24012 11336 24064
rect 11388 24052 11394 24064
rect 16850 24052 16856 24064
rect 11388 24024 16856 24052
rect 11388 24012 11394 24024
rect 16850 24012 16856 24024
rect 16908 24012 16914 24064
rect 16945 24055 17003 24061
rect 16945 24021 16957 24055
rect 16991 24052 17003 24055
rect 17034 24052 17040 24064
rect 16991 24024 17040 24052
rect 16991 24021 17003 24024
rect 16945 24015 17003 24021
rect 17034 24012 17040 24024
rect 17092 24012 17098 24064
rect 17405 24055 17463 24061
rect 17405 24021 17417 24055
rect 17451 24052 17463 24055
rect 17770 24052 17776 24064
rect 17451 24024 17776 24052
rect 17451 24021 17463 24024
rect 17405 24015 17463 24021
rect 17770 24012 17776 24024
rect 17828 24012 17834 24064
rect 17954 24012 17960 24064
rect 18012 24052 18018 24064
rect 18509 24055 18567 24061
rect 18509 24052 18521 24055
rect 18012 24024 18521 24052
rect 18012 24012 18018 24024
rect 18509 24021 18521 24024
rect 18555 24021 18567 24055
rect 18509 24015 18567 24021
rect 18601 24055 18659 24061
rect 18601 24021 18613 24055
rect 18647 24052 18659 24055
rect 19242 24052 19248 24064
rect 18647 24024 19248 24052
rect 18647 24021 18659 24024
rect 18601 24015 18659 24021
rect 19242 24012 19248 24024
rect 19300 24012 19306 24064
rect 19334 24012 19340 24064
rect 19392 24052 19398 24064
rect 19429 24055 19487 24061
rect 19429 24052 19441 24055
rect 19392 24024 19441 24052
rect 19392 24012 19398 24024
rect 19429 24021 19441 24024
rect 19475 24021 19487 24055
rect 19429 24015 19487 24021
rect 20990 24012 20996 24064
rect 21048 24052 21054 24064
rect 21085 24055 21143 24061
rect 21085 24052 21097 24055
rect 21048 24024 21097 24052
rect 21048 24012 21054 24024
rect 21085 24021 21097 24024
rect 21131 24021 21143 24055
rect 21085 24015 21143 24021
rect 21358 24012 21364 24064
rect 21416 24052 21422 24064
rect 21453 24055 21511 24061
rect 21453 24052 21465 24055
rect 21416 24024 21465 24052
rect 21416 24012 21422 24024
rect 21453 24021 21465 24024
rect 21499 24021 21511 24055
rect 21453 24015 21511 24021
rect 21818 24012 21824 24064
rect 21876 24052 21882 24064
rect 21913 24055 21971 24061
rect 21913 24052 21925 24055
rect 21876 24024 21925 24052
rect 21876 24012 21882 24024
rect 21913 24021 21925 24024
rect 21959 24021 21971 24055
rect 22572 24052 22600 24083
rect 23952 24064 23980 24092
rect 24596 24092 25044 24120
rect 23566 24052 23572 24064
rect 22572 24024 23572 24052
rect 21913 24015 21971 24021
rect 23566 24012 23572 24024
rect 23624 24012 23630 24064
rect 23934 24012 23940 24064
rect 23992 24012 23998 24064
rect 24029 24055 24087 24061
rect 24029 24021 24041 24055
rect 24075 24052 24087 24055
rect 24118 24052 24124 24064
rect 24075 24024 24124 24052
rect 24075 24021 24087 24024
rect 24029 24015 24087 24021
rect 24118 24012 24124 24024
rect 24176 24012 24182 24064
rect 24596 24061 24624 24092
rect 25038 24080 25044 24092
rect 25096 24080 25102 24132
rect 24581 24055 24639 24061
rect 24581 24021 24593 24055
rect 24627 24021 24639 24055
rect 24581 24015 24639 24021
rect 24949 24055 25007 24061
rect 24949 24021 24961 24055
rect 24995 24052 25007 24055
rect 25240 24052 25268 24364
rect 24995 24024 25268 24052
rect 24995 24021 25007 24024
rect 24949 24015 25007 24021
rect 1104 23962 25852 23984
rect 1104 23910 7950 23962
rect 8002 23910 8014 23962
rect 8066 23910 8078 23962
rect 8130 23910 8142 23962
rect 8194 23910 8206 23962
rect 8258 23910 17950 23962
rect 18002 23910 18014 23962
rect 18066 23910 18078 23962
rect 18130 23910 18142 23962
rect 18194 23910 18206 23962
rect 18258 23910 25852 23962
rect 1104 23888 25852 23910
rect 4890 23808 4896 23860
rect 4948 23848 4954 23860
rect 4948 23820 7972 23848
rect 4948 23808 4954 23820
rect 3973 23783 4031 23789
rect 3973 23749 3985 23783
rect 4019 23780 4031 23783
rect 5350 23780 5356 23792
rect 4019 23752 5356 23780
rect 4019 23749 4031 23752
rect 3973 23743 4031 23749
rect 5350 23740 5356 23752
rect 5408 23740 5414 23792
rect 5813 23783 5871 23789
rect 5813 23749 5825 23783
rect 5859 23780 5871 23783
rect 7374 23780 7380 23792
rect 5859 23752 7380 23780
rect 5859 23749 5871 23752
rect 5813 23743 5871 23749
rect 7374 23740 7380 23752
rect 7432 23740 7438 23792
rect 1118 23672 1124 23724
rect 1176 23712 1182 23724
rect 1486 23712 1492 23724
rect 1176 23684 1492 23712
rect 1176 23672 1182 23684
rect 1486 23672 1492 23684
rect 1544 23712 1550 23724
rect 1673 23715 1731 23721
rect 1673 23712 1685 23715
rect 1544 23684 1685 23712
rect 1544 23672 1550 23684
rect 1673 23681 1685 23684
rect 1719 23681 1731 23715
rect 1673 23675 1731 23681
rect 2961 23715 3019 23721
rect 2961 23681 2973 23715
rect 3007 23712 3019 23715
rect 3786 23712 3792 23724
rect 3007 23684 3792 23712
rect 3007 23681 3019 23684
rect 2961 23675 3019 23681
rect 3786 23672 3792 23684
rect 3844 23672 3850 23724
rect 7944 23721 7972 23820
rect 9306 23808 9312 23860
rect 9364 23848 9370 23860
rect 11514 23848 11520 23860
rect 9364 23820 11520 23848
rect 9364 23808 9370 23820
rect 11514 23808 11520 23820
rect 11572 23808 11578 23860
rect 13725 23851 13783 23857
rect 13725 23848 13737 23851
rect 11716 23820 13737 23848
rect 9125 23783 9183 23789
rect 9125 23749 9137 23783
rect 9171 23780 9183 23783
rect 10134 23780 10140 23792
rect 9171 23752 10140 23780
rect 9171 23749 9183 23752
rect 9125 23743 9183 23749
rect 10134 23740 10140 23752
rect 10192 23740 10198 23792
rect 10870 23740 10876 23792
rect 10928 23740 10934 23792
rect 11716 23789 11744 23820
rect 13725 23817 13737 23820
rect 13771 23848 13783 23851
rect 13998 23848 14004 23860
rect 13771 23820 14004 23848
rect 13771 23817 13783 23820
rect 13725 23811 13783 23817
rect 13998 23808 14004 23820
rect 14056 23808 14062 23860
rect 14090 23808 14096 23860
rect 14148 23808 14154 23860
rect 14461 23851 14519 23857
rect 14461 23817 14473 23851
rect 14507 23848 14519 23851
rect 15562 23848 15568 23860
rect 14507 23820 15568 23848
rect 14507 23817 14519 23820
rect 14461 23811 14519 23817
rect 15562 23808 15568 23820
rect 15620 23808 15626 23860
rect 15746 23808 15752 23860
rect 15804 23848 15810 23860
rect 16025 23851 16083 23857
rect 16025 23848 16037 23851
rect 15804 23820 16037 23848
rect 15804 23808 15810 23820
rect 16025 23817 16037 23820
rect 16071 23817 16083 23851
rect 16025 23811 16083 23817
rect 16574 23808 16580 23860
rect 16632 23848 16638 23860
rect 19334 23848 19340 23860
rect 16632 23820 19340 23848
rect 16632 23808 16638 23820
rect 19334 23808 19340 23820
rect 19392 23808 19398 23860
rect 20070 23808 20076 23860
rect 20128 23848 20134 23860
rect 20855 23851 20913 23857
rect 20855 23848 20867 23851
rect 20128 23820 20867 23848
rect 20128 23808 20134 23820
rect 20855 23817 20867 23820
rect 20901 23817 20913 23851
rect 20855 23811 20913 23817
rect 22278 23808 22284 23860
rect 22336 23848 22342 23860
rect 23290 23848 23296 23860
rect 22336 23820 23296 23848
rect 22336 23808 22342 23820
rect 23290 23808 23296 23820
rect 23348 23808 23354 23860
rect 11701 23783 11759 23789
rect 11701 23780 11713 23783
rect 11164 23752 11713 23780
rect 4801 23715 4859 23721
rect 4801 23681 4813 23715
rect 4847 23712 4859 23715
rect 7929 23715 7987 23721
rect 4847 23684 7880 23712
rect 4847 23681 4859 23684
rect 4801 23675 4859 23681
rect 6549 23647 6607 23653
rect 6549 23613 6561 23647
rect 6595 23613 6607 23647
rect 6549 23607 6607 23613
rect 6825 23647 6883 23653
rect 6825 23613 6837 23647
rect 6871 23644 6883 23647
rect 7558 23644 7564 23656
rect 6871 23616 7564 23644
rect 6871 23613 6883 23616
rect 6825 23607 6883 23613
rect 1857 23579 1915 23585
rect 1857 23545 1869 23579
rect 1903 23576 1915 23579
rect 6454 23576 6460 23588
rect 1903 23548 6460 23576
rect 1903 23545 1915 23548
rect 1857 23539 1915 23545
rect 6454 23536 6460 23548
rect 6512 23536 6518 23588
rect 6564 23576 6592 23607
rect 7558 23604 7564 23616
rect 7616 23604 7622 23656
rect 7852 23644 7880 23684
rect 7929 23681 7941 23715
rect 7975 23681 7987 23715
rect 7929 23675 7987 23681
rect 8570 23672 8576 23724
rect 8628 23712 8634 23724
rect 9769 23715 9827 23721
rect 9769 23712 9781 23715
rect 8628 23684 9781 23712
rect 8628 23672 8634 23684
rect 9769 23681 9781 23684
rect 9815 23681 9827 23715
rect 9769 23675 9827 23681
rect 9950 23672 9956 23724
rect 10008 23712 10014 23724
rect 11164 23712 11192 23752
rect 11701 23749 11713 23752
rect 11747 23749 11759 23783
rect 11701 23743 11759 23749
rect 11882 23740 11888 23792
rect 11940 23780 11946 23792
rect 18414 23780 18420 23792
rect 11940 23752 18420 23780
rect 11940 23740 11946 23752
rect 18414 23740 18420 23752
rect 18472 23740 18478 23792
rect 18966 23740 18972 23792
rect 19024 23740 19030 23792
rect 19610 23740 19616 23792
rect 19668 23780 19674 23792
rect 22094 23780 22100 23792
rect 19668 23752 22100 23780
rect 19668 23740 19674 23752
rect 22094 23740 22100 23752
rect 22152 23740 22158 23792
rect 12069 23715 12127 23721
rect 12069 23712 12081 23715
rect 10008 23684 11192 23712
rect 11256 23684 12081 23712
rect 10008 23672 10014 23684
rect 11054 23644 11060 23656
rect 7852 23616 11060 23644
rect 11054 23604 11060 23616
rect 11112 23604 11118 23656
rect 7374 23576 7380 23588
rect 6564 23548 7380 23576
rect 7374 23536 7380 23548
rect 7432 23536 7438 23588
rect 2317 23511 2375 23517
rect 2317 23477 2329 23511
rect 2363 23508 2375 23511
rect 2409 23511 2467 23517
rect 2409 23508 2421 23511
rect 2363 23480 2421 23508
rect 2363 23477 2375 23480
rect 2317 23471 2375 23477
rect 2409 23477 2421 23480
rect 2455 23508 2467 23511
rect 7098 23508 7104 23520
rect 2455 23480 7104 23508
rect 2455 23477 2467 23480
rect 2409 23471 2467 23477
rect 7098 23468 7104 23480
rect 7156 23468 7162 23520
rect 9490 23468 9496 23520
rect 9548 23508 9554 23520
rect 11256 23508 11284 23684
rect 12069 23681 12081 23684
rect 12115 23681 12127 23715
rect 12069 23675 12127 23681
rect 14553 23715 14611 23721
rect 14553 23681 14565 23715
rect 14599 23712 14611 23715
rect 15194 23712 15200 23724
rect 14599 23684 15200 23712
rect 14599 23681 14611 23684
rect 14553 23675 14611 23681
rect 15194 23672 15200 23684
rect 15252 23672 15258 23724
rect 15933 23715 15991 23721
rect 15933 23681 15945 23715
rect 15979 23681 15991 23715
rect 15933 23675 15991 23681
rect 17221 23715 17279 23721
rect 17221 23681 17233 23715
rect 17267 23712 17279 23715
rect 17770 23712 17776 23724
rect 17267 23684 17776 23712
rect 17267 23681 17279 23684
rect 17221 23675 17279 23681
rect 11974 23604 11980 23656
rect 12032 23644 12038 23656
rect 12529 23647 12587 23653
rect 12529 23644 12541 23647
rect 12032 23616 12541 23644
rect 12032 23604 12038 23616
rect 12529 23613 12541 23616
rect 12575 23613 12587 23647
rect 12529 23607 12587 23613
rect 14734 23604 14740 23656
rect 14792 23604 14798 23656
rect 15470 23604 15476 23656
rect 15528 23644 15534 23656
rect 15746 23644 15752 23656
rect 15528 23616 15752 23644
rect 15528 23604 15534 23616
rect 15746 23604 15752 23616
rect 15804 23604 15810 23656
rect 11514 23536 11520 23588
rect 11572 23576 11578 23588
rect 14550 23576 14556 23588
rect 11572 23548 14556 23576
rect 11572 23536 11578 23548
rect 14550 23536 14556 23548
rect 14608 23536 14614 23588
rect 15289 23579 15347 23585
rect 15289 23545 15301 23579
rect 15335 23576 15347 23579
rect 15654 23576 15660 23588
rect 15335 23548 15660 23576
rect 15335 23545 15347 23548
rect 15289 23539 15347 23545
rect 15654 23536 15660 23548
rect 15712 23536 15718 23588
rect 15838 23536 15844 23588
rect 15896 23576 15902 23588
rect 15948 23576 15976 23675
rect 17770 23672 17776 23684
rect 17828 23672 17834 23724
rect 22296 23721 22324 23808
rect 24026 23780 24032 23792
rect 23782 23752 24032 23780
rect 24026 23740 24032 23752
rect 24084 23780 24090 23792
rect 24305 23783 24363 23789
rect 24305 23780 24317 23783
rect 24084 23752 24317 23780
rect 24084 23740 24090 23752
rect 24305 23749 24317 23752
rect 24351 23780 24363 23783
rect 24673 23783 24731 23789
rect 24673 23780 24685 23783
rect 24351 23752 24685 23780
rect 24351 23749 24363 23752
rect 24305 23743 24363 23749
rect 24673 23749 24685 23752
rect 24719 23749 24731 23783
rect 24673 23743 24731 23749
rect 24949 23783 25007 23789
rect 24949 23749 24961 23783
rect 24995 23780 25007 23783
rect 25130 23780 25136 23792
rect 24995 23752 25136 23780
rect 24995 23749 25007 23752
rect 24949 23743 25007 23749
rect 25130 23740 25136 23752
rect 25188 23740 25194 23792
rect 22281 23715 22339 23721
rect 22281 23681 22293 23715
rect 22327 23681 22339 23715
rect 22281 23675 22339 23681
rect 16209 23647 16267 23653
rect 16209 23613 16221 23647
rect 16255 23644 16267 23647
rect 16298 23644 16304 23656
rect 16255 23616 16304 23644
rect 16255 23613 16267 23616
rect 16209 23607 16267 23613
rect 16298 23604 16304 23616
rect 16356 23604 16362 23656
rect 17310 23604 17316 23656
rect 17368 23604 17374 23656
rect 17497 23647 17555 23653
rect 17497 23613 17509 23647
rect 17543 23613 17555 23647
rect 17497 23607 17555 23613
rect 15896 23548 15976 23576
rect 15896 23536 15902 23548
rect 9548 23480 11284 23508
rect 9548 23468 9554 23480
rect 11698 23468 11704 23520
rect 11756 23508 11762 23520
rect 14918 23508 14924 23520
rect 11756 23480 14924 23508
rect 11756 23468 11762 23480
rect 14918 23468 14924 23480
rect 14976 23468 14982 23520
rect 15565 23511 15623 23517
rect 15565 23477 15577 23511
rect 15611 23508 15623 23511
rect 16758 23508 16764 23520
rect 15611 23480 16764 23508
rect 15611 23477 15623 23480
rect 15565 23471 15623 23477
rect 16758 23468 16764 23480
rect 16816 23468 16822 23520
rect 16850 23468 16856 23520
rect 16908 23468 16914 23520
rect 17512 23508 17540 23607
rect 18046 23604 18052 23656
rect 18104 23604 18110 23656
rect 18325 23647 18383 23653
rect 18325 23644 18337 23647
rect 18156 23616 18337 23644
rect 17954 23536 17960 23588
rect 18012 23576 18018 23588
rect 18156 23576 18184 23616
rect 18325 23613 18337 23616
rect 18371 23613 18383 23647
rect 18325 23607 18383 23613
rect 18414 23604 18420 23656
rect 18472 23644 18478 23656
rect 19334 23644 19340 23656
rect 18472 23616 19340 23644
rect 18472 23604 18478 23616
rect 19334 23604 19340 23616
rect 19392 23604 19398 23656
rect 20622 23604 20628 23656
rect 20680 23604 20686 23656
rect 22554 23604 22560 23656
rect 22612 23604 22618 23656
rect 24302 23604 24308 23656
rect 24360 23644 24366 23656
rect 24489 23647 24547 23653
rect 24489 23644 24501 23647
rect 24360 23616 24501 23644
rect 24360 23604 24366 23616
rect 24489 23613 24501 23616
rect 24535 23613 24547 23647
rect 24489 23607 24547 23613
rect 18012 23548 18184 23576
rect 19720 23548 21956 23576
rect 18012 23536 18018 23548
rect 19720 23508 19748 23548
rect 17512 23480 19748 23508
rect 19794 23468 19800 23520
rect 19852 23468 19858 23520
rect 19886 23468 19892 23520
rect 19944 23508 19950 23520
rect 20073 23511 20131 23517
rect 20073 23508 20085 23511
rect 19944 23480 20085 23508
rect 19944 23468 19950 23480
rect 20073 23477 20085 23480
rect 20119 23508 20131 23511
rect 20257 23511 20315 23517
rect 20257 23508 20269 23511
rect 20119 23480 20269 23508
rect 20119 23477 20131 23480
rect 20073 23471 20131 23477
rect 20257 23477 20269 23480
rect 20303 23477 20315 23511
rect 20257 23471 20315 23477
rect 20438 23468 20444 23520
rect 20496 23508 20502 23520
rect 21821 23511 21879 23517
rect 21821 23508 21833 23511
rect 20496 23480 21833 23508
rect 20496 23468 20502 23480
rect 21821 23477 21833 23480
rect 21867 23477 21879 23511
rect 21928 23508 21956 23548
rect 23566 23536 23572 23588
rect 23624 23576 23630 23588
rect 24029 23579 24087 23585
rect 24029 23576 24041 23579
rect 23624 23548 24041 23576
rect 23624 23536 23630 23548
rect 24029 23545 24041 23548
rect 24075 23576 24087 23579
rect 25406 23576 25412 23588
rect 24075 23548 25412 23576
rect 24075 23545 24087 23548
rect 24029 23539 24087 23545
rect 25406 23536 25412 23548
rect 25464 23536 25470 23588
rect 24118 23508 24124 23520
rect 21928 23480 24124 23508
rect 21821 23471 21879 23477
rect 24118 23468 24124 23480
rect 24176 23468 24182 23520
rect 25130 23468 25136 23520
rect 25188 23508 25194 23520
rect 25225 23511 25283 23517
rect 25225 23508 25237 23511
rect 25188 23480 25237 23508
rect 25188 23468 25194 23480
rect 25225 23477 25237 23480
rect 25271 23477 25283 23511
rect 25225 23471 25283 23477
rect 1104 23418 25852 23440
rect 1104 23366 2950 23418
rect 3002 23366 3014 23418
rect 3066 23366 3078 23418
rect 3130 23366 3142 23418
rect 3194 23366 3206 23418
rect 3258 23366 12950 23418
rect 13002 23366 13014 23418
rect 13066 23366 13078 23418
rect 13130 23366 13142 23418
rect 13194 23366 13206 23418
rect 13258 23366 22950 23418
rect 23002 23366 23014 23418
rect 23066 23366 23078 23418
rect 23130 23366 23142 23418
rect 23194 23366 23206 23418
rect 23258 23366 25852 23418
rect 1104 23344 25852 23366
rect 1486 23264 1492 23316
rect 1544 23264 1550 23316
rect 1765 23307 1823 23313
rect 1765 23273 1777 23307
rect 1811 23304 1823 23307
rect 6730 23304 6736 23316
rect 1811 23276 6736 23304
rect 1811 23273 1823 23276
rect 1765 23267 1823 23273
rect 6730 23264 6736 23276
rect 6788 23264 6794 23316
rect 7374 23264 7380 23316
rect 7432 23304 7438 23316
rect 11974 23304 11980 23316
rect 7432 23276 11980 23304
rect 7432 23264 7438 23276
rect 11974 23264 11980 23276
rect 12032 23264 12038 23316
rect 12342 23264 12348 23316
rect 12400 23304 12406 23316
rect 12434 23304 12440 23316
rect 12400 23276 12440 23304
rect 12400 23264 12406 23276
rect 12434 23264 12440 23276
rect 12492 23264 12498 23316
rect 12894 23264 12900 23316
rect 12952 23304 12958 23316
rect 13814 23304 13820 23316
rect 12952 23276 13820 23304
rect 12952 23264 12958 23276
rect 13814 23264 13820 23276
rect 13872 23264 13878 23316
rect 13906 23264 13912 23316
rect 13964 23304 13970 23316
rect 16482 23304 16488 23316
rect 13964 23276 16488 23304
rect 13964 23264 13970 23276
rect 16482 23264 16488 23276
rect 16540 23264 16546 23316
rect 16574 23264 16580 23316
rect 16632 23304 16638 23316
rect 16761 23307 16819 23313
rect 16761 23304 16773 23307
rect 16632 23276 16773 23304
rect 16632 23264 16638 23276
rect 16761 23273 16773 23276
rect 16807 23304 16819 23307
rect 17678 23304 17684 23316
rect 16807 23276 17684 23304
rect 16807 23273 16819 23276
rect 16761 23267 16819 23273
rect 17678 23264 17684 23276
rect 17736 23264 17742 23316
rect 17954 23264 17960 23316
rect 18012 23304 18018 23316
rect 18782 23304 18788 23316
rect 18012 23276 18788 23304
rect 18012 23264 18018 23276
rect 18782 23264 18788 23276
rect 18840 23304 18846 23316
rect 21177 23307 21235 23313
rect 21177 23304 21189 23307
rect 18840 23276 21189 23304
rect 18840 23264 18846 23276
rect 21177 23273 21189 23276
rect 21223 23273 21235 23307
rect 21177 23267 21235 23273
rect 22554 23264 22560 23316
rect 22612 23304 22618 23316
rect 23385 23307 23443 23313
rect 23385 23304 23397 23307
rect 22612 23276 23397 23304
rect 22612 23264 22618 23276
rect 23385 23273 23397 23276
rect 23431 23273 23443 23307
rect 23385 23267 23443 23273
rect 9398 23236 9404 23248
rect 8312 23208 9404 23236
rect 3237 23171 3295 23177
rect 3237 23137 3249 23171
rect 3283 23168 3295 23171
rect 4614 23168 4620 23180
rect 3283 23140 4620 23168
rect 3283 23137 3295 23140
rect 3237 23131 3295 23137
rect 4614 23128 4620 23140
rect 4672 23128 4678 23180
rect 6549 23171 6607 23177
rect 6549 23137 6561 23171
rect 6595 23168 6607 23171
rect 7650 23168 7656 23180
rect 6595 23140 7656 23168
rect 6595 23137 6607 23140
rect 6549 23131 6607 23137
rect 7650 23128 7656 23140
rect 7708 23128 7714 23180
rect 8312 23177 8340 23208
rect 9398 23196 9404 23208
rect 9456 23196 9462 23248
rect 11698 23236 11704 23248
rect 9508 23208 11704 23236
rect 8297 23171 8355 23177
rect 8297 23137 8309 23171
rect 8343 23137 8355 23171
rect 8297 23131 8355 23137
rect 8570 23128 8576 23180
rect 8628 23168 8634 23180
rect 9508 23168 9536 23208
rect 11698 23196 11704 23208
rect 11756 23196 11762 23248
rect 13538 23196 13544 23248
rect 13596 23196 13602 23248
rect 17126 23196 17132 23248
rect 17184 23236 17190 23248
rect 18874 23236 18880 23248
rect 17184 23208 18880 23236
rect 17184 23196 17190 23208
rect 18874 23196 18880 23208
rect 18932 23196 18938 23248
rect 18966 23196 18972 23248
rect 19024 23236 19030 23248
rect 19426 23236 19432 23248
rect 19024 23208 19432 23236
rect 19024 23196 19030 23208
rect 19426 23196 19432 23208
rect 19484 23196 19490 23248
rect 8628 23140 9536 23168
rect 8628 23128 8634 23140
rect 10502 23128 10508 23180
rect 10560 23128 10566 23180
rect 11606 23128 11612 23180
rect 11664 23168 11670 23180
rect 12161 23171 12219 23177
rect 12161 23168 12173 23171
rect 11664 23140 12173 23168
rect 11664 23128 11670 23140
rect 12161 23137 12173 23140
rect 12207 23137 12219 23171
rect 14182 23168 14188 23180
rect 12161 23131 12219 23137
rect 12636 23140 14188 23168
rect 2222 23060 2228 23112
rect 2280 23060 2286 23112
rect 3418 23060 3424 23112
rect 3476 23100 3482 23112
rect 4065 23103 4123 23109
rect 4065 23100 4077 23103
rect 3476 23072 4077 23100
rect 3476 23060 3482 23072
rect 4065 23069 4077 23072
rect 4111 23069 4123 23103
rect 4065 23063 4123 23069
rect 5442 23060 5448 23112
rect 5500 23060 5506 23112
rect 7006 23060 7012 23112
rect 7064 23100 7070 23112
rect 7193 23103 7251 23109
rect 7193 23100 7205 23103
rect 7064 23072 7205 23100
rect 7064 23060 7070 23072
rect 7193 23069 7205 23072
rect 7239 23069 7251 23103
rect 9401 23103 9459 23109
rect 9401 23100 9413 23103
rect 7193 23063 7251 23069
rect 7300 23072 9413 23100
rect 4249 23035 4307 23041
rect 4249 23001 4261 23035
rect 4295 23032 4307 23035
rect 5626 23032 5632 23044
rect 4295 23004 5632 23032
rect 4295 23001 4307 23004
rect 4249 22995 4307 23001
rect 5626 22992 5632 23004
rect 5684 22992 5690 23044
rect 6362 22992 6368 23044
rect 6420 23032 6426 23044
rect 7300 23032 7328 23072
rect 9401 23069 9413 23072
rect 9447 23069 9459 23103
rect 9401 23063 9459 23069
rect 9861 23103 9919 23109
rect 9861 23069 9873 23103
rect 9907 23069 9919 23103
rect 9861 23063 9919 23069
rect 11701 23103 11759 23109
rect 11701 23069 11713 23103
rect 11747 23069 11759 23103
rect 11701 23063 11759 23069
rect 6420 23004 7328 23032
rect 6420 22992 6426 23004
rect 7558 22992 7564 23044
rect 7616 23032 7622 23044
rect 9876 23032 9904 23063
rect 7616 23004 9904 23032
rect 7616 22992 7622 23004
rect 4706 22924 4712 22976
rect 4764 22924 4770 22976
rect 9217 22967 9275 22973
rect 9217 22933 9229 22967
rect 9263 22964 9275 22967
rect 11716 22964 11744 23063
rect 11974 22992 11980 23044
rect 12032 23032 12038 23044
rect 12636 23032 12664 23140
rect 14182 23128 14188 23140
rect 14240 23128 14246 23180
rect 15289 23171 15347 23177
rect 15289 23137 15301 23171
rect 15335 23168 15347 23171
rect 17773 23171 17831 23177
rect 17773 23168 17785 23171
rect 15335 23140 17785 23168
rect 15335 23137 15347 23140
rect 15289 23131 15347 23137
rect 17773 23137 17785 23140
rect 17819 23168 17831 23171
rect 18598 23168 18604 23180
rect 17819 23140 18604 23168
rect 17819 23137 17831 23140
rect 17773 23131 17831 23137
rect 18598 23128 18604 23140
rect 18656 23128 18662 23180
rect 18693 23171 18751 23177
rect 18693 23137 18705 23171
rect 18739 23168 18751 23171
rect 19058 23168 19064 23180
rect 18739 23140 19064 23168
rect 18739 23137 18751 23140
rect 18693 23131 18751 23137
rect 19058 23128 19064 23140
rect 19116 23128 19122 23180
rect 19705 23171 19763 23177
rect 19705 23137 19717 23171
rect 19751 23168 19763 23171
rect 20714 23168 20720 23180
rect 19751 23140 20720 23168
rect 19751 23137 19763 23140
rect 19705 23131 19763 23137
rect 20714 23128 20720 23140
rect 20772 23128 20778 23180
rect 21637 23171 21695 23177
rect 21637 23137 21649 23171
rect 21683 23168 21695 23171
rect 22278 23168 22284 23180
rect 21683 23140 22284 23168
rect 21683 23137 21695 23140
rect 21637 23131 21695 23137
rect 22278 23128 22284 23140
rect 22336 23128 22342 23180
rect 24762 23128 24768 23180
rect 24820 23168 24826 23180
rect 25133 23171 25191 23177
rect 25133 23168 25145 23171
rect 24820 23140 25145 23168
rect 24820 23128 24826 23140
rect 25133 23137 25145 23140
rect 25179 23137 25191 23171
rect 25133 23131 25191 23137
rect 12710 23060 12716 23112
rect 12768 23096 12774 23112
rect 13630 23100 13636 23112
rect 12820 23096 13636 23100
rect 12768 23072 13636 23096
rect 12768 23068 12848 23072
rect 12768 23060 12774 23068
rect 13630 23060 13636 23072
rect 13688 23060 13694 23112
rect 13722 23060 13728 23112
rect 13780 23060 13786 23112
rect 13814 23060 13820 23112
rect 13872 23100 13878 23112
rect 15013 23103 15071 23109
rect 15013 23100 15025 23103
rect 13872 23072 15025 23100
rect 13872 23060 13878 23072
rect 15013 23069 15025 23072
rect 15059 23069 15071 23103
rect 15013 23063 15071 23069
rect 16758 23060 16764 23112
rect 16816 23100 16822 23112
rect 17589 23103 17647 23109
rect 17589 23100 17601 23103
rect 16816 23072 17601 23100
rect 16816 23060 16822 23072
rect 17589 23069 17601 23072
rect 17635 23069 17647 23103
rect 17589 23063 17647 23069
rect 18046 23060 18052 23112
rect 18104 23100 18110 23112
rect 19334 23100 19340 23112
rect 18104 23072 19340 23100
rect 18104 23060 18110 23072
rect 19334 23060 19340 23072
rect 19392 23100 19398 23112
rect 19429 23103 19487 23109
rect 19429 23100 19441 23103
rect 19392 23072 19441 23100
rect 19392 23060 19398 23072
rect 19429 23069 19441 23072
rect 19475 23069 19487 23103
rect 19429 23063 19487 23069
rect 12032 23004 12664 23032
rect 12032 22992 12038 23004
rect 12986 22992 12992 23044
rect 13044 23032 13050 23044
rect 14369 23035 14427 23041
rect 14369 23032 14381 23035
rect 13044 23004 14381 23032
rect 13044 22992 13050 23004
rect 14369 23001 14381 23004
rect 14415 23001 14427 23035
rect 14369 22995 14427 23001
rect 14550 22992 14556 23044
rect 14608 23032 14614 23044
rect 15562 23032 15568 23044
rect 14608 23004 15568 23032
rect 14608 22992 14614 23004
rect 15562 22992 15568 23004
rect 15620 23032 15626 23044
rect 18506 23041 18512 23044
rect 17681 23035 17739 23041
rect 17681 23032 17693 23035
rect 15620 23004 15778 23032
rect 16592 23004 17693 23032
rect 15620 22992 15626 23004
rect 9263 22936 11744 22964
rect 9263 22933 9275 22936
rect 9217 22927 9275 22933
rect 11882 22924 11888 22976
rect 11940 22964 11946 22976
rect 14461 22967 14519 22973
rect 14461 22964 14473 22967
rect 11940 22936 14473 22964
rect 11940 22924 11946 22936
rect 14461 22933 14473 22936
rect 14507 22933 14519 22967
rect 14461 22927 14519 22933
rect 15010 22924 15016 22976
rect 15068 22964 15074 22976
rect 16592 22964 16620 23004
rect 17681 23001 17693 23004
rect 17727 23001 17739 23035
rect 17681 22995 17739 23001
rect 18473 23035 18512 23041
rect 18473 23001 18485 23035
rect 18473 22995 18512 23001
rect 18506 22992 18512 22995
rect 18564 22992 18570 23044
rect 18690 22992 18696 23044
rect 18748 23032 18754 23044
rect 18966 23032 18972 23044
rect 18748 23004 18972 23032
rect 18748 22992 18754 23004
rect 18966 22992 18972 23004
rect 19024 22992 19030 23044
rect 19150 22992 19156 23044
rect 19208 23032 19214 23044
rect 19208 23004 19472 23032
rect 19208 22992 19214 23004
rect 15068 22936 16620 22964
rect 15068 22924 15074 22936
rect 16758 22924 16764 22976
rect 16816 22964 16822 22976
rect 17221 22967 17279 22973
rect 17221 22964 17233 22967
rect 16816 22936 17233 22964
rect 16816 22924 16822 22936
rect 17221 22933 17233 22936
rect 17267 22933 17279 22967
rect 17221 22927 17279 22933
rect 17310 22924 17316 22976
rect 17368 22964 17374 22976
rect 18046 22964 18052 22976
rect 17368 22936 18052 22964
rect 17368 22924 17374 22936
rect 18046 22924 18052 22936
rect 18104 22924 18110 22976
rect 19058 22924 19064 22976
rect 19116 22924 19122 22976
rect 19444 22964 19472 23004
rect 19978 22992 19984 23044
rect 20036 23032 20042 23044
rect 21913 23035 21971 23041
rect 20036 23004 20194 23032
rect 20036 22992 20042 23004
rect 21913 23001 21925 23035
rect 21959 23032 21971 23035
rect 22186 23032 22192 23044
rect 21959 23004 22192 23032
rect 21959 23001 21971 23004
rect 21913 22995 21971 23001
rect 22186 22992 22192 23004
rect 22244 22992 22250 23044
rect 22370 22992 22376 23044
rect 22428 22992 22434 23044
rect 25041 23035 25099 23041
rect 25041 23032 25053 23035
rect 23308 23004 25053 23032
rect 23308 22964 23336 23004
rect 25041 23001 25053 23004
rect 25087 23001 25099 23035
rect 25041 22995 25099 23001
rect 19444 22936 23336 22964
rect 23845 22967 23903 22973
rect 23845 22933 23857 22967
rect 23891 22964 23903 22967
rect 23934 22964 23940 22976
rect 23891 22936 23940 22964
rect 23891 22933 23903 22936
rect 23845 22927 23903 22933
rect 23934 22924 23940 22936
rect 23992 22924 23998 22976
rect 24578 22924 24584 22976
rect 24636 22924 24642 22976
rect 24946 22924 24952 22976
rect 25004 22924 25010 22976
rect 1104 22874 25852 22896
rect 1104 22822 7950 22874
rect 8002 22822 8014 22874
rect 8066 22822 8078 22874
rect 8130 22822 8142 22874
rect 8194 22822 8206 22874
rect 8258 22822 17950 22874
rect 18002 22822 18014 22874
rect 18066 22822 18078 22874
rect 18130 22822 18142 22874
rect 18194 22822 18206 22874
rect 18258 22822 25852 22874
rect 1104 22800 25852 22822
rect 2222 22720 2228 22772
rect 2280 22760 2286 22772
rect 2280 22732 4660 22760
rect 2280 22720 2286 22732
rect 2317 22695 2375 22701
rect 2317 22661 2329 22695
rect 2363 22692 2375 22695
rect 3418 22692 3424 22704
rect 2363 22664 3424 22692
rect 2363 22661 2375 22664
rect 2317 22655 2375 22661
rect 3418 22652 3424 22664
rect 3476 22652 3482 22704
rect 3973 22695 4031 22701
rect 3973 22661 3985 22695
rect 4019 22692 4031 22695
rect 4246 22692 4252 22704
rect 4019 22664 4252 22692
rect 4019 22661 4031 22664
rect 3973 22655 4031 22661
rect 4246 22652 4252 22664
rect 4304 22652 4310 22704
rect 4632 22692 4660 22732
rect 4706 22720 4712 22772
rect 4764 22760 4770 22772
rect 12069 22763 12127 22769
rect 12069 22760 12081 22763
rect 4764 22732 12081 22760
rect 4764 22720 4770 22732
rect 12069 22729 12081 22732
rect 12115 22729 12127 22763
rect 13081 22763 13139 22769
rect 13081 22760 13093 22763
rect 12069 22723 12127 22729
rect 12406 22732 13093 22760
rect 4632 22664 4752 22692
rect 1210 22584 1216 22636
rect 1268 22624 1274 22636
rect 1670 22624 1676 22636
rect 1268 22596 1676 22624
rect 1268 22584 1274 22596
rect 1670 22584 1676 22596
rect 1728 22584 1734 22636
rect 2961 22627 3019 22633
rect 2961 22593 2973 22627
rect 3007 22624 3019 22627
rect 3007 22596 3832 22624
rect 3007 22593 3019 22596
rect 2961 22587 3019 22593
rect 2501 22559 2559 22565
rect 2501 22525 2513 22559
rect 2547 22556 2559 22559
rect 3234 22556 3240 22568
rect 2547 22528 3240 22556
rect 2547 22525 2559 22528
rect 2501 22519 2559 22525
rect 3234 22516 3240 22528
rect 3292 22516 3298 22568
rect 3418 22516 3424 22568
rect 3476 22556 3482 22568
rect 3694 22556 3700 22568
rect 3476 22528 3700 22556
rect 3476 22516 3482 22528
rect 3694 22516 3700 22528
rect 3752 22516 3758 22568
rect 3804 22432 3832 22596
rect 4724 22488 4752 22664
rect 5718 22652 5724 22704
rect 5776 22652 5782 22704
rect 7285 22695 7343 22701
rect 7285 22661 7297 22695
rect 7331 22692 7343 22695
rect 7374 22692 7380 22704
rect 7331 22664 7380 22692
rect 7331 22661 7343 22664
rect 7285 22655 7343 22661
rect 7374 22652 7380 22664
rect 7432 22652 7438 22704
rect 8754 22652 8760 22704
rect 8812 22652 8818 22704
rect 9674 22692 9680 22704
rect 8864 22664 9680 22692
rect 4801 22627 4859 22633
rect 4801 22593 4813 22627
rect 4847 22624 4859 22627
rect 5810 22624 5816 22636
rect 4847 22596 5816 22624
rect 4847 22593 4859 22596
rect 4801 22587 4859 22593
rect 5810 22584 5816 22596
rect 5868 22584 5874 22636
rect 6641 22627 6699 22633
rect 6641 22593 6653 22627
rect 6687 22624 6699 22627
rect 6730 22624 6736 22636
rect 6687 22596 6736 22624
rect 6687 22593 6699 22596
rect 6641 22587 6699 22593
rect 6730 22584 6736 22596
rect 6788 22584 6794 22636
rect 7561 22627 7619 22633
rect 7561 22593 7573 22627
rect 7607 22593 7619 22627
rect 7561 22587 7619 22593
rect 6178 22516 6184 22568
rect 6236 22556 6242 22568
rect 7576 22556 7604 22587
rect 6236 22528 7604 22556
rect 6236 22516 6242 22528
rect 8864 22488 8892 22664
rect 9674 22652 9680 22664
rect 9732 22652 9738 22704
rect 9766 22652 9772 22704
rect 9824 22692 9830 22704
rect 9950 22692 9956 22704
rect 9824 22664 9956 22692
rect 9824 22652 9830 22664
rect 9950 22652 9956 22664
rect 10008 22692 10014 22704
rect 10008 22664 10166 22692
rect 10008 22652 10014 22664
rect 11054 22652 11060 22704
rect 11112 22692 11118 22704
rect 12406 22692 12434 22732
rect 13081 22729 13093 22732
rect 13127 22729 13139 22763
rect 14550 22760 14556 22772
rect 13081 22723 13139 22729
rect 14292 22732 14556 22760
rect 13814 22692 13820 22704
rect 11112 22664 12434 22692
rect 13648 22664 13820 22692
rect 11112 22652 11118 22664
rect 12161 22627 12219 22633
rect 12161 22593 12173 22627
rect 12207 22624 12219 22627
rect 12207 22596 12434 22624
rect 12207 22593 12219 22596
rect 12161 22587 12219 22593
rect 9030 22516 9036 22568
rect 9088 22556 9094 22568
rect 9401 22559 9459 22565
rect 9401 22556 9413 22559
rect 9088 22528 9413 22556
rect 9088 22516 9094 22528
rect 9401 22525 9413 22528
rect 9447 22525 9459 22559
rect 9401 22519 9459 22525
rect 9677 22559 9735 22565
rect 9677 22525 9689 22559
rect 9723 22556 9735 22559
rect 12253 22559 12311 22565
rect 12253 22556 12265 22559
rect 9723 22528 12265 22556
rect 9723 22525 9735 22528
rect 9677 22519 9735 22525
rect 12253 22525 12265 22528
rect 12299 22525 12311 22559
rect 12406 22556 12434 22596
rect 12710 22584 12716 22636
rect 12768 22624 12774 22636
rect 13648 22633 13676 22664
rect 13814 22652 13820 22664
rect 13872 22652 13878 22704
rect 13998 22652 14004 22704
rect 14056 22692 14062 22704
rect 14292 22692 14320 22732
rect 14550 22720 14556 22732
rect 14608 22720 14614 22772
rect 14734 22720 14740 22772
rect 14792 22760 14798 22772
rect 15381 22763 15439 22769
rect 15381 22760 15393 22763
rect 14792 22732 15393 22760
rect 14792 22720 14798 22732
rect 15381 22729 15393 22732
rect 15427 22729 15439 22763
rect 15381 22723 15439 22729
rect 15562 22720 15568 22772
rect 15620 22760 15626 22772
rect 16393 22763 16451 22769
rect 16393 22760 16405 22763
rect 15620 22732 16405 22760
rect 15620 22720 15626 22732
rect 16393 22729 16405 22732
rect 16439 22760 16451 22763
rect 16850 22760 16856 22772
rect 16439 22732 16856 22760
rect 16439 22729 16451 22732
rect 16393 22723 16451 22729
rect 16850 22720 16856 22732
rect 16908 22760 16914 22772
rect 16908 22732 17356 22760
rect 16908 22720 16914 22732
rect 16574 22692 16580 22704
rect 14056 22664 14398 22692
rect 15856 22664 16580 22692
rect 14056 22652 14062 22664
rect 12989 22627 13047 22633
rect 12989 22624 13001 22627
rect 12768 22596 13001 22624
rect 12768 22584 12774 22596
rect 12989 22593 13001 22596
rect 13035 22593 13047 22627
rect 12989 22587 13047 22593
rect 13633 22627 13691 22633
rect 13633 22593 13645 22627
rect 13679 22593 13691 22627
rect 15856 22624 15884 22664
rect 16574 22652 16580 22664
rect 16632 22652 16638 22704
rect 17126 22692 17132 22704
rect 16868 22664 17132 22692
rect 13633 22587 13691 22593
rect 15580 22596 15884 22624
rect 13909 22559 13967 22565
rect 12406 22528 13768 22556
rect 12253 22519 12311 22525
rect 12066 22488 12072 22500
rect 4724 22460 8892 22488
rect 10704 22460 12072 22488
rect 1762 22380 1768 22432
rect 1820 22380 1826 22432
rect 3786 22380 3792 22432
rect 3844 22380 3850 22432
rect 5534 22380 5540 22432
rect 5592 22420 5598 22432
rect 6733 22423 6791 22429
rect 6733 22420 6745 22423
rect 5592 22392 6745 22420
rect 5592 22380 5598 22392
rect 6733 22389 6745 22392
rect 6779 22389 6791 22423
rect 6733 22383 6791 22389
rect 9398 22380 9404 22432
rect 9456 22420 9462 22432
rect 10704 22420 10732 22460
rect 12066 22448 12072 22460
rect 12124 22448 12130 22500
rect 12268 22488 12296 22519
rect 12434 22488 12440 22500
rect 12268 22460 12440 22488
rect 12434 22448 12440 22460
rect 12492 22448 12498 22500
rect 12618 22448 12624 22500
rect 12676 22488 12682 22500
rect 12986 22488 12992 22500
rect 12676 22460 12992 22488
rect 12676 22448 12682 22460
rect 12986 22448 12992 22460
rect 13044 22448 13050 22500
rect 9456 22392 10732 22420
rect 9456 22380 9462 22392
rect 11146 22380 11152 22432
rect 11204 22380 11210 22432
rect 11238 22380 11244 22432
rect 11296 22420 11302 22432
rect 11701 22423 11759 22429
rect 11701 22420 11713 22423
rect 11296 22392 11713 22420
rect 11296 22380 11302 22392
rect 11701 22389 11713 22392
rect 11747 22389 11759 22423
rect 11701 22383 11759 22389
rect 12526 22380 12532 22432
rect 12584 22420 12590 22432
rect 12894 22420 12900 22432
rect 12584 22392 12900 22420
rect 12584 22380 12590 22392
rect 12894 22380 12900 22392
rect 12952 22380 12958 22432
rect 13740 22420 13768 22528
rect 13909 22525 13921 22559
rect 13955 22556 13967 22559
rect 15580 22556 15608 22596
rect 15930 22584 15936 22636
rect 15988 22584 15994 22636
rect 16868 22633 16896 22664
rect 17126 22652 17132 22664
rect 17184 22652 17190 22704
rect 17328 22692 17356 22732
rect 18598 22720 18604 22772
rect 18656 22720 18662 22772
rect 20898 22720 20904 22772
rect 20956 22760 20962 22772
rect 23842 22760 23848 22772
rect 20956 22732 23848 22760
rect 20956 22720 20962 22732
rect 23842 22720 23848 22732
rect 23900 22720 23906 22772
rect 19794 22692 19800 22704
rect 17328 22664 17618 22692
rect 18616 22664 19800 22692
rect 16853 22627 16911 22633
rect 16853 22593 16865 22627
rect 16899 22593 16911 22627
rect 16853 22587 16911 22593
rect 13955 22528 15608 22556
rect 13955 22525 13967 22528
rect 13909 22519 13967 22525
rect 15654 22516 15660 22568
rect 15712 22556 15718 22568
rect 16298 22556 16304 22568
rect 15712 22528 16304 22556
rect 15712 22516 15718 22528
rect 16298 22516 16304 22528
rect 16356 22556 16362 22568
rect 17129 22559 17187 22565
rect 17129 22556 17141 22559
rect 16356 22528 17141 22556
rect 16356 22516 16362 22528
rect 17129 22525 17141 22528
rect 17175 22556 17187 22559
rect 18616 22556 18644 22664
rect 19794 22652 19800 22664
rect 19852 22652 19858 22704
rect 22278 22692 22284 22704
rect 22020 22664 22284 22692
rect 19153 22627 19211 22633
rect 19153 22593 19165 22627
rect 19199 22593 19211 22627
rect 19153 22587 19211 22593
rect 17175 22528 18644 22556
rect 17175 22525 17187 22528
rect 17129 22519 17187 22525
rect 15286 22448 15292 22500
rect 15344 22488 15350 22500
rect 15344 22460 16344 22488
rect 15344 22448 15350 22460
rect 16316 22432 16344 22460
rect 15838 22420 15844 22432
rect 13740 22392 15844 22420
rect 15838 22380 15844 22392
rect 15896 22380 15902 22432
rect 16022 22380 16028 22432
rect 16080 22380 16086 22432
rect 16298 22380 16304 22432
rect 16356 22380 16362 22432
rect 16482 22380 16488 22432
rect 16540 22420 16546 22432
rect 19168 22420 19196 22587
rect 19426 22584 19432 22636
rect 19484 22624 19490 22636
rect 19613 22627 19671 22633
rect 19613 22624 19625 22627
rect 19484 22596 19625 22624
rect 19484 22584 19490 22596
rect 19613 22593 19625 22596
rect 19659 22624 19671 22627
rect 19886 22624 19892 22636
rect 19659 22596 19892 22624
rect 19659 22593 19671 22596
rect 19613 22587 19671 22593
rect 19886 22584 19892 22596
rect 19944 22584 19950 22636
rect 20254 22584 20260 22636
rect 20312 22584 20318 22636
rect 22020 22633 22048 22664
rect 22278 22652 22284 22664
rect 22336 22652 22342 22704
rect 24026 22692 24032 22704
rect 22388 22664 24032 22692
rect 22388 22636 22416 22664
rect 24026 22652 24032 22664
rect 24084 22652 24090 22704
rect 22005 22627 22063 22633
rect 22005 22593 22017 22627
rect 22051 22593 22063 22627
rect 22370 22624 22376 22636
rect 22005 22587 22063 22593
rect 22204 22596 22376 22624
rect 19904 22556 19932 22584
rect 20533 22559 20591 22565
rect 20533 22556 20545 22559
rect 19904 22528 20545 22556
rect 20533 22525 20545 22528
rect 20579 22556 20591 22559
rect 20806 22556 20812 22568
rect 20579 22528 20812 22556
rect 20579 22525 20591 22528
rect 20533 22519 20591 22525
rect 20806 22516 20812 22528
rect 20864 22556 20870 22568
rect 22204 22556 22232 22596
rect 22370 22584 22376 22596
rect 22428 22584 22434 22636
rect 20864 22528 22232 22556
rect 22281 22559 22339 22565
rect 20864 22516 20870 22528
rect 22281 22525 22293 22559
rect 22327 22556 22339 22559
rect 22554 22556 22560 22568
rect 22327 22528 22560 22556
rect 22327 22525 22339 22528
rect 22281 22519 22339 22525
rect 22554 22516 22560 22528
rect 22612 22516 22618 22568
rect 23290 22516 23296 22568
rect 23348 22516 23354 22568
rect 23569 22559 23627 22565
rect 23569 22525 23581 22559
rect 23615 22556 23627 22559
rect 24118 22556 24124 22568
rect 23615 22528 24124 22556
rect 23615 22525 23627 22528
rect 23569 22519 23627 22525
rect 24118 22516 24124 22528
rect 24176 22556 24182 22568
rect 25866 22556 25872 22568
rect 24176 22528 25872 22556
rect 24176 22516 24182 22528
rect 25866 22516 25872 22528
rect 25924 22516 25930 22568
rect 19337 22491 19395 22497
rect 19337 22457 19349 22491
rect 19383 22488 19395 22491
rect 19426 22488 19432 22500
rect 19383 22460 19432 22488
rect 19383 22457 19395 22460
rect 19337 22451 19395 22457
rect 19426 22448 19432 22460
rect 19484 22448 19490 22500
rect 16540 22392 19196 22420
rect 16540 22380 16546 22392
rect 20254 22380 20260 22432
rect 20312 22420 20318 22432
rect 21082 22420 21088 22432
rect 20312 22392 21088 22420
rect 20312 22380 20318 22392
rect 21082 22380 21088 22392
rect 21140 22380 21146 22432
rect 23658 22380 23664 22432
rect 23716 22420 23722 22432
rect 24762 22420 24768 22432
rect 23716 22392 24768 22420
rect 23716 22380 23722 22392
rect 24762 22380 24768 22392
rect 24820 22420 24826 22432
rect 25041 22423 25099 22429
rect 25041 22420 25053 22423
rect 24820 22392 25053 22420
rect 24820 22380 24826 22392
rect 25041 22389 25053 22392
rect 25087 22389 25099 22423
rect 25041 22383 25099 22389
rect 25409 22423 25467 22429
rect 25409 22389 25421 22423
rect 25455 22420 25467 22423
rect 25498 22420 25504 22432
rect 25455 22392 25504 22420
rect 25455 22389 25467 22392
rect 25409 22383 25467 22389
rect 25498 22380 25504 22392
rect 25556 22380 25562 22432
rect 1104 22330 25852 22352
rect 1104 22278 2950 22330
rect 3002 22278 3014 22330
rect 3066 22278 3078 22330
rect 3130 22278 3142 22330
rect 3194 22278 3206 22330
rect 3258 22278 12950 22330
rect 13002 22278 13014 22330
rect 13066 22278 13078 22330
rect 13130 22278 13142 22330
rect 13194 22278 13206 22330
rect 13258 22278 22950 22330
rect 23002 22278 23014 22330
rect 23066 22278 23078 22330
rect 23130 22278 23142 22330
rect 23194 22278 23206 22330
rect 23258 22278 25852 22330
rect 1104 22256 25852 22278
rect 1670 22176 1676 22228
rect 1728 22176 1734 22228
rect 10594 22216 10600 22228
rect 2746 22188 10600 22216
rect 1762 22108 1768 22160
rect 1820 22148 1826 22160
rect 2746 22148 2774 22188
rect 10594 22176 10600 22188
rect 10652 22176 10658 22228
rect 10952 22219 11010 22225
rect 10952 22185 10964 22219
rect 10998 22216 11010 22219
rect 12802 22216 12808 22228
rect 10998 22188 12808 22216
rect 10998 22185 11010 22188
rect 10952 22179 11010 22185
rect 12802 22176 12808 22188
rect 12860 22176 12866 22228
rect 14540 22219 14598 22225
rect 14540 22185 14552 22219
rect 14586 22216 14598 22219
rect 14734 22216 14740 22228
rect 14586 22188 14740 22216
rect 14586 22185 14598 22188
rect 14540 22179 14598 22185
rect 14734 22176 14740 22188
rect 14792 22176 14798 22228
rect 15580 22188 16896 22216
rect 1820 22120 2774 22148
rect 1820 22108 1826 22120
rect 3602 22108 3608 22160
rect 3660 22148 3666 22160
rect 3786 22148 3792 22160
rect 3660 22120 3792 22148
rect 3660 22108 3666 22120
rect 3786 22108 3792 22120
rect 3844 22108 3850 22160
rect 9398 22148 9404 22160
rect 8864 22120 9404 22148
rect 2866 22040 2872 22092
rect 2924 22040 2930 22092
rect 6086 22040 6092 22092
rect 6144 22040 6150 22092
rect 8294 22040 8300 22092
rect 8352 22040 8358 22092
rect 2225 22015 2283 22021
rect 2225 21981 2237 22015
rect 2271 21981 2283 22015
rect 2225 21975 2283 21981
rect 3973 22015 4031 22021
rect 3973 21981 3985 22015
rect 4019 21981 4031 22015
rect 3973 21975 4031 21981
rect 4249 22015 4307 22021
rect 4249 21981 4261 22015
rect 4295 22012 4307 22015
rect 4522 22012 4528 22024
rect 4295 21984 4528 22012
rect 4295 21981 4307 21984
rect 4249 21975 4307 21981
rect 2240 21876 2268 21975
rect 3988 21944 4016 21975
rect 4522 21972 4528 21984
rect 4580 21972 4586 22024
rect 5442 21972 5448 22024
rect 5500 21972 5506 22024
rect 7377 22015 7435 22021
rect 7377 21981 7389 22015
rect 7423 22012 7435 22015
rect 7834 22012 7840 22024
rect 7423 21984 7840 22012
rect 7423 21981 7435 21984
rect 7377 21975 7435 21981
rect 7834 21972 7840 21984
rect 7892 21972 7898 22024
rect 8294 21944 8300 21956
rect 3988 21916 8300 21944
rect 8294 21904 8300 21916
rect 8352 21944 8358 21956
rect 8864 21944 8892 22120
rect 9398 22108 9404 22120
rect 9456 22108 9462 22160
rect 12250 22108 12256 22160
rect 12308 22148 12314 22160
rect 13446 22148 13452 22160
rect 12308 22120 13452 22148
rect 12308 22108 12314 22120
rect 13446 22108 13452 22120
rect 13504 22108 13510 22160
rect 13556 22120 14412 22148
rect 9030 22040 9036 22092
rect 9088 22080 9094 22092
rect 10689 22083 10747 22089
rect 10689 22080 10701 22083
rect 9088 22052 10701 22080
rect 9088 22040 9094 22052
rect 10689 22049 10701 22052
rect 10735 22080 10747 22083
rect 11054 22080 11060 22092
rect 10735 22052 11060 22080
rect 10735 22049 10747 22052
rect 10689 22043 10747 22049
rect 11054 22040 11060 22052
rect 11112 22040 11118 22092
rect 11698 22040 11704 22092
rect 11756 22080 11762 22092
rect 11756 22052 12388 22080
rect 11756 22040 11762 22052
rect 8941 22015 8999 22021
rect 8941 21981 8953 22015
rect 8987 22012 8999 22015
rect 9493 22015 9551 22021
rect 9493 22012 9505 22015
rect 8987 21984 9505 22012
rect 8987 21981 8999 21984
rect 8941 21975 8999 21981
rect 9493 21981 9505 21984
rect 9539 22012 9551 22015
rect 12360 22012 12388 22052
rect 12434 22040 12440 22092
rect 12492 22040 12498 22092
rect 13170 22040 13176 22092
rect 13228 22080 13234 22092
rect 13556 22080 13584 22120
rect 13228 22052 13584 22080
rect 13228 22040 13234 22052
rect 13814 22040 13820 22092
rect 13872 22080 13878 22092
rect 14277 22083 14335 22089
rect 14277 22080 14289 22083
rect 13872 22052 14289 22080
rect 13872 22040 13878 22052
rect 14277 22049 14289 22052
rect 14323 22049 14335 22083
rect 14384 22080 14412 22120
rect 15580 22080 15608 22188
rect 15838 22108 15844 22160
rect 15896 22148 15902 22160
rect 16485 22151 16543 22157
rect 16485 22148 16497 22151
rect 15896 22120 16497 22148
rect 15896 22108 15902 22120
rect 16485 22117 16497 22120
rect 16531 22117 16543 22151
rect 16485 22111 16543 22117
rect 14384 22052 15608 22080
rect 16868 22094 16896 22188
rect 17126 22176 17132 22228
rect 17184 22216 17190 22228
rect 18877 22219 18935 22225
rect 18877 22216 18889 22219
rect 17184 22188 18889 22216
rect 17184 22176 17190 22188
rect 18877 22185 18889 22188
rect 18923 22216 18935 22219
rect 18966 22216 18972 22228
rect 18923 22188 18972 22216
rect 18923 22185 18935 22188
rect 18877 22179 18935 22185
rect 18966 22176 18972 22188
rect 19024 22176 19030 22228
rect 19058 22176 19064 22228
rect 19116 22216 19122 22228
rect 21818 22216 21824 22228
rect 19116 22188 21824 22216
rect 19116 22176 19122 22188
rect 21818 22176 21824 22188
rect 21876 22176 21882 22228
rect 22278 22176 22284 22228
rect 22336 22216 22342 22228
rect 25774 22216 25780 22228
rect 22336 22188 25780 22216
rect 22336 22176 22342 22188
rect 25774 22176 25780 22188
rect 25832 22176 25838 22228
rect 17678 22108 17684 22160
rect 17736 22148 17742 22160
rect 20254 22148 20260 22160
rect 17736 22120 20260 22148
rect 17736 22108 17742 22120
rect 20254 22108 20260 22120
rect 20312 22108 20318 22160
rect 21634 22108 21640 22160
rect 21692 22148 21698 22160
rect 22738 22148 22744 22160
rect 21692 22120 22744 22148
rect 21692 22108 21698 22120
rect 22738 22108 22744 22120
rect 22796 22108 22802 22160
rect 25314 22148 25320 22160
rect 25240 22120 25320 22148
rect 16868 22089 17080 22094
rect 16868 22083 17095 22089
rect 16868 22066 17049 22083
rect 14277 22043 14335 22049
rect 17037 22049 17049 22066
rect 17083 22049 17095 22083
rect 17037 22043 17095 22049
rect 17218 22040 17224 22092
rect 17276 22080 17282 22092
rect 18138 22080 18144 22092
rect 17276 22052 18144 22080
rect 17276 22040 17282 22052
rect 18138 22040 18144 22052
rect 18196 22040 18202 22092
rect 18233 22083 18291 22089
rect 18233 22049 18245 22083
rect 18279 22049 18291 22083
rect 19981 22083 20039 22089
rect 19981 22080 19993 22083
rect 18233 22043 18291 22049
rect 18340 22052 19993 22080
rect 12989 22015 13047 22021
rect 12989 22012 13001 22015
rect 9539 21984 10272 22012
rect 12360 21984 13001 22012
rect 9539 21981 9551 21984
rect 9493 21975 9551 21981
rect 8352 21916 8892 21944
rect 8352 21904 8358 21916
rect 4982 21876 4988 21888
rect 2240 21848 4988 21876
rect 4982 21836 4988 21848
rect 5040 21836 5046 21888
rect 9306 21836 9312 21888
rect 9364 21836 9370 21888
rect 10042 21836 10048 21888
rect 10100 21836 10106 21888
rect 10244 21876 10272 21984
rect 12989 21981 13001 21984
rect 13035 22012 13047 22015
rect 13354 22012 13360 22024
rect 13035 21984 13360 22012
rect 13035 21981 13047 21984
rect 12989 21975 13047 21981
rect 13354 21972 13360 21984
rect 13412 21972 13418 22024
rect 14182 22012 14188 22024
rect 13464 21984 14188 22012
rect 11698 21904 11704 21956
rect 11756 21904 11762 21956
rect 12434 21904 12440 21956
rect 12492 21944 12498 21956
rect 13464 21944 13492 21984
rect 14182 21972 14188 21984
rect 14240 21972 14246 22024
rect 18248 22012 18276 22043
rect 16040 21984 18276 22012
rect 12492 21916 13492 21944
rect 12492 21904 12498 21916
rect 13538 21904 13544 21956
rect 13596 21904 13602 21956
rect 13998 21904 14004 21956
rect 14056 21944 14062 21956
rect 14056 21916 15042 21944
rect 14056 21904 14062 21916
rect 12250 21876 12256 21888
rect 10244 21848 12256 21876
rect 12250 21836 12256 21848
rect 12308 21836 12314 21888
rect 12894 21836 12900 21888
rect 12952 21836 12958 21888
rect 13170 21836 13176 21888
rect 13228 21876 13234 21888
rect 13633 21879 13691 21885
rect 13633 21876 13645 21879
rect 13228 21848 13645 21876
rect 13228 21836 13234 21848
rect 13633 21845 13645 21848
rect 13679 21845 13691 21879
rect 13633 21839 13691 21845
rect 15286 21836 15292 21888
rect 15344 21876 15350 21888
rect 16040 21885 16068 21984
rect 16853 21947 16911 21953
rect 16853 21913 16865 21947
rect 16899 21944 16911 21947
rect 17310 21944 17316 21956
rect 16899 21916 17316 21944
rect 16899 21913 16911 21916
rect 16853 21907 16911 21913
rect 17310 21904 17316 21916
rect 17368 21904 17374 21956
rect 17494 21904 17500 21956
rect 17552 21944 17558 21956
rect 18340 21944 18368 22052
rect 19981 22049 19993 22052
rect 20027 22049 20039 22083
rect 19981 22043 20039 22049
rect 20162 22040 20168 22092
rect 20220 22080 20226 22092
rect 20220 22052 22094 22080
rect 20220 22040 20226 22052
rect 19058 22012 19064 22024
rect 17552 21916 18368 21944
rect 18616 21984 19064 22012
rect 17552 21904 17558 21916
rect 16025 21879 16083 21885
rect 16025 21876 16037 21879
rect 15344 21848 16037 21876
rect 15344 21836 15350 21848
rect 16025 21845 16037 21848
rect 16071 21845 16083 21879
rect 16025 21839 16083 21845
rect 16758 21836 16764 21888
rect 16816 21876 16822 21888
rect 16945 21879 17003 21885
rect 16945 21876 16957 21879
rect 16816 21848 16957 21876
rect 16816 21836 16822 21848
rect 16945 21845 16957 21848
rect 16991 21876 17003 21879
rect 17126 21876 17132 21888
rect 16991 21848 17132 21876
rect 16991 21845 17003 21848
rect 16945 21839 17003 21845
rect 17126 21836 17132 21848
rect 17184 21836 17190 21888
rect 17678 21836 17684 21888
rect 17736 21836 17742 21888
rect 17770 21836 17776 21888
rect 17828 21876 17834 21888
rect 18049 21879 18107 21885
rect 18049 21876 18061 21879
rect 17828 21848 18061 21876
rect 17828 21836 17834 21848
rect 18049 21845 18061 21848
rect 18095 21845 18107 21879
rect 18049 21839 18107 21845
rect 18138 21836 18144 21888
rect 18196 21876 18202 21888
rect 18616 21876 18644 21984
rect 19058 21972 19064 21984
rect 19116 21972 19122 22024
rect 19334 21972 19340 22024
rect 19392 22012 19398 22024
rect 20349 22015 20407 22021
rect 20349 22012 20361 22015
rect 19392 21984 20361 22012
rect 19392 21972 19398 21984
rect 20349 21981 20361 21984
rect 20395 21981 20407 22015
rect 22066 22012 22094 22052
rect 22186 22040 22192 22092
rect 22244 22080 22250 22092
rect 22244 22052 23612 22080
rect 22244 22040 22250 22052
rect 22741 22015 22799 22021
rect 22741 22012 22753 22015
rect 22066 21984 22753 22012
rect 20349 21975 20407 21981
rect 22741 21981 22753 21984
rect 22787 21981 22799 22015
rect 22741 21975 22799 21981
rect 22830 21972 22836 22024
rect 22888 22012 22894 22024
rect 23198 22012 23204 22024
rect 22888 21984 23204 22012
rect 22888 21972 22894 21984
rect 23198 21972 23204 21984
rect 23256 21972 23262 22024
rect 23474 21972 23480 22024
rect 23532 21972 23538 22024
rect 23584 22012 23612 22052
rect 24854 22040 24860 22092
rect 24912 22080 24918 22092
rect 25130 22080 25136 22092
rect 24912 22052 25136 22080
rect 24912 22040 24918 22052
rect 25130 22040 25136 22052
rect 25188 22040 25194 22092
rect 25240 22089 25268 22120
rect 25314 22108 25320 22120
rect 25372 22108 25378 22160
rect 25225 22083 25283 22089
rect 25225 22049 25237 22083
rect 25271 22080 25283 22083
rect 25271 22052 25305 22080
rect 25271 22049 25283 22052
rect 25225 22043 25283 22049
rect 25958 22012 25964 22024
rect 23584 21984 25964 22012
rect 25958 21972 25964 21984
rect 26016 21972 26022 22024
rect 19518 21904 19524 21956
rect 19576 21904 19582 21956
rect 20625 21947 20683 21953
rect 20625 21913 20637 21947
rect 20671 21944 20683 21947
rect 20898 21944 20904 21956
rect 20671 21916 20904 21944
rect 20671 21913 20683 21916
rect 20625 21907 20683 21913
rect 20898 21904 20904 21916
rect 20956 21904 20962 21956
rect 23842 21944 23848 21956
rect 21008 21916 21114 21944
rect 22296 21916 23848 21944
rect 18196 21848 18644 21876
rect 18196 21836 18202 21848
rect 18690 21836 18696 21888
rect 18748 21836 18754 21888
rect 19610 21836 19616 21888
rect 19668 21836 19674 21888
rect 20806 21836 20812 21888
rect 20864 21876 20870 21888
rect 21008 21876 21036 21916
rect 22296 21888 22324 21916
rect 23842 21904 23848 21916
rect 23900 21904 23906 21956
rect 24026 21904 24032 21956
rect 24084 21944 24090 21956
rect 24949 21947 25007 21953
rect 24949 21944 24961 21947
rect 24084 21916 24961 21944
rect 24084 21904 24090 21916
rect 24949 21913 24961 21916
rect 24995 21913 25007 21947
rect 24949 21907 25007 21913
rect 20864 21848 21036 21876
rect 20864 21836 20870 21848
rect 21266 21836 21272 21888
rect 21324 21876 21330 21888
rect 21450 21876 21456 21888
rect 21324 21848 21456 21876
rect 21324 21836 21330 21848
rect 21450 21836 21456 21848
rect 21508 21836 21514 21888
rect 22097 21879 22155 21885
rect 22097 21845 22109 21879
rect 22143 21876 22155 21879
rect 22186 21876 22192 21888
rect 22143 21848 22192 21876
rect 22143 21845 22155 21848
rect 22097 21839 22155 21845
rect 22186 21836 22192 21848
rect 22244 21836 22250 21888
rect 22278 21836 22284 21888
rect 22336 21836 22342 21888
rect 22557 21879 22615 21885
rect 22557 21845 22569 21879
rect 22603 21876 22615 21879
rect 23566 21876 23572 21888
rect 22603 21848 23572 21876
rect 22603 21845 22615 21848
rect 22557 21839 22615 21845
rect 23566 21836 23572 21848
rect 23624 21836 23630 21888
rect 23750 21836 23756 21888
rect 23808 21876 23814 21888
rect 24581 21879 24639 21885
rect 24581 21876 24593 21879
rect 23808 21848 24593 21876
rect 23808 21836 23814 21848
rect 24581 21845 24593 21848
rect 24627 21845 24639 21879
rect 24581 21839 24639 21845
rect 25041 21879 25099 21885
rect 25041 21845 25053 21879
rect 25087 21876 25099 21879
rect 26234 21876 26240 21888
rect 25087 21848 26240 21876
rect 25087 21845 25099 21848
rect 25041 21839 25099 21845
rect 26234 21836 26240 21848
rect 26292 21836 26298 21888
rect 1104 21786 25852 21808
rect 1104 21734 7950 21786
rect 8002 21734 8014 21786
rect 8066 21734 8078 21786
rect 8130 21734 8142 21786
rect 8194 21734 8206 21786
rect 8258 21734 17950 21786
rect 18002 21734 18014 21786
rect 18066 21734 18078 21786
rect 18130 21734 18142 21786
rect 18194 21734 18206 21786
rect 18258 21734 25852 21786
rect 1104 21712 25852 21734
rect 2133 21675 2191 21681
rect 2133 21641 2145 21675
rect 2179 21672 2191 21675
rect 3418 21672 3424 21684
rect 2179 21644 3424 21672
rect 2179 21641 2191 21644
rect 2133 21635 2191 21641
rect 1673 21607 1731 21613
rect 1673 21573 1685 21607
rect 1719 21604 1731 21607
rect 2148 21604 2176 21635
rect 3418 21632 3424 21644
rect 3476 21632 3482 21684
rect 6454 21632 6460 21684
rect 6512 21672 6518 21684
rect 8202 21672 8208 21684
rect 6512 21644 8208 21672
rect 6512 21632 6518 21644
rect 8202 21632 8208 21644
rect 8260 21672 8266 21684
rect 8478 21672 8484 21684
rect 8260 21644 8484 21672
rect 8260 21632 8266 21644
rect 8478 21632 8484 21644
rect 8536 21632 8542 21684
rect 10042 21632 10048 21684
rect 10100 21672 10106 21684
rect 12621 21675 12679 21681
rect 12621 21672 12633 21675
rect 10100 21644 12633 21672
rect 10100 21632 10106 21644
rect 12621 21641 12633 21644
rect 12667 21641 12679 21675
rect 12621 21635 12679 21641
rect 13446 21632 13452 21684
rect 13504 21632 13510 21684
rect 16206 21672 16212 21684
rect 13556 21644 16212 21672
rect 5534 21604 5540 21616
rect 1719 21576 2176 21604
rect 2976 21576 5540 21604
rect 1719 21573 1731 21576
rect 1673 21567 1731 21573
rect 2976 21545 3004 21576
rect 5534 21564 5540 21576
rect 5592 21564 5598 21616
rect 9398 21604 9404 21616
rect 6748 21576 9404 21604
rect 2961 21539 3019 21545
rect 2961 21505 2973 21539
rect 3007 21505 3019 21539
rect 2961 21499 3019 21505
rect 4798 21496 4804 21548
rect 4856 21496 4862 21548
rect 6748 21545 6776 21576
rect 9398 21564 9404 21576
rect 9456 21564 9462 21616
rect 9766 21564 9772 21616
rect 9824 21564 9830 21616
rect 11793 21607 11851 21613
rect 11793 21573 11805 21607
rect 11839 21604 11851 21607
rect 13556 21604 13584 21644
rect 16206 21632 16212 21644
rect 16264 21672 16270 21684
rect 20162 21672 20168 21684
rect 16264 21644 20168 21672
rect 16264 21632 16270 21644
rect 20162 21632 20168 21644
rect 20220 21632 20226 21684
rect 20438 21632 20444 21684
rect 20496 21632 20502 21684
rect 20732 21644 21496 21672
rect 11839 21576 13584 21604
rect 14277 21607 14335 21613
rect 11839 21573 11851 21576
rect 11793 21567 11851 21573
rect 14277 21573 14289 21607
rect 14323 21604 14335 21607
rect 17678 21604 17684 21616
rect 14323 21576 17684 21604
rect 14323 21573 14335 21576
rect 14277 21567 14335 21573
rect 17678 21564 17684 21576
rect 17736 21564 17742 21616
rect 18233 21607 18291 21613
rect 18233 21573 18245 21607
rect 18279 21604 18291 21607
rect 18506 21604 18512 21616
rect 18279 21576 18512 21604
rect 18279 21573 18291 21576
rect 18233 21567 18291 21573
rect 18506 21564 18512 21576
rect 18564 21604 18570 21616
rect 20732 21604 20760 21644
rect 18564 21576 20760 21604
rect 18564 21564 18570 21576
rect 21468 21548 21496 21644
rect 21542 21632 21548 21684
rect 21600 21672 21606 21684
rect 22005 21675 22063 21681
rect 22005 21672 22017 21675
rect 21600 21644 22017 21672
rect 21600 21632 21606 21644
rect 22005 21641 22017 21644
rect 22051 21641 22063 21675
rect 22005 21635 22063 21641
rect 22094 21632 22100 21684
rect 22152 21672 22158 21684
rect 24670 21672 24676 21684
rect 22152 21644 24676 21672
rect 22152 21632 22158 21644
rect 24670 21632 24676 21644
rect 24728 21632 24734 21684
rect 23658 21564 23664 21616
rect 23716 21564 23722 21616
rect 24118 21564 24124 21616
rect 24176 21564 24182 21616
rect 6733 21539 6791 21545
rect 6733 21505 6745 21539
rect 6779 21505 6791 21539
rect 6733 21499 6791 21505
rect 7374 21496 7380 21548
rect 7432 21496 7438 21548
rect 9030 21496 9036 21548
rect 9088 21496 9094 21548
rect 11146 21496 11152 21548
rect 11204 21536 11210 21548
rect 13262 21536 13268 21548
rect 11204 21508 13268 21536
rect 11204 21496 11210 21508
rect 13262 21496 13268 21508
rect 13320 21496 13326 21548
rect 13357 21539 13415 21545
rect 13357 21505 13369 21539
rect 13403 21536 13415 21539
rect 14090 21536 14096 21548
rect 13403 21508 14096 21536
rect 13403 21505 13415 21508
rect 13357 21499 13415 21505
rect 14090 21496 14096 21508
rect 14148 21496 14154 21548
rect 14182 21496 14188 21548
rect 14240 21496 14246 21548
rect 14826 21496 14832 21548
rect 14884 21536 14890 21548
rect 15381 21539 15439 21545
rect 15381 21536 15393 21539
rect 14884 21508 15393 21536
rect 14884 21496 14890 21508
rect 15381 21505 15393 21508
rect 15427 21505 15439 21539
rect 15381 21499 15439 21505
rect 15473 21539 15531 21545
rect 15473 21505 15485 21539
rect 15519 21536 15531 21539
rect 15562 21536 15568 21548
rect 15519 21508 15568 21536
rect 15519 21505 15531 21508
rect 15473 21499 15531 21505
rect 15562 21496 15568 21508
rect 15620 21536 15626 21548
rect 16206 21536 16212 21548
rect 15620 21508 16212 21536
rect 15620 21496 15626 21508
rect 16206 21496 16212 21508
rect 16264 21496 16270 21548
rect 16298 21496 16304 21548
rect 16356 21536 16362 21548
rect 16850 21536 16856 21548
rect 16356 21508 16856 21536
rect 16356 21496 16362 21508
rect 16850 21496 16856 21508
rect 16908 21536 16914 21548
rect 17218 21536 17224 21548
rect 16908 21508 17224 21536
rect 16908 21496 16914 21508
rect 17218 21496 17224 21508
rect 17276 21496 17282 21548
rect 17402 21496 17408 21548
rect 17460 21536 17466 21548
rect 17862 21536 17868 21548
rect 17460 21508 17868 21536
rect 17460 21496 17466 21508
rect 17862 21496 17868 21508
rect 17920 21496 17926 21548
rect 20806 21496 20812 21548
rect 20864 21496 20870 21548
rect 21450 21496 21456 21548
rect 21508 21496 21514 21548
rect 22186 21496 22192 21548
rect 22244 21536 22250 21548
rect 22373 21539 22431 21545
rect 22373 21536 22385 21539
rect 22244 21508 22385 21536
rect 22244 21496 22250 21508
rect 22373 21505 22385 21508
rect 22419 21505 22431 21539
rect 22373 21499 22431 21505
rect 23290 21496 23296 21548
rect 23348 21536 23354 21548
rect 23385 21539 23443 21545
rect 23385 21536 23397 21539
rect 23348 21508 23397 21536
rect 23348 21496 23354 21508
rect 23385 21505 23397 21508
rect 23431 21505 23443 21539
rect 23385 21499 23443 21505
rect 3510 21428 3516 21480
rect 3568 21428 3574 21480
rect 5074 21428 5080 21480
rect 5132 21428 5138 21480
rect 7282 21428 7288 21480
rect 7340 21468 7346 21480
rect 7653 21471 7711 21477
rect 7653 21468 7665 21471
rect 7340 21440 7665 21468
rect 7340 21428 7346 21440
rect 7653 21437 7665 21440
rect 7699 21437 7711 21471
rect 7653 21431 7711 21437
rect 9309 21471 9367 21477
rect 9309 21437 9321 21471
rect 9355 21468 9367 21471
rect 11164 21468 11192 21496
rect 12526 21468 12532 21480
rect 9355 21440 11192 21468
rect 11256 21440 12532 21468
rect 9355 21437 9367 21440
rect 9309 21431 9367 21437
rect 10686 21360 10692 21412
rect 10744 21400 10750 21412
rect 11256 21400 11284 21440
rect 12526 21428 12532 21440
rect 12584 21428 12590 21480
rect 12713 21471 12771 21477
rect 12713 21437 12725 21471
rect 12759 21437 12771 21471
rect 12713 21431 12771 21437
rect 10744 21372 11284 21400
rect 10744 21360 10750 21372
rect 11422 21360 11428 21412
rect 11480 21400 11486 21412
rect 12728 21400 12756 21431
rect 12894 21428 12900 21480
rect 12952 21428 12958 21480
rect 13630 21428 13636 21480
rect 13688 21468 13694 21480
rect 14369 21471 14427 21477
rect 14369 21468 14381 21471
rect 13688 21440 14381 21468
rect 13688 21428 13694 21440
rect 14369 21437 14381 21440
rect 14415 21437 14427 21471
rect 14369 21431 14427 21437
rect 15654 21428 15660 21480
rect 15712 21428 15718 21480
rect 16114 21428 16120 21480
rect 16172 21468 16178 21480
rect 16172 21440 16712 21468
rect 16172 21428 16178 21440
rect 16574 21400 16580 21412
rect 11480 21372 12664 21400
rect 12728 21372 13216 21400
rect 11480 21360 11486 21372
rect 1762 21292 1768 21344
rect 1820 21292 1826 21344
rect 6549 21335 6607 21341
rect 6549 21301 6561 21335
rect 6595 21332 6607 21335
rect 7834 21332 7840 21344
rect 6595 21304 7840 21332
rect 6595 21301 6607 21304
rect 6549 21295 6607 21301
rect 7834 21292 7840 21304
rect 7892 21292 7898 21344
rect 10502 21292 10508 21344
rect 10560 21332 10566 21344
rect 10781 21335 10839 21341
rect 10781 21332 10793 21335
rect 10560 21304 10793 21332
rect 10560 21292 10566 21304
rect 10781 21301 10793 21304
rect 10827 21301 10839 21335
rect 10781 21295 10839 21301
rect 11146 21292 11152 21344
rect 11204 21332 11210 21344
rect 11241 21335 11299 21341
rect 11241 21332 11253 21335
rect 11204 21304 11253 21332
rect 11204 21292 11210 21304
rect 11241 21301 11253 21304
rect 11287 21332 11299 21335
rect 11517 21335 11575 21341
rect 11517 21332 11529 21335
rect 11287 21304 11529 21332
rect 11287 21301 11299 21304
rect 11241 21295 11299 21301
rect 11517 21301 11529 21304
rect 11563 21332 11575 21335
rect 11698 21332 11704 21344
rect 11563 21304 11704 21332
rect 11563 21301 11575 21304
rect 11517 21295 11575 21301
rect 11698 21292 11704 21304
rect 11756 21332 11762 21344
rect 11885 21335 11943 21341
rect 11885 21332 11897 21335
rect 11756 21304 11897 21332
rect 11756 21292 11762 21304
rect 11885 21301 11897 21304
rect 11931 21301 11943 21335
rect 11885 21295 11943 21301
rect 11974 21292 11980 21344
rect 12032 21332 12038 21344
rect 12253 21335 12311 21341
rect 12253 21332 12265 21335
rect 12032 21304 12265 21332
rect 12032 21292 12038 21304
rect 12253 21301 12265 21304
rect 12299 21301 12311 21335
rect 12636 21332 12664 21372
rect 12894 21332 12900 21344
rect 12636 21304 12900 21332
rect 12253 21295 12311 21301
rect 12894 21292 12900 21304
rect 12952 21292 12958 21344
rect 13188 21332 13216 21372
rect 13372 21372 16580 21400
rect 13372 21332 13400 21372
rect 16574 21360 16580 21372
rect 16632 21360 16638 21412
rect 16684 21400 16712 21440
rect 17494 21428 17500 21480
rect 17552 21428 17558 21480
rect 17678 21428 17684 21480
rect 17736 21428 17742 21480
rect 18414 21428 18420 21480
rect 18472 21468 18478 21480
rect 18966 21468 18972 21480
rect 18472 21440 18972 21468
rect 18472 21428 18478 21440
rect 18966 21428 18972 21440
rect 19024 21468 19030 21480
rect 20901 21471 20959 21477
rect 20901 21468 20913 21471
rect 19024 21440 20913 21468
rect 19024 21428 19030 21440
rect 20901 21437 20913 21440
rect 20947 21468 20959 21471
rect 20990 21468 20996 21480
rect 20947 21440 20996 21468
rect 20947 21437 20959 21440
rect 20901 21431 20959 21437
rect 20990 21428 20996 21440
rect 21048 21428 21054 21480
rect 21082 21428 21088 21480
rect 21140 21428 21146 21480
rect 22462 21428 22468 21480
rect 22520 21428 22526 21480
rect 22646 21428 22652 21480
rect 22704 21428 22710 21480
rect 22738 21428 22744 21480
rect 22796 21468 22802 21480
rect 23017 21471 23075 21477
rect 23017 21468 23029 21471
rect 22796 21440 23029 21468
rect 22796 21428 22802 21440
rect 23017 21437 23029 21440
rect 23063 21437 23075 21471
rect 23017 21431 23075 21437
rect 23198 21428 23204 21480
rect 23256 21468 23262 21480
rect 25682 21468 25688 21480
rect 23256 21440 25688 21468
rect 23256 21428 23262 21440
rect 25682 21428 25688 21440
rect 25740 21428 25746 21480
rect 16684 21372 19656 21400
rect 13188 21304 13400 21332
rect 13817 21335 13875 21341
rect 13817 21301 13829 21335
rect 13863 21332 13875 21335
rect 13906 21332 13912 21344
rect 13863 21304 13912 21332
rect 13863 21301 13875 21304
rect 13817 21295 13875 21301
rect 13906 21292 13912 21304
rect 13964 21292 13970 21344
rect 15010 21292 15016 21344
rect 15068 21292 15074 21344
rect 15838 21292 15844 21344
rect 15896 21332 15902 21344
rect 16025 21335 16083 21341
rect 16025 21332 16037 21335
rect 15896 21304 16037 21332
rect 15896 21292 15902 21304
rect 16025 21301 16037 21304
rect 16071 21301 16083 21335
rect 16025 21295 16083 21301
rect 16206 21292 16212 21344
rect 16264 21332 16270 21344
rect 16393 21335 16451 21341
rect 16393 21332 16405 21335
rect 16264 21304 16405 21332
rect 16264 21292 16270 21304
rect 16393 21301 16405 21304
rect 16439 21301 16451 21335
rect 16393 21295 16451 21301
rect 16666 21292 16672 21344
rect 16724 21292 16730 21344
rect 17037 21335 17095 21341
rect 17037 21301 17049 21335
rect 17083 21332 17095 21335
rect 19058 21332 19064 21344
rect 17083 21304 19064 21332
rect 17083 21301 17095 21304
rect 17037 21295 17095 21301
rect 19058 21292 19064 21304
rect 19116 21292 19122 21344
rect 19334 21292 19340 21344
rect 19392 21332 19398 21344
rect 19521 21335 19579 21341
rect 19521 21332 19533 21335
rect 19392 21304 19533 21332
rect 19392 21292 19398 21304
rect 19521 21301 19533 21304
rect 19567 21301 19579 21335
rect 19628 21332 19656 21372
rect 19978 21360 19984 21412
rect 20036 21400 20042 21412
rect 21542 21400 21548 21412
rect 20036 21372 21548 21400
rect 20036 21360 20042 21372
rect 21542 21360 21548 21372
rect 21600 21360 21606 21412
rect 22278 21400 22284 21412
rect 21652 21372 22284 21400
rect 21652 21332 21680 21372
rect 22278 21360 22284 21372
rect 22336 21360 22342 21412
rect 24854 21360 24860 21412
rect 24912 21400 24918 21412
rect 25409 21403 25467 21409
rect 25409 21400 25421 21403
rect 24912 21372 25421 21400
rect 24912 21360 24918 21372
rect 25409 21369 25421 21372
rect 25455 21369 25467 21403
rect 25409 21363 25467 21369
rect 19628 21304 21680 21332
rect 19521 21295 19579 21301
rect 21818 21292 21824 21344
rect 21876 21332 21882 21344
rect 22830 21332 22836 21344
rect 21876 21304 22836 21332
rect 21876 21292 21882 21304
rect 22830 21292 22836 21304
rect 22888 21292 22894 21344
rect 23842 21292 23848 21344
rect 23900 21332 23906 21344
rect 25133 21335 25191 21341
rect 25133 21332 25145 21335
rect 23900 21304 25145 21332
rect 23900 21292 23906 21304
rect 25133 21301 25145 21304
rect 25179 21301 25191 21335
rect 25133 21295 25191 21301
rect 1104 21242 25852 21264
rect 1104 21190 2950 21242
rect 3002 21190 3014 21242
rect 3066 21190 3078 21242
rect 3130 21190 3142 21242
rect 3194 21190 3206 21242
rect 3258 21190 12950 21242
rect 13002 21190 13014 21242
rect 13066 21190 13078 21242
rect 13130 21190 13142 21242
rect 13194 21190 13206 21242
rect 13258 21190 22950 21242
rect 23002 21190 23014 21242
rect 23066 21190 23078 21242
rect 23130 21190 23142 21242
rect 23194 21190 23206 21242
rect 23258 21190 25852 21242
rect 1104 21168 25852 21190
rect 1762 21088 1768 21140
rect 1820 21128 1826 21140
rect 10318 21128 10324 21140
rect 1820 21100 10324 21128
rect 1820 21088 1826 21100
rect 10318 21088 10324 21100
rect 10376 21088 10382 21140
rect 10428 21100 12756 21128
rect 6365 21063 6423 21069
rect 6365 21029 6377 21063
rect 6411 21060 6423 21063
rect 8294 21060 8300 21072
rect 6411 21032 8300 21060
rect 6411 21029 6423 21032
rect 6365 21023 6423 21029
rect 8294 21020 8300 21032
rect 8352 21020 8358 21072
rect 8478 21020 8484 21072
rect 8536 21060 8542 21072
rect 9953 21063 10011 21069
rect 9953 21060 9965 21063
rect 8536 21032 9965 21060
rect 8536 21020 8542 21032
rect 9953 21029 9965 21032
rect 9999 21029 10011 21063
rect 9953 21023 10011 21029
rect 2774 20952 2780 21004
rect 2832 20952 2838 21004
rect 4154 20952 4160 21004
rect 4212 20992 4218 21004
rect 4433 20995 4491 21001
rect 4433 20992 4445 20995
rect 4212 20964 4445 20992
rect 4212 20952 4218 20964
rect 4433 20961 4445 20964
rect 4479 20961 4491 20995
rect 4433 20955 4491 20961
rect 5626 20952 5632 21004
rect 5684 20992 5690 21004
rect 5684 20964 5856 20992
rect 5684 20952 5690 20964
rect 2225 20927 2283 20933
rect 2225 20893 2237 20927
rect 2271 20893 2283 20927
rect 2225 20887 2283 20893
rect 4065 20927 4123 20933
rect 4065 20893 4077 20927
rect 4111 20924 4123 20927
rect 5718 20924 5724 20936
rect 4111 20896 5724 20924
rect 4111 20893 4123 20896
rect 4065 20887 4123 20893
rect 2240 20788 2268 20887
rect 5718 20884 5724 20896
rect 5776 20884 5782 20936
rect 5828 20924 5856 20964
rect 6914 20952 6920 21004
rect 6972 20992 6978 21004
rect 7377 20995 7435 21001
rect 7377 20992 7389 20995
rect 6972 20964 7389 20992
rect 6972 20952 6978 20964
rect 7377 20961 7389 20964
rect 7423 20961 7435 20995
rect 7377 20955 7435 20961
rect 8202 20952 8208 21004
rect 8260 20992 8266 21004
rect 10428 21001 10456 21100
rect 12452 21032 12664 21060
rect 8665 20995 8723 21001
rect 8665 20992 8677 20995
rect 8260 20964 8677 20992
rect 8260 20952 8266 20964
rect 8665 20961 8677 20964
rect 8711 20961 8723 20995
rect 8665 20955 8723 20961
rect 10413 20995 10471 21001
rect 10413 20961 10425 20995
rect 10459 20961 10471 20995
rect 10413 20955 10471 20961
rect 10502 20952 10508 21004
rect 10560 20952 10566 21004
rect 11054 20952 11060 21004
rect 11112 20992 11118 21004
rect 11149 20995 11207 21001
rect 11149 20992 11161 20995
rect 11112 20964 11161 20992
rect 11112 20952 11118 20964
rect 11149 20961 11161 20964
rect 11195 20961 11207 20995
rect 11149 20955 11207 20961
rect 11422 20952 11428 21004
rect 11480 20992 11486 21004
rect 12452 20992 12480 21032
rect 11480 20964 12480 20992
rect 11480 20952 11486 20964
rect 5997 20927 6055 20933
rect 5997 20924 6009 20927
rect 5828 20896 6009 20924
rect 5997 20893 6009 20896
rect 6043 20893 6055 20927
rect 5997 20887 6055 20893
rect 7098 20884 7104 20936
rect 7156 20884 7162 20936
rect 7742 20884 7748 20936
rect 7800 20924 7806 20936
rect 10321 20927 10379 20933
rect 10321 20924 10333 20927
rect 7800 20896 10333 20924
rect 7800 20884 7806 20896
rect 10321 20893 10333 20896
rect 10367 20893 10379 20927
rect 12636 20924 12664 21032
rect 12728 20992 12756 21100
rect 12802 21088 12808 21140
rect 12860 21128 12866 21140
rect 12897 21131 12955 21137
rect 12897 21128 12909 21131
rect 12860 21100 12909 21128
rect 12860 21088 12866 21100
rect 12897 21097 12909 21100
rect 12943 21097 12955 21131
rect 12897 21091 12955 21097
rect 13446 21088 13452 21140
rect 13504 21128 13510 21140
rect 13504 21100 16068 21128
rect 13504 21088 13510 21100
rect 13722 21020 13728 21072
rect 13780 21060 13786 21072
rect 15378 21060 15384 21072
rect 13780 21032 15384 21060
rect 13780 21020 13786 21032
rect 15378 21020 15384 21032
rect 15436 21020 15442 21072
rect 15473 21063 15531 21069
rect 15473 21029 15485 21063
rect 15519 21029 15531 21063
rect 15473 21023 15531 21029
rect 15488 20992 15516 21023
rect 12728 20964 15516 20992
rect 15838 20952 15844 21004
rect 15896 20992 15902 21004
rect 16040 21001 16068 21100
rect 16574 21088 16580 21140
rect 16632 21128 16638 21140
rect 16669 21131 16727 21137
rect 16669 21128 16681 21131
rect 16632 21100 16681 21128
rect 16632 21088 16638 21100
rect 16669 21097 16681 21100
rect 16715 21097 16727 21131
rect 24581 21131 24639 21137
rect 24581 21128 24593 21131
rect 16669 21091 16727 21097
rect 18340 21100 24593 21128
rect 16942 21020 16948 21072
rect 17000 21060 17006 21072
rect 18230 21060 18236 21072
rect 17000 21032 18236 21060
rect 17000 21020 17006 21032
rect 18230 21020 18236 21032
rect 18288 21020 18294 21072
rect 15933 20995 15991 21001
rect 15933 20992 15945 20995
rect 15896 20964 15945 20992
rect 15896 20952 15902 20964
rect 15933 20961 15945 20964
rect 15979 20961 15991 20995
rect 15933 20955 15991 20961
rect 16025 20995 16083 21001
rect 16025 20961 16037 20995
rect 16071 20961 16083 20995
rect 16025 20955 16083 20961
rect 16206 20952 16212 21004
rect 16264 20992 16270 21004
rect 18340 21001 18368 21100
rect 24581 21097 24593 21100
rect 24627 21097 24639 21131
rect 24581 21091 24639 21097
rect 18598 21020 18604 21072
rect 18656 21060 18662 21072
rect 18877 21063 18935 21069
rect 18877 21060 18889 21063
rect 18656 21032 18889 21060
rect 18656 21020 18662 21032
rect 18877 21029 18889 21032
rect 18923 21029 18935 21063
rect 18877 21023 18935 21029
rect 20714 21020 20720 21072
rect 20772 21060 20778 21072
rect 21174 21060 21180 21072
rect 20772 21032 21180 21060
rect 20772 21020 20778 21032
rect 21174 21020 21180 21032
rect 21232 21020 21238 21072
rect 21637 21063 21695 21069
rect 21637 21029 21649 21063
rect 21683 21060 21695 21063
rect 22278 21060 22284 21072
rect 21683 21032 22284 21060
rect 21683 21029 21695 21032
rect 21637 21023 21695 21029
rect 22278 21020 22284 21032
rect 22336 21020 22342 21072
rect 22646 21020 22652 21072
rect 22704 21060 22710 21072
rect 22704 21032 23428 21060
rect 22704 21020 22710 21032
rect 17129 20995 17187 21001
rect 17129 20992 17141 20995
rect 16264 20964 17141 20992
rect 16264 20952 16270 20964
rect 17129 20961 17141 20964
rect 17175 20961 17187 20995
rect 17129 20955 17187 20961
rect 17221 20995 17279 21001
rect 17221 20961 17233 20995
rect 17267 20961 17279 20995
rect 17221 20955 17279 20961
rect 18325 20995 18383 21001
rect 18325 20961 18337 20995
rect 18371 20961 18383 20995
rect 18325 20955 18383 20961
rect 18509 20995 18567 21001
rect 18509 20961 18521 20995
rect 18555 20992 18567 20995
rect 18690 20992 18696 21004
rect 18555 20964 18696 20992
rect 18555 20961 18567 20964
rect 18509 20955 18567 20961
rect 13354 20924 13360 20936
rect 12636 20896 13360 20924
rect 10321 20887 10379 20893
rect 13354 20884 13360 20896
rect 13412 20884 13418 20936
rect 14369 20927 14427 20933
rect 14369 20893 14381 20927
rect 14415 20924 14427 20927
rect 14458 20924 14464 20936
rect 14415 20896 14464 20924
rect 14415 20893 14427 20896
rect 14369 20887 14427 20893
rect 14458 20884 14464 20896
rect 14516 20884 14522 20936
rect 14550 20884 14556 20936
rect 14608 20924 14614 20936
rect 17236 20924 17264 20955
rect 18690 20952 18696 20964
rect 18748 20992 18754 21004
rect 19705 20995 19763 21001
rect 19705 20992 19717 20995
rect 18748 20964 19717 20992
rect 18748 20952 18754 20964
rect 19705 20961 19717 20964
rect 19751 20961 19763 20995
rect 21542 20992 21548 21004
rect 19705 20955 19763 20961
rect 20824 20964 21548 20992
rect 14608 20896 17264 20924
rect 14608 20884 14614 20896
rect 19334 20884 19340 20936
rect 19392 20924 19398 20936
rect 19429 20927 19487 20933
rect 19429 20924 19441 20927
rect 19392 20896 19441 20924
rect 19392 20884 19398 20896
rect 19429 20893 19441 20896
rect 19475 20893 19487 20927
rect 19429 20887 19487 20893
rect 20714 20884 20720 20936
rect 20772 20924 20778 20936
rect 20824 20924 20852 20964
rect 21542 20952 21548 20964
rect 21600 20952 21606 21004
rect 22002 20952 22008 21004
rect 22060 20992 22066 21004
rect 22189 20995 22247 21001
rect 22189 20992 22201 20995
rect 22060 20964 22201 20992
rect 22060 20952 22066 20964
rect 22189 20961 22201 20964
rect 22235 20961 22247 20995
rect 22189 20955 22247 20961
rect 22830 20952 22836 21004
rect 22888 20992 22894 21004
rect 23400 21001 23428 21032
rect 23658 21020 23664 21072
rect 23716 21060 23722 21072
rect 23937 21063 23995 21069
rect 23937 21060 23949 21063
rect 23716 21032 23949 21060
rect 23716 21020 23722 21032
rect 23937 21029 23949 21032
rect 23983 21060 23995 21063
rect 24118 21060 24124 21072
rect 23983 21032 24124 21060
rect 23983 21029 23995 21032
rect 23937 21023 23995 21029
rect 24118 21020 24124 21032
rect 24176 21020 24182 21072
rect 23293 20995 23351 21001
rect 23293 20992 23305 20995
rect 22888 20964 23305 20992
rect 22888 20952 22894 20964
rect 23293 20961 23305 20964
rect 23339 20961 23351 20995
rect 23293 20955 23351 20961
rect 23385 20995 23443 21001
rect 23385 20961 23397 20995
rect 23431 20961 23443 20995
rect 23385 20955 23443 20961
rect 25130 20952 25136 21004
rect 25188 20952 25194 21004
rect 20772 20910 20852 20924
rect 20772 20896 20838 20910
rect 20772 20884 20778 20896
rect 20990 20884 20996 20936
rect 21048 20924 21054 20936
rect 21048 20896 22968 20924
rect 21048 20884 21054 20896
rect 8294 20856 8300 20868
rect 2746 20828 8300 20856
rect 2746 20788 2774 20828
rect 8294 20816 8300 20828
rect 8352 20816 8358 20868
rect 8754 20856 8760 20868
rect 8588 20828 8760 20856
rect 2240 20760 2774 20788
rect 5813 20791 5871 20797
rect 5813 20757 5825 20791
rect 5859 20788 5871 20791
rect 6178 20788 6184 20800
rect 5859 20760 6184 20788
rect 5859 20757 5871 20760
rect 5813 20751 5871 20757
rect 6178 20748 6184 20760
rect 6236 20748 6242 20800
rect 6641 20791 6699 20797
rect 6641 20757 6653 20791
rect 6687 20788 6699 20791
rect 8588 20788 8616 20828
rect 8754 20816 8760 20828
rect 8812 20816 8818 20868
rect 9309 20859 9367 20865
rect 9309 20825 9321 20859
rect 9355 20856 9367 20859
rect 9355 20828 10916 20856
rect 9355 20825 9367 20828
rect 9309 20819 9367 20825
rect 6687 20760 8616 20788
rect 6687 20757 6699 20760
rect 6641 20751 6699 20757
rect 8938 20748 8944 20800
rect 8996 20748 9002 20800
rect 10888 20788 10916 20828
rect 11882 20816 11888 20868
rect 11940 20816 11946 20868
rect 13541 20859 13599 20865
rect 13541 20825 13553 20859
rect 13587 20856 13599 20859
rect 13998 20856 14004 20868
rect 13587 20828 14004 20856
rect 13587 20825 13599 20828
rect 13541 20819 13599 20825
rect 13998 20816 14004 20828
rect 14056 20816 14062 20868
rect 14090 20816 14096 20868
rect 14148 20856 14154 20868
rect 15286 20856 15292 20868
rect 14148 20828 15292 20856
rect 14148 20816 14154 20828
rect 15286 20816 15292 20828
rect 15344 20816 15350 20868
rect 15378 20816 15384 20868
rect 15436 20856 15442 20868
rect 18233 20859 18291 20865
rect 15436 20828 17908 20856
rect 15436 20816 15442 20828
rect 12434 20788 12440 20800
rect 10888 20760 12440 20788
rect 12434 20748 12440 20760
rect 12492 20748 12498 20800
rect 12802 20748 12808 20800
rect 12860 20788 12866 20800
rect 13633 20791 13691 20797
rect 13633 20788 13645 20791
rect 12860 20760 13645 20788
rect 12860 20748 12866 20760
rect 13633 20757 13645 20760
rect 13679 20757 13691 20791
rect 13633 20751 13691 20757
rect 13722 20748 13728 20800
rect 13780 20788 13786 20800
rect 14461 20791 14519 20797
rect 14461 20788 14473 20791
rect 13780 20760 14473 20788
rect 13780 20748 13786 20760
rect 14461 20757 14473 20760
rect 14507 20757 14519 20791
rect 14461 20751 14519 20757
rect 14826 20748 14832 20800
rect 14884 20788 14890 20800
rect 15013 20791 15071 20797
rect 15013 20788 15025 20791
rect 14884 20760 15025 20788
rect 14884 20748 14890 20760
rect 15013 20757 15025 20760
rect 15059 20757 15071 20791
rect 15013 20751 15071 20757
rect 15838 20748 15844 20800
rect 15896 20748 15902 20800
rect 17034 20748 17040 20800
rect 17092 20748 17098 20800
rect 17880 20797 17908 20828
rect 18233 20825 18245 20859
rect 18279 20856 18291 20859
rect 18966 20856 18972 20868
rect 18279 20828 18972 20856
rect 18279 20825 18291 20828
rect 18233 20819 18291 20825
rect 18966 20816 18972 20828
rect 19024 20816 19030 20868
rect 22940 20856 22968 20896
rect 23198 20884 23204 20936
rect 23256 20884 23262 20936
rect 25041 20859 25099 20865
rect 25041 20856 25053 20859
rect 21100 20828 22876 20856
rect 22940 20828 25053 20856
rect 17865 20791 17923 20797
rect 17865 20757 17877 20791
rect 17911 20757 17923 20791
rect 17865 20751 17923 20757
rect 19242 20748 19248 20800
rect 19300 20788 19306 20800
rect 21100 20788 21128 20828
rect 19300 20760 21128 20788
rect 19300 20748 19306 20760
rect 21174 20748 21180 20800
rect 21232 20788 21238 20800
rect 21910 20788 21916 20800
rect 21232 20760 21916 20788
rect 21232 20748 21238 20760
rect 21910 20748 21916 20760
rect 21968 20788 21974 20800
rect 22005 20791 22063 20797
rect 22005 20788 22017 20791
rect 21968 20760 22017 20788
rect 21968 20748 21974 20760
rect 22005 20757 22017 20760
rect 22051 20757 22063 20791
rect 22005 20751 22063 20757
rect 22094 20748 22100 20800
rect 22152 20748 22158 20800
rect 22848 20797 22876 20828
rect 25041 20825 25053 20828
rect 25087 20825 25099 20859
rect 25041 20819 25099 20825
rect 22833 20791 22891 20797
rect 22833 20757 22845 20791
rect 22879 20757 22891 20791
rect 22833 20751 22891 20757
rect 24949 20791 25007 20797
rect 24949 20757 24961 20791
rect 24995 20788 25007 20791
rect 26050 20788 26056 20800
rect 24995 20760 26056 20788
rect 24995 20757 25007 20760
rect 24949 20751 25007 20757
rect 26050 20748 26056 20760
rect 26108 20748 26114 20800
rect 1104 20698 25852 20720
rect 1104 20646 7950 20698
rect 8002 20646 8014 20698
rect 8066 20646 8078 20698
rect 8130 20646 8142 20698
rect 8194 20646 8206 20698
rect 8258 20646 17950 20698
rect 18002 20646 18014 20698
rect 18066 20646 18078 20698
rect 18130 20646 18142 20698
rect 18194 20646 18206 20698
rect 18258 20646 25852 20698
rect 1104 20624 25852 20646
rect 2225 20587 2283 20593
rect 2225 20553 2237 20587
rect 2271 20584 2283 20587
rect 3970 20584 3976 20596
rect 2271 20556 3976 20584
rect 2271 20553 2283 20556
rect 2225 20547 2283 20553
rect 3970 20544 3976 20556
rect 4028 20544 4034 20596
rect 4706 20544 4712 20596
rect 4764 20584 4770 20596
rect 4801 20587 4859 20593
rect 4801 20584 4813 20587
rect 4764 20556 4813 20584
rect 4764 20544 4770 20556
rect 4801 20553 4813 20556
rect 4847 20553 4859 20587
rect 4801 20547 4859 20553
rect 5166 20544 5172 20596
rect 5224 20544 5230 20596
rect 6546 20544 6552 20596
rect 6604 20544 6610 20596
rect 6825 20587 6883 20593
rect 6825 20553 6837 20587
rect 6871 20584 6883 20587
rect 7190 20584 7196 20596
rect 6871 20556 7196 20584
rect 6871 20553 6883 20556
rect 6825 20547 6883 20553
rect 7190 20544 7196 20556
rect 7248 20544 7254 20596
rect 7742 20544 7748 20596
rect 7800 20544 7806 20596
rect 10134 20584 10140 20596
rect 8588 20556 10140 20584
rect 5350 20516 5356 20528
rect 1780 20488 5356 20516
rect 1780 20457 1808 20488
rect 5350 20476 5356 20488
rect 5408 20476 5414 20528
rect 7208 20516 7236 20544
rect 7208 20488 8524 20516
rect 1765 20451 1823 20457
rect 1765 20417 1777 20451
rect 1811 20417 1823 20451
rect 1765 20411 1823 20417
rect 2409 20451 2467 20457
rect 2409 20417 2421 20451
rect 2455 20417 2467 20451
rect 2409 20411 2467 20417
rect 3053 20451 3111 20457
rect 3053 20417 3065 20451
rect 3099 20448 3111 20451
rect 5534 20448 5540 20460
rect 3099 20420 5540 20448
rect 3099 20417 3111 20420
rect 3053 20411 3111 20417
rect 2424 20312 2452 20411
rect 5534 20408 5540 20420
rect 5592 20408 5598 20460
rect 5997 20451 6055 20457
rect 5997 20417 6009 20451
rect 6043 20448 6055 20451
rect 7190 20448 7196 20460
rect 6043 20420 7196 20448
rect 6043 20417 6055 20420
rect 5997 20411 6055 20417
rect 7190 20408 7196 20420
rect 7248 20408 7254 20460
rect 7285 20451 7343 20457
rect 7285 20417 7297 20451
rect 7331 20417 7343 20451
rect 7285 20411 7343 20417
rect 3326 20340 3332 20392
rect 3384 20340 3390 20392
rect 6546 20380 6552 20392
rect 3988 20352 6552 20380
rect 3988 20312 4016 20352
rect 6546 20340 6552 20352
rect 6604 20340 6610 20392
rect 7006 20340 7012 20392
rect 7064 20380 7070 20392
rect 7300 20380 7328 20411
rect 7064 20352 7328 20380
rect 7064 20340 7070 20352
rect 7742 20340 7748 20392
rect 7800 20380 7806 20392
rect 8386 20380 8392 20392
rect 7800 20352 8392 20380
rect 7800 20340 7806 20352
rect 8386 20340 8392 20352
rect 8444 20340 8450 20392
rect 8496 20380 8524 20488
rect 8588 20457 8616 20556
rect 10134 20544 10140 20556
rect 10192 20544 10198 20596
rect 10318 20544 10324 20596
rect 10376 20584 10382 20596
rect 10376 20556 10732 20584
rect 10376 20544 10382 20556
rect 8938 20476 8944 20528
rect 8996 20516 9002 20528
rect 9766 20516 9772 20528
rect 8996 20488 9772 20516
rect 8996 20476 9002 20488
rect 9766 20476 9772 20488
rect 9824 20476 9830 20528
rect 8573 20451 8631 20457
rect 8573 20417 8585 20451
rect 8619 20417 8631 20451
rect 8573 20411 8631 20417
rect 9030 20408 9036 20460
rect 9088 20408 9094 20460
rect 10704 20448 10732 20556
rect 10778 20544 10784 20596
rect 10836 20584 10842 20596
rect 12342 20584 12348 20596
rect 10836 20556 12348 20584
rect 10836 20544 10842 20556
rect 12342 20544 12348 20556
rect 12400 20544 12406 20596
rect 12434 20544 12440 20596
rect 12492 20544 12498 20596
rect 12526 20544 12532 20596
rect 12584 20584 12590 20596
rect 12802 20584 12808 20596
rect 12584 20556 12808 20584
rect 12584 20544 12590 20556
rect 12802 20544 12808 20556
rect 12860 20544 12866 20596
rect 14826 20584 14832 20596
rect 13188 20556 14832 20584
rect 11146 20476 11152 20528
rect 11204 20516 11210 20528
rect 11333 20519 11391 20525
rect 11333 20516 11345 20519
rect 11204 20488 11345 20516
rect 11204 20476 11210 20488
rect 11333 20485 11345 20488
rect 11379 20516 11391 20519
rect 11609 20519 11667 20525
rect 11609 20516 11621 20519
rect 11379 20488 11621 20516
rect 11379 20485 11391 20488
rect 11333 20479 11391 20485
rect 11609 20485 11621 20488
rect 11655 20516 11667 20519
rect 11882 20516 11888 20528
rect 11655 20488 11888 20516
rect 11655 20485 11667 20488
rect 11609 20479 11667 20485
rect 11882 20476 11888 20488
rect 11940 20476 11946 20528
rect 13188 20457 13216 20556
rect 14826 20544 14832 20556
rect 14884 20584 14890 20596
rect 15378 20584 15384 20596
rect 14884 20556 15384 20584
rect 14884 20544 14890 20556
rect 15378 20544 15384 20556
rect 15436 20544 15442 20596
rect 18598 20584 18604 20596
rect 17604 20556 18604 20584
rect 13817 20519 13875 20525
rect 13817 20485 13829 20519
rect 13863 20516 13875 20519
rect 14090 20516 14096 20528
rect 13863 20488 14096 20516
rect 13863 20485 13875 20488
rect 13817 20479 13875 20485
rect 14090 20476 14096 20488
rect 14148 20476 14154 20528
rect 15286 20516 15292 20528
rect 15042 20488 15292 20516
rect 15286 20476 15292 20488
rect 15344 20516 15350 20528
rect 16301 20519 16359 20525
rect 16301 20516 16313 20519
rect 15344 20488 16313 20516
rect 15344 20476 15350 20488
rect 16301 20485 16313 20488
rect 16347 20485 16359 20519
rect 16301 20479 16359 20485
rect 16758 20476 16764 20528
rect 16816 20516 16822 20528
rect 17604 20516 17632 20556
rect 16816 20488 17710 20516
rect 16816 20476 16822 20488
rect 18340 20460 18368 20556
rect 18598 20544 18604 20556
rect 18656 20544 18662 20596
rect 18690 20544 18696 20596
rect 18748 20544 18754 20596
rect 18800 20556 20852 20584
rect 13173 20451 13231 20457
rect 13173 20448 13185 20451
rect 10704 20420 13185 20448
rect 13173 20417 13185 20420
rect 13219 20417 13231 20451
rect 13173 20411 13231 20417
rect 13541 20451 13599 20457
rect 13541 20417 13553 20451
rect 13587 20417 13599 20451
rect 13541 20411 13599 20417
rect 8938 20380 8944 20392
rect 8496 20352 8944 20380
rect 8938 20340 8944 20352
rect 8996 20340 9002 20392
rect 9309 20383 9367 20389
rect 9309 20349 9321 20383
rect 9355 20380 9367 20383
rect 10502 20380 10508 20392
rect 9355 20352 10508 20380
rect 9355 20349 9367 20352
rect 9309 20343 9367 20349
rect 10502 20340 10508 20352
rect 10560 20340 10566 20392
rect 11793 20383 11851 20389
rect 10704 20352 11652 20380
rect 5166 20312 5172 20324
rect 2424 20284 4016 20312
rect 4080 20284 5172 20312
rect 1581 20247 1639 20253
rect 1581 20213 1593 20247
rect 1627 20244 1639 20247
rect 4080 20244 4108 20284
rect 5166 20272 5172 20284
rect 5224 20272 5230 20324
rect 1627 20216 4108 20244
rect 1627 20213 1639 20216
rect 1581 20207 1639 20213
rect 4154 20204 4160 20256
rect 4212 20244 4218 20256
rect 5813 20247 5871 20253
rect 5813 20244 5825 20247
rect 4212 20216 5825 20244
rect 4212 20204 4218 20216
rect 5813 20213 5825 20216
rect 5859 20213 5871 20247
rect 5813 20207 5871 20213
rect 6822 20204 6828 20256
rect 6880 20244 6886 20256
rect 7101 20247 7159 20253
rect 7101 20244 7113 20247
rect 6880 20216 7113 20244
rect 6880 20204 6886 20216
rect 7101 20213 7113 20216
rect 7147 20213 7159 20247
rect 7101 20207 7159 20213
rect 8386 20204 8392 20256
rect 8444 20204 8450 20256
rect 9398 20204 9404 20256
rect 9456 20244 9462 20256
rect 10704 20244 10732 20352
rect 9456 20216 10732 20244
rect 9456 20204 9462 20216
rect 10778 20204 10784 20256
rect 10836 20204 10842 20256
rect 11624 20244 11652 20352
rect 11793 20349 11805 20383
rect 11839 20380 11851 20383
rect 12158 20380 12164 20392
rect 11839 20352 12164 20380
rect 11839 20349 11851 20352
rect 11793 20343 11851 20349
rect 12158 20340 12164 20352
rect 12216 20340 12222 20392
rect 12529 20383 12587 20389
rect 12529 20380 12541 20383
rect 12452 20352 12541 20380
rect 12452 20312 12480 20352
rect 12529 20349 12541 20352
rect 12575 20349 12587 20383
rect 12529 20343 12587 20349
rect 12713 20383 12771 20389
rect 12713 20349 12725 20383
rect 12759 20380 12771 20383
rect 12802 20380 12808 20392
rect 12759 20352 12808 20380
rect 12759 20349 12771 20352
rect 12713 20343 12771 20349
rect 12802 20340 12808 20352
rect 12860 20340 12866 20392
rect 13556 20380 13584 20411
rect 15838 20408 15844 20460
rect 15896 20408 15902 20460
rect 18322 20408 18328 20460
rect 18380 20408 18386 20460
rect 13814 20380 13820 20392
rect 13556 20352 13820 20380
rect 13446 20312 13452 20324
rect 12452 20284 13452 20312
rect 13446 20272 13452 20284
rect 13504 20272 13510 20324
rect 12069 20247 12127 20253
rect 12069 20244 12081 20247
rect 11624 20216 12081 20244
rect 12069 20213 12081 20216
rect 12115 20213 12127 20247
rect 12069 20207 12127 20213
rect 12250 20204 12256 20256
rect 12308 20244 12314 20256
rect 13556 20244 13584 20352
rect 13814 20340 13820 20352
rect 13872 20380 13878 20392
rect 16482 20380 16488 20392
rect 13872 20352 16488 20380
rect 13872 20340 13878 20352
rect 16482 20340 16488 20352
rect 16540 20380 16546 20392
rect 16945 20383 17003 20389
rect 16945 20380 16957 20383
rect 16540 20352 16957 20380
rect 16540 20340 16546 20352
rect 16945 20349 16957 20352
rect 16991 20349 17003 20383
rect 16945 20343 17003 20349
rect 17218 20340 17224 20392
rect 17276 20380 17282 20392
rect 18800 20380 18828 20556
rect 20824 20516 20852 20556
rect 20898 20544 20904 20596
rect 20956 20584 20962 20596
rect 20993 20587 21051 20593
rect 20993 20584 21005 20587
rect 20956 20556 21005 20584
rect 20956 20544 20962 20556
rect 20993 20553 21005 20556
rect 21039 20553 21051 20587
rect 25130 20584 25136 20596
rect 20993 20547 21051 20553
rect 21100 20556 25136 20584
rect 21100 20516 21128 20556
rect 25130 20544 25136 20556
rect 25188 20544 25194 20596
rect 20824 20488 21128 20516
rect 22462 20476 22468 20528
rect 22520 20476 22526 20528
rect 23201 20519 23259 20525
rect 23201 20485 23213 20519
rect 23247 20516 23259 20519
rect 23658 20516 23664 20528
rect 23247 20488 23664 20516
rect 23247 20485 23259 20488
rect 23201 20479 23259 20485
rect 23658 20476 23664 20488
rect 23716 20476 23722 20528
rect 23753 20519 23811 20525
rect 23753 20485 23765 20519
rect 23799 20516 23811 20519
rect 23842 20516 23848 20528
rect 23799 20488 23848 20516
rect 23799 20485 23811 20488
rect 23753 20479 23811 20485
rect 23842 20476 23848 20488
rect 23900 20476 23906 20528
rect 24210 20476 24216 20528
rect 24268 20476 24274 20528
rect 20622 20408 20628 20460
rect 20680 20408 20686 20460
rect 22557 20451 22615 20457
rect 22557 20417 22569 20451
rect 22603 20448 22615 20451
rect 22603 20420 23244 20448
rect 22603 20417 22615 20420
rect 22557 20411 22615 20417
rect 17276 20352 18828 20380
rect 17276 20340 17282 20352
rect 19242 20340 19248 20392
rect 19300 20340 19306 20392
rect 19521 20383 19579 20389
rect 19521 20349 19533 20383
rect 19567 20380 19579 20383
rect 19886 20380 19892 20392
rect 19567 20352 19892 20380
rect 19567 20349 19579 20352
rect 19521 20343 19579 20349
rect 19886 20340 19892 20352
rect 19944 20340 19950 20392
rect 20806 20340 20812 20392
rect 20864 20380 20870 20392
rect 20864 20352 21588 20380
rect 20864 20340 20870 20352
rect 14826 20272 14832 20324
rect 14884 20312 14890 20324
rect 14884 20284 16068 20312
rect 14884 20272 14890 20284
rect 12308 20216 13584 20244
rect 12308 20204 12314 20216
rect 13630 20204 13636 20256
rect 13688 20244 13694 20256
rect 15289 20247 15347 20253
rect 15289 20244 15301 20247
rect 13688 20216 15301 20244
rect 13688 20204 13694 20216
rect 15289 20213 15301 20216
rect 15335 20213 15347 20247
rect 15289 20207 15347 20213
rect 15930 20204 15936 20256
rect 15988 20204 15994 20256
rect 16040 20244 16068 20284
rect 20898 20272 20904 20324
rect 20956 20312 20962 20324
rect 21453 20315 21511 20321
rect 21453 20312 21465 20315
rect 20956 20284 21465 20312
rect 20956 20272 20962 20284
rect 21453 20281 21465 20284
rect 21499 20281 21511 20315
rect 21560 20312 21588 20352
rect 22646 20340 22652 20392
rect 22704 20340 22710 20392
rect 23216 20380 23244 20420
rect 23290 20408 23296 20460
rect 23348 20448 23354 20460
rect 23477 20451 23535 20457
rect 23477 20448 23489 20451
rect 23348 20420 23489 20448
rect 23348 20408 23354 20420
rect 23477 20417 23489 20420
rect 23523 20417 23535 20451
rect 23477 20411 23535 20417
rect 24118 20380 24124 20392
rect 23216 20352 24124 20380
rect 24118 20340 24124 20352
rect 24176 20380 24182 20392
rect 24762 20380 24768 20392
rect 24176 20352 24768 20380
rect 24176 20340 24182 20352
rect 24762 20340 24768 20352
rect 24820 20340 24826 20392
rect 21560 20284 22968 20312
rect 21453 20275 21511 20281
rect 18598 20244 18604 20256
rect 16040 20216 18604 20244
rect 18598 20204 18604 20216
rect 18656 20204 18662 20256
rect 19610 20204 19616 20256
rect 19668 20244 19674 20256
rect 20530 20244 20536 20256
rect 19668 20216 20536 20244
rect 19668 20204 19674 20216
rect 20530 20204 20536 20216
rect 20588 20244 20594 20256
rect 21269 20247 21327 20253
rect 21269 20244 21281 20247
rect 20588 20216 21281 20244
rect 20588 20204 20594 20216
rect 21269 20213 21281 20216
rect 21315 20213 21327 20247
rect 21269 20207 21327 20213
rect 22097 20247 22155 20253
rect 22097 20213 22109 20247
rect 22143 20244 22155 20247
rect 22830 20244 22836 20256
rect 22143 20216 22836 20244
rect 22143 20213 22155 20216
rect 22097 20207 22155 20213
rect 22830 20204 22836 20216
rect 22888 20204 22894 20256
rect 22940 20244 22968 20284
rect 23934 20244 23940 20256
rect 22940 20216 23940 20244
rect 23934 20204 23940 20216
rect 23992 20204 23998 20256
rect 25222 20204 25228 20256
rect 25280 20204 25286 20256
rect 1104 20154 25852 20176
rect 1104 20102 2950 20154
rect 3002 20102 3014 20154
rect 3066 20102 3078 20154
rect 3130 20102 3142 20154
rect 3194 20102 3206 20154
rect 3258 20102 12950 20154
rect 13002 20102 13014 20154
rect 13066 20102 13078 20154
rect 13130 20102 13142 20154
rect 13194 20102 13206 20154
rect 13258 20102 22950 20154
rect 23002 20102 23014 20154
rect 23066 20102 23078 20154
rect 23130 20102 23142 20154
rect 23194 20102 23206 20154
rect 23258 20102 25852 20154
rect 1104 20080 25852 20102
rect 3970 20000 3976 20052
rect 4028 20040 4034 20052
rect 4028 20012 7144 20040
rect 4028 20000 4034 20012
rect 4525 19975 4583 19981
rect 4525 19941 4537 19975
rect 4571 19972 4583 19975
rect 4571 19944 7052 19972
rect 4571 19941 4583 19944
rect 4525 19935 4583 19941
rect 2038 19864 2044 19916
rect 2096 19904 2102 19916
rect 2501 19907 2559 19913
rect 2501 19904 2513 19907
rect 2096 19876 2513 19904
rect 2096 19864 2102 19876
rect 2501 19873 2513 19876
rect 2547 19873 2559 19907
rect 2501 19867 2559 19873
rect 5258 19864 5264 19916
rect 5316 19904 5322 19916
rect 5445 19907 5503 19913
rect 5445 19904 5457 19907
rect 5316 19876 5457 19904
rect 5316 19864 5322 19876
rect 5445 19873 5457 19876
rect 5491 19873 5503 19907
rect 5445 19867 5503 19873
rect 2225 19839 2283 19845
rect 2225 19805 2237 19839
rect 2271 19805 2283 19839
rect 2225 19799 2283 19805
rect 2240 19768 2268 19799
rect 4706 19796 4712 19848
rect 4764 19796 4770 19848
rect 5169 19839 5227 19845
rect 5169 19805 5181 19839
rect 5215 19836 5227 19839
rect 5810 19836 5816 19848
rect 5215 19808 5816 19836
rect 5215 19805 5227 19808
rect 5169 19799 5227 19805
rect 5810 19796 5816 19808
rect 5868 19796 5874 19848
rect 6638 19796 6644 19848
rect 6696 19796 6702 19848
rect 7024 19836 7052 19944
rect 7116 19913 7144 20012
rect 7190 20000 7196 20052
rect 7248 20040 7254 20052
rect 10413 20043 10471 20049
rect 10413 20040 10425 20043
rect 7248 20012 10425 20040
rect 7248 20000 7254 20012
rect 10413 20009 10425 20012
rect 10459 20009 10471 20043
rect 14921 20043 14979 20049
rect 14921 20040 14933 20043
rect 10413 20003 10471 20009
rect 10888 20012 14933 20040
rect 7101 19907 7159 19913
rect 7101 19873 7113 19907
rect 7147 19873 7159 19907
rect 7101 19867 7159 19873
rect 7377 19907 7435 19913
rect 7377 19873 7389 19907
rect 7423 19904 7435 19907
rect 7466 19904 7472 19916
rect 7423 19876 7472 19904
rect 7423 19873 7435 19876
rect 7377 19867 7435 19873
rect 7466 19864 7472 19876
rect 7524 19864 7530 19916
rect 10888 19913 10916 20012
rect 14921 20009 14933 20012
rect 14967 20009 14979 20043
rect 14921 20003 14979 20009
rect 15194 20000 15200 20052
rect 15252 20040 15258 20052
rect 17129 20043 17187 20049
rect 17129 20040 17141 20043
rect 15252 20012 17141 20040
rect 15252 20000 15258 20012
rect 17129 20009 17141 20012
rect 17175 20009 17187 20043
rect 17129 20003 17187 20009
rect 18322 20000 18328 20052
rect 18380 20040 18386 20052
rect 20622 20040 20628 20052
rect 18380 20012 20628 20040
rect 18380 20000 18386 20012
rect 20622 20000 20628 20012
rect 20680 20000 20686 20052
rect 20717 20043 20775 20049
rect 20717 20009 20729 20043
rect 20763 20040 20775 20043
rect 21082 20040 21088 20052
rect 20763 20012 21088 20040
rect 20763 20009 20775 20012
rect 20717 20003 20775 20009
rect 21082 20000 21088 20012
rect 21140 20000 21146 20052
rect 23382 20040 23388 20052
rect 21192 20012 23388 20040
rect 13354 19932 13360 19984
rect 13412 19932 13418 19984
rect 13446 19932 13452 19984
rect 13504 19972 13510 19984
rect 17681 19975 17739 19981
rect 17681 19972 17693 19975
rect 13504 19944 17693 19972
rect 13504 19932 13510 19944
rect 17681 19941 17693 19944
rect 17727 19941 17739 19975
rect 17681 19935 17739 19941
rect 17788 19944 18368 19972
rect 10873 19907 10931 19913
rect 10873 19873 10885 19907
rect 10919 19873 10931 19907
rect 10873 19867 10931 19873
rect 10962 19864 10968 19916
rect 11020 19864 11026 19916
rect 11609 19907 11667 19913
rect 11609 19873 11621 19907
rect 11655 19904 11667 19907
rect 12250 19904 12256 19916
rect 11655 19876 12256 19904
rect 11655 19873 11667 19876
rect 11609 19867 11667 19873
rect 12250 19864 12256 19876
rect 12308 19864 12314 19916
rect 12342 19864 12348 19916
rect 12400 19904 12406 19916
rect 15473 19907 15531 19913
rect 15473 19904 15485 19907
rect 12400 19876 15485 19904
rect 12400 19864 12406 19876
rect 15473 19873 15485 19876
rect 15519 19873 15531 19907
rect 15473 19867 15531 19873
rect 15654 19864 15660 19916
rect 15712 19904 15718 19916
rect 17788 19904 17816 19944
rect 15712 19876 17816 19904
rect 15712 19864 15718 19876
rect 17954 19864 17960 19916
rect 18012 19904 18018 19916
rect 18233 19907 18291 19913
rect 18233 19904 18245 19907
rect 18012 19876 18245 19904
rect 18012 19864 18018 19876
rect 18233 19873 18245 19876
rect 18279 19873 18291 19907
rect 18340 19904 18368 19944
rect 18598 19932 18604 19984
rect 18656 19972 18662 19984
rect 21192 19972 21220 20012
rect 23382 20000 23388 20012
rect 23440 20000 23446 20052
rect 23934 20000 23940 20052
rect 23992 20040 23998 20052
rect 24210 20040 24216 20052
rect 23992 20012 24216 20040
rect 23992 20000 23998 20012
rect 24210 20000 24216 20012
rect 24268 20000 24274 20052
rect 18656 19944 21220 19972
rect 18656 19932 18662 19944
rect 20073 19907 20131 19913
rect 20073 19904 20085 19907
rect 18340 19876 20085 19904
rect 18233 19867 18291 19873
rect 20073 19873 20085 19876
rect 20119 19904 20131 19907
rect 20898 19904 20904 19916
rect 20119 19876 20904 19904
rect 20119 19873 20131 19876
rect 20073 19867 20131 19873
rect 20898 19864 20904 19876
rect 20956 19864 20962 19916
rect 21085 19907 21143 19913
rect 21085 19873 21097 19907
rect 21131 19904 21143 19907
rect 23290 19904 23296 19916
rect 21131 19876 23296 19904
rect 21131 19873 21143 19876
rect 21085 19867 21143 19873
rect 23290 19864 23296 19876
rect 23348 19864 23354 19916
rect 23937 19907 23995 19913
rect 23937 19873 23949 19907
rect 23983 19904 23995 19907
rect 24486 19904 24492 19916
rect 23983 19876 24492 19904
rect 23983 19873 23995 19876
rect 23937 19867 23995 19873
rect 24486 19864 24492 19876
rect 24544 19864 24550 19916
rect 25038 19864 25044 19916
rect 25096 19864 25102 19916
rect 25225 19907 25283 19913
rect 25225 19873 25237 19907
rect 25271 19904 25283 19907
rect 25958 19904 25964 19916
rect 25271 19876 25964 19904
rect 25271 19873 25283 19876
rect 25225 19867 25283 19873
rect 25958 19864 25964 19876
rect 26016 19864 26022 19916
rect 11054 19836 11060 19848
rect 7024 19808 11060 19836
rect 11054 19796 11060 19808
rect 11112 19796 11118 19848
rect 13909 19839 13967 19845
rect 13909 19836 13921 19839
rect 13018 19808 13921 19836
rect 13909 19805 13921 19808
rect 13955 19836 13967 19839
rect 14090 19836 14096 19848
rect 13955 19808 14096 19836
rect 13955 19805 13967 19808
rect 13909 19799 13967 19805
rect 14090 19796 14096 19808
rect 14148 19796 14154 19848
rect 14182 19796 14188 19848
rect 14240 19836 14246 19848
rect 14277 19839 14335 19845
rect 14277 19836 14289 19839
rect 14240 19808 14289 19836
rect 14240 19796 14246 19808
rect 14277 19805 14289 19808
rect 14323 19805 14335 19839
rect 14277 19799 14335 19805
rect 15102 19796 15108 19848
rect 15160 19836 15166 19848
rect 18414 19836 18420 19848
rect 15160 19808 18420 19836
rect 15160 19796 15166 19808
rect 18414 19796 18420 19808
rect 18472 19796 18478 19848
rect 18874 19796 18880 19848
rect 18932 19796 18938 19848
rect 19702 19796 19708 19848
rect 19760 19836 19766 19848
rect 20441 19839 20499 19845
rect 20441 19836 20453 19839
rect 19760 19808 20453 19836
rect 19760 19796 19766 19808
rect 20441 19805 20453 19808
rect 20487 19805 20499 19839
rect 20441 19799 20499 19805
rect 23661 19839 23719 19845
rect 23661 19805 23673 19839
rect 23707 19836 23719 19839
rect 24026 19836 24032 19848
rect 23707 19808 24032 19836
rect 23707 19805 23719 19808
rect 23661 19799 23719 19805
rect 24026 19796 24032 19808
rect 24084 19796 24090 19848
rect 8294 19768 8300 19780
rect 2240 19740 8300 19768
rect 8294 19728 8300 19740
rect 8352 19728 8358 19780
rect 8389 19771 8447 19777
rect 8389 19737 8401 19771
rect 8435 19768 8447 19771
rect 10781 19771 10839 19777
rect 10781 19768 10793 19771
rect 8435 19740 10793 19768
rect 8435 19737 8447 19740
rect 8389 19731 8447 19737
rect 10781 19737 10793 19740
rect 10827 19737 10839 19771
rect 10781 19731 10839 19737
rect 11892 19771 11950 19777
rect 11892 19737 11904 19771
rect 11938 19737 11950 19771
rect 11892 19731 11950 19737
rect 13633 19771 13691 19777
rect 13633 19737 13645 19771
rect 13679 19768 13691 19771
rect 13722 19768 13728 19780
rect 13679 19740 13728 19768
rect 13679 19737 13691 19740
rect 13633 19731 13691 19737
rect 5534 19660 5540 19712
rect 5592 19700 5598 19712
rect 6457 19703 6515 19709
rect 6457 19700 6469 19703
rect 5592 19672 6469 19700
rect 5592 19660 5598 19672
rect 6457 19669 6469 19672
rect 6503 19669 6515 19703
rect 6457 19663 6515 19669
rect 7006 19660 7012 19712
rect 7064 19700 7070 19712
rect 7466 19700 7472 19712
rect 7064 19672 7472 19700
rect 7064 19660 7070 19672
rect 7466 19660 7472 19672
rect 7524 19660 7530 19712
rect 9122 19660 9128 19712
rect 9180 19660 9186 19712
rect 9769 19703 9827 19709
rect 9769 19669 9781 19703
rect 9815 19700 9827 19703
rect 10870 19700 10876 19712
rect 9815 19672 10876 19700
rect 9815 19669 9827 19672
rect 9769 19663 9827 19669
rect 10870 19660 10876 19672
rect 10928 19660 10934 19712
rect 11514 19660 11520 19712
rect 11572 19700 11578 19712
rect 11790 19700 11796 19712
rect 11572 19672 11796 19700
rect 11572 19660 11578 19672
rect 11790 19660 11796 19672
rect 11848 19660 11854 19712
rect 11907 19700 11935 19731
rect 13722 19728 13728 19740
rect 13780 19728 13786 19780
rect 14550 19768 14556 19780
rect 13832 19740 14556 19768
rect 13832 19700 13860 19740
rect 14550 19728 14556 19740
rect 14608 19728 14614 19780
rect 14642 19728 14648 19780
rect 14700 19768 14706 19780
rect 14826 19768 14832 19780
rect 14700 19740 14832 19768
rect 14700 19728 14706 19740
rect 14826 19728 14832 19740
rect 14884 19728 14890 19780
rect 15010 19728 15016 19780
rect 15068 19768 15074 19780
rect 15378 19768 15384 19780
rect 15068 19740 15384 19768
rect 15068 19728 15074 19740
rect 15378 19728 15384 19740
rect 15436 19728 15442 19780
rect 16206 19728 16212 19780
rect 16264 19728 16270 19780
rect 16758 19728 16764 19780
rect 16816 19768 16822 19780
rect 17037 19771 17095 19777
rect 17037 19768 17049 19771
rect 16816 19740 17049 19768
rect 16816 19728 16822 19740
rect 17037 19737 17049 19740
rect 17083 19737 17095 19771
rect 17037 19731 17095 19737
rect 18141 19771 18199 19777
rect 18141 19737 18153 19771
rect 18187 19768 18199 19771
rect 18230 19768 18236 19780
rect 18187 19740 18236 19768
rect 18187 19737 18199 19740
rect 18141 19731 18199 19737
rect 18230 19728 18236 19740
rect 18288 19728 18294 19780
rect 19797 19771 19855 19777
rect 19797 19737 19809 19771
rect 19843 19768 19855 19771
rect 20530 19768 20536 19780
rect 19843 19740 20536 19768
rect 19843 19737 19855 19740
rect 19797 19731 19855 19737
rect 20530 19728 20536 19740
rect 20588 19728 20594 19780
rect 21358 19728 21364 19780
rect 21416 19728 21422 19780
rect 21634 19728 21640 19780
rect 21692 19768 21698 19780
rect 23753 19771 23811 19777
rect 21692 19740 21850 19768
rect 21692 19728 21698 19740
rect 23753 19737 23765 19771
rect 23799 19768 23811 19771
rect 24302 19768 24308 19780
rect 23799 19740 24308 19768
rect 23799 19737 23811 19740
rect 23753 19731 23811 19737
rect 24302 19728 24308 19740
rect 24360 19728 24366 19780
rect 11907 19672 13860 19700
rect 13906 19660 13912 19712
rect 13964 19700 13970 19712
rect 15289 19703 15347 19709
rect 15289 19700 15301 19703
rect 13964 19672 15301 19700
rect 13964 19660 13970 19672
rect 15289 19669 15301 19672
rect 15335 19669 15347 19703
rect 15289 19663 15347 19669
rect 16298 19660 16304 19712
rect 16356 19660 16362 19712
rect 16574 19660 16580 19712
rect 16632 19700 16638 19712
rect 18049 19703 18107 19709
rect 18049 19700 18061 19703
rect 16632 19672 18061 19700
rect 16632 19660 16638 19672
rect 18049 19669 18061 19672
rect 18095 19669 18107 19703
rect 18248 19700 18276 19728
rect 18414 19700 18420 19712
rect 18248 19672 18420 19700
rect 18049 19663 18107 19669
rect 18414 19660 18420 19672
rect 18472 19660 18478 19712
rect 18598 19660 18604 19712
rect 18656 19700 18662 19712
rect 18693 19703 18751 19709
rect 18693 19700 18705 19703
rect 18656 19672 18705 19700
rect 18656 19660 18662 19672
rect 18693 19669 18705 19672
rect 18739 19669 18751 19703
rect 18693 19663 18751 19669
rect 18782 19660 18788 19712
rect 18840 19700 18846 19712
rect 19429 19703 19487 19709
rect 19429 19700 19441 19703
rect 18840 19672 19441 19700
rect 18840 19660 18846 19672
rect 19429 19669 19441 19672
rect 19475 19669 19487 19703
rect 19429 19663 19487 19669
rect 19518 19660 19524 19712
rect 19576 19700 19582 19712
rect 19889 19703 19947 19709
rect 19889 19700 19901 19703
rect 19576 19672 19901 19700
rect 19576 19660 19582 19672
rect 19889 19669 19901 19672
rect 19935 19669 19947 19703
rect 19889 19663 19947 19669
rect 20714 19660 20720 19712
rect 20772 19700 20778 19712
rect 22002 19700 22008 19712
rect 20772 19672 22008 19700
rect 20772 19660 20778 19672
rect 22002 19660 22008 19672
rect 22060 19700 22066 19712
rect 22833 19703 22891 19709
rect 22833 19700 22845 19703
rect 22060 19672 22845 19700
rect 22060 19660 22066 19672
rect 22833 19669 22845 19672
rect 22879 19669 22891 19703
rect 22833 19663 22891 19669
rect 23293 19703 23351 19709
rect 23293 19669 23305 19703
rect 23339 19700 23351 19703
rect 23566 19700 23572 19712
rect 23339 19672 23572 19700
rect 23339 19669 23351 19672
rect 23293 19663 23351 19669
rect 23566 19660 23572 19672
rect 23624 19660 23630 19712
rect 24578 19660 24584 19712
rect 24636 19660 24642 19712
rect 24854 19660 24860 19712
rect 24912 19700 24918 19712
rect 24949 19703 25007 19709
rect 24949 19700 24961 19703
rect 24912 19672 24961 19700
rect 24912 19660 24918 19672
rect 24949 19669 24961 19672
rect 24995 19700 25007 19703
rect 25958 19700 25964 19712
rect 24995 19672 25964 19700
rect 24995 19669 25007 19672
rect 24949 19663 25007 19669
rect 25958 19660 25964 19672
rect 26016 19660 26022 19712
rect 1104 19610 25852 19632
rect 1104 19558 7950 19610
rect 8002 19558 8014 19610
rect 8066 19558 8078 19610
rect 8130 19558 8142 19610
rect 8194 19558 8206 19610
rect 8258 19558 17950 19610
rect 18002 19558 18014 19610
rect 18066 19558 18078 19610
rect 18130 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 25852 19610
rect 1104 19536 25852 19558
rect 3878 19456 3884 19508
rect 3936 19456 3942 19508
rect 5810 19456 5816 19508
rect 5868 19456 5874 19508
rect 6730 19456 6736 19508
rect 6788 19496 6794 19508
rect 8389 19499 8447 19505
rect 8389 19496 8401 19499
rect 6788 19468 8401 19496
rect 6788 19456 6794 19468
rect 8389 19465 8401 19468
rect 8435 19465 8447 19499
rect 8389 19459 8447 19465
rect 12158 19456 12164 19508
rect 12216 19496 12222 19508
rect 12342 19496 12348 19508
rect 12216 19468 12348 19496
rect 12216 19456 12222 19468
rect 12342 19456 12348 19468
rect 12400 19456 12406 19508
rect 13354 19456 13360 19508
rect 13412 19496 13418 19508
rect 14366 19496 14372 19508
rect 13412 19468 14372 19496
rect 13412 19456 13418 19468
rect 14366 19456 14372 19468
rect 14424 19456 14430 19508
rect 14461 19499 14519 19505
rect 14461 19465 14473 19499
rect 14507 19496 14519 19499
rect 14550 19496 14556 19508
rect 14507 19468 14556 19496
rect 14507 19465 14519 19468
rect 14461 19459 14519 19465
rect 14550 19456 14556 19468
rect 14608 19456 14614 19508
rect 14826 19456 14832 19508
rect 14884 19496 14890 19508
rect 14921 19499 14979 19505
rect 14921 19496 14933 19499
rect 14884 19468 14933 19496
rect 14884 19456 14890 19468
rect 14921 19465 14933 19468
rect 14967 19465 14979 19499
rect 14921 19459 14979 19465
rect 15289 19499 15347 19505
rect 15289 19465 15301 19499
rect 15335 19496 15347 19499
rect 18690 19496 18696 19508
rect 15335 19468 18696 19496
rect 15335 19465 15347 19468
rect 15289 19459 15347 19465
rect 18690 19456 18696 19468
rect 18748 19456 18754 19508
rect 18785 19499 18843 19505
rect 18785 19465 18797 19499
rect 18831 19465 18843 19499
rect 18785 19459 18843 19465
rect 19245 19499 19303 19505
rect 19245 19465 19257 19499
rect 19291 19496 19303 19499
rect 19334 19496 19340 19508
rect 19291 19468 19340 19496
rect 19291 19465 19303 19468
rect 19245 19459 19303 19465
rect 8294 19428 8300 19440
rect 4080 19400 8300 19428
rect 1949 19363 2007 19369
rect 1949 19329 1961 19363
rect 1995 19360 2007 19363
rect 3786 19360 3792 19372
rect 1995 19332 3792 19360
rect 1995 19329 2007 19332
rect 1949 19323 2007 19329
rect 3786 19320 3792 19332
rect 3844 19320 3850 19372
rect 4080 19369 4108 19400
rect 8294 19388 8300 19400
rect 8352 19388 8358 19440
rect 9214 19428 9220 19440
rect 8588 19400 9220 19428
rect 4065 19363 4123 19369
rect 4065 19329 4077 19363
rect 4111 19329 4123 19363
rect 4065 19323 4123 19329
rect 4801 19363 4859 19369
rect 4801 19329 4813 19363
rect 4847 19360 4859 19363
rect 4890 19360 4896 19372
rect 4847 19332 4896 19360
rect 4847 19329 4859 19332
rect 4801 19323 4859 19329
rect 4890 19320 4896 19332
rect 4948 19320 4954 19372
rect 5994 19320 6000 19372
rect 6052 19320 6058 19372
rect 7285 19363 7343 19369
rect 7285 19360 7297 19363
rect 6748 19332 7297 19360
rect 1854 19252 1860 19304
rect 1912 19292 1918 19304
rect 2225 19295 2283 19301
rect 2225 19292 2237 19295
rect 1912 19264 2237 19292
rect 1912 19252 1918 19264
rect 2225 19261 2237 19264
rect 2271 19261 2283 19295
rect 2225 19255 2283 19261
rect 3326 19252 3332 19304
rect 3384 19292 3390 19304
rect 4525 19295 4583 19301
rect 4525 19292 4537 19295
rect 3384 19264 4537 19292
rect 3384 19252 3390 19264
rect 4525 19261 4537 19264
rect 4571 19261 4583 19295
rect 4525 19255 4583 19261
rect 6454 19252 6460 19304
rect 6512 19252 6518 19304
rect 6641 19295 6699 19301
rect 6641 19261 6653 19295
rect 6687 19292 6699 19295
rect 6748 19292 6776 19332
rect 7285 19329 7297 19332
rect 7331 19360 7343 19363
rect 7742 19360 7748 19372
rect 7331 19332 7748 19360
rect 7331 19329 7343 19332
rect 7285 19323 7343 19329
rect 7742 19320 7748 19332
rect 7800 19320 7806 19372
rect 8588 19369 8616 19400
rect 9214 19388 9220 19400
rect 9272 19388 9278 19440
rect 9766 19388 9772 19440
rect 9824 19388 9830 19440
rect 14274 19388 14280 19440
rect 14332 19428 14338 19440
rect 15381 19431 15439 19437
rect 15381 19428 15393 19431
rect 14332 19400 15393 19428
rect 14332 19388 14338 19400
rect 15381 19397 15393 19400
rect 15427 19397 15439 19431
rect 16666 19428 16672 19440
rect 15381 19391 15439 19397
rect 16316 19400 16672 19428
rect 7929 19363 7987 19369
rect 7929 19360 7941 19363
rect 7852 19332 7941 19360
rect 6687 19264 6776 19292
rect 6825 19295 6883 19301
rect 6687 19261 6699 19264
rect 6641 19255 6699 19261
rect 6825 19261 6837 19295
rect 6871 19292 6883 19295
rect 7190 19292 7196 19304
rect 6871 19264 7196 19292
rect 6871 19261 6883 19264
rect 6825 19255 6883 19261
rect 7190 19252 7196 19264
rect 7248 19292 7254 19304
rect 7650 19292 7656 19304
rect 7248 19264 7656 19292
rect 7248 19252 7254 19264
rect 7650 19252 7656 19264
rect 7708 19252 7714 19304
rect 6914 19184 6920 19236
rect 6972 19224 6978 19236
rect 7745 19227 7803 19233
rect 7745 19224 7757 19227
rect 6972 19196 7757 19224
rect 6972 19184 6978 19196
rect 7745 19193 7757 19196
rect 7791 19193 7803 19227
rect 7745 19187 7803 19193
rect 5350 19116 5356 19168
rect 5408 19156 5414 19168
rect 7006 19156 7012 19168
rect 5408 19128 7012 19156
rect 5408 19116 5414 19128
rect 7006 19116 7012 19128
rect 7064 19116 7070 19168
rect 7101 19159 7159 19165
rect 7101 19125 7113 19159
rect 7147 19156 7159 19159
rect 7282 19156 7288 19168
rect 7147 19128 7288 19156
rect 7147 19125 7159 19128
rect 7101 19119 7159 19125
rect 7282 19116 7288 19128
rect 7340 19116 7346 19168
rect 7650 19116 7656 19168
rect 7708 19156 7714 19168
rect 7852 19156 7880 19332
rect 7929 19329 7941 19332
rect 7975 19329 7987 19363
rect 7929 19323 7987 19329
rect 8573 19363 8631 19369
rect 8573 19329 8585 19363
rect 8619 19329 8631 19363
rect 8573 19323 8631 19329
rect 9030 19320 9036 19372
rect 9088 19320 9094 19372
rect 12250 19320 12256 19372
rect 12308 19360 12314 19372
rect 12713 19363 12771 19369
rect 12713 19360 12725 19363
rect 12308 19332 12725 19360
rect 12308 19320 12314 19332
rect 12713 19329 12725 19332
rect 12759 19329 12771 19363
rect 12713 19323 12771 19329
rect 14090 19320 14096 19372
rect 14148 19360 14154 19372
rect 15286 19360 15292 19372
rect 14148 19332 15292 19360
rect 14148 19320 14154 19332
rect 15286 19320 15292 19332
rect 15344 19320 15350 19372
rect 15654 19360 15660 19372
rect 15396 19332 15660 19360
rect 9309 19295 9367 19301
rect 9309 19261 9321 19295
rect 9355 19292 9367 19295
rect 10778 19292 10784 19304
rect 9355 19264 10784 19292
rect 9355 19261 9367 19264
rect 9309 19255 9367 19261
rect 10778 19252 10784 19264
rect 10836 19252 10842 19304
rect 12066 19252 12072 19304
rect 12124 19252 12130 19304
rect 12989 19295 13047 19301
rect 12989 19261 13001 19295
rect 13035 19292 13047 19295
rect 13630 19292 13636 19304
rect 13035 19264 13636 19292
rect 13035 19261 13047 19264
rect 12989 19255 13047 19261
rect 13630 19252 13636 19264
rect 13688 19252 13694 19304
rect 15102 19252 15108 19304
rect 15160 19292 15166 19304
rect 15396 19292 15424 19332
rect 15654 19320 15660 19332
rect 15712 19320 15718 19372
rect 16316 19369 16344 19400
rect 16666 19388 16672 19400
rect 16724 19388 16730 19440
rect 18322 19388 18328 19440
rect 18380 19388 18386 19440
rect 18800 19428 18828 19459
rect 19334 19456 19340 19468
rect 19392 19456 19398 19508
rect 19613 19499 19671 19505
rect 19613 19465 19625 19499
rect 19659 19496 19671 19499
rect 20441 19499 20499 19505
rect 20441 19496 20453 19499
rect 19659 19468 20453 19496
rect 19659 19465 19671 19468
rect 19613 19459 19671 19465
rect 20441 19465 20453 19468
rect 20487 19465 20499 19499
rect 20441 19459 20499 19465
rect 20806 19456 20812 19508
rect 20864 19456 20870 19508
rect 21266 19456 21272 19508
rect 21324 19496 21330 19508
rect 22005 19499 22063 19505
rect 22005 19496 22017 19499
rect 21324 19468 22017 19496
rect 21324 19456 21330 19468
rect 22005 19465 22017 19468
rect 22051 19465 22063 19499
rect 22005 19459 22063 19465
rect 22094 19456 22100 19508
rect 22152 19496 22158 19508
rect 22373 19499 22431 19505
rect 22373 19496 22385 19499
rect 22152 19468 22385 19496
rect 22152 19456 22158 19468
rect 22373 19465 22385 19468
rect 22419 19496 22431 19499
rect 22462 19496 22468 19508
rect 22419 19468 22468 19496
rect 22419 19465 22431 19468
rect 22373 19459 22431 19465
rect 22462 19456 22468 19468
rect 22520 19456 22526 19508
rect 23842 19496 23848 19508
rect 23216 19468 23848 19496
rect 19886 19428 19892 19440
rect 18800 19400 19892 19428
rect 19886 19388 19892 19400
rect 19944 19388 19950 19440
rect 23014 19428 23020 19440
rect 20456 19400 23020 19428
rect 20456 19372 20484 19400
rect 23014 19388 23020 19400
rect 23072 19388 23078 19440
rect 16301 19363 16359 19369
rect 16301 19329 16313 19363
rect 16347 19329 16359 19363
rect 16301 19323 16359 19329
rect 16482 19320 16488 19372
rect 16540 19360 16546 19372
rect 17037 19363 17095 19369
rect 17037 19360 17049 19363
rect 16540 19332 17049 19360
rect 16540 19320 16546 19332
rect 17037 19329 17049 19332
rect 17083 19329 17095 19363
rect 17037 19323 17095 19329
rect 19058 19320 19064 19372
rect 19116 19360 19122 19372
rect 19705 19363 19763 19369
rect 19705 19360 19717 19363
rect 19116 19332 19717 19360
rect 19116 19320 19122 19332
rect 19705 19329 19717 19332
rect 19751 19329 19763 19363
rect 19705 19323 19763 19329
rect 19812 19332 20024 19360
rect 15160 19264 15424 19292
rect 15565 19295 15623 19301
rect 15160 19252 15166 19264
rect 15565 19261 15577 19295
rect 15611 19292 15623 19295
rect 16022 19292 16028 19304
rect 15611 19264 16028 19292
rect 15611 19261 15623 19264
rect 15565 19255 15623 19261
rect 16022 19252 16028 19264
rect 16080 19252 16086 19304
rect 17313 19295 17371 19301
rect 17313 19292 17325 19295
rect 17052 19264 17325 19292
rect 17052 19236 17080 19264
rect 17313 19261 17325 19264
rect 17359 19292 17371 19295
rect 17678 19292 17684 19304
rect 17359 19264 17684 19292
rect 17359 19261 17371 19264
rect 17313 19255 17371 19261
rect 17678 19252 17684 19264
rect 17736 19292 17742 19304
rect 19812 19292 19840 19332
rect 17736 19264 19840 19292
rect 17736 19252 17742 19264
rect 19886 19252 19892 19304
rect 19944 19252 19950 19304
rect 19996 19292 20024 19332
rect 20438 19320 20444 19372
rect 20496 19320 20502 19372
rect 20898 19320 20904 19372
rect 20956 19320 20962 19372
rect 21358 19320 21364 19372
rect 21416 19360 21422 19372
rect 23216 19360 23244 19468
rect 23842 19456 23848 19468
rect 23900 19456 23906 19508
rect 23934 19456 23940 19508
rect 23992 19456 23998 19508
rect 25038 19456 25044 19508
rect 25096 19456 25102 19508
rect 23952 19428 23980 19456
rect 23952 19400 24058 19428
rect 21416 19332 23244 19360
rect 21416 19320 21422 19332
rect 23290 19320 23296 19372
rect 23348 19320 23354 19372
rect 20993 19295 21051 19301
rect 20993 19292 21005 19295
rect 19996 19264 21005 19292
rect 20993 19261 21005 19264
rect 21039 19261 21051 19295
rect 20993 19255 21051 19261
rect 21545 19295 21603 19301
rect 21545 19261 21557 19295
rect 21591 19292 21603 19295
rect 21634 19292 21640 19304
rect 21591 19264 21640 19292
rect 21591 19261 21603 19264
rect 21545 19255 21603 19261
rect 21634 19252 21640 19264
rect 21692 19252 21698 19304
rect 22465 19295 22523 19301
rect 22465 19261 22477 19295
rect 22511 19261 22523 19295
rect 22465 19255 22523 19261
rect 8202 19184 8208 19236
rect 8260 19224 8266 19236
rect 8662 19224 8668 19236
rect 8260 19196 8668 19224
rect 8260 19184 8266 19196
rect 8662 19184 8668 19196
rect 8720 19184 8726 19236
rect 10318 19184 10324 19236
rect 10376 19224 10382 19236
rect 11057 19227 11115 19233
rect 11057 19224 11069 19227
rect 10376 19196 11069 19224
rect 10376 19184 10382 19196
rect 11057 19193 11069 19196
rect 11103 19224 11115 19227
rect 11422 19224 11428 19236
rect 11103 19196 11428 19224
rect 11103 19193 11115 19196
rect 11057 19187 11115 19193
rect 11422 19184 11428 19196
rect 11480 19224 11486 19236
rect 11517 19227 11575 19233
rect 11517 19224 11529 19227
rect 11480 19196 11529 19224
rect 11480 19184 11486 19196
rect 11517 19193 11529 19196
rect 11563 19193 11575 19227
rect 11517 19187 11575 19193
rect 14366 19184 14372 19236
rect 14424 19224 14430 19236
rect 14734 19224 14740 19236
rect 14424 19196 14740 19224
rect 14424 19184 14430 19196
rect 14734 19184 14740 19196
rect 14792 19184 14798 19236
rect 16669 19227 16727 19233
rect 16669 19224 16681 19227
rect 15580 19196 16681 19224
rect 15580 19168 15608 19196
rect 16669 19193 16681 19196
rect 16715 19193 16727 19227
rect 16669 19187 16727 19193
rect 17034 19184 17040 19236
rect 17092 19184 17098 19236
rect 18414 19184 18420 19236
rect 18472 19224 18478 19236
rect 22094 19224 22100 19236
rect 18472 19196 22100 19224
rect 18472 19184 18478 19196
rect 22094 19184 22100 19196
rect 22152 19184 22158 19236
rect 7708 19128 7880 19156
rect 7708 19116 7714 19128
rect 7926 19116 7932 19168
rect 7984 19156 7990 19168
rect 9490 19156 9496 19168
rect 7984 19128 9496 19156
rect 7984 19116 7990 19128
rect 9490 19116 9496 19128
rect 9548 19116 9554 19168
rect 10778 19116 10784 19168
rect 10836 19156 10842 19168
rect 10962 19156 10968 19168
rect 10836 19128 10968 19156
rect 10836 19116 10842 19128
rect 10962 19116 10968 19128
rect 11020 19116 11026 19168
rect 11238 19116 11244 19168
rect 11296 19116 11302 19168
rect 11790 19116 11796 19168
rect 11848 19116 11854 19168
rect 11882 19116 11888 19168
rect 11940 19156 11946 19168
rect 13354 19156 13360 19168
rect 11940 19128 13360 19156
rect 11940 19116 11946 19128
rect 13354 19116 13360 19128
rect 13412 19116 13418 19168
rect 13722 19116 13728 19168
rect 13780 19156 13786 19168
rect 14826 19156 14832 19168
rect 13780 19128 14832 19156
rect 13780 19116 13786 19128
rect 14826 19116 14832 19128
rect 14884 19156 14890 19168
rect 15562 19156 15568 19168
rect 14884 19128 15568 19156
rect 14884 19116 14890 19128
rect 15562 19116 15568 19128
rect 15620 19116 15626 19168
rect 16114 19116 16120 19168
rect 16172 19116 16178 19168
rect 17126 19116 17132 19168
rect 17184 19156 17190 19168
rect 18782 19156 18788 19168
rect 17184 19128 18788 19156
rect 17184 19116 17190 19128
rect 18782 19116 18788 19128
rect 18840 19116 18846 19168
rect 20714 19116 20720 19168
rect 20772 19156 20778 19168
rect 20990 19156 20996 19168
rect 20772 19128 20996 19156
rect 20772 19116 20778 19128
rect 20990 19116 20996 19128
rect 21048 19116 21054 19168
rect 21910 19116 21916 19168
rect 21968 19156 21974 19168
rect 22480 19156 22508 19255
rect 22554 19252 22560 19304
rect 22612 19252 22618 19304
rect 23569 19295 23627 19301
rect 23569 19261 23581 19295
rect 23615 19292 23627 19295
rect 25222 19292 25228 19304
rect 23615 19264 25228 19292
rect 23615 19261 23627 19264
rect 23569 19255 23627 19261
rect 25222 19252 25228 19264
rect 25280 19252 25286 19304
rect 21968 19128 22508 19156
rect 21968 19116 21974 19128
rect 24026 19116 24032 19168
rect 24084 19156 24090 19168
rect 24670 19156 24676 19168
rect 24084 19128 24676 19156
rect 24084 19116 24090 19128
rect 24670 19116 24676 19128
rect 24728 19156 24734 19168
rect 25317 19159 25375 19165
rect 25317 19156 25329 19159
rect 24728 19128 25329 19156
rect 24728 19116 24734 19128
rect 25317 19125 25329 19128
rect 25363 19125 25375 19159
rect 25317 19119 25375 19125
rect 1104 19066 25852 19088
rect 1104 19014 2950 19066
rect 3002 19014 3014 19066
rect 3066 19014 3078 19066
rect 3130 19014 3142 19066
rect 3194 19014 3206 19066
rect 3258 19014 12950 19066
rect 13002 19014 13014 19066
rect 13066 19014 13078 19066
rect 13130 19014 13142 19066
rect 13194 19014 13206 19066
rect 13258 19014 22950 19066
rect 23002 19014 23014 19066
rect 23066 19014 23078 19066
rect 23130 19014 23142 19066
rect 23194 19014 23206 19066
rect 23258 19014 25852 19066
rect 1104 18992 25852 19014
rect 1946 18912 1952 18964
rect 2004 18912 2010 18964
rect 5813 18955 5871 18961
rect 5813 18921 5825 18955
rect 5859 18952 5871 18955
rect 5902 18952 5908 18964
rect 5859 18924 5908 18952
rect 5859 18921 5871 18924
rect 5813 18915 5871 18921
rect 5902 18912 5908 18924
rect 5960 18912 5966 18964
rect 6457 18955 6515 18961
rect 6457 18921 6469 18955
rect 6503 18952 6515 18955
rect 6730 18952 6736 18964
rect 6503 18924 6736 18952
rect 6503 18921 6515 18924
rect 6457 18915 6515 18921
rect 6730 18912 6736 18924
rect 6788 18912 6794 18964
rect 7006 18912 7012 18964
rect 7064 18952 7070 18964
rect 7064 18924 8248 18952
rect 7064 18912 7070 18924
rect 2590 18844 2596 18896
rect 2648 18844 2654 18896
rect 3237 18887 3295 18893
rect 3237 18853 3249 18887
rect 3283 18853 3295 18887
rect 3237 18847 3295 18853
rect 5169 18887 5227 18893
rect 5169 18853 5181 18887
rect 5215 18884 5227 18887
rect 8110 18884 8116 18896
rect 5215 18856 8116 18884
rect 5215 18853 5227 18856
rect 5169 18847 5227 18853
rect 3252 18816 3280 18847
rect 8110 18844 8116 18856
rect 8168 18844 8174 18896
rect 8220 18884 8248 18924
rect 8294 18912 8300 18964
rect 8352 18952 8358 18964
rect 8389 18955 8447 18961
rect 8389 18952 8401 18955
rect 8352 18924 8401 18952
rect 8352 18912 8358 18924
rect 8389 18921 8401 18924
rect 8435 18921 8447 18955
rect 9217 18955 9275 18961
rect 9217 18952 9229 18955
rect 8389 18915 8447 18921
rect 8496 18924 9229 18952
rect 8496 18884 8524 18924
rect 9217 18921 9229 18924
rect 9263 18921 9275 18955
rect 9217 18915 9275 18921
rect 9674 18912 9680 18964
rect 9732 18952 9738 18964
rect 12989 18955 13047 18961
rect 12989 18952 13001 18955
rect 9732 18924 13001 18952
rect 9732 18912 9738 18924
rect 12989 18921 13001 18924
rect 13035 18921 13047 18955
rect 12989 18915 13047 18921
rect 14274 18912 14280 18964
rect 14332 18912 14338 18964
rect 15580 18924 18736 18952
rect 8220 18856 8524 18884
rect 9490 18844 9496 18896
rect 9548 18884 9554 18896
rect 11882 18884 11888 18896
rect 9548 18856 11888 18884
rect 9548 18844 9554 18856
rect 11882 18844 11888 18856
rect 11940 18844 11946 18896
rect 15580 18884 15608 18924
rect 11992 18856 15608 18884
rect 6086 18816 6092 18828
rect 3252 18788 6092 18816
rect 6086 18776 6092 18788
rect 6144 18776 6150 18828
rect 7377 18819 7435 18825
rect 7377 18785 7389 18819
rect 7423 18816 7435 18819
rect 7558 18816 7564 18828
rect 7423 18788 7564 18816
rect 7423 18785 7435 18788
rect 7377 18779 7435 18785
rect 7558 18776 7564 18788
rect 7616 18776 7622 18828
rect 9861 18819 9919 18825
rect 9861 18785 9873 18819
rect 9907 18816 9919 18819
rect 10042 18816 10048 18828
rect 9907 18788 10048 18816
rect 9907 18785 9919 18788
rect 9861 18779 9919 18785
rect 10042 18776 10048 18788
rect 10100 18776 10106 18828
rect 11146 18776 11152 18828
rect 11204 18816 11210 18828
rect 11992 18816 12020 18856
rect 17218 18844 17224 18896
rect 17276 18844 17282 18896
rect 12618 18816 12624 18828
rect 11204 18788 12020 18816
rect 12084 18788 12624 18816
rect 11204 18776 11210 18788
rect 1673 18751 1731 18757
rect 1673 18717 1685 18751
rect 1719 18748 1731 18751
rect 2130 18748 2136 18760
rect 1719 18720 2136 18748
rect 1719 18717 1731 18720
rect 1673 18711 1731 18717
rect 2130 18708 2136 18720
rect 2188 18708 2194 18760
rect 2777 18751 2835 18757
rect 2777 18717 2789 18751
rect 2823 18717 2835 18751
rect 2777 18711 2835 18717
rect 3421 18751 3479 18757
rect 3421 18717 3433 18751
rect 3467 18748 3479 18751
rect 4154 18748 4160 18760
rect 3467 18720 4160 18748
rect 3467 18717 3479 18720
rect 3421 18711 3479 18717
rect 2792 18680 2820 18711
rect 4154 18708 4160 18720
rect 4212 18708 4218 18760
rect 4249 18751 4307 18757
rect 4249 18717 4261 18751
rect 4295 18748 4307 18751
rect 4706 18748 4712 18760
rect 4295 18720 4712 18748
rect 4295 18717 4307 18720
rect 4249 18711 4307 18717
rect 4706 18708 4712 18720
rect 4764 18708 4770 18760
rect 5353 18751 5411 18757
rect 5353 18717 5365 18751
rect 5399 18717 5411 18751
rect 5353 18711 5411 18717
rect 3878 18680 3884 18692
rect 2792 18652 3884 18680
rect 3878 18640 3884 18652
rect 3936 18640 3942 18692
rect 4065 18683 4123 18689
rect 4065 18649 4077 18683
rect 4111 18680 4123 18683
rect 5368 18680 5396 18711
rect 5994 18708 6000 18760
rect 6052 18708 6058 18760
rect 6454 18708 6460 18760
rect 6512 18748 6518 18760
rect 6641 18751 6699 18757
rect 6641 18748 6653 18751
rect 6512 18720 6653 18748
rect 6512 18708 6518 18720
rect 6641 18717 6653 18720
rect 6687 18717 6699 18751
rect 6641 18711 6699 18717
rect 7101 18751 7159 18757
rect 7101 18717 7113 18751
rect 7147 18748 7159 18751
rect 8386 18748 8392 18760
rect 7147 18720 8392 18748
rect 7147 18717 7159 18720
rect 7101 18711 7159 18717
rect 8386 18708 8392 18720
rect 8444 18708 8450 18760
rect 8581 18751 8639 18757
rect 8581 18717 8593 18751
rect 8627 18748 8639 18751
rect 8627 18720 9076 18748
rect 8627 18717 8639 18720
rect 8581 18711 8639 18717
rect 7926 18680 7932 18692
rect 4111 18652 7932 18680
rect 4111 18649 4123 18652
rect 4065 18643 4123 18649
rect 7926 18640 7932 18652
rect 7984 18640 7990 18692
rect 9048 18680 9076 18720
rect 9122 18708 9128 18760
rect 9180 18748 9186 18760
rect 9585 18751 9643 18757
rect 9585 18748 9597 18751
rect 9180 18720 9597 18748
rect 9180 18708 9186 18720
rect 9585 18717 9597 18720
rect 9631 18717 9643 18751
rect 9585 18711 9643 18717
rect 9766 18708 9772 18760
rect 9824 18748 9830 18760
rect 10318 18748 10324 18760
rect 9824 18720 10324 18748
rect 9824 18708 9830 18720
rect 10318 18708 10324 18720
rect 10376 18708 10382 18760
rect 10413 18751 10471 18757
rect 10413 18717 10425 18751
rect 10459 18748 10471 18751
rect 11790 18748 11796 18760
rect 10459 18720 11796 18748
rect 10459 18717 10471 18720
rect 10413 18711 10471 18717
rect 11790 18708 11796 18720
rect 11848 18708 11854 18760
rect 11882 18708 11888 18760
rect 11940 18748 11946 18760
rect 12084 18748 12112 18788
rect 12618 18776 12624 18788
rect 12676 18776 12682 18828
rect 12710 18776 12716 18828
rect 12768 18816 12774 18828
rect 13446 18816 13452 18828
rect 12768 18788 13452 18816
rect 12768 18776 12774 18788
rect 13446 18776 13452 18788
rect 13504 18776 13510 18828
rect 13630 18776 13636 18828
rect 13688 18776 13694 18828
rect 14550 18816 14556 18828
rect 13740 18788 14556 18816
rect 13740 18748 13768 18788
rect 14550 18776 14556 18788
rect 14608 18776 14614 18828
rect 14734 18776 14740 18828
rect 14792 18776 14798 18828
rect 14829 18819 14887 18825
rect 14829 18785 14841 18819
rect 14875 18816 14887 18819
rect 15102 18816 15108 18828
rect 14875 18788 15108 18816
rect 14875 18785 14887 18788
rect 14829 18779 14887 18785
rect 15102 18776 15108 18788
rect 15160 18776 15166 18828
rect 15286 18776 15292 18828
rect 15344 18816 15350 18828
rect 16482 18816 16488 18828
rect 15344 18788 16488 18816
rect 15344 18776 15350 18788
rect 16482 18776 16488 18788
rect 16540 18816 16546 18828
rect 16540 18788 16896 18816
rect 16540 18776 16546 18788
rect 11940 18720 12112 18748
rect 12406 18720 13768 18748
rect 11940 18708 11946 18720
rect 9306 18680 9312 18692
rect 9048 18652 9312 18680
rect 9306 18640 9312 18652
rect 9364 18640 9370 18692
rect 9677 18683 9735 18689
rect 9677 18649 9689 18683
rect 9723 18680 9735 18683
rect 12406 18680 12434 18720
rect 13814 18708 13820 18760
rect 13872 18748 13878 18760
rect 14918 18748 14924 18760
rect 13872 18720 14924 18748
rect 13872 18708 13878 18720
rect 14918 18708 14924 18720
rect 14976 18748 14982 18760
rect 15473 18751 15531 18757
rect 15473 18748 15485 18751
rect 14976 18720 15485 18748
rect 14976 18708 14982 18720
rect 15473 18717 15485 18720
rect 15519 18717 15531 18751
rect 16868 18748 16896 18788
rect 17862 18776 17868 18828
rect 17920 18816 17926 18828
rect 18322 18816 18328 18828
rect 17920 18788 18328 18816
rect 17920 18776 17926 18788
rect 18322 18776 18328 18788
rect 18380 18776 18386 18828
rect 18601 18819 18659 18825
rect 18601 18785 18613 18819
rect 18647 18785 18659 18819
rect 18708 18816 18736 18924
rect 18782 18912 18788 18964
rect 18840 18952 18846 18964
rect 18840 18924 21680 18952
rect 18840 18912 18846 18924
rect 21652 18884 21680 18924
rect 21818 18912 21824 18964
rect 21876 18952 21882 18964
rect 24397 18955 24455 18961
rect 24397 18952 24409 18955
rect 21876 18924 24409 18952
rect 21876 18912 21882 18924
rect 24397 18921 24409 18924
rect 24443 18952 24455 18955
rect 24443 18924 25084 18952
rect 24443 18921 24455 18924
rect 24397 18915 24455 18921
rect 24854 18884 24860 18896
rect 21652 18856 24860 18884
rect 24854 18844 24860 18856
rect 24912 18844 24918 18896
rect 22922 18816 22928 18828
rect 18708 18788 22928 18816
rect 18601 18779 18659 18785
rect 17497 18751 17555 18757
rect 17497 18748 17509 18751
rect 16868 18734 17509 18748
rect 16882 18720 17509 18734
rect 15473 18711 15531 18717
rect 17497 18717 17509 18720
rect 17543 18717 17555 18751
rect 17497 18711 17555 18717
rect 18414 18708 18420 18760
rect 18472 18708 18478 18760
rect 18616 18748 18644 18779
rect 22922 18776 22928 18788
rect 22980 18776 22986 18828
rect 25056 18825 25084 18924
rect 23109 18819 23167 18825
rect 23109 18785 23121 18819
rect 23155 18785 23167 18819
rect 23109 18779 23167 18785
rect 25041 18819 25099 18825
rect 25041 18785 25053 18819
rect 25087 18785 25099 18819
rect 25041 18779 25099 18785
rect 18782 18748 18788 18760
rect 18616 18720 18788 18748
rect 18782 18708 18788 18720
rect 18840 18708 18846 18760
rect 19610 18708 19616 18760
rect 19668 18708 19674 18760
rect 20349 18751 20407 18757
rect 20349 18717 20361 18751
rect 20395 18717 20407 18751
rect 20349 18711 20407 18717
rect 9723 18652 12434 18680
rect 13357 18683 13415 18689
rect 9723 18649 9735 18652
rect 9677 18643 9735 18649
rect 13357 18649 13369 18683
rect 13403 18680 13415 18683
rect 13722 18680 13728 18692
rect 13403 18652 13728 18680
rect 13403 18649 13415 18652
rect 13357 18643 13415 18649
rect 13722 18640 13728 18652
rect 13780 18640 13786 18692
rect 15194 18680 15200 18692
rect 13832 18652 15200 18680
rect 4525 18615 4583 18621
rect 4525 18581 4537 18615
rect 4571 18612 4583 18615
rect 8846 18612 8852 18624
rect 4571 18584 8852 18612
rect 4571 18581 4583 18584
rect 4525 18575 4583 18581
rect 8846 18572 8852 18584
rect 8904 18572 8910 18624
rect 9490 18572 9496 18624
rect 9548 18612 9554 18624
rect 10502 18612 10508 18624
rect 9548 18584 10508 18612
rect 9548 18572 9554 18584
rect 10502 18572 10508 18584
rect 10560 18572 10566 18624
rect 11698 18572 11704 18624
rect 11756 18572 11762 18624
rect 12529 18615 12587 18621
rect 12529 18581 12541 18615
rect 12575 18612 12587 18615
rect 12618 18612 12624 18624
rect 12575 18584 12624 18612
rect 12575 18581 12587 18584
rect 12529 18575 12587 18581
rect 12618 18572 12624 18584
rect 12676 18572 12682 18624
rect 12710 18572 12716 18624
rect 12768 18572 12774 18624
rect 13446 18572 13452 18624
rect 13504 18572 13510 18624
rect 13630 18572 13636 18624
rect 13688 18612 13694 18624
rect 13832 18612 13860 18652
rect 15194 18640 15200 18652
rect 15252 18640 15258 18692
rect 15749 18683 15807 18689
rect 15749 18649 15761 18683
rect 15795 18680 15807 18683
rect 16022 18680 16028 18692
rect 15795 18652 16028 18680
rect 15795 18649 15807 18652
rect 15749 18643 15807 18649
rect 16022 18640 16028 18652
rect 16080 18640 16086 18692
rect 17126 18640 17132 18692
rect 17184 18680 17190 18692
rect 17954 18680 17960 18692
rect 17184 18652 17960 18680
rect 17184 18640 17190 18652
rect 17954 18640 17960 18652
rect 18012 18640 18018 18692
rect 18322 18640 18328 18692
rect 18380 18680 18386 18692
rect 19242 18680 19248 18692
rect 18380 18652 19248 18680
rect 18380 18640 18386 18652
rect 19242 18640 19248 18652
rect 19300 18680 19306 18692
rect 20364 18680 20392 18711
rect 22370 18708 22376 18760
rect 22428 18748 22434 18760
rect 23124 18748 23152 18779
rect 25222 18776 25228 18828
rect 25280 18776 25286 18828
rect 22428 18720 23152 18748
rect 22428 18708 22434 18720
rect 23474 18708 23480 18760
rect 23532 18748 23538 18760
rect 24121 18751 24179 18757
rect 24121 18748 24133 18751
rect 23532 18720 24133 18748
rect 23532 18708 23538 18720
rect 24121 18717 24133 18720
rect 24167 18748 24179 18751
rect 24949 18751 25007 18757
rect 24949 18748 24961 18751
rect 24167 18720 24961 18748
rect 24167 18717 24179 18720
rect 24121 18711 24179 18717
rect 24949 18717 24961 18720
rect 24995 18717 25007 18751
rect 24949 18711 25007 18717
rect 19300 18652 20392 18680
rect 19300 18640 19306 18652
rect 20622 18640 20628 18692
rect 20680 18640 20686 18692
rect 21634 18640 21640 18692
rect 21692 18640 21698 18692
rect 22462 18680 22468 18692
rect 21928 18652 22468 18680
rect 13688 18584 13860 18612
rect 14645 18615 14703 18621
rect 13688 18572 13694 18584
rect 14645 18581 14657 18615
rect 14691 18612 14703 18615
rect 15010 18612 15016 18624
rect 14691 18584 15016 18612
rect 14691 18581 14703 18584
rect 14645 18575 14703 18581
rect 15010 18572 15016 18584
rect 15068 18612 15074 18624
rect 17678 18612 17684 18624
rect 15068 18584 17684 18612
rect 15068 18572 15074 18584
rect 17678 18572 17684 18584
rect 17736 18572 17742 18624
rect 18049 18615 18107 18621
rect 18049 18581 18061 18615
rect 18095 18612 18107 18615
rect 18414 18612 18420 18624
rect 18095 18584 18420 18612
rect 18095 18581 18107 18584
rect 18049 18575 18107 18581
rect 18414 18572 18420 18584
rect 18472 18572 18478 18624
rect 18509 18615 18567 18621
rect 18509 18581 18521 18615
rect 18555 18612 18567 18615
rect 19429 18615 19487 18621
rect 19429 18612 19441 18615
rect 18555 18584 19441 18612
rect 18555 18581 18567 18584
rect 18509 18575 18567 18581
rect 19429 18581 19441 18584
rect 19475 18581 19487 18615
rect 19429 18575 19487 18581
rect 19518 18572 19524 18624
rect 19576 18612 19582 18624
rect 19889 18615 19947 18621
rect 19889 18612 19901 18615
rect 19576 18584 19901 18612
rect 19576 18572 19582 18584
rect 19889 18581 19901 18584
rect 19935 18581 19947 18615
rect 19889 18575 19947 18581
rect 20438 18572 20444 18624
rect 20496 18612 20502 18624
rect 20898 18612 20904 18624
rect 20496 18584 20904 18612
rect 20496 18572 20502 18584
rect 20898 18572 20904 18584
rect 20956 18612 20962 18624
rect 21928 18612 21956 18652
rect 22462 18640 22468 18652
rect 22520 18680 22526 18692
rect 22520 18652 22692 18680
rect 22520 18640 22526 18652
rect 20956 18584 21956 18612
rect 22097 18615 22155 18621
rect 20956 18572 20962 18584
rect 22097 18581 22109 18615
rect 22143 18612 22155 18615
rect 22186 18612 22192 18624
rect 22143 18584 22192 18612
rect 22143 18581 22155 18584
rect 22097 18575 22155 18581
rect 22186 18572 22192 18584
rect 22244 18572 22250 18624
rect 22554 18572 22560 18624
rect 22612 18572 22618 18624
rect 22664 18612 22692 18652
rect 22738 18640 22744 18692
rect 22796 18680 22802 18692
rect 23017 18683 23075 18689
rect 23017 18680 23029 18683
rect 22796 18652 23029 18680
rect 22796 18640 22802 18652
rect 23017 18649 23029 18652
rect 23063 18649 23075 18683
rect 23017 18643 23075 18649
rect 23845 18683 23903 18689
rect 23845 18649 23857 18683
rect 23891 18680 23903 18683
rect 23934 18680 23940 18692
rect 23891 18652 23940 18680
rect 23891 18649 23903 18652
rect 23845 18643 23903 18649
rect 23934 18640 23940 18652
rect 23992 18640 23998 18692
rect 24029 18683 24087 18689
rect 24029 18649 24041 18683
rect 24075 18680 24087 18683
rect 25498 18680 25504 18692
rect 24075 18652 25504 18680
rect 24075 18649 24087 18652
rect 24029 18643 24087 18649
rect 25498 18640 25504 18652
rect 25556 18640 25562 18692
rect 22925 18615 22983 18621
rect 22925 18612 22937 18615
rect 22664 18584 22937 18612
rect 22925 18581 22937 18584
rect 22971 18612 22983 18615
rect 23198 18612 23204 18624
rect 22971 18584 23204 18612
rect 22971 18581 22983 18584
rect 22925 18575 22983 18581
rect 23198 18572 23204 18584
rect 23256 18572 23262 18624
rect 24578 18572 24584 18624
rect 24636 18572 24642 18624
rect 1104 18522 25852 18544
rect 1104 18470 7950 18522
rect 8002 18470 8014 18522
rect 8066 18470 8078 18522
rect 8130 18470 8142 18522
rect 8194 18470 8206 18522
rect 8258 18470 17950 18522
rect 18002 18470 18014 18522
rect 18066 18470 18078 18522
rect 18130 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 25852 18522
rect 1104 18448 25852 18470
rect 1581 18411 1639 18417
rect 1581 18377 1593 18411
rect 1627 18408 1639 18411
rect 3510 18408 3516 18420
rect 1627 18380 3516 18408
rect 1627 18377 1639 18380
rect 1581 18371 1639 18377
rect 3510 18368 3516 18380
rect 3568 18368 3574 18420
rect 3694 18368 3700 18420
rect 3752 18408 3758 18420
rect 3881 18411 3939 18417
rect 3881 18408 3893 18411
rect 3752 18380 3893 18408
rect 3752 18368 3758 18380
rect 3881 18377 3893 18380
rect 3927 18377 3939 18411
rect 3881 18371 3939 18377
rect 4982 18368 4988 18420
rect 5040 18408 5046 18420
rect 5169 18411 5227 18417
rect 5169 18408 5181 18411
rect 5040 18380 5181 18408
rect 5040 18368 5046 18380
rect 5169 18377 5181 18380
rect 5215 18377 5227 18411
rect 5169 18371 5227 18377
rect 5718 18368 5724 18420
rect 5776 18408 5782 18420
rect 5813 18411 5871 18417
rect 5813 18408 5825 18411
rect 5776 18380 5825 18408
rect 5776 18368 5782 18380
rect 5813 18377 5825 18380
rect 5859 18377 5871 18411
rect 5813 18371 5871 18377
rect 5994 18368 6000 18420
rect 6052 18408 6058 18420
rect 8297 18411 8355 18417
rect 8297 18408 8309 18411
rect 6052 18380 8309 18408
rect 6052 18368 6058 18380
rect 8297 18377 8309 18380
rect 8343 18377 8355 18411
rect 10778 18408 10784 18420
rect 8297 18371 8355 18377
rect 9232 18380 10784 18408
rect 2222 18300 2228 18352
rect 2280 18300 2286 18352
rect 2777 18343 2835 18349
rect 2777 18309 2789 18343
rect 2823 18340 2835 18343
rect 4614 18340 4620 18352
rect 2823 18312 4620 18340
rect 2823 18309 2835 18312
rect 2777 18303 2835 18309
rect 1765 18275 1823 18281
rect 1765 18241 1777 18275
rect 1811 18272 1823 18275
rect 2884 18272 2912 18312
rect 4614 18300 4620 18312
rect 4672 18300 4678 18352
rect 6822 18340 6828 18352
rect 4724 18312 6828 18340
rect 4724 18281 4752 18312
rect 6822 18300 6828 18312
rect 6880 18300 6886 18352
rect 8570 18340 8576 18352
rect 7852 18312 8576 18340
rect 1811 18244 2912 18272
rect 2961 18275 3019 18281
rect 1811 18241 1823 18244
rect 1765 18235 1823 18241
rect 2961 18241 2973 18275
rect 3007 18272 3019 18275
rect 3421 18275 3479 18281
rect 3421 18272 3433 18275
rect 3007 18244 3433 18272
rect 3007 18241 3019 18244
rect 2961 18235 3019 18241
rect 3421 18241 3433 18244
rect 3467 18241 3479 18275
rect 3421 18235 3479 18241
rect 4709 18275 4767 18281
rect 4709 18241 4721 18275
rect 4755 18241 4767 18275
rect 4709 18235 4767 18241
rect 5353 18275 5411 18281
rect 5353 18241 5365 18275
rect 5399 18272 5411 18275
rect 5534 18272 5540 18284
rect 5399 18244 5540 18272
rect 5399 18241 5411 18244
rect 5353 18235 5411 18241
rect 3436 18204 3464 18235
rect 5534 18232 5540 18244
rect 5592 18232 5598 18284
rect 5997 18275 6055 18281
rect 5997 18241 6009 18275
rect 6043 18272 6055 18275
rect 6914 18272 6920 18284
rect 6043 18244 6920 18272
rect 6043 18241 6055 18244
rect 5997 18235 6055 18241
rect 6914 18232 6920 18244
rect 6972 18232 6978 18284
rect 7190 18232 7196 18284
rect 7248 18232 7254 18284
rect 7852 18281 7880 18312
rect 8570 18300 8576 18312
rect 8628 18300 8634 18352
rect 9232 18349 9260 18380
rect 10778 18368 10784 18380
rect 10836 18368 10842 18420
rect 10962 18368 10968 18420
rect 11020 18408 11026 18420
rect 11882 18408 11888 18420
rect 11020 18380 11888 18408
rect 11020 18368 11026 18380
rect 11882 18368 11888 18380
rect 11940 18368 11946 18420
rect 12066 18368 12072 18420
rect 12124 18408 12130 18420
rect 12161 18411 12219 18417
rect 12161 18408 12173 18411
rect 12124 18380 12173 18408
rect 12124 18368 12130 18380
rect 12161 18377 12173 18380
rect 12207 18377 12219 18411
rect 12161 18371 12219 18377
rect 13814 18368 13820 18420
rect 13872 18408 13878 18420
rect 14277 18411 14335 18417
rect 14277 18408 14289 18411
rect 13872 18380 14289 18408
rect 13872 18368 13878 18380
rect 14277 18377 14289 18380
rect 14323 18377 14335 18411
rect 14277 18371 14335 18377
rect 14550 18368 14556 18420
rect 14608 18408 14614 18420
rect 15197 18411 15255 18417
rect 15197 18408 15209 18411
rect 14608 18380 15209 18408
rect 14608 18368 14614 18380
rect 15197 18377 15209 18380
rect 15243 18377 15255 18411
rect 15197 18371 15255 18377
rect 15562 18368 15568 18420
rect 15620 18408 15626 18420
rect 15657 18411 15715 18417
rect 15657 18408 15669 18411
rect 15620 18380 15669 18408
rect 15620 18368 15626 18380
rect 15657 18377 15669 18380
rect 15703 18377 15715 18411
rect 15657 18371 15715 18377
rect 16301 18411 16359 18417
rect 16301 18377 16313 18411
rect 16347 18408 16359 18411
rect 18506 18408 18512 18420
rect 16347 18380 18512 18408
rect 16347 18377 16359 18380
rect 16301 18371 16359 18377
rect 9217 18343 9275 18349
rect 9217 18309 9229 18343
rect 9263 18309 9275 18343
rect 9217 18303 9275 18309
rect 9766 18300 9772 18352
rect 9824 18300 9830 18352
rect 10594 18300 10600 18352
rect 10652 18340 10658 18352
rect 11057 18343 11115 18349
rect 11057 18340 11069 18343
rect 10652 18312 11069 18340
rect 10652 18300 10658 18312
rect 11057 18309 11069 18312
rect 11103 18309 11115 18343
rect 11057 18303 11115 18309
rect 11790 18300 11796 18352
rect 11848 18340 11854 18352
rect 12989 18343 13047 18349
rect 12989 18340 13001 18343
rect 11848 18312 13001 18340
rect 11848 18300 11854 18312
rect 12989 18309 13001 18312
rect 13035 18340 13047 18343
rect 16316 18340 16344 18371
rect 18506 18368 18512 18380
rect 18564 18368 18570 18420
rect 19702 18368 19708 18420
rect 19760 18368 19766 18420
rect 20070 18368 20076 18420
rect 20128 18408 20134 18420
rect 21545 18411 21603 18417
rect 21545 18408 21557 18411
rect 20128 18380 21557 18408
rect 20128 18368 20134 18380
rect 21545 18377 21557 18380
rect 21591 18377 21603 18411
rect 21545 18371 21603 18377
rect 21634 18368 21640 18420
rect 21692 18408 21698 18420
rect 23014 18408 23020 18420
rect 21692 18380 23020 18408
rect 21692 18368 21698 18380
rect 23014 18368 23020 18380
rect 23072 18368 23078 18420
rect 23106 18368 23112 18420
rect 23164 18408 23170 18420
rect 23290 18408 23296 18420
rect 23164 18380 23296 18408
rect 23164 18368 23170 18380
rect 23290 18368 23296 18380
rect 23348 18368 23354 18420
rect 24305 18411 24363 18417
rect 24305 18377 24317 18411
rect 24351 18408 24363 18411
rect 24670 18408 24676 18420
rect 24351 18380 24676 18408
rect 24351 18377 24363 18380
rect 24305 18371 24363 18377
rect 24670 18368 24676 18380
rect 24728 18368 24734 18420
rect 24854 18368 24860 18420
rect 24912 18408 24918 18420
rect 25041 18411 25099 18417
rect 25041 18408 25053 18411
rect 24912 18380 25053 18408
rect 24912 18368 24918 18380
rect 25041 18377 25053 18380
rect 25087 18377 25099 18411
rect 25041 18371 25099 18377
rect 13035 18312 16344 18340
rect 13035 18309 13047 18312
rect 12989 18303 13047 18309
rect 16482 18300 16488 18352
rect 16540 18300 16546 18352
rect 17126 18300 17132 18352
rect 17184 18340 17190 18352
rect 20622 18340 20628 18352
rect 17184 18312 20628 18340
rect 17184 18300 17190 18312
rect 20622 18300 20628 18312
rect 20680 18300 20686 18352
rect 20901 18343 20959 18349
rect 20901 18309 20913 18343
rect 20947 18340 20959 18343
rect 21082 18340 21088 18352
rect 20947 18312 21088 18340
rect 20947 18309 20959 18312
rect 20901 18303 20959 18309
rect 21082 18300 21088 18312
rect 21140 18300 21146 18352
rect 21450 18300 21456 18352
rect 21508 18340 21514 18352
rect 22005 18343 22063 18349
rect 22005 18340 22017 18343
rect 21508 18312 22017 18340
rect 21508 18300 21514 18312
rect 22005 18309 22017 18312
rect 22051 18340 22063 18343
rect 24029 18343 24087 18349
rect 24029 18340 24041 18343
rect 22051 18312 24041 18340
rect 22051 18309 22063 18312
rect 22005 18303 22063 18309
rect 24029 18309 24041 18312
rect 24075 18309 24087 18343
rect 24029 18303 24087 18309
rect 24949 18343 25007 18349
rect 24949 18309 24961 18343
rect 24995 18340 25007 18343
rect 25590 18340 25596 18352
rect 24995 18312 25596 18340
rect 24995 18309 25007 18312
rect 24949 18303 25007 18309
rect 25590 18300 25596 18312
rect 25648 18300 25654 18352
rect 7837 18275 7895 18281
rect 7837 18241 7849 18275
rect 7883 18241 7895 18275
rect 7837 18235 7895 18241
rect 6270 18204 6276 18216
rect 3436 18176 6276 18204
rect 6270 18164 6276 18176
rect 6328 18164 6334 18216
rect 6733 18207 6791 18213
rect 6733 18173 6745 18207
rect 6779 18204 6791 18207
rect 7852 18204 7880 18235
rect 8478 18232 8484 18284
rect 8536 18232 8542 18284
rect 8938 18232 8944 18284
rect 8996 18232 9002 18284
rect 10502 18232 10508 18284
rect 10560 18272 10566 18284
rect 15565 18275 15623 18281
rect 15565 18272 15577 18275
rect 10560 18244 15577 18272
rect 10560 18232 10566 18244
rect 15565 18241 15577 18244
rect 15611 18241 15623 18275
rect 15565 18235 15623 18241
rect 15672 18244 15884 18272
rect 6779 18176 7880 18204
rect 6779 18173 6791 18176
rect 6733 18167 6791 18173
rect 9306 18164 9312 18216
rect 9364 18204 9370 18216
rect 12253 18207 12311 18213
rect 9364 18176 11836 18204
rect 9364 18164 9370 18176
rect 3602 18096 3608 18148
rect 3660 18136 3666 18148
rect 4525 18139 4583 18145
rect 4525 18136 4537 18139
rect 3660 18108 4537 18136
rect 3660 18096 3666 18108
rect 4525 18105 4537 18108
rect 4571 18105 4583 18139
rect 4525 18099 4583 18105
rect 4614 18096 4620 18148
rect 4672 18136 4678 18148
rect 6362 18136 6368 18148
rect 4672 18108 6368 18136
rect 4672 18096 4678 18108
rect 6362 18096 6368 18108
rect 6420 18096 6426 18148
rect 7006 18096 7012 18148
rect 7064 18096 7070 18148
rect 11808 18145 11836 18176
rect 12253 18173 12265 18207
rect 12299 18173 12311 18207
rect 12253 18167 12311 18173
rect 11793 18139 11851 18145
rect 10704 18108 11376 18136
rect 3237 18071 3295 18077
rect 3237 18037 3249 18071
rect 3283 18068 3295 18071
rect 4062 18068 4068 18080
rect 3283 18040 4068 18068
rect 3283 18037 3295 18040
rect 3237 18031 3295 18037
rect 4062 18028 4068 18040
rect 4120 18028 4126 18080
rect 6549 18071 6607 18077
rect 6549 18037 6561 18071
rect 6595 18068 6607 18071
rect 7282 18068 7288 18080
rect 6595 18040 7288 18068
rect 6595 18037 6607 18040
rect 6549 18031 6607 18037
rect 7282 18028 7288 18040
rect 7340 18028 7346 18080
rect 7650 18028 7656 18080
rect 7708 18028 7714 18080
rect 9766 18028 9772 18080
rect 9824 18068 9830 18080
rect 10704 18077 10732 18108
rect 10689 18071 10747 18077
rect 10689 18068 10701 18071
rect 9824 18040 10701 18068
rect 9824 18028 9830 18040
rect 10689 18037 10701 18040
rect 10735 18037 10747 18071
rect 10689 18031 10747 18037
rect 11146 18028 11152 18080
rect 11204 18068 11210 18080
rect 11241 18071 11299 18077
rect 11241 18068 11253 18071
rect 11204 18040 11253 18068
rect 11204 18028 11210 18040
rect 11241 18037 11253 18040
rect 11287 18037 11299 18071
rect 11348 18068 11376 18108
rect 11793 18105 11805 18139
rect 11839 18105 11851 18139
rect 12268 18136 12296 18167
rect 12342 18164 12348 18216
rect 12400 18164 12406 18216
rect 12618 18164 12624 18216
rect 12676 18204 12682 18216
rect 15102 18204 15108 18216
rect 12676 18176 15108 18204
rect 12676 18164 12682 18176
rect 15102 18164 15108 18176
rect 15160 18164 15166 18216
rect 15672 18136 15700 18244
rect 15749 18207 15807 18213
rect 15749 18173 15761 18207
rect 15795 18173 15807 18207
rect 15749 18167 15807 18173
rect 12268 18108 15700 18136
rect 11793 18099 11851 18105
rect 15764 18068 15792 18167
rect 15856 18136 15884 18244
rect 16850 18232 16856 18284
rect 16908 18232 16914 18284
rect 17218 18232 17224 18284
rect 17276 18232 17282 18284
rect 17494 18232 17500 18284
rect 17552 18272 17558 18284
rect 18417 18275 18475 18281
rect 18417 18272 18429 18275
rect 17552 18244 18429 18272
rect 17552 18232 17558 18244
rect 18417 18241 18429 18244
rect 18463 18272 18475 18275
rect 19518 18272 19524 18284
rect 18463 18244 19524 18272
rect 18463 18241 18475 18244
rect 18417 18235 18475 18241
rect 19518 18232 19524 18244
rect 19576 18232 19582 18284
rect 19613 18275 19671 18281
rect 19613 18241 19625 18275
rect 19659 18272 19671 18275
rect 20438 18272 20444 18284
rect 19659 18244 20444 18272
rect 19659 18241 19671 18244
rect 19613 18235 19671 18241
rect 20438 18232 20444 18244
rect 20496 18232 20502 18284
rect 20806 18232 20812 18284
rect 20864 18272 20870 18284
rect 21174 18272 21180 18284
rect 20864 18244 21180 18272
rect 20864 18232 20870 18244
rect 21174 18232 21180 18244
rect 21232 18232 21238 18284
rect 22554 18232 22560 18284
rect 22612 18272 22618 18284
rect 25314 18272 25320 18284
rect 22612 18244 25320 18272
rect 22612 18232 22618 18244
rect 25314 18232 25320 18244
rect 25372 18232 25378 18284
rect 16868 18204 16896 18232
rect 17313 18207 17371 18213
rect 17313 18204 17325 18207
rect 16868 18176 17325 18204
rect 17313 18173 17325 18176
rect 17359 18173 17371 18207
rect 17313 18167 17371 18173
rect 16853 18139 16911 18145
rect 16853 18136 16865 18139
rect 15856 18108 16865 18136
rect 16853 18105 16865 18108
rect 16899 18105 16911 18139
rect 17328 18136 17356 18167
rect 17402 18164 17408 18216
rect 17460 18164 17466 18216
rect 18230 18164 18236 18216
rect 18288 18204 18294 18216
rect 18509 18207 18567 18213
rect 18509 18204 18521 18207
rect 18288 18176 18521 18204
rect 18288 18164 18294 18176
rect 18509 18173 18521 18176
rect 18555 18173 18567 18207
rect 18509 18167 18567 18173
rect 18690 18164 18696 18216
rect 18748 18164 18754 18216
rect 19426 18204 19432 18216
rect 19260 18176 19432 18204
rect 19058 18136 19064 18148
rect 17328 18108 19064 18136
rect 16853 18099 16911 18105
rect 19058 18096 19064 18108
rect 19116 18136 19122 18148
rect 19260 18136 19288 18176
rect 19426 18164 19432 18176
rect 19484 18164 19490 18216
rect 19794 18164 19800 18216
rect 19852 18213 19858 18216
rect 19852 18207 19901 18213
rect 19852 18173 19855 18207
rect 19889 18173 19901 18207
rect 19852 18167 19901 18173
rect 20993 18207 21051 18213
rect 20993 18173 21005 18207
rect 21039 18173 21051 18207
rect 20993 18167 21051 18173
rect 19852 18164 19858 18167
rect 19116 18108 19288 18136
rect 19116 18096 19122 18108
rect 20806 18096 20812 18148
rect 20864 18136 20870 18148
rect 21008 18136 21036 18167
rect 21910 18164 21916 18216
rect 21968 18204 21974 18216
rect 22094 18204 22100 18216
rect 21968 18176 22100 18204
rect 21968 18164 21974 18176
rect 22094 18164 22100 18176
rect 22152 18164 22158 18216
rect 22462 18164 22468 18216
rect 22520 18204 22526 18216
rect 23934 18204 23940 18216
rect 22520 18176 23940 18204
rect 22520 18164 22526 18176
rect 23934 18164 23940 18176
rect 23992 18164 23998 18216
rect 25225 18207 25283 18213
rect 25225 18173 25237 18207
rect 25271 18204 25283 18207
rect 25406 18204 25412 18216
rect 25271 18176 25412 18204
rect 25271 18173 25283 18176
rect 25225 18167 25283 18173
rect 25406 18164 25412 18176
rect 25464 18164 25470 18216
rect 20864 18108 21036 18136
rect 20864 18096 20870 18108
rect 21174 18096 21180 18148
rect 21232 18136 21238 18148
rect 24581 18139 24639 18145
rect 24581 18136 24593 18139
rect 21232 18108 24593 18136
rect 21232 18096 21238 18108
rect 24581 18105 24593 18108
rect 24627 18105 24639 18139
rect 24581 18099 24639 18105
rect 11348 18040 15792 18068
rect 11241 18031 11299 18037
rect 17494 18028 17500 18080
rect 17552 18068 17558 18080
rect 18049 18071 18107 18077
rect 18049 18068 18061 18071
rect 17552 18040 18061 18068
rect 17552 18028 17558 18040
rect 18049 18037 18061 18040
rect 18095 18037 18107 18071
rect 18049 18031 18107 18037
rect 19245 18071 19303 18077
rect 19245 18037 19257 18071
rect 19291 18068 19303 18071
rect 19886 18068 19892 18080
rect 19291 18040 19892 18068
rect 19291 18037 19303 18040
rect 19245 18031 19303 18037
rect 19886 18028 19892 18040
rect 19944 18028 19950 18080
rect 20438 18028 20444 18080
rect 20496 18028 20502 18080
rect 22554 18028 22560 18080
rect 22612 18068 22618 18080
rect 23106 18068 23112 18080
rect 22612 18040 23112 18068
rect 22612 18028 22618 18040
rect 23106 18028 23112 18040
rect 23164 18028 23170 18080
rect 1104 17978 25852 18000
rect 1104 17926 2950 17978
rect 3002 17926 3014 17978
rect 3066 17926 3078 17978
rect 3130 17926 3142 17978
rect 3194 17926 3206 17978
rect 3258 17926 12950 17978
rect 13002 17926 13014 17978
rect 13066 17926 13078 17978
rect 13130 17926 13142 17978
rect 13194 17926 13206 17978
rect 13258 17926 22950 17978
rect 23002 17926 23014 17978
rect 23066 17926 23078 17978
rect 23130 17926 23142 17978
rect 23194 17926 23206 17978
rect 23258 17926 25852 17978
rect 1104 17904 25852 17926
rect 3237 17867 3295 17873
rect 3237 17833 3249 17867
rect 3283 17864 3295 17867
rect 3326 17864 3332 17876
rect 3283 17836 3332 17864
rect 3283 17833 3295 17836
rect 3237 17827 3295 17833
rect 3326 17824 3332 17836
rect 3384 17824 3390 17876
rect 5442 17824 5448 17876
rect 5500 17864 5506 17876
rect 6457 17867 6515 17873
rect 6457 17864 6469 17867
rect 5500 17836 6469 17864
rect 5500 17824 5506 17836
rect 6457 17833 6469 17836
rect 6503 17833 6515 17867
rect 6457 17827 6515 17833
rect 7098 17824 7104 17876
rect 7156 17864 7162 17876
rect 7745 17867 7803 17873
rect 7745 17864 7757 17867
rect 7156 17836 7757 17864
rect 7156 17824 7162 17836
rect 7745 17833 7757 17836
rect 7791 17833 7803 17867
rect 7745 17827 7803 17833
rect 7852 17836 13400 17864
rect 6914 17796 6920 17808
rect 5184 17768 6920 17796
rect 5184 17737 5212 17768
rect 6914 17756 6920 17768
rect 6972 17756 6978 17808
rect 7190 17756 7196 17808
rect 7248 17796 7254 17808
rect 7852 17796 7880 17836
rect 9674 17796 9680 17808
rect 7248 17768 7880 17796
rect 8588 17768 9680 17796
rect 7248 17756 7254 17768
rect 5169 17731 5227 17737
rect 5169 17697 5181 17731
rect 5215 17697 5227 17731
rect 5169 17691 5227 17697
rect 3418 17620 3424 17672
rect 3476 17620 3482 17672
rect 4065 17663 4123 17669
rect 4065 17629 4077 17663
rect 4111 17660 4123 17663
rect 4709 17663 4767 17669
rect 4709 17660 4721 17663
rect 4111 17632 4721 17660
rect 4111 17629 4123 17632
rect 4065 17623 4123 17629
rect 4709 17629 4721 17632
rect 4755 17629 4767 17663
rect 4709 17623 4767 17629
rect 4724 17592 4752 17623
rect 5442 17620 5448 17672
rect 5500 17620 5506 17672
rect 6178 17620 6184 17672
rect 6236 17660 6242 17672
rect 6641 17663 6699 17669
rect 6641 17660 6653 17663
rect 6236 17632 6653 17660
rect 6236 17620 6242 17632
rect 6641 17629 6653 17632
rect 6687 17629 6699 17663
rect 6641 17623 6699 17629
rect 7282 17620 7288 17672
rect 7340 17620 7346 17672
rect 7834 17620 7840 17672
rect 7892 17660 7898 17672
rect 8588 17669 8616 17768
rect 9674 17756 9680 17768
rect 9732 17756 9738 17808
rect 11238 17756 11244 17808
rect 11296 17796 11302 17808
rect 11882 17796 11888 17808
rect 11296 17768 11888 17796
rect 11296 17756 11302 17768
rect 11882 17756 11888 17768
rect 11940 17756 11946 17808
rect 13372 17796 13400 17836
rect 13446 17824 13452 17876
rect 13504 17864 13510 17876
rect 17129 17867 17187 17873
rect 17129 17864 17141 17867
rect 13504 17836 17141 17864
rect 13504 17824 13510 17836
rect 17129 17833 17141 17836
rect 17175 17833 17187 17867
rect 20622 17864 20628 17876
rect 17129 17827 17187 17833
rect 17236 17836 20628 17864
rect 13906 17796 13912 17808
rect 13372 17768 13912 17796
rect 13906 17756 13912 17768
rect 13964 17756 13970 17808
rect 17236 17796 17264 17836
rect 20622 17824 20628 17836
rect 20680 17824 20686 17876
rect 20980 17867 21038 17873
rect 20980 17833 20992 17867
rect 21026 17864 21038 17867
rect 22186 17864 22192 17876
rect 21026 17836 22192 17864
rect 21026 17833 21038 17836
rect 20980 17827 21038 17833
rect 22186 17824 22192 17836
rect 22244 17824 22250 17876
rect 22465 17867 22523 17873
rect 22465 17833 22477 17867
rect 22511 17864 22523 17867
rect 22646 17864 22652 17876
rect 22511 17836 22652 17864
rect 22511 17833 22523 17836
rect 22465 17827 22523 17833
rect 22646 17824 22652 17836
rect 22704 17824 22710 17876
rect 24581 17867 24639 17873
rect 24581 17833 24593 17867
rect 24627 17864 24639 17867
rect 24946 17864 24952 17876
rect 24627 17836 24952 17864
rect 24627 17833 24639 17836
rect 24581 17827 24639 17833
rect 24946 17824 24952 17836
rect 25004 17824 25010 17876
rect 16224 17768 17264 17796
rect 8938 17688 8944 17740
rect 8996 17728 9002 17740
rect 9769 17731 9827 17737
rect 9769 17728 9781 17731
rect 8996 17700 9781 17728
rect 8996 17688 9002 17700
rect 9769 17697 9781 17700
rect 9815 17728 9827 17731
rect 11698 17728 11704 17740
rect 9815 17700 11704 17728
rect 9815 17697 9827 17700
rect 9769 17691 9827 17697
rect 11698 17688 11704 17700
rect 11756 17728 11762 17740
rect 11977 17731 12035 17737
rect 11977 17728 11989 17731
rect 11756 17700 11989 17728
rect 11756 17688 11762 17700
rect 11977 17697 11989 17700
rect 12023 17697 12035 17731
rect 11977 17691 12035 17697
rect 12253 17731 12311 17737
rect 12253 17697 12265 17731
rect 12299 17728 12311 17731
rect 12802 17728 12808 17740
rect 12299 17700 12808 17728
rect 12299 17697 12311 17700
rect 12253 17691 12311 17697
rect 12802 17688 12808 17700
rect 12860 17728 12866 17740
rect 13262 17728 13268 17740
rect 12860 17700 13268 17728
rect 12860 17688 12866 17700
rect 13262 17688 13268 17700
rect 13320 17688 13326 17740
rect 13722 17688 13728 17740
rect 13780 17728 13786 17740
rect 14277 17731 14335 17737
rect 14277 17728 14289 17731
rect 13780 17700 14289 17728
rect 13780 17688 13786 17700
rect 14277 17697 14289 17700
rect 14323 17697 14335 17731
rect 14277 17691 14335 17697
rect 14918 17688 14924 17740
rect 14976 17688 14982 17740
rect 15746 17688 15752 17740
rect 15804 17728 15810 17740
rect 16224 17728 16252 17768
rect 17862 17756 17868 17808
rect 17920 17796 17926 17808
rect 18141 17799 18199 17805
rect 18141 17796 18153 17799
rect 17920 17768 18153 17796
rect 17920 17756 17926 17768
rect 18141 17765 18153 17768
rect 18187 17765 18199 17799
rect 18141 17759 18199 17765
rect 19426 17756 19432 17808
rect 19484 17796 19490 17808
rect 20162 17796 20168 17808
rect 19484 17768 20168 17796
rect 19484 17756 19490 17768
rect 20162 17756 20168 17768
rect 20220 17756 20226 17808
rect 22554 17796 22560 17808
rect 22066 17768 22560 17796
rect 15804 17700 16252 17728
rect 16669 17731 16727 17737
rect 15804 17688 15810 17700
rect 16669 17697 16681 17731
rect 16715 17697 16727 17731
rect 16669 17691 16727 17697
rect 7929 17663 7987 17669
rect 7929 17660 7941 17663
rect 7892 17632 7941 17660
rect 7892 17620 7898 17632
rect 7929 17629 7941 17632
rect 7975 17629 7987 17663
rect 7929 17623 7987 17629
rect 8573 17663 8631 17669
rect 8573 17629 8585 17663
rect 8619 17629 8631 17663
rect 8573 17623 8631 17629
rect 9309 17663 9367 17669
rect 9309 17629 9321 17663
rect 9355 17629 9367 17663
rect 9309 17623 9367 17629
rect 8294 17592 8300 17604
rect 4724 17564 8300 17592
rect 8294 17552 8300 17564
rect 8352 17552 8358 17604
rect 9324 17592 9352 17623
rect 16298 17620 16304 17672
rect 16356 17660 16362 17672
rect 16482 17660 16488 17672
rect 16356 17632 16488 17660
rect 16356 17620 16362 17632
rect 16482 17620 16488 17632
rect 16540 17620 16546 17672
rect 16684 17660 16712 17691
rect 16850 17688 16856 17740
rect 16908 17728 16914 17740
rect 17681 17731 17739 17737
rect 17681 17728 17693 17731
rect 16908 17700 17693 17728
rect 16908 17688 16914 17700
rect 17681 17697 17693 17700
rect 17727 17697 17739 17731
rect 17681 17691 17739 17697
rect 19794 17688 19800 17740
rect 19852 17728 19858 17740
rect 19981 17731 20039 17737
rect 19981 17728 19993 17731
rect 19852 17700 19993 17728
rect 19852 17688 19858 17700
rect 19981 17697 19993 17700
rect 20027 17697 20039 17731
rect 19981 17691 20039 17697
rect 20717 17731 20775 17737
rect 20717 17697 20729 17731
rect 20763 17728 20775 17731
rect 22066 17728 22094 17768
rect 22554 17756 22560 17768
rect 22612 17756 22618 17808
rect 23290 17756 23296 17808
rect 23348 17796 23354 17808
rect 23348 17768 25084 17796
rect 23348 17756 23354 17768
rect 20763 17700 22094 17728
rect 20763 17697 20775 17700
rect 20717 17691 20775 17697
rect 23750 17688 23756 17740
rect 23808 17688 23814 17740
rect 23842 17688 23848 17740
rect 23900 17688 23906 17740
rect 25056 17737 25084 17768
rect 25041 17731 25099 17737
rect 25041 17697 25053 17731
rect 25087 17697 25099 17731
rect 25041 17691 25099 17697
rect 25225 17731 25283 17737
rect 25225 17697 25237 17731
rect 25271 17728 25283 17731
rect 25866 17728 25872 17740
rect 25271 17700 25872 17728
rect 25271 17697 25283 17700
rect 25225 17691 25283 17697
rect 25866 17688 25872 17700
rect 25924 17688 25930 17740
rect 17034 17660 17040 17672
rect 16684 17632 17040 17660
rect 17034 17620 17040 17632
rect 17092 17620 17098 17672
rect 17497 17663 17555 17669
rect 17497 17629 17509 17663
rect 17543 17660 17555 17663
rect 18598 17660 18604 17672
rect 17543 17632 18604 17660
rect 17543 17629 17555 17632
rect 17497 17623 17555 17629
rect 18598 17620 18604 17632
rect 18656 17620 18662 17672
rect 18785 17663 18843 17669
rect 18785 17629 18797 17663
rect 18831 17660 18843 17663
rect 18874 17660 18880 17672
rect 18831 17632 18880 17660
rect 18831 17629 18843 17632
rect 18785 17623 18843 17629
rect 18874 17620 18880 17632
rect 18932 17620 18938 17672
rect 19889 17663 19947 17669
rect 19889 17629 19901 17663
rect 19935 17660 19947 17663
rect 20070 17660 20076 17672
rect 19935 17632 20076 17660
rect 19935 17629 19947 17632
rect 19889 17623 19947 17629
rect 20070 17620 20076 17632
rect 20128 17620 20134 17672
rect 22738 17620 22744 17672
rect 22796 17660 22802 17672
rect 23661 17663 23719 17669
rect 23661 17660 23673 17663
rect 22796 17632 23673 17660
rect 22796 17620 22802 17632
rect 23661 17629 23673 17632
rect 23707 17629 23719 17663
rect 23661 17623 23719 17629
rect 9950 17592 9956 17604
rect 9324 17564 9956 17592
rect 9950 17552 9956 17564
rect 10008 17552 10014 17604
rect 10042 17552 10048 17604
rect 10100 17552 10106 17604
rect 10318 17552 10324 17604
rect 10376 17592 10382 17604
rect 10502 17592 10508 17604
rect 10376 17564 10508 17592
rect 10376 17552 10382 17564
rect 10502 17552 10508 17564
rect 10560 17552 10566 17604
rect 12158 17592 12164 17604
rect 11348 17564 12164 17592
rect 4246 17484 4252 17536
rect 4304 17484 4310 17536
rect 4525 17527 4583 17533
rect 4525 17493 4537 17527
rect 4571 17524 4583 17527
rect 6822 17524 6828 17536
rect 4571 17496 6828 17524
rect 4571 17493 4583 17496
rect 4525 17487 4583 17493
rect 6822 17484 6828 17496
rect 6880 17484 6886 17536
rect 7098 17484 7104 17536
rect 7156 17484 7162 17536
rect 8386 17484 8392 17536
rect 8444 17484 8450 17536
rect 9122 17484 9128 17536
rect 9180 17484 9186 17536
rect 9306 17484 9312 17536
rect 9364 17524 9370 17536
rect 11348 17524 11376 17564
rect 12158 17552 12164 17564
rect 12216 17552 12222 17604
rect 12710 17552 12716 17604
rect 12768 17552 12774 17604
rect 14550 17552 14556 17604
rect 14608 17592 14614 17604
rect 15102 17592 15108 17604
rect 14608 17564 15108 17592
rect 14608 17552 14614 17564
rect 15102 17552 15108 17564
rect 15160 17552 15166 17604
rect 15194 17552 15200 17604
rect 15252 17552 15258 17604
rect 17402 17592 17408 17604
rect 16500 17564 17408 17592
rect 9364 17496 11376 17524
rect 9364 17484 9370 17496
rect 11422 17484 11428 17536
rect 11480 17524 11486 17536
rect 11517 17527 11575 17533
rect 11517 17524 11529 17527
rect 11480 17496 11529 17524
rect 11480 17484 11486 17496
rect 11517 17493 11529 17496
rect 11563 17493 11575 17527
rect 11517 17487 11575 17493
rect 12250 17484 12256 17536
rect 12308 17524 12314 17536
rect 13725 17527 13783 17533
rect 13725 17524 13737 17527
rect 12308 17496 13737 17524
rect 12308 17484 12314 17496
rect 13725 17493 13737 17496
rect 13771 17524 13783 17527
rect 16500 17524 16528 17564
rect 17402 17552 17408 17564
rect 17460 17552 17466 17604
rect 22462 17592 22468 17604
rect 18616 17564 20668 17592
rect 22218 17564 22468 17592
rect 13771 17496 16528 17524
rect 13771 17493 13783 17496
rect 13725 17487 13783 17493
rect 16574 17484 16580 17536
rect 16632 17524 16638 17536
rect 17589 17527 17647 17533
rect 17589 17524 17601 17527
rect 16632 17496 17601 17524
rect 16632 17484 16638 17496
rect 17589 17493 17601 17496
rect 17635 17524 17647 17527
rect 17678 17524 17684 17536
rect 17635 17496 17684 17524
rect 17635 17493 17647 17496
rect 17589 17487 17647 17493
rect 17678 17484 17684 17496
rect 17736 17484 17742 17536
rect 18616 17533 18644 17564
rect 18601 17527 18659 17533
rect 18601 17493 18613 17527
rect 18647 17493 18659 17527
rect 18601 17487 18659 17493
rect 19429 17527 19487 17533
rect 19429 17493 19441 17527
rect 19475 17524 19487 17527
rect 19518 17524 19524 17536
rect 19475 17496 19524 17524
rect 19475 17493 19487 17496
rect 19429 17487 19487 17493
rect 19518 17484 19524 17496
rect 19576 17484 19582 17536
rect 19797 17527 19855 17533
rect 19797 17493 19809 17527
rect 19843 17524 19855 17527
rect 20254 17524 20260 17536
rect 19843 17496 20260 17524
rect 19843 17493 19855 17496
rect 19797 17487 19855 17493
rect 20254 17484 20260 17496
rect 20312 17484 20318 17536
rect 20640 17524 20668 17564
rect 22462 17552 22468 17564
rect 22520 17592 22526 17604
rect 22833 17595 22891 17601
rect 22833 17592 22845 17595
rect 22520 17564 22845 17592
rect 22520 17552 22526 17564
rect 22833 17561 22845 17564
rect 22879 17592 22891 17595
rect 23017 17595 23075 17601
rect 23017 17592 23029 17595
rect 22879 17564 23029 17592
rect 22879 17561 22891 17564
rect 22833 17555 22891 17561
rect 23017 17561 23029 17564
rect 23063 17592 23075 17595
rect 23750 17592 23756 17604
rect 23063 17564 23756 17592
rect 23063 17561 23075 17564
rect 23017 17555 23075 17561
rect 23750 17552 23756 17564
rect 23808 17592 23814 17604
rect 24670 17592 24676 17604
rect 23808 17564 24676 17592
rect 23808 17552 23814 17564
rect 24670 17552 24676 17564
rect 24728 17552 24734 17604
rect 21910 17524 21916 17536
rect 20640 17496 21916 17524
rect 21910 17484 21916 17496
rect 21968 17484 21974 17536
rect 23293 17527 23351 17533
rect 23293 17493 23305 17527
rect 23339 17524 23351 17527
rect 23382 17524 23388 17536
rect 23339 17496 23388 17524
rect 23339 17493 23351 17496
rect 23293 17487 23351 17493
rect 23382 17484 23388 17496
rect 23440 17484 23446 17536
rect 23842 17484 23848 17536
rect 23900 17524 23906 17536
rect 24397 17527 24455 17533
rect 24397 17524 24409 17527
rect 23900 17496 24409 17524
rect 23900 17484 23906 17496
rect 24397 17493 24409 17496
rect 24443 17524 24455 17527
rect 24949 17527 25007 17533
rect 24949 17524 24961 17527
rect 24443 17496 24961 17524
rect 24443 17493 24455 17496
rect 24397 17487 24455 17493
rect 24949 17493 24961 17496
rect 24995 17493 25007 17527
rect 24949 17487 25007 17493
rect 1104 17434 25852 17456
rect 1104 17382 7950 17434
rect 8002 17382 8014 17434
rect 8066 17382 8078 17434
rect 8130 17382 8142 17434
rect 8194 17382 8206 17434
rect 8258 17382 17950 17434
rect 18002 17382 18014 17434
rect 18066 17382 18078 17434
rect 18130 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 25852 17434
rect 1104 17360 25852 17382
rect 3881 17323 3939 17329
rect 3881 17289 3893 17323
rect 3927 17320 3939 17323
rect 3970 17320 3976 17332
rect 3927 17292 3976 17320
rect 3927 17289 3939 17292
rect 3881 17283 3939 17289
rect 3970 17280 3976 17292
rect 4028 17280 4034 17332
rect 4246 17320 4252 17332
rect 4080 17292 4252 17320
rect 4080 17193 4108 17292
rect 4246 17280 4252 17292
rect 4304 17320 4310 17332
rect 7006 17320 7012 17332
rect 4304 17292 7012 17320
rect 4304 17280 4310 17292
rect 7006 17280 7012 17292
rect 7064 17280 7070 17332
rect 7190 17280 7196 17332
rect 7248 17280 7254 17332
rect 7374 17280 7380 17332
rect 7432 17320 7438 17332
rect 7837 17323 7895 17329
rect 7837 17320 7849 17323
rect 7432 17292 7849 17320
rect 7432 17280 7438 17292
rect 7837 17289 7849 17292
rect 7883 17289 7895 17323
rect 7837 17283 7895 17289
rect 8386 17280 8392 17332
rect 8444 17320 8450 17332
rect 15841 17323 15899 17329
rect 15841 17320 15853 17323
rect 8444 17292 15853 17320
rect 8444 17280 8450 17292
rect 15841 17289 15853 17292
rect 15887 17289 15899 17323
rect 15841 17283 15899 17289
rect 15930 17280 15936 17332
rect 15988 17320 15994 17332
rect 15988 17292 18000 17320
rect 15988 17280 15994 17292
rect 5166 17212 5172 17264
rect 5224 17252 5230 17264
rect 9398 17252 9404 17264
rect 5224 17224 8064 17252
rect 5224 17212 5230 17224
rect 4065 17187 4123 17193
rect 4065 17153 4077 17187
rect 4111 17153 4123 17187
rect 4065 17147 4123 17153
rect 6733 17187 6791 17193
rect 6733 17153 6745 17187
rect 6779 17184 6791 17187
rect 6914 17184 6920 17196
rect 6779 17156 6920 17184
rect 6779 17153 6791 17156
rect 6733 17147 6791 17153
rect 6914 17144 6920 17156
rect 6972 17144 6978 17196
rect 7282 17144 7288 17196
rect 7340 17184 7346 17196
rect 7377 17187 7435 17193
rect 7377 17184 7389 17187
rect 7340 17156 7389 17184
rect 7340 17144 7346 17156
rect 7377 17153 7389 17156
rect 7423 17184 7435 17187
rect 7742 17184 7748 17196
rect 7423 17156 7748 17184
rect 7423 17153 7435 17156
rect 7377 17147 7435 17153
rect 7742 17144 7748 17156
rect 7800 17144 7806 17196
rect 8036 17193 8064 17224
rect 8864 17224 9404 17252
rect 8021 17187 8079 17193
rect 8021 17153 8033 17187
rect 8067 17153 8079 17187
rect 8021 17147 8079 17153
rect 8754 17144 8760 17196
rect 8812 17144 8818 17196
rect 4525 17119 4583 17125
rect 4525 17085 4537 17119
rect 4571 17085 4583 17119
rect 4525 17079 4583 17085
rect 4540 17048 4568 17079
rect 4798 17076 4804 17128
rect 4856 17076 4862 17128
rect 5442 17076 5448 17128
rect 5500 17116 5506 17128
rect 8864 17116 8892 17224
rect 9398 17212 9404 17224
rect 9456 17212 9462 17264
rect 9493 17255 9551 17261
rect 9493 17221 9505 17255
rect 9539 17252 9551 17255
rect 9766 17252 9772 17264
rect 9539 17224 9772 17252
rect 9539 17221 9551 17224
rect 9493 17215 9551 17221
rect 9766 17212 9772 17224
rect 9824 17212 9830 17264
rect 11422 17212 11428 17264
rect 11480 17252 11486 17264
rect 11977 17255 12035 17261
rect 11977 17252 11989 17255
rect 11480 17224 11989 17252
rect 11480 17212 11486 17224
rect 11977 17221 11989 17224
rect 12023 17221 12035 17255
rect 11977 17215 12035 17221
rect 12710 17212 12716 17264
rect 12768 17212 12774 17264
rect 16206 17212 16212 17264
rect 16264 17252 16270 17264
rect 16850 17252 16856 17264
rect 16264 17224 16856 17252
rect 16264 17212 16270 17224
rect 16850 17212 16856 17224
rect 16908 17212 16914 17264
rect 17313 17255 17371 17261
rect 17313 17221 17325 17255
rect 17359 17252 17371 17255
rect 17862 17252 17868 17264
rect 17359 17224 17868 17252
rect 17359 17221 17371 17224
rect 17313 17215 17371 17221
rect 17862 17212 17868 17224
rect 17920 17212 17926 17264
rect 8938 17144 8944 17196
rect 8996 17184 9002 17196
rect 9217 17187 9275 17193
rect 9217 17184 9229 17187
rect 8996 17156 9229 17184
rect 8996 17144 9002 17156
rect 9217 17153 9229 17156
rect 9263 17153 9275 17187
rect 9217 17147 9275 17153
rect 10594 17144 10600 17196
rect 10652 17184 10658 17196
rect 11241 17187 11299 17193
rect 11241 17184 11253 17187
rect 10652 17156 11253 17184
rect 10652 17144 10658 17156
rect 11241 17153 11253 17156
rect 11287 17153 11299 17187
rect 11241 17147 11299 17153
rect 11698 17144 11704 17196
rect 11756 17144 11762 17196
rect 14461 17187 14519 17193
rect 14461 17153 14473 17187
rect 14507 17184 14519 17187
rect 14550 17184 14556 17196
rect 14507 17156 14556 17184
rect 14507 17153 14519 17156
rect 14461 17147 14519 17153
rect 14550 17144 14556 17156
rect 14608 17144 14614 17196
rect 15010 17144 15016 17196
rect 15068 17144 15074 17196
rect 15120 17156 16068 17184
rect 5500 17088 8892 17116
rect 5500 17076 5506 17088
rect 10042 17076 10048 17128
rect 10100 17116 10106 17128
rect 10965 17119 11023 17125
rect 10965 17116 10977 17119
rect 10100 17088 10977 17116
rect 10100 17076 10106 17088
rect 10965 17085 10977 17088
rect 11011 17085 11023 17119
rect 10965 17079 11023 17085
rect 13262 17076 13268 17128
rect 13320 17116 13326 17128
rect 13449 17119 13507 17125
rect 13449 17116 13461 17119
rect 13320 17088 13461 17116
rect 13320 17076 13326 17088
rect 13449 17085 13461 17088
rect 13495 17085 13507 17119
rect 13449 17079 13507 17085
rect 13814 17076 13820 17128
rect 13872 17116 13878 17128
rect 13909 17119 13967 17125
rect 13909 17116 13921 17119
rect 13872 17088 13921 17116
rect 13872 17076 13878 17088
rect 13909 17085 13921 17088
rect 13955 17085 13967 17119
rect 13909 17079 13967 17085
rect 14090 17076 14096 17128
rect 14148 17116 14154 17128
rect 15120 17116 15148 17156
rect 16040 17125 16068 17156
rect 16942 17144 16948 17196
rect 17000 17184 17006 17196
rect 17221 17187 17279 17193
rect 17221 17184 17233 17187
rect 17000 17156 17233 17184
rect 17000 17144 17006 17156
rect 17221 17153 17233 17156
rect 17267 17153 17279 17187
rect 17221 17147 17279 17153
rect 14148 17088 15148 17116
rect 15933 17119 15991 17125
rect 14148 17076 14154 17088
rect 15933 17085 15945 17119
rect 15979 17085 15991 17119
rect 15933 17079 15991 17085
rect 16025 17119 16083 17125
rect 16025 17085 16037 17119
rect 16071 17085 16083 17119
rect 16025 17079 16083 17085
rect 17405 17119 17463 17125
rect 17405 17085 17417 17119
rect 17451 17085 17463 17119
rect 17405 17079 17463 17085
rect 8662 17048 8668 17060
rect 4540 17020 8668 17048
rect 8662 17008 8668 17020
rect 8720 17008 8726 17060
rect 6546 16940 6552 16992
rect 6604 16940 6610 16992
rect 8573 16983 8631 16989
rect 8573 16949 8585 16983
rect 8619 16980 8631 16983
rect 9490 16980 9496 16992
rect 8619 16952 9496 16980
rect 8619 16949 8631 16952
rect 8573 16943 8631 16949
rect 9490 16940 9496 16952
rect 9548 16940 9554 16992
rect 9950 16940 9956 16992
rect 10008 16980 10014 16992
rect 11054 16980 11060 16992
rect 10008 16952 11060 16980
rect 10008 16940 10014 16952
rect 11054 16940 11060 16952
rect 11112 16940 11118 16992
rect 14826 16940 14832 16992
rect 14884 16940 14890 16992
rect 15010 16940 15016 16992
rect 15068 16980 15074 16992
rect 15473 16983 15531 16989
rect 15473 16980 15485 16983
rect 15068 16952 15485 16980
rect 15068 16940 15074 16952
rect 15473 16949 15485 16952
rect 15519 16949 15531 16983
rect 15948 16980 15976 17079
rect 16850 17008 16856 17060
rect 16908 17008 16914 17060
rect 16482 16980 16488 16992
rect 15948 16952 16488 16980
rect 15473 16943 15531 16949
rect 16482 16940 16488 16952
rect 16540 16940 16546 16992
rect 16574 16940 16580 16992
rect 16632 16980 16638 16992
rect 17420 16980 17448 17079
rect 17678 17076 17684 17128
rect 17736 17116 17742 17128
rect 17865 17119 17923 17125
rect 17865 17116 17877 17119
rect 17736 17088 17877 17116
rect 17736 17076 17742 17088
rect 17865 17085 17877 17088
rect 17911 17085 17923 17119
rect 17865 17079 17923 17085
rect 16632 16952 17448 16980
rect 17972 16980 18000 17292
rect 18966 17280 18972 17332
rect 19024 17320 19030 17332
rect 20073 17323 20131 17329
rect 19024 17292 19932 17320
rect 19024 17280 19030 17292
rect 19904 17252 19932 17292
rect 20073 17289 20085 17323
rect 20119 17320 20131 17323
rect 20162 17320 20168 17332
rect 20119 17292 20168 17320
rect 20119 17289 20131 17292
rect 20073 17283 20131 17289
rect 20162 17280 20168 17292
rect 20220 17280 20226 17332
rect 20530 17280 20536 17332
rect 20588 17280 20594 17332
rect 20622 17280 20628 17332
rect 20680 17320 20686 17332
rect 24762 17320 24768 17332
rect 20680 17292 24768 17320
rect 20680 17280 20686 17292
rect 24762 17280 24768 17292
rect 24820 17280 24826 17332
rect 21177 17255 21235 17261
rect 21177 17252 21189 17255
rect 19904 17224 21189 17252
rect 21177 17221 21189 17224
rect 21223 17221 21235 17255
rect 21177 17215 21235 17221
rect 21913 17255 21971 17261
rect 21913 17221 21925 17255
rect 21959 17252 21971 17255
rect 22002 17252 22008 17264
rect 21959 17224 22008 17252
rect 21959 17221 21971 17224
rect 21913 17215 21971 17221
rect 18322 17144 18328 17196
rect 18380 17144 18386 17196
rect 21928 17184 21956 17215
rect 22002 17212 22008 17224
rect 22060 17252 22066 17264
rect 22097 17255 22155 17261
rect 22097 17252 22109 17255
rect 22060 17224 22109 17252
rect 22060 17212 22066 17224
rect 22097 17221 22109 17224
rect 22143 17252 22155 17255
rect 22281 17255 22339 17261
rect 22281 17252 22293 17255
rect 22143 17224 22293 17252
rect 22143 17221 22155 17224
rect 22097 17215 22155 17221
rect 22281 17221 22293 17224
rect 22327 17252 22339 17255
rect 22462 17252 22468 17264
rect 22327 17224 22468 17252
rect 22327 17221 22339 17224
rect 22281 17215 22339 17221
rect 22462 17212 22468 17224
rect 22520 17212 22526 17264
rect 24670 17252 24676 17264
rect 24058 17224 24676 17252
rect 24670 17212 24676 17224
rect 24728 17212 24734 17264
rect 19734 17156 21956 17184
rect 22554 17144 22560 17196
rect 22612 17144 22618 17196
rect 24854 17144 24860 17196
rect 24912 17184 24918 17196
rect 25317 17187 25375 17193
rect 25317 17184 25329 17187
rect 24912 17156 25329 17184
rect 24912 17144 24918 17156
rect 25317 17153 25329 17156
rect 25363 17153 25375 17187
rect 25317 17147 25375 17153
rect 18601 17119 18659 17125
rect 18601 17085 18613 17119
rect 18647 17116 18659 17119
rect 21082 17116 21088 17128
rect 18647 17088 21088 17116
rect 18647 17085 18659 17088
rect 18601 17079 18659 17085
rect 21082 17076 21088 17088
rect 21140 17076 21146 17128
rect 23474 17076 23480 17128
rect 23532 17116 23538 17128
rect 25041 17119 25099 17125
rect 25041 17116 25053 17119
rect 23532 17088 25053 17116
rect 23532 17076 23538 17088
rect 25041 17085 25053 17088
rect 25087 17085 25099 17119
rect 25041 17079 25099 17085
rect 20162 17008 20168 17060
rect 20220 17048 20226 17060
rect 22462 17048 22468 17060
rect 20220 17020 22468 17048
rect 20220 17008 20226 17020
rect 22462 17008 22468 17020
rect 22520 17008 22526 17060
rect 23934 17008 23940 17060
rect 23992 17048 23998 17060
rect 24305 17051 24363 17057
rect 24305 17048 24317 17051
rect 23992 17020 24317 17048
rect 23992 17008 23998 17020
rect 24305 17017 24317 17020
rect 24351 17017 24363 17051
rect 24305 17011 24363 17017
rect 19610 16980 19616 16992
rect 17972 16952 19616 16980
rect 16632 16940 16638 16952
rect 19610 16940 19616 16952
rect 19668 16940 19674 16992
rect 22820 16983 22878 16989
rect 22820 16949 22832 16983
rect 22866 16980 22878 16983
rect 25038 16980 25044 16992
rect 22866 16952 25044 16980
rect 22866 16949 22878 16952
rect 22820 16943 22878 16949
rect 25038 16940 25044 16952
rect 25096 16940 25102 16992
rect 1104 16890 25852 16912
rect 1104 16838 2950 16890
rect 3002 16838 3014 16890
rect 3066 16838 3078 16890
rect 3130 16838 3142 16890
rect 3194 16838 3206 16890
rect 3258 16838 12950 16890
rect 13002 16838 13014 16890
rect 13066 16838 13078 16890
rect 13130 16838 13142 16890
rect 13194 16838 13206 16890
rect 13258 16838 22950 16890
rect 23002 16838 23014 16890
rect 23066 16838 23078 16890
rect 23130 16838 23142 16890
rect 23194 16838 23206 16890
rect 23258 16838 25852 16890
rect 1104 16816 25852 16838
rect 7282 16736 7288 16788
rect 7340 16736 7346 16788
rect 8386 16736 8392 16788
rect 8444 16736 8450 16788
rect 9033 16779 9091 16785
rect 9033 16745 9045 16779
rect 9079 16776 9091 16779
rect 9306 16776 9312 16788
rect 9079 16748 9312 16776
rect 9079 16745 9091 16748
rect 9033 16739 9091 16745
rect 9306 16736 9312 16748
rect 9364 16776 9370 16788
rect 9582 16776 9588 16788
rect 9364 16748 9588 16776
rect 9364 16736 9370 16748
rect 9582 16736 9588 16748
rect 9640 16736 9646 16788
rect 9766 16736 9772 16788
rect 9824 16776 9830 16788
rect 10686 16776 10692 16788
rect 9824 16748 10692 16776
rect 9824 16736 9830 16748
rect 10686 16736 10692 16748
rect 10744 16736 10750 16788
rect 15010 16776 15016 16788
rect 11348 16748 15016 16776
rect 3418 16668 3424 16720
rect 3476 16708 3482 16720
rect 11146 16708 11152 16720
rect 3476 16680 11152 16708
rect 3476 16668 3482 16680
rect 11146 16668 11152 16680
rect 11204 16668 11210 16720
rect 6914 16600 6920 16652
rect 6972 16640 6978 16652
rect 9122 16640 9128 16652
rect 6972 16612 9128 16640
rect 6972 16600 6978 16612
rect 9122 16600 9128 16612
rect 9180 16600 9186 16652
rect 9217 16643 9275 16649
rect 9217 16609 9229 16643
rect 9263 16640 9275 16643
rect 9950 16640 9956 16652
rect 9263 16612 9956 16640
rect 9263 16609 9275 16612
rect 9217 16603 9275 16609
rect 9950 16600 9956 16612
rect 10008 16600 10014 16652
rect 11054 16640 11060 16652
rect 10796 16612 11060 16640
rect 4154 16532 4160 16584
rect 4212 16532 4218 16584
rect 4709 16575 4767 16581
rect 4709 16541 4721 16575
rect 4755 16572 4767 16575
rect 7374 16572 7380 16584
rect 4755 16544 7380 16572
rect 4755 16541 4767 16544
rect 4709 16535 4767 16541
rect 7374 16532 7380 16544
rect 7432 16532 7438 16584
rect 7469 16575 7527 16581
rect 7469 16541 7481 16575
rect 7515 16572 7527 16575
rect 7926 16572 7932 16584
rect 7515 16544 7932 16572
rect 7515 16541 7527 16544
rect 7469 16535 7527 16541
rect 7926 16532 7932 16544
rect 7984 16532 7990 16584
rect 8570 16532 8576 16584
rect 8628 16532 8634 16584
rect 9582 16572 9588 16584
rect 8680 16544 9588 16572
rect 8680 16504 8708 16544
rect 9582 16532 9588 16544
rect 9640 16532 9646 16584
rect 9677 16575 9735 16581
rect 9677 16541 9689 16575
rect 9723 16572 9735 16575
rect 10796 16572 10824 16612
rect 11054 16600 11060 16612
rect 11112 16600 11118 16652
rect 11241 16643 11299 16649
rect 11241 16609 11253 16643
rect 11287 16640 11299 16643
rect 11348 16640 11376 16748
rect 15010 16736 15016 16748
rect 15068 16736 15074 16788
rect 16022 16736 16028 16788
rect 16080 16736 16086 16788
rect 16114 16736 16120 16788
rect 16172 16776 16178 16788
rect 17862 16776 17868 16788
rect 16172 16748 17868 16776
rect 16172 16736 16178 16748
rect 17862 16736 17868 16748
rect 17920 16736 17926 16788
rect 19426 16776 19432 16788
rect 18432 16748 19432 16776
rect 11287 16612 11376 16640
rect 11425 16643 11483 16649
rect 11287 16609 11299 16612
rect 11241 16603 11299 16609
rect 11425 16609 11437 16643
rect 11471 16609 11483 16643
rect 11425 16603 11483 16609
rect 9723 16568 9812 16572
rect 9876 16568 10824 16572
rect 9723 16544 10824 16568
rect 9723 16541 9735 16544
rect 9677 16535 9735 16541
rect 9784 16540 9904 16544
rect 10870 16532 10876 16584
rect 10928 16572 10934 16584
rect 11149 16575 11207 16581
rect 11149 16572 11161 16575
rect 10928 16544 11161 16572
rect 10928 16532 10934 16544
rect 11149 16541 11161 16544
rect 11195 16541 11207 16575
rect 11149 16535 11207 16541
rect 11054 16504 11060 16516
rect 3988 16476 8708 16504
rect 9600 16476 11060 16504
rect 3988 16445 4016 16476
rect 3973 16439 4031 16445
rect 3973 16405 3985 16439
rect 4019 16405 4031 16439
rect 3973 16399 4031 16405
rect 7745 16439 7803 16445
rect 7745 16405 7757 16439
rect 7791 16436 7803 16439
rect 9398 16436 9404 16448
rect 7791 16408 9404 16436
rect 7791 16405 7803 16408
rect 7745 16399 7803 16405
rect 9398 16396 9404 16408
rect 9456 16396 9462 16448
rect 9493 16439 9551 16445
rect 9493 16405 9505 16439
rect 9539 16436 9551 16439
rect 9600 16436 9628 16476
rect 11054 16464 11060 16476
rect 11112 16464 11118 16516
rect 11440 16504 11468 16603
rect 12250 16600 12256 16652
rect 12308 16600 12314 16652
rect 14277 16643 14335 16649
rect 14277 16609 14289 16643
rect 14323 16640 14335 16643
rect 14918 16640 14924 16652
rect 14323 16612 14924 16640
rect 14323 16609 14335 16612
rect 14277 16603 14335 16609
rect 14918 16600 14924 16612
rect 14976 16600 14982 16652
rect 15010 16600 15016 16652
rect 15068 16640 15074 16652
rect 16850 16640 16856 16652
rect 15068 16612 16856 16640
rect 15068 16600 15074 16612
rect 16850 16600 16856 16612
rect 16908 16600 16914 16652
rect 17126 16600 17132 16652
rect 17184 16600 17190 16652
rect 17405 16643 17463 16649
rect 17405 16609 17417 16643
rect 17451 16640 17463 16643
rect 18432 16640 18460 16748
rect 19426 16736 19432 16748
rect 19484 16736 19490 16788
rect 19692 16779 19750 16785
rect 19692 16745 19704 16779
rect 19738 16776 19750 16779
rect 20714 16776 20720 16788
rect 19738 16748 20720 16776
rect 19738 16745 19750 16748
rect 19692 16739 19750 16745
rect 20714 16736 20720 16748
rect 20772 16776 20778 16788
rect 20772 16748 20944 16776
rect 20772 16736 20778 16748
rect 20916 16708 20944 16748
rect 21082 16736 21088 16788
rect 21140 16776 21146 16788
rect 21177 16779 21235 16785
rect 21177 16776 21189 16779
rect 21140 16748 21189 16776
rect 21140 16736 21146 16748
rect 21177 16745 21189 16748
rect 21223 16776 21235 16779
rect 21358 16776 21364 16788
rect 21223 16748 21364 16776
rect 21223 16745 21235 16748
rect 21177 16739 21235 16745
rect 21358 16736 21364 16748
rect 21416 16736 21422 16788
rect 22554 16785 22560 16788
rect 22544 16779 22560 16785
rect 22544 16745 22556 16779
rect 22544 16739 22560 16745
rect 22554 16736 22560 16739
rect 22612 16736 22618 16788
rect 21542 16708 21548 16720
rect 20916 16680 21548 16708
rect 21542 16668 21548 16680
rect 21600 16668 21606 16720
rect 17451 16612 18460 16640
rect 19429 16643 19487 16649
rect 17451 16609 17463 16612
rect 17405 16603 17463 16609
rect 19429 16609 19441 16643
rect 19475 16640 19487 16643
rect 22281 16643 22339 16649
rect 22281 16640 22293 16643
rect 19475 16612 22293 16640
rect 19475 16609 19487 16612
rect 19429 16603 19487 16609
rect 22281 16609 22293 16612
rect 22327 16640 22339 16643
rect 22554 16640 22560 16652
rect 22327 16612 22560 16640
rect 22327 16609 22339 16612
rect 22281 16603 22339 16609
rect 22554 16600 22560 16612
rect 22612 16600 22618 16652
rect 23750 16600 23756 16652
rect 23808 16600 23814 16652
rect 11698 16532 11704 16584
rect 11756 16572 11762 16584
rect 11977 16575 12035 16581
rect 11977 16572 11989 16575
rect 11756 16544 11989 16572
rect 11756 16532 11762 16544
rect 11977 16541 11989 16544
rect 12023 16541 12035 16575
rect 11977 16535 12035 16541
rect 16669 16575 16727 16581
rect 16669 16541 16681 16575
rect 16715 16541 16727 16575
rect 16669 16535 16727 16541
rect 12250 16504 12256 16516
rect 11440 16476 12256 16504
rect 12250 16464 12256 16476
rect 12308 16464 12314 16516
rect 12710 16464 12716 16516
rect 12768 16464 12774 16516
rect 14550 16464 14556 16516
rect 14608 16464 14614 16516
rect 16298 16504 16304 16516
rect 15778 16476 16304 16504
rect 16298 16464 16304 16476
rect 16356 16464 16362 16516
rect 16684 16448 16712 16535
rect 21082 16532 21088 16584
rect 21140 16572 21146 16584
rect 21637 16575 21695 16581
rect 21637 16572 21649 16575
rect 21140 16544 21649 16572
rect 21140 16532 21146 16544
rect 21637 16541 21649 16544
rect 21683 16541 21695 16575
rect 23768 16572 23796 16600
rect 23690 16544 23796 16572
rect 21637 16535 21695 16541
rect 24394 16532 24400 16584
rect 24452 16572 24458 16584
rect 24581 16575 24639 16581
rect 24581 16572 24593 16575
rect 24452 16544 24593 16572
rect 24452 16532 24458 16544
rect 24581 16541 24593 16544
rect 24627 16541 24639 16575
rect 24581 16535 24639 16541
rect 24762 16532 24768 16584
rect 24820 16572 24826 16584
rect 25225 16575 25283 16581
rect 25225 16572 25237 16575
rect 24820 16544 25237 16572
rect 24820 16532 24826 16544
rect 25225 16541 25237 16544
rect 25271 16541 25283 16575
rect 25225 16535 25283 16541
rect 16850 16464 16856 16516
rect 16908 16504 16914 16516
rect 17678 16504 17684 16516
rect 16908 16476 17684 16504
rect 16908 16464 16914 16476
rect 17678 16464 17684 16476
rect 17736 16504 17742 16516
rect 22002 16504 22008 16516
rect 17736 16476 17894 16504
rect 18708 16476 19012 16504
rect 20930 16476 22008 16504
rect 17736 16464 17742 16476
rect 9539 16408 9628 16436
rect 9539 16405 9551 16408
rect 9493 16399 9551 16405
rect 9674 16396 9680 16448
rect 9732 16436 9738 16448
rect 10042 16436 10048 16448
rect 9732 16408 10048 16436
rect 9732 16396 9738 16408
rect 10042 16396 10048 16408
rect 10100 16396 10106 16448
rect 10134 16396 10140 16448
rect 10192 16396 10198 16448
rect 10778 16396 10784 16448
rect 10836 16396 10842 16448
rect 12342 16396 12348 16448
rect 12400 16436 12406 16448
rect 13725 16439 13783 16445
rect 13725 16436 13737 16439
rect 12400 16408 13737 16436
rect 12400 16396 12406 16408
rect 13725 16405 13737 16408
rect 13771 16405 13783 16439
rect 13725 16399 13783 16405
rect 16482 16396 16488 16448
rect 16540 16396 16546 16448
rect 16666 16396 16672 16448
rect 16724 16436 16730 16448
rect 17586 16436 17592 16448
rect 16724 16408 17592 16436
rect 16724 16396 16730 16408
rect 17586 16396 17592 16408
rect 17644 16396 17650 16448
rect 18322 16396 18328 16448
rect 18380 16436 18386 16448
rect 18708 16436 18736 16476
rect 18380 16408 18736 16436
rect 18380 16396 18386 16408
rect 18874 16396 18880 16448
rect 18932 16396 18938 16448
rect 18984 16436 19012 16476
rect 22002 16464 22008 16476
rect 22060 16464 22066 16516
rect 22186 16464 22192 16516
rect 22244 16504 22250 16516
rect 22646 16504 22652 16516
rect 22244 16476 22652 16504
rect 22244 16464 22250 16476
rect 22646 16464 22652 16476
rect 22704 16464 22710 16516
rect 23842 16436 23848 16448
rect 18984 16408 23848 16436
rect 23842 16396 23848 16408
rect 23900 16396 23906 16448
rect 23934 16396 23940 16448
rect 23992 16436 23998 16448
rect 24029 16439 24087 16445
rect 24029 16436 24041 16439
rect 23992 16408 24041 16436
rect 23992 16396 23998 16408
rect 24029 16405 24041 16408
rect 24075 16405 24087 16439
rect 24029 16399 24087 16405
rect 1104 16346 25852 16368
rect 1104 16294 7950 16346
rect 8002 16294 8014 16346
rect 8066 16294 8078 16346
rect 8130 16294 8142 16346
rect 8194 16294 8206 16346
rect 8258 16294 17950 16346
rect 18002 16294 18014 16346
rect 18066 16294 18078 16346
rect 18130 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 25852 16346
rect 1104 16272 25852 16294
rect 4154 16192 4160 16244
rect 4212 16232 4218 16244
rect 4249 16235 4307 16241
rect 4249 16232 4261 16235
rect 4212 16204 4261 16232
rect 4212 16192 4218 16204
rect 4249 16201 4261 16204
rect 4295 16201 4307 16235
rect 4249 16195 4307 16201
rect 8021 16235 8079 16241
rect 8021 16201 8033 16235
rect 8067 16232 8079 16235
rect 8754 16232 8760 16244
rect 8067 16204 8760 16232
rect 8067 16201 8079 16204
rect 8021 16195 8079 16201
rect 8754 16192 8760 16204
rect 8812 16192 8818 16244
rect 9214 16192 9220 16244
rect 9272 16232 9278 16244
rect 9272 16204 10088 16232
rect 9272 16192 9278 16204
rect 5626 16124 5632 16176
rect 5684 16164 5690 16176
rect 5684 16136 9628 16164
rect 5684 16124 5690 16136
rect 8665 16099 8723 16105
rect 8665 16065 8677 16099
rect 8711 16065 8723 16099
rect 8665 16059 8723 16065
rect 8205 16031 8263 16037
rect 8205 15997 8217 16031
rect 8251 16028 8263 16031
rect 8680 16028 8708 16059
rect 9306 16056 9312 16108
rect 9364 16056 9370 16108
rect 9600 16096 9628 16136
rect 9600 16068 9904 16096
rect 9582 16028 9588 16040
rect 8251 16000 9588 16028
rect 8251 15997 8263 16000
rect 8205 15991 8263 15997
rect 9582 15988 9588 16000
rect 9640 15988 9646 16040
rect 9876 16028 9904 16068
rect 9950 16056 9956 16108
rect 10008 16056 10014 16108
rect 10060 16096 10088 16204
rect 10134 16192 10140 16244
rect 10192 16232 10198 16244
rect 10781 16235 10839 16241
rect 10781 16232 10793 16235
rect 10192 16204 10793 16232
rect 10192 16192 10198 16204
rect 10781 16201 10793 16204
rect 10827 16201 10839 16235
rect 10781 16195 10839 16201
rect 10873 16235 10931 16241
rect 10873 16201 10885 16235
rect 10919 16232 10931 16235
rect 15473 16235 15531 16241
rect 15473 16232 15485 16235
rect 10919 16204 15485 16232
rect 10919 16201 10931 16204
rect 10873 16195 10931 16201
rect 15473 16201 15485 16204
rect 15519 16201 15531 16235
rect 15473 16195 15531 16201
rect 15562 16192 15568 16244
rect 15620 16192 15626 16244
rect 15841 16235 15899 16241
rect 15841 16201 15853 16235
rect 15887 16232 15899 16235
rect 15887 16204 15976 16232
rect 15887 16201 15899 16204
rect 15841 16195 15899 16201
rect 12710 16124 12716 16176
rect 12768 16124 12774 16176
rect 15105 16167 15163 16173
rect 15105 16133 15117 16167
rect 15151 16164 15163 16167
rect 15580 16164 15608 16192
rect 15746 16164 15752 16176
rect 15151 16136 15752 16164
rect 15151 16133 15163 16136
rect 15105 16127 15163 16133
rect 15746 16124 15752 16136
rect 15804 16124 15810 16176
rect 11422 16096 11428 16108
rect 10060 16068 11428 16096
rect 11422 16056 11428 16068
rect 11480 16056 11486 16108
rect 13906 16056 13912 16108
rect 13964 16096 13970 16108
rect 14277 16099 14335 16105
rect 14277 16096 14289 16099
rect 13964 16068 14289 16096
rect 13964 16056 13970 16068
rect 14277 16065 14289 16068
rect 14323 16065 14335 16099
rect 15948 16100 15976 16204
rect 16298 16192 16304 16244
rect 16356 16232 16362 16244
rect 16669 16235 16727 16241
rect 16669 16232 16681 16235
rect 16356 16204 16681 16232
rect 16356 16192 16362 16204
rect 16669 16201 16681 16204
rect 16715 16232 16727 16235
rect 16850 16232 16856 16244
rect 16715 16204 16856 16232
rect 16715 16201 16727 16204
rect 16669 16195 16727 16201
rect 16850 16192 16856 16204
rect 16908 16192 16914 16244
rect 17770 16232 17776 16244
rect 17052 16204 17776 16232
rect 15948 16096 16068 16100
rect 17052 16096 17080 16204
rect 17770 16192 17776 16204
rect 17828 16192 17834 16244
rect 18417 16235 18475 16241
rect 18417 16201 18429 16235
rect 18463 16232 18475 16235
rect 18506 16232 18512 16244
rect 18463 16204 18512 16232
rect 18463 16201 18475 16204
rect 18417 16195 18475 16201
rect 18506 16192 18512 16204
rect 18564 16192 18570 16244
rect 19058 16192 19064 16244
rect 19116 16232 19122 16244
rect 19797 16235 19855 16241
rect 19797 16232 19809 16235
rect 19116 16204 19809 16232
rect 19116 16192 19122 16204
rect 19797 16201 19809 16204
rect 19843 16232 19855 16235
rect 20622 16232 20628 16244
rect 19843 16204 20628 16232
rect 19843 16201 19855 16204
rect 19797 16195 19855 16201
rect 20622 16192 20628 16204
rect 20680 16192 20686 16244
rect 20898 16192 20904 16244
rect 20956 16192 20962 16244
rect 21082 16192 21088 16244
rect 21140 16232 21146 16244
rect 21634 16232 21640 16244
rect 21140 16204 21640 16232
rect 21140 16192 21146 16204
rect 21634 16192 21640 16204
rect 21692 16192 21698 16244
rect 22278 16192 22284 16244
rect 22336 16232 22342 16244
rect 22465 16235 22523 16241
rect 22465 16232 22477 16235
rect 22336 16204 22477 16232
rect 22336 16192 22342 16204
rect 22465 16201 22477 16204
rect 22511 16201 22523 16235
rect 22465 16195 22523 16201
rect 24394 16192 24400 16244
rect 24452 16232 24458 16244
rect 25317 16235 25375 16241
rect 25317 16232 25329 16235
rect 24452 16204 25329 16232
rect 24452 16192 24458 16204
rect 25317 16201 25329 16204
rect 25363 16201 25375 16235
rect 25317 16195 25375 16201
rect 17218 16124 17224 16176
rect 17276 16164 17282 16176
rect 23753 16167 23811 16173
rect 17276 16136 22094 16164
rect 17276 16124 17282 16136
rect 15948 16072 17080 16096
rect 16040 16068 17080 16072
rect 17129 16099 17187 16105
rect 14277 16059 14335 16065
rect 17129 16065 17141 16099
rect 17175 16096 17187 16099
rect 18966 16096 18972 16108
rect 17175 16068 18972 16096
rect 17175 16065 17187 16068
rect 17129 16059 17187 16065
rect 18966 16056 18972 16068
rect 19024 16056 19030 16108
rect 19058 16056 19064 16108
rect 19116 16096 19122 16108
rect 19705 16099 19763 16105
rect 19705 16096 19717 16099
rect 19116 16068 19717 16096
rect 19116 16056 19122 16068
rect 19705 16065 19717 16068
rect 19751 16065 19763 16099
rect 19705 16059 19763 16065
rect 20622 16056 20628 16108
rect 20680 16096 20686 16108
rect 21545 16099 21603 16105
rect 21545 16096 21557 16099
rect 20680 16068 21557 16096
rect 20680 16056 20686 16068
rect 21545 16065 21557 16068
rect 21591 16065 21603 16099
rect 21545 16059 21603 16065
rect 10778 16028 10784 16040
rect 9876 16000 10784 16028
rect 10778 15988 10784 16000
rect 10836 15988 10842 16040
rect 11054 15988 11060 16040
rect 11112 15988 11118 16040
rect 11698 15988 11704 16040
rect 11756 15988 11762 16040
rect 11977 16031 12035 16037
rect 11977 15997 11989 16031
rect 12023 16028 12035 16031
rect 12342 16028 12348 16040
rect 12023 16000 12348 16028
rect 12023 15997 12035 16000
rect 11977 15991 12035 15997
rect 12342 15988 12348 16000
rect 12400 15988 12406 16040
rect 12710 15988 12716 16040
rect 12768 16028 12774 16040
rect 12768 16000 13308 16028
rect 12768 15988 12774 16000
rect 7466 15920 7472 15972
rect 7524 15960 7530 15972
rect 7524 15932 8892 15960
rect 7524 15920 7530 15932
rect 8478 15852 8484 15904
rect 8536 15852 8542 15904
rect 8864 15892 8892 15932
rect 9122 15920 9128 15972
rect 9180 15920 9186 15972
rect 9766 15920 9772 15972
rect 9824 15920 9830 15972
rect 13280 15960 13308 16000
rect 13446 15988 13452 16040
rect 13504 16028 13510 16040
rect 14090 16028 14096 16040
rect 13504 16000 14096 16028
rect 13504 15988 13510 16000
rect 14090 15988 14096 16000
rect 14148 15988 14154 16040
rect 14369 16031 14427 16037
rect 14369 15997 14381 16031
rect 14415 15997 14427 16031
rect 14369 15991 14427 15997
rect 14384 15960 14412 15991
rect 14550 15988 14556 16040
rect 14608 15988 14614 16040
rect 15838 15988 15844 16040
rect 15896 16028 15902 16040
rect 15933 16031 15991 16037
rect 15933 16028 15945 16031
rect 15896 16000 15945 16028
rect 15896 15988 15902 16000
rect 15933 15997 15945 16000
rect 15979 15997 15991 16031
rect 15933 15991 15991 15997
rect 16022 15988 16028 16040
rect 16080 15988 16086 16040
rect 16298 15988 16304 16040
rect 16356 16028 16362 16040
rect 19889 16031 19947 16037
rect 16356 16000 19472 16028
rect 16356 15988 16362 16000
rect 19337 15963 19395 15969
rect 19337 15960 19349 15963
rect 13280 15932 14320 15960
rect 14384 15932 16160 15960
rect 10413 15895 10471 15901
rect 10413 15892 10425 15895
rect 8864 15864 10425 15892
rect 10413 15861 10425 15864
rect 10459 15861 10471 15895
rect 10413 15855 10471 15861
rect 13538 15852 13544 15904
rect 13596 15892 13602 15904
rect 13909 15895 13967 15901
rect 13909 15892 13921 15895
rect 13596 15864 13921 15892
rect 13596 15852 13602 15864
rect 13909 15861 13921 15864
rect 13955 15861 13967 15895
rect 14292 15892 14320 15932
rect 14921 15895 14979 15901
rect 14921 15892 14933 15895
rect 14292 15864 14933 15892
rect 13909 15855 13967 15861
rect 14921 15861 14933 15864
rect 14967 15892 14979 15895
rect 15102 15892 15108 15904
rect 14967 15864 15108 15892
rect 14967 15861 14979 15864
rect 14921 15855 14979 15861
rect 15102 15852 15108 15864
rect 15160 15852 15166 15904
rect 15378 15852 15384 15904
rect 15436 15892 15442 15904
rect 16022 15892 16028 15904
rect 15436 15864 16028 15892
rect 15436 15852 15442 15864
rect 16022 15852 16028 15864
rect 16080 15852 16086 15904
rect 16132 15892 16160 15932
rect 16408 15932 19349 15960
rect 16408 15892 16436 15932
rect 19337 15929 19349 15932
rect 19383 15929 19395 15963
rect 19444 15960 19472 16000
rect 19889 15997 19901 16031
rect 19935 15997 19947 16031
rect 19889 15991 19947 15997
rect 19904 15960 19932 15991
rect 20254 15988 20260 16040
rect 20312 16028 20318 16040
rect 20993 16031 21051 16037
rect 20993 16028 21005 16031
rect 20312 16000 21005 16028
rect 20312 15988 20318 16000
rect 20993 15997 21005 16000
rect 21039 15997 21051 16031
rect 20993 15991 21051 15997
rect 19444 15932 19932 15960
rect 21008 15960 21036 15991
rect 21082 15988 21088 16040
rect 21140 15988 21146 16040
rect 22066 16028 22094 16136
rect 23753 16133 23765 16167
rect 23799 16164 23811 16167
rect 23842 16164 23848 16176
rect 23799 16136 23848 16164
rect 23799 16133 23811 16136
rect 23753 16127 23811 16133
rect 23842 16124 23848 16136
rect 23900 16124 23906 16176
rect 22278 16056 22284 16108
rect 22336 16096 22342 16108
rect 22373 16099 22431 16105
rect 22373 16096 22385 16099
rect 22336 16068 22385 16096
rect 22336 16056 22342 16068
rect 22373 16065 22385 16068
rect 22419 16065 22431 16099
rect 24118 16096 24124 16108
rect 22373 16059 22431 16065
rect 22480 16068 24124 16096
rect 22480 16028 22508 16068
rect 24118 16056 24124 16068
rect 24176 16056 24182 16108
rect 24670 16056 24676 16108
rect 24728 16096 24734 16108
rect 25133 16099 25191 16105
rect 25133 16096 25145 16099
rect 24728 16068 25145 16096
rect 24728 16056 24734 16068
rect 25133 16065 25145 16068
rect 25179 16065 25191 16099
rect 25133 16059 25191 16065
rect 22066 16000 22508 16028
rect 22646 15988 22652 16040
rect 22704 15988 22710 16040
rect 22830 15988 22836 16040
rect 22888 16028 22894 16040
rect 23845 16031 23903 16037
rect 23845 16028 23857 16031
rect 22888 16000 23857 16028
rect 22888 15988 22894 16000
rect 23845 15997 23857 16000
rect 23891 15997 23903 16031
rect 23845 15991 23903 15997
rect 23934 15988 23940 16040
rect 23992 15988 23998 16040
rect 25866 15988 25872 16040
rect 25924 16028 25930 16040
rect 26234 16028 26240 16040
rect 25924 16000 26240 16028
rect 25924 15988 25930 16000
rect 26234 15988 26240 16000
rect 26292 15988 26298 16040
rect 23017 15963 23075 15969
rect 23017 15960 23029 15963
rect 21008 15932 23029 15960
rect 19337 15923 19395 15929
rect 23017 15929 23029 15932
rect 23063 15929 23075 15963
rect 23017 15923 23075 15929
rect 24857 15963 24915 15969
rect 24857 15929 24869 15963
rect 24903 15960 24915 15963
rect 24946 15960 24952 15972
rect 24903 15932 24952 15960
rect 24903 15929 24915 15932
rect 24857 15923 24915 15929
rect 24946 15920 24952 15932
rect 25004 15920 25010 15972
rect 16132 15864 16436 15892
rect 16482 15852 16488 15904
rect 16540 15892 16546 15904
rect 20346 15892 20352 15904
rect 16540 15864 20352 15892
rect 16540 15852 16546 15864
rect 20346 15852 20352 15864
rect 20404 15852 20410 15904
rect 20530 15852 20536 15904
rect 20588 15852 20594 15904
rect 22005 15895 22063 15901
rect 22005 15861 22017 15895
rect 22051 15892 22063 15895
rect 22186 15892 22192 15904
rect 22051 15864 22192 15892
rect 22051 15861 22063 15864
rect 22005 15855 22063 15861
rect 22186 15852 22192 15864
rect 22244 15852 22250 15904
rect 23290 15852 23296 15904
rect 23348 15892 23354 15904
rect 23385 15895 23443 15901
rect 23385 15892 23397 15895
rect 23348 15864 23397 15892
rect 23348 15852 23354 15864
rect 23385 15861 23397 15864
rect 23431 15861 23443 15895
rect 23385 15855 23443 15861
rect 1104 15802 25852 15824
rect 1104 15750 2950 15802
rect 3002 15750 3014 15802
rect 3066 15750 3078 15802
rect 3130 15750 3142 15802
rect 3194 15750 3206 15802
rect 3258 15750 12950 15802
rect 13002 15750 13014 15802
rect 13066 15750 13078 15802
rect 13130 15750 13142 15802
rect 13194 15750 13206 15802
rect 13258 15750 22950 15802
rect 23002 15750 23014 15802
rect 23066 15750 23078 15802
rect 23130 15750 23142 15802
rect 23194 15750 23206 15802
rect 23258 15750 25852 15802
rect 1104 15728 25852 15750
rect 9858 15648 9864 15700
rect 9916 15648 9922 15700
rect 10962 15688 10968 15700
rect 10612 15660 10968 15688
rect 9217 15623 9275 15629
rect 9217 15589 9229 15623
rect 9263 15620 9275 15623
rect 10612 15620 10640 15660
rect 10962 15648 10968 15660
rect 11020 15648 11026 15700
rect 11146 15648 11152 15700
rect 11204 15688 11210 15700
rect 12713 15691 12771 15697
rect 12713 15688 12725 15691
rect 11204 15660 12725 15688
rect 11204 15648 11210 15660
rect 12713 15657 12725 15660
rect 12759 15657 12771 15691
rect 13446 15688 13452 15700
rect 12713 15651 12771 15657
rect 13096 15660 13452 15688
rect 9263 15592 10640 15620
rect 9263 15589 9275 15592
rect 9217 15583 9275 15589
rect 12250 15580 12256 15632
rect 12308 15580 12314 15632
rect 10781 15555 10839 15561
rect 10781 15521 10793 15555
rect 10827 15552 10839 15555
rect 13096 15552 13124 15660
rect 13446 15648 13452 15660
rect 13504 15648 13510 15700
rect 13817 15691 13875 15697
rect 13817 15657 13829 15691
rect 13863 15688 13875 15691
rect 13998 15688 14004 15700
rect 13863 15660 14004 15688
rect 13863 15657 13875 15660
rect 13817 15651 13875 15657
rect 13998 15648 14004 15660
rect 14056 15648 14062 15700
rect 15010 15688 15016 15700
rect 14108 15660 15016 15688
rect 14108 15620 14136 15660
rect 15010 15648 15016 15660
rect 15068 15648 15074 15700
rect 15194 15648 15200 15700
rect 15252 15688 15258 15700
rect 16025 15691 16083 15697
rect 16025 15688 16037 15691
rect 15252 15660 16037 15688
rect 15252 15648 15258 15660
rect 16025 15657 16037 15660
rect 16071 15657 16083 15691
rect 16025 15651 16083 15657
rect 16666 15648 16672 15700
rect 16724 15648 16730 15700
rect 18598 15648 18604 15700
rect 18656 15688 18662 15700
rect 18693 15691 18751 15697
rect 18693 15688 18705 15691
rect 18656 15660 18705 15688
rect 18656 15648 18662 15660
rect 18693 15657 18705 15660
rect 18739 15688 18751 15691
rect 19334 15688 19340 15700
rect 18739 15660 19340 15688
rect 18739 15657 18751 15660
rect 18693 15651 18751 15657
rect 19334 15648 19340 15660
rect 19392 15648 19398 15700
rect 23385 15691 23443 15697
rect 23385 15688 23397 15691
rect 19444 15660 23397 15688
rect 13188 15592 14136 15620
rect 16393 15623 16451 15629
rect 13188 15561 13216 15592
rect 16393 15589 16405 15623
rect 16439 15620 16451 15623
rect 16850 15620 16856 15632
rect 16439 15592 16856 15620
rect 16439 15589 16451 15592
rect 16393 15583 16451 15589
rect 16850 15580 16856 15592
rect 16908 15580 16914 15632
rect 19242 15580 19248 15632
rect 19300 15620 19306 15632
rect 19444 15620 19472 15660
rect 23385 15657 23397 15660
rect 23431 15657 23443 15691
rect 23385 15651 23443 15657
rect 24489 15691 24547 15697
rect 24489 15657 24501 15691
rect 24535 15688 24547 15691
rect 24854 15688 24860 15700
rect 24535 15660 24860 15688
rect 24535 15657 24547 15660
rect 24489 15651 24547 15657
rect 19300 15592 19472 15620
rect 20717 15623 20775 15629
rect 19300 15580 19306 15592
rect 20717 15589 20729 15623
rect 20763 15620 20775 15623
rect 21174 15620 21180 15632
rect 20763 15592 21180 15620
rect 20763 15589 20775 15592
rect 20717 15583 20775 15589
rect 21174 15580 21180 15592
rect 21232 15580 21238 15632
rect 24029 15623 24087 15629
rect 24029 15620 24041 15623
rect 21284 15592 24041 15620
rect 10827 15524 13124 15552
rect 13173 15555 13231 15561
rect 10827 15521 10839 15524
rect 10781 15515 10839 15521
rect 13173 15521 13185 15555
rect 13219 15521 13231 15555
rect 13173 15515 13231 15521
rect 13357 15555 13415 15561
rect 13357 15521 13369 15555
rect 13403 15552 13415 15555
rect 14182 15552 14188 15564
rect 13403 15524 14188 15552
rect 13403 15521 13415 15524
rect 13357 15515 13415 15521
rect 14182 15512 14188 15524
rect 14240 15512 14246 15564
rect 14274 15512 14280 15564
rect 14332 15552 14338 15564
rect 17221 15555 17279 15561
rect 14332 15524 15792 15552
rect 14332 15512 14338 15524
rect 8754 15444 8760 15496
rect 8812 15444 8818 15496
rect 9398 15444 9404 15496
rect 9456 15444 9462 15496
rect 10045 15487 10103 15493
rect 10045 15453 10057 15487
rect 10091 15484 10103 15487
rect 10226 15484 10232 15496
rect 10091 15456 10232 15484
rect 10091 15453 10103 15456
rect 10045 15447 10103 15453
rect 10226 15444 10232 15456
rect 10284 15444 10290 15496
rect 10505 15487 10563 15493
rect 10505 15453 10517 15487
rect 10551 15453 10563 15487
rect 10505 15447 10563 15453
rect 13081 15487 13139 15493
rect 13081 15453 13093 15487
rect 13127 15484 13139 15487
rect 13814 15484 13820 15496
rect 13127 15456 13820 15484
rect 13127 15453 13139 15456
rect 13081 15447 13139 15453
rect 10520 15416 10548 15447
rect 13814 15444 13820 15456
rect 13872 15444 13878 15496
rect 15764 15484 15792 15524
rect 17221 15521 17233 15555
rect 17267 15552 17279 15555
rect 18874 15552 18880 15564
rect 17267 15524 18880 15552
rect 17267 15521 17279 15524
rect 17221 15515 17279 15521
rect 18874 15512 18880 15524
rect 18932 15552 18938 15564
rect 20073 15555 20131 15561
rect 20073 15552 20085 15555
rect 18932 15524 20085 15552
rect 18932 15512 18938 15524
rect 20073 15521 20085 15524
rect 20119 15521 20131 15555
rect 20073 15515 20131 15521
rect 20162 15512 20168 15564
rect 20220 15552 20226 15564
rect 21284 15552 21312 15592
rect 20220 15524 21312 15552
rect 20220 15512 20226 15524
rect 21358 15512 21364 15564
rect 21416 15512 21422 15564
rect 16850 15484 16856 15496
rect 15764 15456 16856 15484
rect 16850 15444 16856 15456
rect 16908 15484 16914 15496
rect 16945 15487 17003 15493
rect 16945 15484 16957 15487
rect 16908 15456 16957 15484
rect 16908 15444 16914 15456
rect 16945 15453 16957 15456
rect 16991 15453 17003 15487
rect 16945 15447 17003 15453
rect 19978 15444 19984 15496
rect 20036 15444 20042 15496
rect 21085 15487 21143 15493
rect 21085 15453 21097 15487
rect 21131 15484 21143 15487
rect 21131 15456 21956 15484
rect 21131 15453 21143 15456
rect 21085 15447 21143 15453
rect 10686 15416 10692 15428
rect 10520 15388 10692 15416
rect 10686 15376 10692 15388
rect 10744 15376 10750 15428
rect 12710 15416 12716 15428
rect 12006 15388 12716 15416
rect 12710 15376 12716 15388
rect 12768 15376 12774 15428
rect 13538 15416 13544 15428
rect 13096 15388 13544 15416
rect 7558 15308 7564 15360
rect 7616 15348 7622 15360
rect 11146 15348 11152 15360
rect 7616 15320 11152 15348
rect 7616 15308 7622 15320
rect 11146 15308 11152 15320
rect 11204 15308 11210 15360
rect 11422 15308 11428 15360
rect 11480 15348 11486 15360
rect 13096 15348 13124 15388
rect 13538 15376 13544 15388
rect 13596 15376 13602 15428
rect 14553 15419 14611 15425
rect 14553 15385 14565 15419
rect 14599 15385 14611 15419
rect 14553 15379 14611 15385
rect 11480 15320 13124 15348
rect 14568 15348 14596 15379
rect 15102 15376 15108 15428
rect 15160 15376 15166 15428
rect 17678 15416 17684 15428
rect 17604 15388 17684 15416
rect 16206 15348 16212 15360
rect 14568 15320 16212 15348
rect 11480 15308 11486 15320
rect 16206 15308 16212 15320
rect 16264 15308 16270 15360
rect 17604 15348 17632 15388
rect 17678 15376 17684 15388
rect 17736 15376 17742 15428
rect 19889 15419 19947 15425
rect 19889 15385 19901 15419
rect 19935 15416 19947 15419
rect 21634 15416 21640 15428
rect 19935 15388 21640 15416
rect 19935 15385 19947 15388
rect 19889 15379 19947 15385
rect 21634 15376 21640 15388
rect 21692 15376 21698 15428
rect 21928 15416 21956 15456
rect 22002 15444 22008 15496
rect 22060 15444 22066 15496
rect 22646 15484 22652 15496
rect 22112 15456 22652 15484
rect 22112 15416 22140 15456
rect 22646 15444 22652 15456
rect 22704 15444 22710 15496
rect 22741 15487 22799 15493
rect 22741 15453 22753 15487
rect 22787 15484 22799 15487
rect 22848 15484 22876 15592
rect 24029 15589 24041 15592
rect 24075 15589 24087 15623
rect 24029 15583 24087 15589
rect 22787 15456 22876 15484
rect 23569 15487 23627 15493
rect 22787 15453 22799 15456
rect 22741 15447 22799 15453
rect 23569 15453 23581 15487
rect 23615 15484 23627 15487
rect 24504 15484 24532 15651
rect 24854 15648 24860 15660
rect 24912 15648 24918 15700
rect 25406 15484 25412 15496
rect 23615 15456 24532 15484
rect 24780 15456 25412 15484
rect 23615 15453 23627 15456
rect 23569 15447 23627 15453
rect 21928 15388 22140 15416
rect 22189 15419 22247 15425
rect 22189 15385 22201 15419
rect 22235 15416 22247 15419
rect 22235 15388 22968 15416
rect 22235 15385 22247 15388
rect 22189 15379 22247 15385
rect 18969 15351 19027 15357
rect 18969 15348 18981 15351
rect 17604 15320 18981 15348
rect 18969 15317 18981 15320
rect 19015 15317 19027 15351
rect 18969 15311 19027 15317
rect 19521 15351 19579 15357
rect 19521 15317 19533 15351
rect 19567 15348 19579 15351
rect 19702 15348 19708 15360
rect 19567 15320 19708 15348
rect 19567 15317 19579 15320
rect 19521 15311 19579 15317
rect 19702 15308 19708 15320
rect 19760 15308 19766 15360
rect 21177 15351 21235 15357
rect 21177 15317 21189 15351
rect 21223 15348 21235 15351
rect 21266 15348 21272 15360
rect 21223 15320 21272 15348
rect 21223 15317 21235 15320
rect 21177 15311 21235 15317
rect 21266 15308 21272 15320
rect 21324 15308 21330 15360
rect 22646 15308 22652 15360
rect 22704 15348 22710 15360
rect 22833 15351 22891 15357
rect 22833 15348 22845 15351
rect 22704 15320 22845 15348
rect 22704 15308 22710 15320
rect 22833 15317 22845 15320
rect 22879 15317 22891 15351
rect 22940 15348 22968 15388
rect 23198 15376 23204 15428
rect 23256 15416 23262 15428
rect 23845 15419 23903 15425
rect 23845 15416 23857 15419
rect 23256 15388 23857 15416
rect 23256 15376 23262 15388
rect 23845 15385 23857 15388
rect 23891 15385 23903 15419
rect 23845 15379 23903 15385
rect 24780 15348 24808 15456
rect 25406 15444 25412 15456
rect 25464 15444 25470 15496
rect 24854 15376 24860 15428
rect 24912 15376 24918 15428
rect 25038 15376 25044 15428
rect 25096 15376 25102 15428
rect 22940 15320 24808 15348
rect 24872 15348 24900 15376
rect 25317 15351 25375 15357
rect 25317 15348 25329 15351
rect 24872 15320 25329 15348
rect 22833 15311 22891 15317
rect 25317 15317 25329 15320
rect 25363 15317 25375 15351
rect 25317 15311 25375 15317
rect 1104 15258 25852 15280
rect 1104 15206 7950 15258
rect 8002 15206 8014 15258
rect 8066 15206 8078 15258
rect 8130 15206 8142 15258
rect 8194 15206 8206 15258
rect 8258 15206 17950 15258
rect 18002 15206 18014 15258
rect 18066 15206 18078 15258
rect 18130 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 25852 15258
rect 1104 15184 25852 15206
rect 9398 15104 9404 15156
rect 9456 15104 9462 15156
rect 9677 15147 9735 15153
rect 9677 15113 9689 15147
rect 9723 15144 9735 15147
rect 10226 15144 10232 15156
rect 9723 15116 10232 15144
rect 9723 15113 9735 15116
rect 9677 15107 9735 15113
rect 10226 15104 10232 15116
rect 10284 15104 10290 15156
rect 10962 15104 10968 15156
rect 11020 15104 11026 15156
rect 11054 15104 11060 15156
rect 11112 15144 11118 15156
rect 12066 15144 12072 15156
rect 11112 15116 12072 15144
rect 11112 15104 11118 15116
rect 12066 15104 12072 15116
rect 12124 15144 12130 15156
rect 13449 15147 13507 15153
rect 13449 15144 13461 15147
rect 12124 15116 13461 15144
rect 12124 15104 12130 15116
rect 13449 15113 13461 15116
rect 13495 15113 13507 15147
rect 13449 15107 13507 15113
rect 13906 15104 13912 15156
rect 13964 15104 13970 15156
rect 15286 15104 15292 15156
rect 15344 15144 15350 15156
rect 15473 15147 15531 15153
rect 15473 15144 15485 15147
rect 15344 15116 15485 15144
rect 15344 15104 15350 15116
rect 15473 15113 15485 15116
rect 15519 15113 15531 15147
rect 17034 15144 17040 15156
rect 15473 15107 15531 15113
rect 15948 15116 17040 15144
rect 9861 15079 9919 15085
rect 9861 15045 9873 15079
rect 9907 15076 9919 15079
rect 9907 15048 11192 15076
rect 9907 15045 9919 15048
rect 9861 15039 9919 15045
rect 11164 15020 11192 15048
rect 12710 15036 12716 15088
rect 12768 15036 12774 15088
rect 10502 14968 10508 15020
rect 10560 14968 10566 15020
rect 11146 14968 11152 15020
rect 11204 14968 11210 15020
rect 14553 15011 14611 15017
rect 14553 14977 14565 15011
rect 14599 15008 14611 15011
rect 15013 15011 15071 15017
rect 15013 15008 15025 15011
rect 14599 14980 15025 15008
rect 14599 14977 14611 14980
rect 14553 14971 14611 14977
rect 15013 14977 15025 14980
rect 15059 15008 15071 15011
rect 15948 15008 15976 15116
rect 17034 15104 17040 15116
rect 17092 15104 17098 15156
rect 18598 15144 18604 15156
rect 17144 15116 18604 15144
rect 17144 15085 17172 15116
rect 18598 15104 18604 15116
rect 18656 15104 18662 15156
rect 18966 15104 18972 15156
rect 19024 15104 19030 15156
rect 20622 15104 20628 15156
rect 20680 15144 20686 15156
rect 21085 15147 21143 15153
rect 21085 15144 21097 15147
rect 20680 15116 21097 15144
rect 20680 15104 20686 15116
rect 21085 15113 21097 15116
rect 21131 15113 21143 15147
rect 21085 15107 21143 15113
rect 21450 15104 21456 15156
rect 21508 15104 21514 15156
rect 21637 15147 21695 15153
rect 21637 15113 21649 15147
rect 21683 15144 21695 15147
rect 22094 15144 22100 15156
rect 21683 15116 22100 15144
rect 21683 15113 21695 15116
rect 21637 15107 21695 15113
rect 17129 15079 17187 15085
rect 17129 15045 17141 15079
rect 17175 15045 17187 15079
rect 17129 15039 17187 15045
rect 17678 15036 17684 15088
rect 17736 15036 17742 15088
rect 20898 15076 20904 15088
rect 20838 15048 20904 15076
rect 20898 15036 20904 15048
rect 20956 15076 20962 15088
rect 21652 15076 21680 15107
rect 22094 15104 22100 15116
rect 22152 15104 22158 15156
rect 23934 15144 23940 15156
rect 23124 15116 23940 15144
rect 23124 15085 23152 15116
rect 23934 15104 23940 15116
rect 23992 15104 23998 15156
rect 24486 15104 24492 15156
rect 24544 15144 24550 15156
rect 24581 15147 24639 15153
rect 24581 15144 24593 15147
rect 24544 15116 24593 15144
rect 24544 15104 24550 15116
rect 24581 15113 24593 15116
rect 24627 15113 24639 15147
rect 24581 15107 24639 15113
rect 20956 15048 21680 15076
rect 23109 15079 23167 15085
rect 20956 15036 20962 15048
rect 23109 15045 23121 15079
rect 23155 15045 23167 15079
rect 23109 15039 23167 15045
rect 23750 15036 23756 15088
rect 23808 15036 23814 15088
rect 15059 14980 15976 15008
rect 16853 15011 16911 15017
rect 15059 14977 15071 14980
rect 15013 14971 15071 14977
rect 16853 14977 16865 15011
rect 16899 14977 16911 15011
rect 18874 15008 18880 15020
rect 16853 14971 16911 14977
rect 18340 14980 18880 15008
rect 10686 14900 10692 14952
rect 10744 14940 10750 14952
rect 11698 14940 11704 14952
rect 10744 14912 11704 14940
rect 10744 14900 10750 14912
rect 11698 14900 11704 14912
rect 11756 14900 11762 14952
rect 11977 14943 12035 14949
rect 11977 14909 11989 14943
rect 12023 14940 12035 14943
rect 12434 14940 12440 14952
rect 12023 14912 12440 14940
rect 12023 14909 12035 14912
rect 11977 14903 12035 14909
rect 12434 14900 12440 14912
rect 12492 14940 12498 14952
rect 15378 14940 15384 14952
rect 12492 14912 15384 14940
rect 12492 14900 12498 14912
rect 15378 14900 15384 14912
rect 15436 14900 15442 14952
rect 16114 14900 16120 14952
rect 16172 14900 16178 14952
rect 16482 14940 16488 14952
rect 16316 14912 16488 14940
rect 10321 14875 10379 14881
rect 10321 14841 10333 14875
rect 10367 14872 10379 14875
rect 10367 14844 11376 14872
rect 10367 14841 10379 14844
rect 10321 14835 10379 14841
rect 10042 14764 10048 14816
rect 10100 14764 10106 14816
rect 11348 14804 11376 14844
rect 14090 14832 14096 14884
rect 14148 14872 14154 14884
rect 14734 14872 14740 14884
rect 14148 14844 14740 14872
rect 14148 14832 14154 14844
rect 14734 14832 14740 14844
rect 14792 14832 14798 14884
rect 14829 14875 14887 14881
rect 14829 14841 14841 14875
rect 14875 14872 14887 14875
rect 16316 14872 16344 14912
rect 16482 14900 16488 14912
rect 16540 14900 16546 14952
rect 16666 14872 16672 14884
rect 14875 14844 16344 14872
rect 16408 14844 16672 14872
rect 14875 14841 14887 14844
rect 14829 14835 14887 14841
rect 16408 14804 16436 14844
rect 16666 14832 16672 14844
rect 16724 14832 16730 14884
rect 11348 14776 16436 14804
rect 16482 14764 16488 14816
rect 16540 14804 16546 14816
rect 16868 14804 16896 14971
rect 17862 14900 17868 14952
rect 17920 14940 17926 14952
rect 18340 14940 18368 14980
rect 18874 14968 18880 14980
rect 18932 14968 18938 15020
rect 22097 15011 22155 15017
rect 22097 14977 22109 15011
rect 22143 14977 22155 15011
rect 22097 14971 22155 14977
rect 19334 14940 19340 14952
rect 17920 14912 18368 14940
rect 18432 14912 19340 14940
rect 17920 14900 17926 14912
rect 17126 14804 17132 14816
rect 16540 14776 17132 14804
rect 16540 14764 16546 14776
rect 17126 14764 17132 14776
rect 17184 14804 17190 14816
rect 18432 14804 18460 14912
rect 19334 14900 19340 14912
rect 19392 14900 19398 14952
rect 19613 14943 19671 14949
rect 19613 14909 19625 14943
rect 19659 14940 19671 14943
rect 21266 14940 21272 14952
rect 19659 14912 21272 14940
rect 19659 14909 19671 14912
rect 19613 14903 19671 14909
rect 21266 14900 21272 14912
rect 21324 14900 21330 14952
rect 18874 14832 18880 14884
rect 18932 14872 18938 14884
rect 22112 14872 22140 14971
rect 22554 14900 22560 14952
rect 22612 14940 22618 14952
rect 22833 14943 22891 14949
rect 22833 14940 22845 14943
rect 22612 14912 22845 14940
rect 22612 14900 22618 14912
rect 22833 14909 22845 14912
rect 22879 14909 22891 14943
rect 25041 14943 25099 14949
rect 25041 14940 25053 14943
rect 22833 14903 22891 14909
rect 22940 14912 25053 14940
rect 18932 14844 19472 14872
rect 18932 14832 18938 14844
rect 17184 14776 18460 14804
rect 17184 14764 17190 14776
rect 18598 14764 18604 14816
rect 18656 14764 18662 14816
rect 19444 14804 19472 14844
rect 20640 14844 22140 14872
rect 22281 14875 22339 14881
rect 20640 14804 20668 14844
rect 22281 14841 22293 14875
rect 22327 14872 22339 14875
rect 22462 14872 22468 14884
rect 22327 14844 22468 14872
rect 22327 14841 22339 14844
rect 22281 14835 22339 14841
rect 22462 14832 22468 14844
rect 22520 14832 22526 14884
rect 22738 14832 22744 14884
rect 22796 14872 22802 14884
rect 22940 14872 22968 14912
rect 25041 14909 25053 14912
rect 25087 14909 25099 14943
rect 25041 14903 25099 14909
rect 22796 14844 22968 14872
rect 22796 14832 22802 14844
rect 19444 14776 20668 14804
rect 1104 14714 25852 14736
rect 1104 14662 2950 14714
rect 3002 14662 3014 14714
rect 3066 14662 3078 14714
rect 3130 14662 3142 14714
rect 3194 14662 3206 14714
rect 3258 14662 12950 14714
rect 13002 14662 13014 14714
rect 13066 14662 13078 14714
rect 13130 14662 13142 14714
rect 13194 14662 13206 14714
rect 13258 14662 22950 14714
rect 23002 14662 23014 14714
rect 23066 14662 23078 14714
rect 23130 14662 23142 14714
rect 23194 14662 23206 14714
rect 23258 14662 25852 14714
rect 1104 14640 25852 14662
rect 10413 14603 10471 14609
rect 10413 14569 10425 14603
rect 10459 14600 10471 14603
rect 10502 14600 10508 14612
rect 10459 14572 10508 14600
rect 10459 14569 10471 14572
rect 10413 14563 10471 14569
rect 10502 14560 10508 14572
rect 10560 14560 10566 14612
rect 11146 14560 11152 14612
rect 11204 14600 11210 14612
rect 11204 14572 12388 14600
rect 11204 14560 11210 14572
rect 10965 14467 11023 14473
rect 10965 14433 10977 14467
rect 11011 14464 11023 14467
rect 12250 14464 12256 14476
rect 11011 14436 12256 14464
rect 11011 14433 11023 14436
rect 10965 14427 11023 14433
rect 12250 14424 12256 14436
rect 12308 14424 12314 14476
rect 10686 14356 10692 14408
rect 10744 14356 10750 14408
rect 12360 14328 12388 14572
rect 12434 14560 12440 14612
rect 12492 14560 12498 14612
rect 12897 14603 12955 14609
rect 12897 14569 12909 14603
rect 12943 14600 12955 14603
rect 13354 14600 13360 14612
rect 12943 14572 13360 14600
rect 12943 14569 12955 14572
rect 12897 14563 12955 14569
rect 13354 14560 13360 14572
rect 13412 14560 13418 14612
rect 13449 14603 13507 14609
rect 13449 14569 13461 14603
rect 13495 14600 13507 14603
rect 15930 14600 15936 14612
rect 13495 14572 15936 14600
rect 13495 14569 13507 14572
rect 13449 14563 13507 14569
rect 13556 14473 13584 14572
rect 15930 14560 15936 14572
rect 15988 14560 15994 14612
rect 16114 14560 16120 14612
rect 16172 14600 16178 14612
rect 19429 14603 19487 14609
rect 16172 14572 19380 14600
rect 16172 14560 16178 14572
rect 16025 14535 16083 14541
rect 16025 14501 16037 14535
rect 16071 14532 16083 14535
rect 16206 14532 16212 14544
rect 16071 14504 16212 14532
rect 16071 14501 16083 14504
rect 16025 14495 16083 14501
rect 16206 14492 16212 14504
rect 16264 14492 16270 14544
rect 18233 14535 18291 14541
rect 18233 14501 18245 14535
rect 18279 14532 18291 14535
rect 18690 14532 18696 14544
rect 18279 14504 18696 14532
rect 18279 14501 18291 14504
rect 18233 14495 18291 14501
rect 18690 14492 18696 14504
rect 18748 14492 18754 14544
rect 19352 14532 19380 14572
rect 19429 14569 19441 14603
rect 19475 14600 19487 14603
rect 19978 14600 19984 14612
rect 19475 14572 19984 14600
rect 19475 14569 19487 14572
rect 19429 14563 19487 14569
rect 19978 14560 19984 14572
rect 20036 14560 20042 14612
rect 20254 14560 20260 14612
rect 20312 14600 20318 14612
rect 20441 14603 20499 14609
rect 20441 14600 20453 14603
rect 20312 14572 20453 14600
rect 20312 14560 20318 14572
rect 20441 14569 20453 14572
rect 20487 14600 20499 14603
rect 20898 14600 20904 14612
rect 20487 14572 20904 14600
rect 20487 14569 20499 14572
rect 20441 14563 20499 14569
rect 20898 14560 20904 14572
rect 20956 14560 20962 14612
rect 22094 14560 22100 14612
rect 22152 14600 22158 14612
rect 22554 14600 22560 14612
rect 22152 14572 22560 14600
rect 22152 14560 22158 14572
rect 22554 14560 22560 14572
rect 22612 14560 22618 14612
rect 22925 14603 22983 14609
rect 22925 14569 22937 14603
rect 22971 14600 22983 14603
rect 23750 14600 23756 14612
rect 22971 14572 23756 14600
rect 22971 14569 22983 14572
rect 22925 14563 22983 14569
rect 23750 14560 23756 14572
rect 23808 14560 23814 14612
rect 25130 14560 25136 14612
rect 25188 14600 25194 14612
rect 25225 14603 25283 14609
rect 25225 14600 25237 14603
rect 25188 14572 25237 14600
rect 25188 14560 25194 14572
rect 25225 14569 25237 14572
rect 25271 14600 25283 14603
rect 26142 14600 26148 14612
rect 25271 14572 26148 14600
rect 25271 14569 25283 14572
rect 25225 14563 25283 14569
rect 26142 14560 26148 14572
rect 26200 14560 26206 14612
rect 19352 14504 20484 14532
rect 13541 14467 13599 14473
rect 13541 14433 13553 14467
rect 13587 14433 13599 14467
rect 13541 14427 13599 14433
rect 14274 14424 14280 14476
rect 14332 14424 14338 14476
rect 14550 14424 14556 14476
rect 14608 14424 14614 14476
rect 16761 14467 16819 14473
rect 16761 14433 16773 14467
rect 16807 14464 16819 14467
rect 18598 14464 18604 14476
rect 16807 14436 18604 14464
rect 16807 14433 16819 14436
rect 16761 14427 16819 14433
rect 18598 14424 18604 14436
rect 18656 14464 18662 14476
rect 19981 14467 20039 14473
rect 19981 14464 19993 14467
rect 18656 14436 19993 14464
rect 18656 14424 18662 14436
rect 19981 14433 19993 14436
rect 20027 14433 20039 14467
rect 19981 14427 20039 14433
rect 13081 14399 13139 14405
rect 13081 14365 13093 14399
rect 13127 14396 13139 14399
rect 13998 14396 14004 14408
rect 13127 14368 14004 14396
rect 13127 14365 13139 14368
rect 13081 14359 13139 14365
rect 13998 14356 14004 14368
rect 14056 14356 14062 14408
rect 16482 14356 16488 14408
rect 16540 14356 16546 14408
rect 19886 14356 19892 14408
rect 19944 14356 19950 14408
rect 14090 14328 14096 14340
rect 12190 14300 12296 14328
rect 12360 14300 14096 14328
rect 10042 14220 10048 14272
rect 10100 14260 10106 14272
rect 12268 14260 12296 14300
rect 14090 14288 14096 14300
rect 14148 14288 14154 14340
rect 15010 14288 15016 14340
rect 15068 14288 15074 14340
rect 16666 14288 16672 14340
rect 16724 14328 16730 14340
rect 18693 14331 18751 14337
rect 16724 14300 17250 14328
rect 16724 14288 16730 14300
rect 18693 14297 18705 14331
rect 18739 14328 18751 14331
rect 19797 14331 19855 14337
rect 19797 14328 19809 14331
rect 18739 14300 19809 14328
rect 18739 14297 18751 14300
rect 18693 14291 18751 14297
rect 19797 14297 19809 14300
rect 19843 14297 19855 14331
rect 20456 14328 20484 14504
rect 20530 14492 20536 14544
rect 20588 14532 20594 14544
rect 25409 14535 25467 14541
rect 20588 14504 25268 14532
rect 20588 14492 20594 14504
rect 25240 14476 25268 14504
rect 25409 14501 25421 14535
rect 25455 14532 25467 14535
rect 25590 14532 25596 14544
rect 25455 14504 25596 14532
rect 25455 14501 25467 14504
rect 25409 14495 25467 14501
rect 25590 14492 25596 14504
rect 25648 14492 25654 14544
rect 23382 14464 23388 14476
rect 20548 14436 23388 14464
rect 20548 14408 20576 14436
rect 23382 14424 23388 14436
rect 23440 14424 23446 14476
rect 23566 14424 23572 14476
rect 23624 14464 23630 14476
rect 23753 14467 23811 14473
rect 23753 14464 23765 14467
rect 23624 14436 23765 14464
rect 23624 14424 23630 14436
rect 23753 14433 23765 14436
rect 23799 14433 23811 14467
rect 23753 14427 23811 14433
rect 23937 14467 23995 14473
rect 23937 14433 23949 14467
rect 23983 14464 23995 14467
rect 24578 14464 24584 14476
rect 23983 14436 24584 14464
rect 23983 14433 23995 14436
rect 23937 14427 23995 14433
rect 24578 14424 24584 14436
rect 24636 14424 24642 14476
rect 25222 14424 25228 14476
rect 25280 14424 25286 14476
rect 20530 14356 20536 14408
rect 20588 14356 20594 14408
rect 20809 14399 20867 14405
rect 20809 14365 20821 14399
rect 20855 14396 20867 14399
rect 21450 14396 21456 14408
rect 20855 14368 21456 14396
rect 20855 14365 20867 14368
rect 20809 14359 20867 14365
rect 21450 14356 21456 14368
rect 21508 14356 21514 14408
rect 22066 14368 23336 14396
rect 20456 14300 20576 14328
rect 19797 14291 19855 14297
rect 12710 14260 12716 14272
rect 10100 14232 12716 14260
rect 10100 14220 10106 14232
rect 12710 14220 12716 14232
rect 12768 14220 12774 14272
rect 13630 14220 13636 14272
rect 13688 14260 13694 14272
rect 16758 14260 16764 14272
rect 13688 14232 16764 14260
rect 13688 14220 13694 14232
rect 16758 14220 16764 14232
rect 16816 14220 16822 14272
rect 18598 14220 18604 14272
rect 18656 14260 18662 14272
rect 19150 14260 19156 14272
rect 18656 14232 19156 14260
rect 18656 14220 18662 14232
rect 19150 14220 19156 14232
rect 19208 14220 19214 14272
rect 20548 14260 20576 14300
rect 20622 14288 20628 14340
rect 20680 14328 20686 14340
rect 22066 14328 22094 14368
rect 20680 14300 22094 14328
rect 20680 14288 20686 14300
rect 22554 14288 22560 14340
rect 22612 14288 22618 14340
rect 22830 14288 22836 14340
rect 22888 14288 22894 14340
rect 22848 14260 22876 14288
rect 23308 14269 23336 14368
rect 23658 14356 23664 14408
rect 23716 14396 23722 14408
rect 24673 14399 24731 14405
rect 24673 14396 24685 14399
rect 23716 14368 24685 14396
rect 23716 14356 23722 14368
rect 24673 14365 24685 14368
rect 24719 14365 24731 14399
rect 24673 14359 24731 14365
rect 25590 14356 25596 14408
rect 25648 14396 25654 14408
rect 25866 14396 25872 14408
rect 25648 14368 25872 14396
rect 25648 14356 25654 14368
rect 25866 14356 25872 14368
rect 25924 14356 25930 14408
rect 20548 14232 22876 14260
rect 23293 14263 23351 14269
rect 23293 14229 23305 14263
rect 23339 14229 23351 14263
rect 23293 14223 23351 14229
rect 23658 14220 23664 14272
rect 23716 14220 23722 14272
rect 24302 14220 24308 14272
rect 24360 14260 24366 14272
rect 24765 14263 24823 14269
rect 24765 14260 24777 14263
rect 24360 14232 24777 14260
rect 24360 14220 24366 14232
rect 24765 14229 24777 14232
rect 24811 14229 24823 14263
rect 24765 14223 24823 14229
rect 1104 14170 25852 14192
rect 1104 14118 7950 14170
rect 8002 14118 8014 14170
rect 8066 14118 8078 14170
rect 8130 14118 8142 14170
rect 8194 14118 8206 14170
rect 8258 14118 17950 14170
rect 18002 14118 18014 14170
rect 18066 14118 18078 14170
rect 18130 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 25852 14170
rect 1104 14096 25852 14118
rect 11790 14016 11796 14068
rect 11848 14016 11854 14068
rect 12437 14059 12495 14065
rect 12437 14025 12449 14059
rect 12483 14056 12495 14059
rect 12526 14056 12532 14068
rect 12483 14028 12532 14056
rect 12483 14025 12495 14028
rect 12437 14019 12495 14025
rect 12526 14016 12532 14028
rect 12584 14016 12590 14068
rect 13081 14059 13139 14065
rect 13081 14025 13093 14059
rect 13127 14056 13139 14059
rect 13630 14056 13636 14068
rect 13127 14028 13636 14056
rect 13127 14025 13139 14028
rect 13081 14019 13139 14025
rect 13630 14016 13636 14028
rect 13688 14016 13694 14068
rect 13722 14016 13728 14068
rect 13780 14056 13786 14068
rect 13780 14028 14412 14056
rect 13780 14016 13786 14028
rect 11333 13991 11391 13997
rect 11333 13957 11345 13991
rect 11379 13988 11391 13991
rect 13538 13988 13544 14000
rect 11379 13960 13544 13988
rect 11379 13957 11391 13960
rect 11333 13951 11391 13957
rect 11149 13923 11207 13929
rect 11149 13889 11161 13923
rect 11195 13920 11207 13923
rect 11974 13920 11980 13932
rect 11195 13892 11980 13920
rect 11195 13889 11207 13892
rect 11149 13883 11207 13889
rect 11974 13880 11980 13892
rect 12032 13880 12038 13932
rect 12636 13929 12664 13960
rect 13538 13948 13544 13960
rect 13596 13948 13602 14000
rect 14274 13988 14280 14000
rect 13740 13960 14280 13988
rect 13740 13929 13768 13960
rect 14274 13948 14280 13960
rect 14332 13948 14338 14000
rect 14384 13988 14412 14028
rect 14642 14016 14648 14068
rect 14700 14056 14706 14068
rect 15473 14059 15531 14065
rect 15473 14056 15485 14059
rect 14700 14028 15485 14056
rect 14700 14016 14706 14028
rect 15473 14025 15485 14028
rect 15519 14025 15531 14059
rect 15473 14019 15531 14025
rect 16117 14059 16175 14065
rect 16117 14025 16129 14059
rect 16163 14056 16175 14059
rect 16390 14056 16396 14068
rect 16163 14028 16396 14056
rect 16163 14025 16175 14028
rect 16117 14019 16175 14025
rect 16390 14016 16396 14028
rect 16448 14016 16454 14068
rect 17494 14016 17500 14068
rect 17552 14016 17558 14068
rect 17604 14028 18644 14056
rect 17604 13988 17632 14028
rect 14384 13960 14490 13988
rect 16316 13960 17632 13988
rect 18233 13991 18291 13997
rect 12621 13923 12679 13929
rect 12621 13889 12633 13923
rect 12667 13920 12679 13923
rect 13265 13923 13323 13929
rect 12667 13892 12701 13920
rect 12667 13889 12679 13892
rect 12621 13883 12679 13889
rect 13265 13889 13277 13923
rect 13311 13889 13323 13923
rect 13265 13883 13323 13889
rect 13725 13923 13783 13929
rect 13725 13889 13737 13923
rect 13771 13889 13783 13923
rect 13725 13883 13783 13889
rect 13280 13852 13308 13883
rect 15010 13880 15016 13932
rect 15068 13920 15074 13932
rect 16316 13929 16344 13960
rect 18233 13957 18245 13991
rect 18279 13988 18291 13991
rect 18506 13988 18512 14000
rect 18279 13960 18512 13988
rect 18279 13957 18291 13960
rect 18233 13951 18291 13957
rect 15749 13923 15807 13929
rect 15749 13920 15761 13923
rect 15068 13892 15761 13920
rect 15068 13880 15074 13892
rect 15749 13889 15761 13892
rect 15795 13889 15807 13923
rect 15749 13883 15807 13889
rect 16301 13923 16359 13929
rect 16301 13889 16313 13923
rect 16347 13889 16359 13923
rect 16301 13883 16359 13889
rect 13998 13852 14004 13864
rect 13280 13824 14004 13852
rect 13998 13812 14004 13824
rect 14056 13852 14062 13864
rect 14366 13852 14372 13864
rect 14056 13824 14372 13852
rect 14056 13812 14062 13824
rect 14366 13812 14372 13824
rect 14424 13812 14430 13864
rect 15764 13852 15792 13883
rect 17402 13880 17408 13932
rect 17460 13880 17466 13932
rect 16666 13852 16672 13864
rect 15764 13824 16672 13852
rect 16666 13812 16672 13824
rect 16724 13812 16730 13864
rect 17586 13812 17592 13864
rect 17644 13812 17650 13864
rect 15562 13744 15568 13796
rect 15620 13784 15626 13796
rect 18248 13784 18276 13951
rect 18506 13948 18512 13960
rect 18564 13948 18570 14000
rect 18616 13988 18644 14028
rect 19334 14016 19340 14068
rect 19392 14056 19398 14068
rect 19521 14059 19579 14065
rect 19521 14056 19533 14059
rect 19392 14028 19533 14056
rect 19392 14016 19398 14028
rect 19521 14025 19533 14028
rect 19567 14025 19579 14059
rect 19521 14019 19579 14025
rect 20254 14016 20260 14068
rect 20312 14016 20318 14068
rect 20438 14016 20444 14068
rect 20496 14056 20502 14068
rect 21177 14059 21235 14065
rect 21177 14056 21189 14059
rect 20496 14028 21189 14056
rect 20496 14016 20502 14028
rect 21177 14025 21189 14028
rect 21223 14025 21235 14059
rect 22738 14056 22744 14068
rect 21177 14019 21235 14025
rect 22066 14028 22744 14056
rect 20070 13988 20076 14000
rect 18616 13960 20076 13988
rect 20070 13948 20076 13960
rect 20128 13948 20134 14000
rect 21085 13991 21143 13997
rect 21085 13957 21097 13991
rect 21131 13988 21143 13991
rect 22066 13988 22094 14028
rect 22738 14016 22744 14028
rect 22796 14016 22802 14068
rect 23382 13988 23388 14000
rect 21131 13960 22094 13988
rect 22480 13960 23388 13988
rect 21131 13957 21143 13960
rect 21085 13951 21143 13957
rect 19426 13880 19432 13932
rect 19484 13920 19490 13932
rect 22097 13923 22155 13929
rect 22097 13920 22109 13923
rect 19484 13892 22109 13920
rect 19484 13880 19490 13892
rect 22097 13889 22109 13892
rect 22143 13920 22155 13923
rect 22480 13920 22508 13960
rect 23382 13948 23388 13960
rect 23440 13948 23446 14000
rect 23750 13948 23756 14000
rect 23808 13948 23814 14000
rect 25130 13948 25136 14000
rect 25188 13948 25194 14000
rect 22143 13892 22508 13920
rect 22143 13889 22155 13892
rect 22097 13883 22155 13889
rect 22554 13880 22560 13932
rect 22612 13920 22618 13932
rect 22833 13923 22891 13929
rect 22833 13920 22845 13923
rect 22612 13892 22845 13920
rect 22612 13880 22618 13892
rect 22833 13889 22845 13892
rect 22879 13889 22891 13923
rect 22833 13883 22891 13889
rect 19242 13812 19248 13864
rect 19300 13852 19306 13864
rect 20254 13852 20260 13864
rect 19300 13824 20260 13852
rect 19300 13812 19306 13824
rect 20254 13812 20260 13824
rect 20312 13812 20318 13864
rect 21266 13812 21272 13864
rect 21324 13812 21330 13864
rect 22278 13812 22284 13864
rect 22336 13812 22342 13864
rect 23109 13855 23167 13861
rect 23109 13821 23121 13855
rect 23155 13852 23167 13855
rect 24486 13852 24492 13864
rect 23155 13824 24492 13852
rect 23155 13821 23167 13824
rect 23109 13815 23167 13821
rect 24486 13812 24492 13824
rect 24544 13812 24550 13864
rect 24578 13812 24584 13864
rect 24636 13812 24642 13864
rect 25317 13855 25375 13861
rect 25317 13821 25329 13855
rect 25363 13852 25375 13855
rect 25866 13852 25872 13864
rect 25363 13824 25872 13852
rect 25363 13821 25375 13824
rect 25317 13815 25375 13821
rect 25866 13812 25872 13824
rect 25924 13812 25930 13864
rect 15620 13756 18276 13784
rect 15620 13744 15626 13756
rect 13988 13719 14046 13725
rect 13988 13685 14000 13719
rect 14034 13716 14046 13719
rect 15194 13716 15200 13728
rect 14034 13688 15200 13716
rect 14034 13685 14046 13688
rect 13988 13679 14046 13685
rect 15194 13676 15200 13688
rect 15252 13676 15258 13728
rect 17034 13676 17040 13728
rect 17092 13676 17098 13728
rect 19886 13676 19892 13728
rect 19944 13716 19950 13728
rect 20070 13716 20076 13728
rect 19944 13688 20076 13716
rect 19944 13676 19950 13688
rect 20070 13676 20076 13688
rect 20128 13676 20134 13728
rect 20714 13676 20720 13728
rect 20772 13676 20778 13728
rect 1104 13626 25852 13648
rect 1104 13574 2950 13626
rect 3002 13574 3014 13626
rect 3066 13574 3078 13626
rect 3130 13574 3142 13626
rect 3194 13574 3206 13626
rect 3258 13574 12950 13626
rect 13002 13574 13014 13626
rect 13066 13574 13078 13626
rect 13130 13574 13142 13626
rect 13194 13574 13206 13626
rect 13258 13574 22950 13626
rect 23002 13574 23014 13626
rect 23066 13574 23078 13626
rect 23130 13574 23142 13626
rect 23194 13574 23206 13626
rect 23258 13574 25852 13626
rect 1104 13552 25852 13574
rect 12710 13472 12716 13524
rect 12768 13512 12774 13524
rect 13722 13512 13728 13524
rect 12768 13484 13728 13512
rect 12768 13472 12774 13484
rect 13722 13472 13728 13484
rect 13780 13512 13786 13524
rect 13817 13515 13875 13521
rect 13817 13512 13829 13515
rect 13780 13484 13829 13512
rect 13780 13472 13786 13484
rect 13817 13481 13829 13484
rect 13863 13481 13875 13515
rect 13817 13475 13875 13481
rect 15194 13472 15200 13524
rect 15252 13512 15258 13524
rect 16025 13515 16083 13521
rect 16025 13512 16037 13515
rect 15252 13484 16037 13512
rect 15252 13472 15258 13484
rect 16025 13481 16037 13484
rect 16071 13512 16083 13515
rect 16298 13512 16304 13524
rect 16071 13484 16304 13512
rect 16071 13481 16083 13484
rect 16025 13475 16083 13481
rect 16298 13472 16304 13484
rect 16356 13472 16362 13524
rect 16574 13472 16580 13524
rect 16632 13472 16638 13524
rect 18693 13515 18751 13521
rect 18693 13481 18705 13515
rect 18739 13512 18751 13515
rect 19058 13512 19064 13524
rect 18739 13484 19064 13512
rect 18739 13481 18751 13484
rect 18693 13475 18751 13481
rect 19058 13472 19064 13484
rect 19116 13472 19122 13524
rect 19610 13512 19616 13524
rect 19352 13484 19616 13512
rect 13354 13404 13360 13456
rect 13412 13444 13418 13456
rect 13541 13447 13599 13453
rect 13541 13444 13553 13447
rect 13412 13416 13553 13444
rect 13412 13404 13418 13416
rect 13541 13413 13553 13416
rect 13587 13444 13599 13447
rect 16592 13444 16620 13472
rect 13587 13416 14412 13444
rect 13587 13413 13599 13416
rect 13541 13407 13599 13413
rect 12066 13336 12072 13388
rect 12124 13336 12130 13388
rect 14274 13336 14280 13388
rect 14332 13336 14338 13388
rect 14384 13376 14412 13416
rect 15580 13416 16620 13444
rect 15580 13376 15608 13416
rect 14384 13348 15608 13376
rect 16482 13336 16488 13388
rect 16540 13336 16546 13388
rect 16761 13379 16819 13385
rect 16761 13345 16773 13379
rect 16807 13376 16819 13379
rect 18690 13376 18696 13388
rect 16807 13348 18696 13376
rect 16807 13345 16819 13348
rect 16761 13339 16819 13345
rect 18690 13336 18696 13348
rect 18748 13336 18754 13388
rect 11793 13311 11851 13317
rect 11793 13277 11805 13311
rect 11839 13277 11851 13311
rect 11793 13271 11851 13277
rect 18877 13311 18935 13317
rect 18877 13277 18889 13311
rect 18923 13308 18935 13311
rect 19352 13308 19380 13484
rect 19610 13472 19616 13484
rect 19668 13512 19674 13524
rect 20530 13512 20536 13524
rect 19668 13484 20536 13512
rect 19668 13472 19674 13484
rect 20530 13472 20536 13484
rect 20588 13472 20594 13524
rect 21266 13472 21272 13524
rect 21324 13512 21330 13524
rect 21453 13515 21511 13521
rect 21453 13512 21465 13515
rect 21324 13484 21465 13512
rect 21324 13472 21330 13484
rect 21453 13481 21465 13484
rect 21499 13481 21511 13515
rect 21453 13475 21511 13481
rect 22176 13515 22234 13521
rect 22176 13481 22188 13515
rect 22222 13512 22234 13515
rect 23198 13512 23204 13524
rect 22222 13484 23204 13512
rect 22222 13481 22234 13484
rect 22176 13475 22234 13481
rect 23198 13472 23204 13484
rect 23256 13472 23262 13524
rect 23474 13472 23480 13524
rect 23532 13512 23538 13524
rect 23937 13515 23995 13521
rect 23937 13512 23949 13515
rect 23532 13484 23949 13512
rect 23532 13472 23538 13484
rect 23937 13481 23949 13484
rect 23983 13481 23995 13515
rect 23937 13475 23995 13481
rect 23750 13404 23756 13456
rect 23808 13444 23814 13456
rect 24121 13447 24179 13453
rect 24121 13444 24133 13447
rect 23808 13416 24133 13444
rect 23808 13404 23814 13416
rect 24121 13413 24133 13416
rect 24167 13413 24179 13447
rect 24121 13407 24179 13413
rect 21910 13376 21916 13388
rect 19720 13348 21916 13376
rect 18923 13280 19380 13308
rect 18923 13277 18935 13280
rect 18877 13271 18935 13277
rect 9585 13243 9643 13249
rect 9585 13209 9597 13243
rect 9631 13240 9643 13243
rect 11514 13240 11520 13252
rect 9631 13212 11520 13240
rect 9631 13209 9643 13212
rect 9585 13203 9643 13209
rect 11514 13200 11520 13212
rect 11572 13200 11578 13252
rect 10042 13132 10048 13184
rect 10100 13172 10106 13184
rect 10686 13172 10692 13184
rect 10100 13144 10692 13172
rect 10100 13132 10106 13144
rect 10686 13132 10692 13144
rect 10744 13172 10750 13184
rect 10873 13175 10931 13181
rect 10873 13172 10885 13175
rect 10744 13144 10885 13172
rect 10744 13132 10750 13144
rect 10873 13141 10885 13144
rect 10919 13172 10931 13175
rect 11808 13172 11836 13271
rect 19426 13268 19432 13320
rect 19484 13308 19490 13320
rect 19720 13317 19748 13348
rect 21910 13336 21916 13348
rect 21968 13336 21974 13388
rect 22646 13336 22652 13388
rect 22704 13376 22710 13388
rect 22830 13376 22836 13388
rect 22704 13348 22836 13376
rect 22704 13336 22710 13348
rect 22830 13336 22836 13348
rect 22888 13336 22894 13388
rect 23198 13336 23204 13388
rect 23256 13376 23262 13388
rect 25133 13379 25191 13385
rect 25133 13376 25145 13379
rect 23256 13348 25145 13376
rect 23256 13336 23262 13348
rect 25133 13345 25145 13348
rect 25179 13345 25191 13379
rect 25133 13339 25191 13345
rect 19705 13311 19763 13317
rect 19705 13308 19717 13311
rect 19484 13280 19717 13308
rect 19484 13268 19490 13280
rect 19705 13277 19717 13280
rect 19751 13277 19763 13311
rect 19705 13271 19763 13277
rect 25041 13311 25099 13317
rect 25041 13277 25053 13311
rect 25087 13308 25099 13311
rect 25314 13308 25320 13320
rect 25087 13280 25320 13308
rect 25087 13277 25099 13280
rect 25041 13271 25099 13277
rect 25314 13268 25320 13280
rect 25372 13268 25378 13320
rect 12710 13200 12716 13252
rect 12768 13200 12774 13252
rect 14182 13200 14188 13252
rect 14240 13240 14246 13252
rect 14550 13240 14556 13252
rect 14240 13212 14556 13240
rect 14240 13200 14246 13212
rect 14550 13200 14556 13212
rect 14608 13200 14614 13252
rect 15010 13240 15016 13252
rect 14660 13212 15016 13240
rect 10919 13144 11836 13172
rect 10919 13141 10931 13144
rect 10873 13135 10931 13141
rect 13722 13132 13728 13184
rect 13780 13172 13786 13184
rect 14660 13172 14688 13212
rect 15010 13200 15016 13212
rect 15068 13200 15074 13252
rect 16482 13200 16488 13252
rect 16540 13240 16546 13252
rect 17218 13240 17224 13252
rect 16540 13212 17224 13240
rect 16540 13200 16546 13212
rect 17218 13200 17224 13212
rect 17276 13200 17282 13252
rect 19337 13243 19395 13249
rect 19337 13209 19349 13243
rect 19383 13240 19395 13243
rect 19886 13240 19892 13252
rect 19383 13212 19892 13240
rect 19383 13209 19395 13212
rect 19337 13203 19395 13209
rect 19886 13200 19892 13212
rect 19944 13200 19950 13252
rect 19981 13243 20039 13249
rect 19981 13209 19993 13243
rect 20027 13209 20039 13243
rect 19981 13203 20039 13209
rect 13780 13144 14688 13172
rect 13780 13132 13786 13144
rect 16298 13132 16304 13184
rect 16356 13172 16362 13184
rect 17586 13172 17592 13184
rect 16356 13144 17592 13172
rect 16356 13132 16362 13144
rect 17586 13132 17592 13144
rect 17644 13172 17650 13184
rect 18233 13175 18291 13181
rect 18233 13172 18245 13175
rect 17644 13144 18245 13172
rect 17644 13132 17650 13144
rect 18233 13141 18245 13144
rect 18279 13141 18291 13175
rect 19996 13172 20024 13203
rect 20254 13200 20260 13252
rect 20312 13240 20318 13252
rect 23750 13240 23756 13252
rect 20312 13212 20470 13240
rect 23414 13212 23756 13240
rect 20312 13200 20318 13212
rect 23750 13200 23756 13212
rect 23808 13200 23814 13252
rect 24026 13200 24032 13252
rect 24084 13240 24090 13252
rect 24397 13243 24455 13249
rect 24397 13240 24409 13243
rect 24084 13212 24409 13240
rect 24084 13200 24090 13212
rect 24397 13209 24409 13212
rect 24443 13240 24455 13243
rect 24949 13243 25007 13249
rect 24949 13240 24961 13243
rect 24443 13212 24961 13240
rect 24443 13209 24455 13212
rect 24397 13203 24455 13209
rect 24949 13209 24961 13212
rect 24995 13209 25007 13243
rect 24949 13203 25007 13209
rect 20806 13172 20812 13184
rect 19996 13144 20812 13172
rect 18233 13135 18291 13141
rect 20806 13132 20812 13144
rect 20864 13172 20870 13184
rect 23661 13175 23719 13181
rect 23661 13172 23673 13175
rect 20864 13144 23673 13172
rect 20864 13132 20870 13144
rect 23661 13141 23673 13144
rect 23707 13141 23719 13175
rect 23661 13135 23719 13141
rect 24486 13132 24492 13184
rect 24544 13172 24550 13184
rect 24581 13175 24639 13181
rect 24581 13172 24593 13175
rect 24544 13144 24593 13172
rect 24544 13132 24550 13144
rect 24581 13141 24593 13144
rect 24627 13141 24639 13175
rect 24581 13135 24639 13141
rect 1104 13082 25852 13104
rect 1104 13030 7950 13082
rect 8002 13030 8014 13082
rect 8066 13030 8078 13082
rect 8130 13030 8142 13082
rect 8194 13030 8206 13082
rect 8258 13030 17950 13082
rect 18002 13030 18014 13082
rect 18066 13030 18078 13082
rect 18130 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 25852 13082
rect 1104 13008 25852 13030
rect 11514 12928 11520 12980
rect 11572 12968 11578 12980
rect 12621 12971 12679 12977
rect 11572 12940 12434 12968
rect 11572 12928 11578 12940
rect 12406 12900 12434 12940
rect 12621 12937 12633 12971
rect 12667 12968 12679 12971
rect 12710 12968 12716 12980
rect 12667 12940 12716 12968
rect 12667 12937 12679 12940
rect 12621 12931 12679 12937
rect 12710 12928 12716 12940
rect 12768 12928 12774 12980
rect 13814 12928 13820 12980
rect 13872 12968 13878 12980
rect 14274 12968 14280 12980
rect 13872 12940 14280 12968
rect 13872 12928 13878 12940
rect 14274 12928 14280 12940
rect 14332 12928 14338 12980
rect 15010 12928 15016 12980
rect 15068 12968 15074 12980
rect 16301 12971 16359 12977
rect 16301 12968 16313 12971
rect 15068 12940 16313 12968
rect 15068 12928 15074 12940
rect 16301 12937 16313 12940
rect 16347 12968 16359 12971
rect 16482 12968 16488 12980
rect 16347 12940 16488 12968
rect 16347 12937 16359 12940
rect 16301 12931 16359 12937
rect 16482 12928 16488 12940
rect 16540 12928 16546 12980
rect 17862 12968 17868 12980
rect 17144 12940 17868 12968
rect 12989 12903 13047 12909
rect 12989 12900 13001 12903
rect 12406 12872 13001 12900
rect 12989 12869 13001 12872
rect 13035 12900 13047 12903
rect 15562 12900 15568 12912
rect 13035 12872 15568 12900
rect 13035 12869 13047 12872
rect 12989 12863 13047 12869
rect 15562 12860 15568 12872
rect 15620 12860 15626 12912
rect 17144 12909 17172 12940
rect 17862 12928 17868 12940
rect 17920 12968 17926 12980
rect 18690 12968 18696 12980
rect 17920 12940 18696 12968
rect 17920 12928 17926 12940
rect 18690 12928 18696 12940
rect 18748 12928 18754 12980
rect 19518 12928 19524 12980
rect 19576 12968 19582 12980
rect 20717 12971 20775 12977
rect 20717 12968 20729 12971
rect 19576 12940 20729 12968
rect 19576 12928 19582 12940
rect 20717 12937 20729 12940
rect 20763 12937 20775 12971
rect 20717 12931 20775 12937
rect 21361 12971 21419 12977
rect 21361 12937 21373 12971
rect 21407 12968 21419 12971
rect 21450 12968 21456 12980
rect 21407 12940 21456 12968
rect 21407 12937 21419 12940
rect 21361 12931 21419 12937
rect 21450 12928 21456 12940
rect 21508 12928 21514 12980
rect 23198 12928 23204 12980
rect 23256 12968 23262 12980
rect 23753 12971 23811 12977
rect 23753 12968 23765 12971
rect 23256 12940 23765 12968
rect 23256 12928 23262 12940
rect 23753 12937 23765 12940
rect 23799 12937 23811 12971
rect 23753 12931 23811 12937
rect 25501 12971 25559 12977
rect 25501 12937 25513 12971
rect 25547 12968 25559 12971
rect 25682 12968 25688 12980
rect 25547 12940 25688 12968
rect 25547 12937 25559 12940
rect 25501 12931 25559 12937
rect 25682 12928 25688 12940
rect 25740 12928 25746 12980
rect 17129 12903 17187 12909
rect 17129 12869 17141 12903
rect 17175 12869 17187 12903
rect 17129 12863 17187 12869
rect 17218 12860 17224 12912
rect 17276 12900 17282 12912
rect 17586 12900 17592 12912
rect 17276 12872 17592 12900
rect 17276 12860 17282 12872
rect 17586 12860 17592 12872
rect 17644 12860 17650 12912
rect 18782 12860 18788 12912
rect 18840 12900 18846 12912
rect 22370 12900 22376 12912
rect 18840 12872 22376 12900
rect 18840 12860 18846 12872
rect 22370 12860 22376 12872
rect 22428 12860 22434 12912
rect 25041 12903 25099 12909
rect 25041 12900 25053 12903
rect 24228 12872 25053 12900
rect 24228 12844 24256 12872
rect 25041 12869 25053 12872
rect 25087 12869 25099 12903
rect 25041 12863 25099 12869
rect 25317 12903 25375 12909
rect 25317 12869 25329 12903
rect 25363 12900 25375 12903
rect 25958 12900 25964 12912
rect 25363 12872 25964 12900
rect 25363 12869 25375 12872
rect 25317 12863 25375 12869
rect 25958 12860 25964 12872
rect 26016 12860 26022 12912
rect 16850 12792 16856 12844
rect 16908 12792 16914 12844
rect 18506 12792 18512 12844
rect 18564 12832 18570 12844
rect 19429 12835 19487 12841
rect 19429 12832 19441 12835
rect 18564 12804 19441 12832
rect 18564 12792 18570 12804
rect 19429 12801 19441 12804
rect 19475 12801 19487 12835
rect 19429 12795 19487 12801
rect 20622 12792 20628 12844
rect 20680 12792 20686 12844
rect 21453 12835 21511 12841
rect 21453 12832 21465 12835
rect 20732 12804 21465 12832
rect 15194 12724 15200 12776
rect 15252 12724 15258 12776
rect 15473 12767 15531 12773
rect 15473 12733 15485 12767
rect 15519 12764 15531 12767
rect 16666 12764 16672 12776
rect 15519 12736 16672 12764
rect 15519 12733 15531 12736
rect 15473 12727 15531 12733
rect 16666 12724 16672 12736
rect 16724 12724 16730 12776
rect 17586 12724 17592 12776
rect 17644 12764 17650 12776
rect 17862 12764 17868 12776
rect 17644 12736 17868 12764
rect 17644 12724 17650 12736
rect 17862 12724 17868 12736
rect 17920 12724 17926 12776
rect 18414 12724 18420 12776
rect 18472 12764 18478 12776
rect 19521 12767 19579 12773
rect 19521 12764 19533 12767
rect 18472 12736 19533 12764
rect 18472 12724 18478 12736
rect 19521 12733 19533 12736
rect 19567 12733 19579 12767
rect 19521 12727 19579 12733
rect 19613 12767 19671 12773
rect 19613 12733 19625 12767
rect 19659 12733 19671 12767
rect 19613 12727 19671 12733
rect 18598 12656 18604 12708
rect 18656 12696 18662 12708
rect 19628 12696 19656 12727
rect 20254 12724 20260 12776
rect 20312 12764 20318 12776
rect 20732 12764 20760 12804
rect 21453 12801 21465 12804
rect 21499 12801 21511 12835
rect 21453 12795 21511 12801
rect 21910 12792 21916 12844
rect 21968 12832 21974 12844
rect 22005 12835 22063 12841
rect 22005 12832 22017 12835
rect 21968 12804 22017 12832
rect 21968 12792 21974 12804
rect 22005 12801 22017 12804
rect 22051 12801 22063 12835
rect 23750 12832 23756 12844
rect 23414 12804 23756 12832
rect 22005 12795 22063 12801
rect 23750 12792 23756 12804
rect 23808 12832 23814 12844
rect 24029 12835 24087 12841
rect 24029 12832 24041 12835
rect 23808 12804 24041 12832
rect 23808 12792 23814 12804
rect 24029 12801 24041 12804
rect 24075 12832 24087 12835
rect 24210 12832 24216 12844
rect 24075 12804 24216 12832
rect 24075 12801 24087 12804
rect 24029 12795 24087 12801
rect 24210 12792 24216 12804
rect 24268 12792 24274 12844
rect 24394 12792 24400 12844
rect 24452 12832 24458 12844
rect 24765 12835 24823 12841
rect 24765 12832 24777 12835
rect 24452 12804 24777 12832
rect 24452 12792 24458 12804
rect 24765 12801 24777 12804
rect 24811 12801 24823 12835
rect 24765 12795 24823 12801
rect 20312 12736 20760 12764
rect 20809 12767 20867 12773
rect 20312 12724 20318 12736
rect 20809 12733 20821 12767
rect 20855 12733 20867 12767
rect 20809 12727 20867 12733
rect 18656 12668 19656 12696
rect 18656 12656 18662 12668
rect 20438 12656 20444 12708
rect 20496 12696 20502 12708
rect 20824 12696 20852 12727
rect 20990 12724 20996 12776
rect 21048 12764 21054 12776
rect 21542 12764 21548 12776
rect 21048 12736 21548 12764
rect 21048 12724 21054 12736
rect 21542 12724 21548 12736
rect 21600 12724 21606 12776
rect 22278 12724 22284 12776
rect 22336 12724 22342 12776
rect 20496 12668 20852 12696
rect 20496 12656 20502 12668
rect 23474 12656 23480 12708
rect 23532 12696 23538 12708
rect 24581 12699 24639 12705
rect 24581 12696 24593 12699
rect 23532 12668 24593 12696
rect 23532 12656 23538 12668
rect 24581 12665 24593 12668
rect 24627 12665 24639 12699
rect 24581 12659 24639 12665
rect 19061 12631 19119 12637
rect 19061 12597 19073 12631
rect 19107 12628 19119 12631
rect 19794 12628 19800 12640
rect 19107 12600 19800 12628
rect 19107 12597 19119 12600
rect 19061 12591 19119 12597
rect 19794 12588 19800 12600
rect 19852 12588 19858 12640
rect 20254 12588 20260 12640
rect 20312 12588 20318 12640
rect 1104 12538 25852 12560
rect 1104 12486 2950 12538
rect 3002 12486 3014 12538
rect 3066 12486 3078 12538
rect 3130 12486 3142 12538
rect 3194 12486 3206 12538
rect 3258 12486 12950 12538
rect 13002 12486 13014 12538
rect 13066 12486 13078 12538
rect 13130 12486 13142 12538
rect 13194 12486 13206 12538
rect 13258 12486 22950 12538
rect 23002 12486 23014 12538
rect 23066 12486 23078 12538
rect 23130 12486 23142 12538
rect 23194 12486 23206 12538
rect 23258 12486 25852 12538
rect 1104 12464 25852 12486
rect 4062 12384 4068 12436
rect 4120 12424 4126 12436
rect 4120 12396 6914 12424
rect 4120 12384 4126 12396
rect 6886 12220 6914 12396
rect 8570 12384 8576 12436
rect 8628 12424 8634 12436
rect 13449 12427 13507 12433
rect 13449 12424 13461 12427
rect 8628 12396 13461 12424
rect 8628 12384 8634 12396
rect 13449 12393 13461 12396
rect 13495 12393 13507 12427
rect 13449 12387 13507 12393
rect 13464 12288 13492 12387
rect 13722 12384 13728 12436
rect 13780 12384 13786 12436
rect 13909 12427 13967 12433
rect 13909 12393 13921 12427
rect 13955 12424 13967 12427
rect 13998 12424 14004 12436
rect 13955 12396 14004 12424
rect 13955 12393 13967 12396
rect 13909 12387 13967 12393
rect 13998 12384 14004 12396
rect 14056 12384 14062 12436
rect 15473 12427 15531 12433
rect 15473 12393 15485 12427
rect 15519 12424 15531 12427
rect 15562 12424 15568 12436
rect 15519 12396 15568 12424
rect 15519 12393 15531 12396
rect 15473 12387 15531 12393
rect 15562 12384 15568 12396
rect 15620 12384 15626 12436
rect 17497 12427 17555 12433
rect 17497 12393 17509 12427
rect 17543 12424 17555 12427
rect 17586 12424 17592 12436
rect 17543 12396 17592 12424
rect 17543 12393 17555 12396
rect 17497 12387 17555 12393
rect 17586 12384 17592 12396
rect 17644 12384 17650 12436
rect 22738 12384 22744 12436
rect 22796 12424 22802 12436
rect 22796 12396 25084 12424
rect 22796 12384 22802 12396
rect 24210 12316 24216 12368
rect 24268 12356 24274 12368
rect 24397 12359 24455 12365
rect 24397 12356 24409 12359
rect 24268 12328 24409 12356
rect 24268 12316 24274 12328
rect 24397 12325 24409 12328
rect 24443 12356 24455 12359
rect 24673 12359 24731 12365
rect 24673 12356 24685 12359
rect 24443 12328 24685 12356
rect 24443 12325 24455 12328
rect 24397 12319 24455 12325
rect 24673 12325 24685 12328
rect 24719 12325 24731 12359
rect 24673 12319 24731 12325
rect 14277 12291 14335 12297
rect 14277 12288 14289 12291
rect 13464 12260 14289 12288
rect 14277 12257 14289 12260
rect 14323 12257 14335 12291
rect 14277 12251 14335 12257
rect 15749 12291 15807 12297
rect 15749 12257 15761 12291
rect 15795 12288 15807 12291
rect 16758 12288 16764 12300
rect 15795 12260 16764 12288
rect 15795 12257 15807 12260
rect 15749 12251 15807 12257
rect 16758 12248 16764 12260
rect 16816 12248 16822 12300
rect 17402 12248 17408 12300
rect 17460 12288 17466 12300
rect 17957 12291 18015 12297
rect 17957 12288 17969 12291
rect 17460 12260 17969 12288
rect 17460 12248 17466 12260
rect 17957 12257 17969 12260
rect 18003 12257 18015 12291
rect 17957 12251 18015 12257
rect 19794 12248 19800 12300
rect 19852 12288 19858 12300
rect 20438 12288 20444 12300
rect 19852 12260 20444 12288
rect 19852 12248 19858 12260
rect 20438 12248 20444 12260
rect 20496 12288 20502 12300
rect 21177 12291 21235 12297
rect 21177 12288 21189 12291
rect 20496 12260 21189 12288
rect 20496 12248 20502 12260
rect 21177 12257 21189 12260
rect 21223 12257 21235 12291
rect 21177 12251 21235 12257
rect 21358 12248 21364 12300
rect 21416 12288 21422 12300
rect 21910 12288 21916 12300
rect 21416 12260 21916 12288
rect 21416 12248 21422 12260
rect 21910 12248 21916 12260
rect 21968 12288 21974 12300
rect 22281 12291 22339 12297
rect 22281 12288 22293 12291
rect 21968 12260 22293 12288
rect 21968 12248 21974 12260
rect 22281 12257 22293 12260
rect 22327 12257 22339 12291
rect 22281 12251 22339 12257
rect 22557 12291 22615 12297
rect 22557 12257 22569 12291
rect 22603 12288 22615 12291
rect 24578 12288 24584 12300
rect 22603 12260 24584 12288
rect 22603 12257 22615 12260
rect 22557 12251 22615 12257
rect 24578 12248 24584 12260
rect 24636 12248 24642 12300
rect 25056 12297 25084 12396
rect 25041 12291 25099 12297
rect 25041 12257 25053 12291
rect 25087 12257 25099 12291
rect 25041 12251 25099 12257
rect 14553 12223 14611 12229
rect 6886 12192 12434 12220
rect 12406 12152 12434 12192
rect 14553 12189 14565 12223
rect 14599 12220 14611 12223
rect 15562 12220 15568 12232
rect 14599 12192 15568 12220
rect 14599 12189 14611 12192
rect 14553 12183 14611 12189
rect 15562 12180 15568 12192
rect 15620 12180 15626 12232
rect 19334 12180 19340 12232
rect 19392 12220 19398 12232
rect 19429 12223 19487 12229
rect 19429 12220 19441 12223
rect 19392 12192 19441 12220
rect 19392 12180 19398 12192
rect 19429 12189 19441 12192
rect 19475 12189 19487 12223
rect 19429 12183 19487 12189
rect 16025 12155 16083 12161
rect 12406 12124 15976 12152
rect 15948 12084 15976 12124
rect 16025 12121 16037 12155
rect 16071 12152 16083 12155
rect 16298 12152 16304 12164
rect 16071 12124 16304 12152
rect 16071 12121 16083 12124
rect 16025 12115 16083 12121
rect 16298 12112 16304 12124
rect 16356 12112 16362 12164
rect 16482 12112 16488 12164
rect 16540 12112 16546 12164
rect 18693 12155 18751 12161
rect 18693 12121 18705 12155
rect 18739 12152 18751 12155
rect 19610 12152 19616 12164
rect 18739 12124 19616 12152
rect 18739 12121 18751 12124
rect 18693 12115 18751 12121
rect 18708 12084 18736 12115
rect 19610 12112 19616 12124
rect 19668 12112 19674 12164
rect 19702 12112 19708 12164
rect 19760 12112 19766 12164
rect 20162 12112 20168 12164
rect 20220 12112 20226 12164
rect 21637 12155 21695 12161
rect 21637 12152 21649 12155
rect 21100 12124 21649 12152
rect 15948 12056 18736 12084
rect 18785 12087 18843 12093
rect 18785 12053 18797 12087
rect 18831 12084 18843 12087
rect 19978 12084 19984 12096
rect 18831 12056 19984 12084
rect 18831 12053 18843 12056
rect 18785 12047 18843 12053
rect 19978 12044 19984 12056
rect 20036 12044 20042 12096
rect 20622 12044 20628 12096
rect 20680 12084 20686 12096
rect 21100 12084 21128 12124
rect 21637 12121 21649 12124
rect 21683 12121 21695 12155
rect 24210 12152 24216 12164
rect 23782 12124 24216 12152
rect 21637 12115 21695 12121
rect 24210 12112 24216 12124
rect 24268 12112 24274 12164
rect 20680 12056 21128 12084
rect 20680 12044 20686 12056
rect 22370 12044 22376 12096
rect 22428 12084 22434 12096
rect 24029 12087 24087 12093
rect 24029 12084 24041 12087
rect 22428 12056 24041 12084
rect 22428 12044 22434 12056
rect 24029 12053 24041 12056
rect 24075 12053 24087 12087
rect 24029 12047 24087 12053
rect 1104 11994 25852 12016
rect 1104 11942 7950 11994
rect 8002 11942 8014 11994
rect 8066 11942 8078 11994
rect 8130 11942 8142 11994
rect 8194 11942 8206 11994
rect 8258 11942 17950 11994
rect 18002 11942 18014 11994
rect 18066 11942 18078 11994
rect 18130 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 25852 11994
rect 1104 11920 25852 11942
rect 13814 11880 13820 11892
rect 12820 11852 13820 11880
rect 12820 11753 12848 11852
rect 13814 11840 13820 11852
rect 13872 11840 13878 11892
rect 14550 11840 14556 11892
rect 14608 11840 14614 11892
rect 15105 11883 15163 11889
rect 15105 11849 15117 11883
rect 15151 11880 15163 11883
rect 15657 11883 15715 11889
rect 15151 11852 15240 11880
rect 15151 11849 15163 11852
rect 15105 11843 15163 11849
rect 13081 11815 13139 11821
rect 13081 11781 13093 11815
rect 13127 11812 13139 11815
rect 13354 11812 13360 11824
rect 13127 11784 13360 11812
rect 13127 11781 13139 11784
rect 13081 11775 13139 11781
rect 13354 11772 13360 11784
rect 13412 11772 13418 11824
rect 13722 11772 13728 11824
rect 13780 11772 13786 11824
rect 12805 11747 12863 11753
rect 12805 11713 12817 11747
rect 12851 11713 12863 11747
rect 12805 11707 12863 11713
rect 15212 11676 15240 11852
rect 15657 11849 15669 11883
rect 15703 11880 15715 11883
rect 15746 11880 15752 11892
rect 15703 11852 15752 11880
rect 15703 11849 15715 11852
rect 15657 11843 15715 11849
rect 15289 11747 15347 11753
rect 15289 11713 15301 11747
rect 15335 11744 15347 11747
rect 15672 11744 15700 11843
rect 15746 11840 15752 11852
rect 15804 11840 15810 11892
rect 19334 11880 19340 11892
rect 17052 11852 19340 11880
rect 15335 11716 15700 11744
rect 16301 11747 16359 11753
rect 15335 11713 15347 11716
rect 15289 11707 15347 11713
rect 16301 11713 16313 11747
rect 16347 11744 16359 11747
rect 16758 11744 16764 11756
rect 16347 11716 16764 11744
rect 16347 11713 16359 11716
rect 16301 11707 16359 11713
rect 16758 11704 16764 11716
rect 16816 11704 16822 11756
rect 16850 11676 16856 11688
rect 15212 11648 16856 11676
rect 16850 11636 16856 11648
rect 16908 11636 16914 11688
rect 17052 11676 17080 11852
rect 19334 11840 19340 11852
rect 19392 11840 19398 11892
rect 21453 11883 21511 11889
rect 21453 11880 21465 11883
rect 19444 11852 21465 11880
rect 17678 11772 17684 11824
rect 17736 11812 17742 11824
rect 17736 11784 17894 11812
rect 17736 11772 17742 11784
rect 19150 11772 19156 11824
rect 19208 11812 19214 11824
rect 19444 11812 19472 11852
rect 21453 11849 21465 11852
rect 21499 11849 21511 11883
rect 21453 11843 21511 11849
rect 19208 11784 19472 11812
rect 19705 11815 19763 11821
rect 19208 11772 19214 11784
rect 19705 11781 19717 11815
rect 19751 11812 19763 11815
rect 19794 11812 19800 11824
rect 19751 11784 19800 11812
rect 19751 11781 19763 11784
rect 19705 11775 19763 11781
rect 19794 11772 19800 11784
rect 19852 11772 19858 11824
rect 20162 11772 20168 11824
rect 20220 11772 20226 11824
rect 23293 11815 23351 11821
rect 23293 11781 23305 11815
rect 23339 11812 23351 11815
rect 24854 11812 24860 11824
rect 23339 11784 24860 11812
rect 23339 11781 23351 11784
rect 23293 11775 23351 11781
rect 24854 11772 24860 11784
rect 24912 11772 24918 11824
rect 25130 11772 25136 11824
rect 25188 11772 25194 11824
rect 19426 11704 19432 11756
rect 19484 11704 19490 11756
rect 22186 11704 22192 11756
rect 22244 11704 22250 11756
rect 23937 11747 23995 11753
rect 23937 11713 23949 11747
rect 23983 11713 23995 11747
rect 23937 11707 23995 11713
rect 17129 11679 17187 11685
rect 17129 11676 17141 11679
rect 17052 11648 17141 11676
rect 17129 11645 17141 11648
rect 17175 11645 17187 11679
rect 17129 11639 17187 11645
rect 17405 11679 17463 11685
rect 17405 11645 17417 11679
rect 17451 11676 17463 11679
rect 18598 11676 18604 11688
rect 17451 11648 18604 11676
rect 17451 11645 17463 11648
rect 17405 11639 17463 11645
rect 18598 11636 18604 11648
rect 18656 11636 18662 11688
rect 19536 11648 20852 11676
rect 14458 11568 14464 11620
rect 14516 11608 14522 11620
rect 16117 11611 16175 11617
rect 16117 11608 16129 11611
rect 14516 11580 16129 11608
rect 14516 11568 14522 11580
rect 16117 11577 16129 11580
rect 16163 11577 16175 11611
rect 16117 11571 16175 11577
rect 18506 11568 18512 11620
rect 18564 11608 18570 11620
rect 19536 11608 19564 11648
rect 20824 11620 20852 11648
rect 20898 11636 20904 11688
rect 20956 11676 20962 11688
rect 23952 11676 23980 11707
rect 20956 11648 23980 11676
rect 20956 11636 20962 11648
rect 18564 11580 19564 11608
rect 18564 11568 18570 11580
rect 20806 11568 20812 11620
rect 20864 11568 20870 11620
rect 21082 11568 21088 11620
rect 21140 11608 21146 11620
rect 21177 11611 21235 11617
rect 21177 11608 21189 11611
rect 21140 11580 21189 11608
rect 21140 11568 21146 11580
rect 21177 11577 21189 11580
rect 21223 11608 21235 11611
rect 21634 11608 21640 11620
rect 21223 11580 21640 11608
rect 21223 11577 21235 11580
rect 21177 11571 21235 11577
rect 21634 11568 21640 11580
rect 21692 11568 21698 11620
rect 14642 11500 14648 11552
rect 14700 11540 14706 11552
rect 15749 11543 15807 11549
rect 15749 11540 15761 11543
rect 14700 11512 15761 11540
rect 14700 11500 14706 11512
rect 15749 11509 15761 11512
rect 15795 11509 15807 11543
rect 15749 11503 15807 11509
rect 16758 11500 16764 11552
rect 16816 11540 16822 11552
rect 18782 11540 18788 11552
rect 16816 11512 18788 11540
rect 16816 11500 16822 11512
rect 18782 11500 18788 11512
rect 18840 11500 18846 11552
rect 18877 11543 18935 11549
rect 18877 11509 18889 11543
rect 18923 11540 18935 11543
rect 19702 11540 19708 11552
rect 18923 11512 19708 11540
rect 18923 11509 18935 11512
rect 18877 11503 18935 11509
rect 19702 11500 19708 11512
rect 19760 11500 19766 11552
rect 20824 11540 20852 11568
rect 21266 11540 21272 11552
rect 20824 11512 21272 11540
rect 21266 11500 21272 11512
rect 21324 11500 21330 11552
rect 21542 11500 21548 11552
rect 21600 11540 21606 11552
rect 24486 11540 24492 11552
rect 21600 11512 24492 11540
rect 21600 11500 21606 11512
rect 24486 11500 24492 11512
rect 24544 11500 24550 11552
rect 1104 11450 25852 11472
rect 1104 11398 2950 11450
rect 3002 11398 3014 11450
rect 3066 11398 3078 11450
rect 3130 11398 3142 11450
rect 3194 11398 3206 11450
rect 3258 11398 12950 11450
rect 13002 11398 13014 11450
rect 13066 11398 13078 11450
rect 13130 11398 13142 11450
rect 13194 11398 13206 11450
rect 13258 11398 22950 11450
rect 23002 11398 23014 11450
rect 23066 11398 23078 11450
rect 23130 11398 23142 11450
rect 23194 11398 23206 11450
rect 23258 11398 25852 11450
rect 1104 11376 25852 11398
rect 12526 11296 12532 11348
rect 12584 11336 12590 11348
rect 13722 11336 13728 11348
rect 12584 11308 13728 11336
rect 12584 11296 12590 11308
rect 13722 11296 13728 11308
rect 13780 11336 13786 11348
rect 14642 11336 14648 11348
rect 13780 11308 14648 11336
rect 13780 11296 13786 11308
rect 14642 11296 14648 11308
rect 14700 11296 14706 11348
rect 15470 11296 15476 11348
rect 15528 11296 15534 11348
rect 16114 11296 16120 11348
rect 16172 11296 16178 11348
rect 16761 11339 16819 11345
rect 16761 11305 16773 11339
rect 16807 11336 16819 11339
rect 16942 11336 16948 11348
rect 16807 11308 16948 11336
rect 16807 11305 16819 11308
rect 16761 11299 16819 11305
rect 16942 11296 16948 11308
rect 17000 11296 17006 11348
rect 17405 11339 17463 11345
rect 17405 11305 17417 11339
rect 17451 11336 17463 11339
rect 17494 11336 17500 11348
rect 17451 11308 17500 11336
rect 17451 11305 17463 11308
rect 17405 11299 17463 11305
rect 17494 11296 17500 11308
rect 17552 11296 17558 11348
rect 19242 11296 19248 11348
rect 19300 11296 19306 11348
rect 19518 11296 19524 11348
rect 19576 11296 19582 11348
rect 19610 11296 19616 11348
rect 19668 11336 19674 11348
rect 20441 11339 20499 11345
rect 20441 11336 20453 11339
rect 19668 11308 20453 11336
rect 19668 11296 19674 11308
rect 20441 11305 20453 11308
rect 20487 11305 20499 11339
rect 20441 11299 20499 11305
rect 20806 11296 20812 11348
rect 20864 11296 20870 11348
rect 21177 11339 21235 11345
rect 21177 11305 21189 11339
rect 21223 11336 21235 11339
rect 23382 11336 23388 11348
rect 21223 11308 23388 11336
rect 21223 11305 21235 11308
rect 21177 11299 21235 11305
rect 23382 11296 23388 11308
rect 23440 11296 23446 11348
rect 24578 11296 24584 11348
rect 24636 11296 24642 11348
rect 24762 11296 24768 11348
rect 24820 11336 24826 11348
rect 25225 11339 25283 11345
rect 25225 11336 25237 11339
rect 24820 11308 25237 11336
rect 24820 11296 24826 11308
rect 25225 11305 25237 11308
rect 25271 11305 25283 11339
rect 25225 11299 25283 11305
rect 25501 11339 25559 11345
rect 25501 11305 25513 11339
rect 25547 11336 25559 11339
rect 25682 11336 25688 11348
rect 25547 11308 25688 11336
rect 25547 11305 25559 11308
rect 25501 11299 25559 11305
rect 25682 11296 25688 11308
rect 25740 11296 25746 11348
rect 18693 11271 18751 11277
rect 18693 11237 18705 11271
rect 18739 11268 18751 11271
rect 19794 11268 19800 11280
rect 18739 11240 19800 11268
rect 18739 11237 18751 11240
rect 18693 11231 18751 11237
rect 19794 11228 19800 11240
rect 19852 11228 19858 11280
rect 20254 11228 20260 11280
rect 20312 11268 20318 11280
rect 22005 11271 22063 11277
rect 22005 11268 22017 11271
rect 20312 11240 22017 11268
rect 20312 11228 20318 11240
rect 22005 11237 22017 11240
rect 22051 11237 22063 11271
rect 22005 11231 22063 11237
rect 22370 11228 22376 11280
rect 22428 11268 22434 11280
rect 22646 11268 22652 11280
rect 22428 11240 22652 11268
rect 22428 11228 22434 11240
rect 22646 11228 22652 11240
rect 22704 11228 22710 11280
rect 25133 11271 25191 11277
rect 25133 11237 25145 11271
rect 25179 11268 25191 11271
rect 25958 11268 25964 11280
rect 25179 11240 25964 11268
rect 25179 11237 25191 11240
rect 25133 11231 25191 11237
rect 25958 11228 25964 11240
rect 26016 11228 26022 11280
rect 18049 11203 18107 11209
rect 18049 11169 18061 11203
rect 18095 11200 18107 11203
rect 18414 11200 18420 11212
rect 18095 11172 18420 11200
rect 18095 11169 18107 11172
rect 18049 11163 18107 11169
rect 18414 11160 18420 11172
rect 18472 11160 18478 11212
rect 21542 11200 21548 11212
rect 18892 11172 21548 11200
rect 15654 11092 15660 11144
rect 15712 11092 15718 11144
rect 16022 11092 16028 11144
rect 16080 11132 16086 11144
rect 16301 11135 16359 11141
rect 16301 11132 16313 11135
rect 16080 11104 16313 11132
rect 16080 11092 16086 11104
rect 16301 11101 16313 11104
rect 16347 11101 16359 11135
rect 16301 11095 16359 11101
rect 16945 11135 17003 11141
rect 16945 11101 16957 11135
rect 16991 11132 17003 11135
rect 17126 11132 17132 11144
rect 16991 11104 17132 11132
rect 16991 11101 17003 11104
rect 16945 11095 17003 11101
rect 17126 11092 17132 11104
rect 17184 11092 17190 11144
rect 17589 11135 17647 11141
rect 17589 11101 17601 11135
rect 17635 11132 17647 11135
rect 18506 11132 18512 11144
rect 17635 11104 18512 11132
rect 17635 11101 17647 11104
rect 17589 11095 17647 11101
rect 18506 11092 18512 11104
rect 18564 11092 18570 11144
rect 18892 11141 18920 11172
rect 21542 11160 21548 11172
rect 21600 11160 21606 11212
rect 23845 11203 23903 11209
rect 23845 11169 23857 11203
rect 23891 11200 23903 11203
rect 24854 11200 24860 11212
rect 23891 11172 24860 11200
rect 23891 11169 23903 11172
rect 23845 11163 23903 11169
rect 24854 11160 24860 11172
rect 24912 11160 24918 11212
rect 18877 11135 18935 11141
rect 18877 11101 18889 11135
rect 18923 11101 18935 11135
rect 18877 11095 18935 11101
rect 19150 11092 19156 11144
rect 19208 11132 19214 11144
rect 19981 11135 20039 11141
rect 19981 11132 19993 11135
rect 19208 11104 19993 11132
rect 19208 11092 19214 11104
rect 19981 11101 19993 11104
rect 20027 11101 20039 11135
rect 19981 11095 20039 11101
rect 20070 11092 20076 11144
rect 20128 11132 20134 11144
rect 21361 11135 21419 11141
rect 21361 11132 21373 11135
rect 20128 11104 21373 11132
rect 20128 11092 20134 11104
rect 21361 11101 21373 11104
rect 21407 11101 21419 11135
rect 21361 11095 21419 11101
rect 22189 11135 22247 11141
rect 22189 11101 22201 11135
rect 22235 11132 22247 11135
rect 22278 11132 22284 11144
rect 22235 11104 22284 11132
rect 22235 11101 22247 11104
rect 22189 11095 22247 11101
rect 22278 11092 22284 11104
rect 22336 11092 22342 11144
rect 22646 11092 22652 11144
rect 22704 11092 22710 11144
rect 24762 11092 24768 11144
rect 24820 11092 24826 11144
rect 15562 11024 15568 11076
rect 15620 11064 15626 11076
rect 23934 11064 23940 11076
rect 15620 11036 23940 11064
rect 15620 11024 15626 11036
rect 23934 11024 23940 11036
rect 23992 11024 23998 11076
rect 20070 10956 20076 11008
rect 20128 10956 20134 11008
rect 20162 10956 20168 11008
rect 20220 10996 20226 11008
rect 20625 10999 20683 11005
rect 20625 10996 20637 10999
rect 20220 10968 20637 10996
rect 20220 10956 20226 10968
rect 20625 10965 20637 10968
rect 20671 10996 20683 10999
rect 21082 10996 21088 11008
rect 20671 10968 21088 10996
rect 20671 10965 20683 10968
rect 20625 10959 20683 10965
rect 21082 10956 21088 10968
rect 21140 10956 21146 11008
rect 21266 10956 21272 11008
rect 21324 10996 21330 11008
rect 21637 10999 21695 11005
rect 21637 10996 21649 10999
rect 21324 10968 21649 10996
rect 21324 10956 21330 10968
rect 21637 10965 21649 10968
rect 21683 10996 21695 10999
rect 21726 10996 21732 11008
rect 21683 10968 21732 10996
rect 21683 10965 21695 10968
rect 21637 10959 21695 10965
rect 21726 10956 21732 10968
rect 21784 10956 21790 11008
rect 1104 10906 25852 10928
rect 1104 10854 7950 10906
rect 8002 10854 8014 10906
rect 8066 10854 8078 10906
rect 8130 10854 8142 10906
rect 8194 10854 8206 10906
rect 8258 10854 17950 10906
rect 18002 10854 18014 10906
rect 18066 10854 18078 10906
rect 18130 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 25852 10906
rect 1104 10832 25852 10854
rect 15654 10752 15660 10804
rect 15712 10792 15718 10804
rect 15749 10795 15807 10801
rect 15749 10792 15761 10795
rect 15712 10764 15761 10792
rect 15712 10752 15718 10764
rect 15749 10761 15761 10764
rect 15795 10761 15807 10795
rect 15749 10755 15807 10761
rect 16022 10752 16028 10804
rect 16080 10792 16086 10804
rect 16393 10795 16451 10801
rect 16393 10792 16405 10795
rect 16080 10764 16405 10792
rect 16080 10752 16086 10764
rect 16393 10761 16405 10764
rect 16439 10761 16451 10795
rect 16393 10755 16451 10761
rect 17126 10752 17132 10804
rect 17184 10752 17190 10804
rect 17313 10795 17371 10801
rect 17313 10761 17325 10795
rect 17359 10792 17371 10795
rect 17405 10795 17463 10801
rect 17405 10792 17417 10795
rect 17359 10764 17417 10792
rect 17359 10761 17371 10764
rect 17313 10755 17371 10761
rect 17405 10761 17417 10764
rect 17451 10792 17463 10795
rect 17862 10792 17868 10804
rect 17451 10764 17868 10792
rect 17451 10761 17463 10764
rect 17405 10755 17463 10761
rect 17862 10752 17868 10764
rect 17920 10752 17926 10804
rect 18049 10795 18107 10801
rect 18049 10761 18061 10795
rect 18095 10792 18107 10795
rect 18322 10792 18328 10804
rect 18095 10764 18328 10792
rect 18095 10761 18107 10764
rect 18049 10755 18107 10761
rect 18322 10752 18328 10764
rect 18380 10752 18386 10804
rect 19337 10795 19395 10801
rect 19337 10761 19349 10795
rect 19383 10792 19395 10795
rect 20990 10792 20996 10804
rect 19383 10764 20996 10792
rect 19383 10761 19395 10764
rect 19337 10755 19395 10761
rect 20990 10752 20996 10764
rect 21048 10752 21054 10804
rect 21082 10752 21088 10804
rect 21140 10792 21146 10804
rect 21910 10792 21916 10804
rect 21140 10764 21916 10792
rect 21140 10752 21146 10764
rect 21910 10752 21916 10764
rect 21968 10752 21974 10804
rect 20530 10724 20536 10736
rect 19536 10696 20536 10724
rect 16945 10659 17003 10665
rect 16945 10625 16957 10659
rect 16991 10656 17003 10659
rect 18233 10659 18291 10665
rect 18233 10656 18245 10659
rect 16991 10628 18245 10656
rect 16991 10625 17003 10628
rect 16945 10619 17003 10625
rect 18233 10625 18245 10628
rect 18279 10656 18291 10659
rect 18690 10656 18696 10668
rect 18279 10628 18696 10656
rect 18279 10625 18291 10628
rect 18233 10619 18291 10625
rect 18690 10616 18696 10628
rect 18748 10616 18754 10668
rect 19536 10665 19564 10696
rect 20530 10684 20536 10696
rect 20588 10684 20594 10736
rect 23293 10727 23351 10733
rect 20640 10696 22140 10724
rect 18877 10659 18935 10665
rect 18877 10625 18889 10659
rect 18923 10625 18935 10659
rect 18877 10619 18935 10625
rect 19521 10659 19579 10665
rect 19521 10625 19533 10659
rect 19567 10625 19579 10659
rect 19521 10619 19579 10625
rect 18892 10588 18920 10619
rect 20162 10616 20168 10668
rect 20220 10616 20226 10668
rect 20438 10616 20444 10668
rect 20496 10656 20502 10668
rect 20640 10656 20668 10696
rect 20496 10628 20668 10656
rect 20496 10616 20502 10628
rect 20714 10616 20720 10668
rect 20772 10656 20778 10668
rect 22112 10665 22140 10696
rect 23293 10693 23305 10727
rect 23339 10724 23351 10727
rect 24854 10724 24860 10736
rect 23339 10696 24860 10724
rect 23339 10693 23351 10696
rect 23293 10687 23351 10693
rect 24854 10684 24860 10696
rect 24912 10684 24918 10736
rect 20809 10659 20867 10665
rect 20809 10656 20821 10659
rect 20772 10628 20821 10656
rect 20772 10616 20778 10628
rect 20809 10625 20821 10628
rect 20855 10625 20867 10659
rect 20809 10619 20867 10625
rect 21453 10659 21511 10665
rect 21453 10625 21465 10659
rect 21499 10625 21511 10659
rect 21453 10619 21511 10625
rect 22097 10659 22155 10665
rect 22097 10625 22109 10659
rect 22143 10625 22155 10659
rect 22097 10619 22155 10625
rect 21266 10588 21272 10600
rect 18892 10560 21272 10588
rect 21266 10548 21272 10560
rect 21324 10548 21330 10600
rect 21468 10588 21496 10619
rect 23934 10616 23940 10668
rect 23992 10616 23998 10668
rect 23290 10588 23296 10600
rect 21468 10560 23296 10588
rect 23290 10548 23296 10560
rect 23348 10548 23354 10600
rect 24670 10548 24676 10600
rect 24728 10548 24734 10600
rect 17310 10480 17316 10532
rect 17368 10520 17374 10532
rect 18693 10523 18751 10529
rect 18693 10520 18705 10523
rect 17368 10492 18705 10520
rect 17368 10480 17374 10492
rect 18693 10489 18705 10492
rect 18739 10489 18751 10523
rect 18693 10483 18751 10489
rect 19981 10523 20039 10529
rect 19981 10489 19993 10523
rect 20027 10520 20039 10523
rect 23934 10520 23940 10532
rect 20027 10492 23940 10520
rect 20027 10489 20039 10492
rect 19981 10483 20039 10489
rect 23934 10480 23940 10492
rect 23992 10480 23998 10532
rect 16666 10412 16672 10464
rect 16724 10452 16730 10464
rect 20438 10452 20444 10464
rect 16724 10424 20444 10452
rect 16724 10412 16730 10424
rect 20438 10412 20444 10424
rect 20496 10412 20502 10464
rect 20625 10455 20683 10461
rect 20625 10421 20637 10455
rect 20671 10452 20683 10455
rect 20806 10452 20812 10464
rect 20671 10424 20812 10452
rect 20671 10421 20683 10424
rect 20625 10415 20683 10421
rect 20806 10412 20812 10424
rect 20864 10412 20870 10464
rect 21266 10412 21272 10464
rect 21324 10412 21330 10464
rect 21542 10412 21548 10464
rect 21600 10452 21606 10464
rect 22094 10452 22100 10464
rect 21600 10424 22100 10452
rect 21600 10412 21606 10424
rect 22094 10412 22100 10424
rect 22152 10412 22158 10464
rect 1104 10362 25852 10384
rect 1104 10310 2950 10362
rect 3002 10310 3014 10362
rect 3066 10310 3078 10362
rect 3130 10310 3142 10362
rect 3194 10310 3206 10362
rect 3258 10310 12950 10362
rect 13002 10310 13014 10362
rect 13066 10310 13078 10362
rect 13130 10310 13142 10362
rect 13194 10310 13206 10362
rect 13258 10310 22950 10362
rect 23002 10310 23014 10362
rect 23066 10310 23078 10362
rect 23130 10310 23142 10362
rect 23194 10310 23206 10362
rect 23258 10310 25852 10362
rect 1104 10288 25852 10310
rect 17405 10251 17463 10257
rect 17405 10217 17417 10251
rect 17451 10248 17463 10251
rect 20162 10248 20168 10260
rect 17451 10220 20168 10248
rect 17451 10217 17463 10220
rect 17405 10211 17463 10217
rect 20162 10208 20168 10220
rect 20220 10208 20226 10260
rect 20714 10208 20720 10260
rect 20772 10208 20778 10260
rect 21726 10208 21732 10260
rect 21784 10248 21790 10260
rect 24581 10251 24639 10257
rect 24581 10248 24593 10251
rect 21784 10220 24593 10248
rect 21784 10208 21790 10220
rect 24581 10217 24593 10220
rect 24627 10217 24639 10251
rect 24581 10211 24639 10217
rect 19426 10140 19432 10192
rect 19484 10140 19490 10192
rect 18049 10115 18107 10121
rect 18049 10081 18061 10115
rect 18095 10112 18107 10115
rect 21266 10112 21272 10124
rect 18095 10084 21272 10112
rect 18095 10081 18107 10084
rect 18049 10075 18107 10081
rect 21266 10072 21272 10084
rect 21324 10072 21330 10124
rect 21358 10072 21364 10124
rect 21416 10072 21422 10124
rect 21634 10072 21640 10124
rect 21692 10072 21698 10124
rect 23658 10072 23664 10124
rect 23716 10112 23722 10124
rect 23845 10115 23903 10121
rect 23845 10112 23857 10115
rect 23716 10084 23857 10112
rect 23716 10072 23722 10084
rect 23845 10081 23857 10084
rect 23891 10081 23903 10115
rect 23845 10075 23903 10081
rect 25133 10115 25191 10121
rect 25133 10081 25145 10115
rect 25179 10081 25191 10115
rect 25133 10075 25191 10081
rect 17586 10004 17592 10056
rect 17644 10004 17650 10056
rect 18325 10047 18383 10053
rect 18325 10013 18337 10047
rect 18371 10013 18383 10047
rect 18325 10007 18383 10013
rect 19613 10047 19671 10053
rect 19613 10013 19625 10047
rect 19659 10044 19671 10047
rect 20714 10044 20720 10056
rect 19659 10016 20720 10044
rect 19659 10013 19671 10016
rect 19613 10007 19671 10013
rect 18340 9908 18368 10007
rect 20714 10004 20720 10016
rect 20772 10004 20778 10056
rect 20901 10047 20959 10053
rect 20901 10013 20913 10047
rect 20947 10044 20959 10047
rect 20947 10016 21404 10044
rect 20947 10013 20959 10016
rect 20901 10007 20959 10013
rect 20073 9979 20131 9985
rect 20073 9945 20085 9979
rect 20119 9976 20131 9979
rect 21376 9976 21404 10016
rect 23106 10004 23112 10056
rect 23164 10044 23170 10056
rect 25148 10044 25176 10075
rect 23164 10016 25176 10044
rect 23164 10004 23170 10016
rect 21542 9976 21548 9988
rect 20119 9948 21128 9976
rect 21376 9948 21548 9976
rect 20119 9945 20131 9948
rect 20073 9939 20131 9945
rect 20438 9908 20444 9920
rect 18340 9880 20444 9908
rect 20438 9868 20444 9880
rect 20496 9868 20502 9920
rect 21100 9908 21128 9948
rect 21542 9936 21548 9948
rect 21600 9936 21606 9988
rect 21634 9936 21640 9988
rect 21692 9976 21698 9988
rect 21910 9976 21916 9988
rect 21692 9948 21916 9976
rect 21692 9936 21698 9948
rect 21910 9936 21916 9948
rect 21968 9976 21974 9988
rect 24949 9979 25007 9985
rect 24949 9976 24961 9979
rect 21968 9948 22126 9976
rect 22940 9948 24961 9976
rect 21968 9936 21974 9948
rect 22940 9908 22968 9948
rect 24949 9945 24961 9948
rect 24995 9945 25007 9979
rect 24949 9939 25007 9945
rect 25041 9979 25099 9985
rect 25041 9945 25053 9979
rect 25087 9976 25099 9979
rect 25222 9976 25228 9988
rect 25087 9948 25228 9976
rect 25087 9945 25099 9948
rect 25041 9939 25099 9945
rect 25222 9936 25228 9948
rect 25280 9936 25286 9988
rect 21100 9880 22968 9908
rect 23106 9868 23112 9920
rect 23164 9868 23170 9920
rect 1104 9818 25852 9840
rect 1104 9766 7950 9818
rect 8002 9766 8014 9818
rect 8066 9766 8078 9818
rect 8130 9766 8142 9818
rect 8194 9766 8206 9818
rect 8258 9766 17950 9818
rect 18002 9766 18014 9818
rect 18066 9766 18078 9818
rect 18130 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 25852 9818
rect 1104 9744 25852 9766
rect 19352 9676 20392 9704
rect 17034 9596 17040 9648
rect 17092 9636 17098 9648
rect 19352 9636 19380 9676
rect 17092 9608 19380 9636
rect 17092 9596 17098 9608
rect 8478 9528 8484 9580
rect 8536 9568 8542 9580
rect 18233 9571 18291 9577
rect 18233 9568 18245 9571
rect 8536 9540 18245 9568
rect 8536 9528 8542 9540
rect 18233 9537 18245 9540
rect 18279 9537 18291 9571
rect 18233 9531 18291 9537
rect 18877 9571 18935 9577
rect 18877 9537 18889 9571
rect 18923 9568 18935 9571
rect 19058 9568 19064 9580
rect 18923 9540 19064 9568
rect 18923 9537 18935 9540
rect 18877 9531 18935 9537
rect 19058 9528 19064 9540
rect 19116 9528 19122 9580
rect 19518 9528 19524 9580
rect 19576 9528 19582 9580
rect 20165 9571 20223 9577
rect 20165 9537 20177 9571
rect 20211 9568 20223 9571
rect 20254 9568 20260 9580
rect 20211 9540 20260 9568
rect 20211 9537 20223 9540
rect 20165 9531 20223 9537
rect 20254 9528 20260 9540
rect 20312 9528 20318 9580
rect 20364 9568 20392 9676
rect 20622 9664 20628 9716
rect 20680 9704 20686 9716
rect 23106 9704 23112 9716
rect 20680 9676 23112 9704
rect 20680 9664 20686 9676
rect 23106 9664 23112 9676
rect 23164 9664 23170 9716
rect 20438 9596 20444 9648
rect 20496 9636 20502 9648
rect 20496 9608 22140 9636
rect 20496 9596 20502 9608
rect 20901 9571 20959 9577
rect 20901 9568 20913 9571
rect 20364 9540 20913 9568
rect 20901 9537 20913 9540
rect 20947 9537 20959 9571
rect 20901 9531 20959 9537
rect 21266 9528 21272 9580
rect 21324 9528 21330 9580
rect 21453 9571 21511 9577
rect 21453 9537 21465 9571
rect 21499 9568 21511 9571
rect 21545 9571 21603 9577
rect 21545 9568 21557 9571
rect 21499 9540 21557 9568
rect 21499 9537 21511 9540
rect 21453 9531 21511 9537
rect 21545 9537 21557 9540
rect 21591 9568 21603 9571
rect 21634 9568 21640 9580
rect 21591 9540 21640 9568
rect 21591 9537 21603 9540
rect 21545 9531 21603 9537
rect 21634 9528 21640 9540
rect 21692 9528 21698 9580
rect 22112 9577 22140 9608
rect 23290 9596 23296 9648
rect 23348 9596 23354 9648
rect 22097 9571 22155 9577
rect 22097 9537 22109 9571
rect 22143 9537 22155 9571
rect 22097 9531 22155 9537
rect 23934 9528 23940 9580
rect 23992 9528 23998 9580
rect 22646 9500 22652 9512
rect 18064 9472 22652 9500
rect 18064 9441 18092 9472
rect 22646 9460 22652 9472
rect 22704 9460 22710 9512
rect 24762 9460 24768 9512
rect 24820 9460 24826 9512
rect 18049 9435 18107 9441
rect 18049 9401 18061 9435
rect 18095 9401 18107 9435
rect 18049 9395 18107 9401
rect 19334 9392 19340 9444
rect 19392 9392 19398 9444
rect 17770 9324 17776 9376
rect 17828 9364 17834 9376
rect 18693 9367 18751 9373
rect 18693 9364 18705 9367
rect 17828 9336 18705 9364
rect 17828 9324 17834 9336
rect 18693 9333 18705 9336
rect 18739 9333 18751 9367
rect 18693 9327 18751 9333
rect 19981 9367 20039 9373
rect 19981 9333 19993 9367
rect 20027 9364 20039 9367
rect 20530 9364 20536 9376
rect 20027 9336 20536 9364
rect 20027 9333 20039 9336
rect 19981 9327 20039 9333
rect 20530 9324 20536 9336
rect 20588 9324 20594 9376
rect 20714 9324 20720 9376
rect 20772 9324 20778 9376
rect 1104 9274 25852 9296
rect 1104 9222 2950 9274
rect 3002 9222 3014 9274
rect 3066 9222 3078 9274
rect 3130 9222 3142 9274
rect 3194 9222 3206 9274
rect 3258 9222 12950 9274
rect 13002 9222 13014 9274
rect 13066 9222 13078 9274
rect 13130 9222 13142 9274
rect 13194 9222 13206 9274
rect 13258 9222 22950 9274
rect 23002 9222 23014 9274
rect 23066 9222 23078 9274
rect 23130 9222 23142 9274
rect 23194 9222 23206 9274
rect 23258 9222 25852 9274
rect 1104 9200 25852 9222
rect 11793 9163 11851 9169
rect 11793 9129 11805 9163
rect 11839 9160 11851 9163
rect 14734 9160 14740 9172
rect 11839 9132 14740 9160
rect 11839 9129 11851 9132
rect 11793 9123 11851 9129
rect 14734 9120 14740 9132
rect 14792 9120 14798 9172
rect 19058 9120 19064 9172
rect 19116 9120 19122 9172
rect 19518 9120 19524 9172
rect 19576 9160 19582 9172
rect 20993 9163 21051 9169
rect 20993 9160 21005 9163
rect 19576 9132 21005 9160
rect 19576 9120 19582 9132
rect 20993 9129 21005 9132
rect 21039 9160 21051 9163
rect 21358 9160 21364 9172
rect 21039 9132 21364 9160
rect 21039 9129 21051 9132
rect 20993 9123 21051 9129
rect 21358 9120 21364 9132
rect 21416 9120 21422 9172
rect 22002 9120 22008 9172
rect 22060 9160 22066 9172
rect 23842 9160 23848 9172
rect 22060 9132 23848 9160
rect 22060 9120 22066 9132
rect 23842 9120 23848 9132
rect 23900 9120 23906 9172
rect 25409 9163 25467 9169
rect 25409 9129 25421 9163
rect 25455 9160 25467 9163
rect 25774 9160 25780 9172
rect 25455 9132 25780 9160
rect 25455 9129 25467 9132
rect 25409 9123 25467 9129
rect 25774 9120 25780 9132
rect 25832 9120 25838 9172
rect 21269 9095 21327 9101
rect 21269 9092 21281 9095
rect 19444 9064 21281 9092
rect 10042 8984 10048 9036
rect 10100 8984 10106 9036
rect 19444 9033 19472 9064
rect 21269 9061 21281 9064
rect 21315 9061 21327 9095
rect 21269 9055 21327 9061
rect 22094 9052 22100 9104
rect 22152 9092 22158 9104
rect 22830 9092 22836 9104
rect 22152 9064 22836 9092
rect 22152 9052 22158 9064
rect 22830 9052 22836 9064
rect 22888 9052 22894 9104
rect 19429 9027 19487 9033
rect 19429 8993 19441 9027
rect 19475 8993 19487 9027
rect 19429 8987 19487 8993
rect 19705 9027 19763 9033
rect 19705 8993 19717 9027
rect 19751 9024 19763 9027
rect 22738 9024 22744 9036
rect 19751 8996 22744 9024
rect 19751 8993 19763 8996
rect 19705 8987 19763 8993
rect 22738 8984 22744 8996
rect 22796 8984 22802 9036
rect 23845 9027 23903 9033
rect 23845 8993 23857 9027
rect 23891 9024 23903 9027
rect 24854 9024 24860 9036
rect 23891 8996 24860 9024
rect 23891 8993 23903 8996
rect 23845 8987 23903 8993
rect 24854 8984 24860 8996
rect 24912 8984 24918 9036
rect 21174 8916 21180 8968
rect 21232 8956 21238 8968
rect 21453 8959 21511 8965
rect 21453 8956 21465 8959
rect 21232 8928 21465 8956
rect 21232 8916 21238 8928
rect 21453 8925 21465 8928
rect 21499 8925 21511 8959
rect 21453 8919 21511 8925
rect 21542 8916 21548 8968
rect 21600 8956 21606 8968
rect 22649 8959 22707 8965
rect 22649 8956 22661 8959
rect 21600 8928 22661 8956
rect 21600 8916 21606 8928
rect 22649 8925 22661 8928
rect 22695 8925 22707 8959
rect 22649 8919 22707 8925
rect 9306 8848 9312 8900
rect 9364 8888 9370 8900
rect 10321 8891 10379 8897
rect 10321 8888 10333 8891
rect 9364 8860 10333 8888
rect 9364 8848 9370 8860
rect 10321 8857 10333 8860
rect 10367 8857 10379 8891
rect 12069 8891 12127 8897
rect 12069 8888 12081 8891
rect 11546 8860 12081 8888
rect 10321 8851 10379 8857
rect 12069 8857 12081 8860
rect 12115 8888 12127 8891
rect 12526 8888 12532 8900
rect 12115 8860 12532 8888
rect 12115 8857 12127 8860
rect 12069 8851 12127 8857
rect 12526 8848 12532 8860
rect 12584 8848 12590 8900
rect 20714 8848 20720 8900
rect 20772 8888 20778 8900
rect 21634 8888 21640 8900
rect 20772 8860 21640 8888
rect 20772 8848 20778 8860
rect 21634 8848 21640 8860
rect 21692 8848 21698 8900
rect 21910 8848 21916 8900
rect 21968 8888 21974 8900
rect 24673 8891 24731 8897
rect 24673 8888 24685 8891
rect 21968 8860 24685 8888
rect 21968 8848 21974 8860
rect 24673 8857 24685 8860
rect 24719 8857 24731 8891
rect 24673 8851 24731 8857
rect 20530 8780 20536 8832
rect 20588 8820 20594 8832
rect 21358 8820 21364 8832
rect 20588 8792 21364 8820
rect 20588 8780 20594 8792
rect 21358 8780 21364 8792
rect 21416 8780 21422 8832
rect 22002 8780 22008 8832
rect 22060 8780 22066 8832
rect 22278 8780 22284 8832
rect 22336 8820 22342 8832
rect 24765 8823 24823 8829
rect 24765 8820 24777 8823
rect 22336 8792 24777 8820
rect 22336 8780 22342 8792
rect 24765 8789 24777 8792
rect 24811 8789 24823 8823
rect 24765 8783 24823 8789
rect 1104 8730 25852 8752
rect 1104 8678 7950 8730
rect 8002 8678 8014 8730
rect 8066 8678 8078 8730
rect 8130 8678 8142 8730
rect 8194 8678 8206 8730
rect 8258 8678 17950 8730
rect 18002 8678 18014 8730
rect 18066 8678 18078 8730
rect 18130 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 25852 8730
rect 1104 8656 25852 8678
rect 19429 8619 19487 8625
rect 19429 8585 19441 8619
rect 19475 8616 19487 8619
rect 22186 8616 22192 8628
rect 19475 8588 22192 8616
rect 19475 8585 19487 8588
rect 19429 8579 19487 8585
rect 22186 8576 22192 8588
rect 22244 8576 22250 8628
rect 20272 8520 21312 8548
rect 14826 8440 14832 8492
rect 14884 8480 14890 8492
rect 20272 8489 20300 8520
rect 21284 8489 21312 8520
rect 21358 8508 21364 8560
rect 21416 8548 21422 8560
rect 23293 8551 23351 8557
rect 21416 8520 22232 8548
rect 21416 8508 21422 8520
rect 19613 8483 19671 8489
rect 19613 8480 19625 8483
rect 14884 8452 19625 8480
rect 14884 8440 14890 8452
rect 19613 8449 19625 8452
rect 19659 8449 19671 8483
rect 19613 8443 19671 8449
rect 20257 8483 20315 8489
rect 20257 8449 20269 8483
rect 20303 8449 20315 8483
rect 20257 8443 20315 8449
rect 20901 8483 20959 8489
rect 20901 8449 20913 8483
rect 20947 8449 20959 8483
rect 20901 8443 20959 8449
rect 21269 8483 21327 8489
rect 21269 8449 21281 8483
rect 21315 8480 21327 8483
rect 22002 8480 22008 8492
rect 21315 8452 22008 8480
rect 21315 8449 21327 8452
rect 21269 8443 21327 8449
rect 19886 8372 19892 8424
rect 19944 8412 19950 8424
rect 20916 8412 20944 8443
rect 22002 8440 22008 8452
rect 22060 8440 22066 8492
rect 22097 8483 22155 8489
rect 22097 8449 22109 8483
rect 22143 8449 22155 8483
rect 22204 8480 22232 8520
rect 23293 8517 23305 8551
rect 23339 8548 23351 8551
rect 24854 8548 24860 8560
rect 23339 8520 24860 8548
rect 23339 8517 23351 8520
rect 23293 8511 23351 8517
rect 24854 8508 24860 8520
rect 24912 8508 24918 8560
rect 23937 8483 23995 8489
rect 23937 8480 23949 8483
rect 22204 8452 23949 8480
rect 22097 8443 22155 8449
rect 23937 8449 23949 8452
rect 23983 8449 23995 8483
rect 24946 8480 24952 8492
rect 23937 8443 23995 8449
rect 24044 8452 24952 8480
rect 19944 8384 20944 8412
rect 19944 8372 19950 8384
rect 21450 8372 21456 8424
rect 21508 8372 21514 8424
rect 22112 8412 22140 8443
rect 24044 8412 24072 8452
rect 24946 8440 24952 8452
rect 25004 8440 25010 8492
rect 22112 8384 24072 8412
rect 24578 8372 24584 8424
rect 24636 8372 24642 8424
rect 19702 8304 19708 8356
rect 19760 8344 19766 8356
rect 20073 8347 20131 8353
rect 20073 8344 20085 8347
rect 19760 8316 20085 8344
rect 19760 8304 19766 8316
rect 20073 8313 20085 8316
rect 20119 8313 20131 8347
rect 20073 8307 20131 8313
rect 20717 8347 20775 8353
rect 20717 8313 20729 8347
rect 20763 8344 20775 8347
rect 24394 8344 24400 8356
rect 20763 8316 24400 8344
rect 20763 8313 20775 8316
rect 20717 8307 20775 8313
rect 24394 8304 24400 8316
rect 24452 8304 24458 8356
rect 1104 8186 25852 8208
rect 1104 8134 2950 8186
rect 3002 8134 3014 8186
rect 3066 8134 3078 8186
rect 3130 8134 3142 8186
rect 3194 8134 3206 8186
rect 3258 8134 12950 8186
rect 13002 8134 13014 8186
rect 13066 8134 13078 8186
rect 13130 8134 13142 8186
rect 13194 8134 13206 8186
rect 13258 8134 22950 8186
rect 23002 8134 23014 8186
rect 23066 8134 23078 8186
rect 23130 8134 23142 8186
rect 23194 8134 23206 8186
rect 23258 8134 25852 8186
rect 1104 8112 25852 8134
rect 20898 8032 20904 8084
rect 20956 8072 20962 8084
rect 21361 8075 21419 8081
rect 21361 8072 21373 8075
rect 20956 8044 21373 8072
rect 20956 8032 20962 8044
rect 21361 8041 21373 8044
rect 21407 8041 21419 8075
rect 21361 8035 21419 8041
rect 21910 8032 21916 8084
rect 21968 8072 21974 8084
rect 22005 8075 22063 8081
rect 22005 8072 22017 8075
rect 21968 8044 22017 8072
rect 21968 8032 21974 8044
rect 22005 8041 22017 8044
rect 22051 8041 22063 8075
rect 22005 8035 22063 8041
rect 24026 8004 24032 8016
rect 20088 7976 24032 8004
rect 20088 7945 20116 7976
rect 24026 7964 24032 7976
rect 24084 7964 24090 8016
rect 19981 7939 20039 7945
rect 19981 7905 19993 7939
rect 20027 7936 20039 7939
rect 20073 7939 20131 7945
rect 20073 7936 20085 7939
rect 20027 7908 20085 7936
rect 20027 7905 20039 7908
rect 19981 7899 20039 7905
rect 20073 7905 20085 7908
rect 20119 7905 20131 7939
rect 23474 7936 23480 7948
rect 20073 7899 20131 7905
rect 21560 7908 23480 7936
rect 19794 7828 19800 7880
rect 19852 7868 19858 7880
rect 21560 7877 21588 7908
rect 23474 7896 23480 7908
rect 23532 7896 23538 7948
rect 23845 7939 23903 7945
rect 23845 7905 23857 7939
rect 23891 7936 23903 7939
rect 24946 7936 24952 7948
rect 23891 7908 24952 7936
rect 23891 7905 23903 7908
rect 23845 7899 23903 7905
rect 24946 7896 24952 7908
rect 25004 7896 25010 7948
rect 20901 7871 20959 7877
rect 20901 7868 20913 7871
rect 19852 7840 20913 7868
rect 19852 7828 19858 7840
rect 20901 7837 20913 7840
rect 20947 7837 20959 7871
rect 20901 7831 20959 7837
rect 21545 7871 21603 7877
rect 21545 7837 21557 7871
rect 21591 7837 21603 7871
rect 21545 7831 21603 7837
rect 22002 7828 22008 7880
rect 22060 7868 22066 7880
rect 22189 7871 22247 7877
rect 22189 7868 22201 7871
rect 22060 7840 22201 7868
rect 22060 7828 22066 7840
rect 22189 7837 22201 7840
rect 22235 7837 22247 7871
rect 22189 7831 22247 7837
rect 22833 7871 22891 7877
rect 22833 7837 22845 7871
rect 22879 7837 22891 7871
rect 22833 7831 22891 7837
rect 22848 7800 22876 7831
rect 23382 7828 23388 7880
rect 23440 7868 23446 7880
rect 24857 7871 24915 7877
rect 24857 7868 24869 7871
rect 23440 7840 24869 7868
rect 23440 7828 23446 7840
rect 24857 7837 24869 7840
rect 24903 7837 24915 7871
rect 24857 7831 24915 7837
rect 25590 7800 25596 7812
rect 22848 7772 25596 7800
rect 25590 7760 25596 7772
rect 25648 7760 25654 7812
rect 20714 7692 20720 7744
rect 20772 7692 20778 7744
rect 23474 7692 23480 7744
rect 23532 7732 23538 7744
rect 24673 7735 24731 7741
rect 24673 7732 24685 7735
rect 23532 7704 24685 7732
rect 23532 7692 23538 7704
rect 24673 7701 24685 7704
rect 24719 7701 24731 7735
rect 24673 7695 24731 7701
rect 1104 7642 25852 7664
rect 1104 7590 7950 7642
rect 8002 7590 8014 7642
rect 8066 7590 8078 7642
rect 8130 7590 8142 7642
rect 8194 7590 8206 7642
rect 8258 7590 17950 7642
rect 18002 7590 18014 7642
rect 18066 7590 18078 7642
rect 18130 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 25852 7642
rect 1104 7568 25852 7590
rect 21266 7488 21272 7540
rect 21324 7488 21330 7540
rect 20714 7420 20720 7472
rect 20772 7460 20778 7472
rect 23293 7463 23351 7469
rect 20772 7432 22416 7460
rect 20772 7420 20778 7432
rect 20346 7352 20352 7404
rect 20404 7392 20410 7404
rect 20809 7395 20867 7401
rect 20809 7392 20821 7395
rect 20404 7364 20821 7392
rect 20404 7352 20410 7364
rect 20809 7361 20821 7364
rect 20855 7361 20867 7395
rect 20809 7355 20867 7361
rect 21453 7395 21511 7401
rect 21453 7361 21465 7395
rect 21499 7392 21511 7395
rect 21818 7392 21824 7404
rect 21499 7364 21824 7392
rect 21499 7361 21511 7364
rect 21453 7355 21511 7361
rect 21818 7352 21824 7364
rect 21876 7352 21882 7404
rect 22281 7395 22339 7401
rect 22281 7361 22293 7395
rect 22327 7361 22339 7395
rect 22388 7392 22416 7432
rect 23293 7429 23305 7463
rect 23339 7460 23351 7463
rect 24854 7460 24860 7472
rect 23339 7432 24860 7460
rect 23339 7429 23351 7432
rect 23293 7423 23351 7429
rect 24854 7420 24860 7432
rect 24912 7420 24918 7472
rect 23937 7395 23995 7401
rect 23937 7392 23949 7395
rect 22388 7364 23949 7392
rect 22281 7355 22339 7361
rect 23937 7361 23949 7364
rect 23983 7361 23995 7395
rect 25038 7392 25044 7404
rect 23937 7355 23995 7361
rect 24044 7364 25044 7392
rect 22296 7324 22324 7355
rect 24044 7324 24072 7364
rect 25038 7352 25044 7364
rect 25096 7352 25102 7404
rect 22296 7296 24072 7324
rect 24670 7284 24676 7336
rect 24728 7284 24734 7336
rect 20625 7259 20683 7265
rect 20625 7225 20637 7259
rect 20671 7256 20683 7259
rect 20671 7228 22094 7256
rect 20671 7225 20683 7228
rect 20625 7219 20683 7225
rect 22066 7188 22094 7228
rect 23382 7188 23388 7200
rect 22066 7160 23388 7188
rect 23382 7148 23388 7160
rect 23440 7148 23446 7200
rect 1104 7098 25852 7120
rect 1104 7046 2950 7098
rect 3002 7046 3014 7098
rect 3066 7046 3078 7098
rect 3130 7046 3142 7098
rect 3194 7046 3206 7098
rect 3258 7046 12950 7098
rect 13002 7046 13014 7098
rect 13066 7046 13078 7098
rect 13130 7046 13142 7098
rect 13194 7046 13206 7098
rect 13258 7046 22950 7098
rect 23002 7046 23014 7098
rect 23066 7046 23078 7098
rect 23130 7046 23142 7098
rect 23194 7046 23206 7098
rect 23258 7046 25852 7098
rect 1104 7024 25852 7046
rect 20625 6919 20683 6925
rect 20625 6885 20637 6919
rect 20671 6885 20683 6919
rect 20625 6879 20683 6885
rect 20640 6848 20668 6879
rect 23845 6851 23903 6857
rect 20640 6820 22692 6848
rect 20806 6740 20812 6792
rect 20864 6740 20870 6792
rect 20990 6740 20996 6792
rect 21048 6780 21054 6792
rect 21453 6783 21511 6789
rect 21453 6780 21465 6783
rect 21048 6752 21465 6780
rect 21048 6740 21054 6752
rect 21453 6749 21465 6752
rect 21499 6749 21511 6783
rect 21453 6743 21511 6749
rect 21634 6740 21640 6792
rect 21692 6780 21698 6792
rect 21692 6752 22140 6780
rect 21692 6740 21698 6752
rect 15194 6672 15200 6724
rect 15252 6712 15258 6724
rect 22112 6712 22140 6752
rect 22186 6740 22192 6792
rect 22244 6740 22250 6792
rect 22664 6789 22692 6820
rect 23845 6817 23857 6851
rect 23891 6848 23903 6851
rect 24854 6848 24860 6860
rect 23891 6820 24860 6848
rect 23891 6817 23903 6820
rect 23845 6811 23903 6817
rect 24854 6808 24860 6820
rect 24912 6808 24918 6860
rect 22649 6783 22707 6789
rect 22649 6749 22661 6783
rect 22695 6749 22707 6783
rect 22649 6743 22707 6749
rect 24673 6715 24731 6721
rect 24673 6712 24685 6715
rect 15252 6684 22048 6712
rect 22112 6684 24685 6712
rect 15252 6672 15258 6684
rect 21269 6647 21327 6653
rect 21269 6613 21281 6647
rect 21315 6644 21327 6647
rect 21542 6644 21548 6656
rect 21315 6616 21548 6644
rect 21315 6613 21327 6616
rect 21269 6607 21327 6613
rect 21542 6604 21548 6616
rect 21600 6604 21606 6656
rect 22020 6653 22048 6684
rect 24673 6681 24685 6684
rect 24719 6681 24731 6715
rect 24673 6675 24731 6681
rect 24857 6715 24915 6721
rect 24857 6681 24869 6715
rect 24903 6712 24915 6715
rect 25038 6712 25044 6724
rect 24903 6684 25044 6712
rect 24903 6681 24915 6684
rect 24857 6675 24915 6681
rect 25038 6672 25044 6684
rect 25096 6672 25102 6724
rect 22005 6647 22063 6653
rect 22005 6613 22017 6647
rect 22051 6613 22063 6647
rect 22005 6607 22063 6613
rect 1104 6554 25852 6576
rect 1104 6502 7950 6554
rect 8002 6502 8014 6554
rect 8066 6502 8078 6554
rect 8130 6502 8142 6554
rect 8194 6502 8206 6554
rect 8258 6502 17950 6554
rect 18002 6502 18014 6554
rect 18066 6502 18078 6554
rect 18130 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 25852 6554
rect 1104 6480 25852 6502
rect 9306 6400 9312 6452
rect 9364 6400 9370 6452
rect 21637 6443 21695 6449
rect 21637 6409 21649 6443
rect 21683 6440 21695 6443
rect 21818 6440 21824 6452
rect 21683 6412 21824 6440
rect 21683 6409 21695 6412
rect 21637 6403 21695 6409
rect 21818 6400 21824 6412
rect 21876 6400 21882 6452
rect 23293 6375 23351 6381
rect 23293 6341 23305 6375
rect 23339 6372 23351 6375
rect 24854 6372 24860 6384
rect 23339 6344 24860 6372
rect 23339 6341 23351 6344
rect 23293 6335 23351 6341
rect 24854 6332 24860 6344
rect 24912 6332 24918 6384
rect 6822 6264 6828 6316
rect 6880 6304 6886 6316
rect 8665 6307 8723 6313
rect 8665 6304 8677 6307
rect 6880 6276 8677 6304
rect 6880 6264 6886 6276
rect 8665 6273 8677 6276
rect 8711 6273 8723 6307
rect 8665 6267 8723 6273
rect 22278 6264 22284 6316
rect 22336 6264 22342 6316
rect 23658 6264 23664 6316
rect 23716 6304 23722 6316
rect 23937 6307 23995 6313
rect 23937 6304 23949 6307
rect 23716 6276 23949 6304
rect 23716 6264 23722 6276
rect 23937 6273 23949 6276
rect 23983 6273 23995 6307
rect 23937 6267 23995 6273
rect 24762 6196 24768 6248
rect 24820 6196 24826 6248
rect 1104 6010 25852 6032
rect 1104 5958 2950 6010
rect 3002 5958 3014 6010
rect 3066 5958 3078 6010
rect 3130 5958 3142 6010
rect 3194 5958 3206 6010
rect 3258 5958 12950 6010
rect 13002 5958 13014 6010
rect 13066 5958 13078 6010
rect 13130 5958 13142 6010
rect 13194 5958 13206 6010
rect 13258 5958 22950 6010
rect 23002 5958 23014 6010
rect 23066 5958 23078 6010
rect 23130 5958 23142 6010
rect 23194 5958 23206 6010
rect 23258 5958 25852 6010
rect 1104 5936 25852 5958
rect 20530 5856 20536 5908
rect 20588 5896 20594 5908
rect 22005 5899 22063 5905
rect 22005 5896 22017 5899
rect 20588 5868 22017 5896
rect 20588 5856 20594 5868
rect 22005 5865 22017 5868
rect 22051 5865 22063 5899
rect 22005 5859 22063 5865
rect 21361 5831 21419 5837
rect 21361 5797 21373 5831
rect 21407 5828 21419 5831
rect 24578 5828 24584 5840
rect 21407 5800 24584 5828
rect 21407 5797 21419 5800
rect 21361 5791 21419 5797
rect 24578 5788 24584 5800
rect 24636 5788 24642 5840
rect 21545 5695 21603 5701
rect 21545 5661 21557 5695
rect 21591 5692 21603 5695
rect 21726 5692 21732 5704
rect 21591 5664 21732 5692
rect 21591 5661 21603 5664
rect 21545 5655 21603 5661
rect 21726 5652 21732 5664
rect 21784 5652 21790 5704
rect 22189 5695 22247 5701
rect 22189 5661 22201 5695
rect 22235 5692 22247 5695
rect 22370 5692 22376 5704
rect 22235 5664 22376 5692
rect 22235 5661 22247 5664
rect 22189 5655 22247 5661
rect 22370 5652 22376 5664
rect 22428 5652 22434 5704
rect 22833 5695 22891 5701
rect 22833 5661 22845 5695
rect 22879 5692 22891 5695
rect 23474 5692 23480 5704
rect 22879 5664 23480 5692
rect 22879 5661 22891 5664
rect 22833 5655 22891 5661
rect 23474 5652 23480 5664
rect 23532 5652 23538 5704
rect 24394 5652 24400 5704
rect 24452 5692 24458 5704
rect 24857 5695 24915 5701
rect 24857 5692 24869 5695
rect 24452 5664 24869 5692
rect 24452 5652 24458 5664
rect 24857 5661 24869 5664
rect 24903 5661 24915 5695
rect 24857 5655 24915 5661
rect 23845 5627 23903 5633
rect 23845 5593 23857 5627
rect 23891 5624 23903 5627
rect 24946 5624 24952 5636
rect 23891 5596 24952 5624
rect 23891 5593 23903 5596
rect 23845 5587 23903 5593
rect 24946 5584 24952 5596
rect 25004 5584 25010 5636
rect 23474 5516 23480 5568
rect 23532 5556 23538 5568
rect 24673 5559 24731 5565
rect 24673 5556 24685 5559
rect 23532 5528 24685 5556
rect 23532 5516 23538 5528
rect 24673 5525 24685 5528
rect 24719 5525 24731 5559
rect 24673 5519 24731 5525
rect 1104 5466 25852 5488
rect 1104 5414 7950 5466
rect 8002 5414 8014 5466
rect 8066 5414 8078 5466
rect 8130 5414 8142 5466
rect 8194 5414 8206 5466
rect 8258 5414 17950 5466
rect 18002 5414 18014 5466
rect 18066 5414 18078 5466
rect 18130 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 25852 5466
rect 1104 5392 25852 5414
rect 23293 5287 23351 5293
rect 23293 5253 23305 5287
rect 23339 5284 23351 5287
rect 24854 5284 24860 5296
rect 23339 5256 24860 5284
rect 23339 5253 23351 5256
rect 23293 5247 23351 5253
rect 24854 5244 24860 5256
rect 24912 5244 24918 5296
rect 22281 5219 22339 5225
rect 22281 5185 22293 5219
rect 22327 5216 22339 5219
rect 22462 5216 22468 5228
rect 22327 5188 22468 5216
rect 22327 5185 22339 5188
rect 22281 5179 22339 5185
rect 22462 5176 22468 5188
rect 22520 5176 22526 5228
rect 22738 5176 22744 5228
rect 22796 5216 22802 5228
rect 23937 5219 23995 5225
rect 23937 5216 23949 5219
rect 22796 5188 23949 5216
rect 22796 5176 22802 5188
rect 23937 5185 23949 5188
rect 23983 5185 23995 5219
rect 23937 5179 23995 5185
rect 24670 5108 24676 5160
rect 24728 5108 24734 5160
rect 1104 4922 25852 4944
rect 1104 4870 2950 4922
rect 3002 4870 3014 4922
rect 3066 4870 3078 4922
rect 3130 4870 3142 4922
rect 3194 4870 3206 4922
rect 3258 4870 12950 4922
rect 13002 4870 13014 4922
rect 13066 4870 13078 4922
rect 13130 4870 13142 4922
rect 13194 4870 13206 4922
rect 13258 4870 22950 4922
rect 23002 4870 23014 4922
rect 23066 4870 23078 4922
rect 23130 4870 23142 4922
rect 23194 4870 23206 4922
rect 23258 4870 25852 4922
rect 1104 4848 25852 4870
rect 22370 4768 22376 4820
rect 22428 4768 22434 4820
rect 22646 4564 22652 4616
rect 22704 4564 22710 4616
rect 23382 4564 23388 4616
rect 23440 4604 23446 4616
rect 24857 4607 24915 4613
rect 24857 4604 24869 4607
rect 23440 4576 24869 4604
rect 23440 4564 23446 4576
rect 24857 4573 24869 4576
rect 24903 4573 24915 4607
rect 24857 4567 24915 4573
rect 23845 4539 23903 4545
rect 23845 4505 23857 4539
rect 23891 4536 23903 4539
rect 24946 4536 24952 4548
rect 23891 4508 24952 4536
rect 23891 4505 23903 4508
rect 23845 4499 23903 4505
rect 24946 4496 24952 4508
rect 25004 4496 25010 4548
rect 23566 4428 23572 4480
rect 23624 4468 23630 4480
rect 24673 4471 24731 4477
rect 24673 4468 24685 4471
rect 23624 4440 24685 4468
rect 23624 4428 23630 4440
rect 24673 4437 24685 4440
rect 24719 4437 24731 4471
rect 24673 4431 24731 4437
rect 1104 4378 25852 4400
rect 1104 4326 7950 4378
rect 8002 4326 8014 4378
rect 8066 4326 8078 4378
rect 8130 4326 8142 4378
rect 8194 4326 8206 4378
rect 8258 4326 17950 4378
rect 18002 4326 18014 4378
rect 18066 4326 18078 4378
rect 18130 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 25852 4378
rect 1104 4304 25852 4326
rect 20254 4088 20260 4140
rect 20312 4088 20318 4140
rect 22281 4131 22339 4137
rect 22281 4097 22293 4131
rect 22327 4128 22339 4131
rect 24121 4131 24179 4137
rect 22327 4100 23244 4128
rect 22327 4097 22339 4100
rect 22281 4091 22339 4097
rect 18966 4020 18972 4072
rect 19024 4060 19030 4072
rect 20162 4060 20168 4072
rect 19024 4032 20168 4060
rect 19024 4020 19030 4032
rect 20162 4020 20168 4032
rect 20220 4020 20226 4072
rect 21269 4063 21327 4069
rect 21269 4029 21281 4063
rect 21315 4060 21327 4063
rect 22094 4060 22100 4072
rect 21315 4032 22100 4060
rect 21315 4029 21327 4032
rect 21269 4023 21327 4029
rect 22094 4020 22100 4032
rect 22152 4020 22158 4072
rect 23216 3924 23244 4100
rect 24121 4097 24133 4131
rect 24167 4128 24179 4131
rect 25130 4128 25136 4140
rect 24167 4100 25136 4128
rect 24167 4097 24179 4100
rect 24121 4091 24179 4097
rect 25130 4088 25136 4100
rect 25188 4088 25194 4140
rect 23293 4063 23351 4069
rect 23293 4029 23305 4063
rect 23339 4029 23351 4063
rect 23293 4023 23351 4029
rect 23308 3992 23336 4023
rect 24762 4020 24768 4072
rect 24820 4020 24826 4072
rect 24946 3992 24952 4004
rect 23308 3964 24952 3992
rect 24946 3952 24952 3964
rect 25004 3952 25010 4004
rect 25038 3924 25044 3936
rect 23216 3896 25044 3924
rect 25038 3884 25044 3896
rect 25096 3884 25102 3936
rect 1104 3834 25852 3856
rect 1104 3782 2950 3834
rect 3002 3782 3014 3834
rect 3066 3782 3078 3834
rect 3130 3782 3142 3834
rect 3194 3782 3206 3834
rect 3258 3782 12950 3834
rect 13002 3782 13014 3834
rect 13066 3782 13078 3834
rect 13130 3782 13142 3834
rect 13194 3782 13206 3834
rect 13258 3782 22950 3834
rect 23002 3782 23014 3834
rect 23066 3782 23078 3834
rect 23130 3782 23142 3834
rect 23194 3782 23206 3834
rect 23258 3782 25852 3834
rect 1104 3760 25852 3782
rect 20070 3476 20076 3528
rect 20128 3516 20134 3528
rect 20809 3519 20867 3525
rect 20809 3516 20821 3519
rect 20128 3488 20821 3516
rect 20128 3476 20134 3488
rect 20809 3485 20821 3488
rect 20855 3485 20867 3519
rect 20809 3479 20867 3485
rect 22833 3519 22891 3525
rect 22833 3485 22845 3519
rect 22879 3516 22891 3519
rect 23474 3516 23480 3528
rect 22879 3488 23480 3516
rect 22879 3485 22891 3488
rect 22833 3479 22891 3485
rect 23474 3476 23480 3488
rect 23532 3476 23538 3528
rect 24578 3476 24584 3528
rect 24636 3516 24642 3528
rect 24765 3519 24823 3525
rect 24765 3516 24777 3519
rect 24636 3488 24777 3516
rect 24636 3476 24642 3488
rect 24765 3485 24777 3488
rect 24811 3485 24823 3519
rect 24765 3479 24823 3485
rect 22002 3408 22008 3460
rect 22060 3408 22066 3460
rect 23845 3451 23903 3457
rect 23845 3417 23857 3451
rect 23891 3448 23903 3451
rect 24946 3448 24952 3460
rect 23891 3420 24952 3448
rect 23891 3417 23903 3420
rect 23845 3411 23903 3417
rect 24946 3408 24952 3420
rect 25004 3408 25010 3460
rect 24578 3340 24584 3392
rect 24636 3340 24642 3392
rect 1104 3290 25852 3312
rect 1104 3238 7950 3290
rect 8002 3238 8014 3290
rect 8066 3238 8078 3290
rect 8130 3238 8142 3290
rect 8194 3238 8206 3290
rect 8258 3238 17950 3290
rect 18002 3238 18014 3290
rect 18066 3238 18078 3290
rect 18130 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 25852 3290
rect 1104 3216 25852 3238
rect 6822 3136 6828 3188
rect 6880 3136 6886 3188
rect 23293 3111 23351 3117
rect 23293 3077 23305 3111
rect 23339 3108 23351 3111
rect 24854 3108 24860 3120
rect 23339 3080 24860 3108
rect 23339 3077 23351 3080
rect 23293 3071 23351 3077
rect 24854 3068 24860 3080
rect 24912 3068 24918 3120
rect 25130 3068 25136 3120
rect 25188 3068 25194 3120
rect 7006 3000 7012 3052
rect 7064 3000 7070 3052
rect 18417 3043 18475 3049
rect 18417 3009 18429 3043
rect 18463 3040 18475 3043
rect 19794 3040 19800 3052
rect 18463 3012 19800 3040
rect 18463 3009 18475 3012
rect 18417 3003 18475 3009
rect 19794 3000 19800 3012
rect 19852 3000 19858 3052
rect 19978 3000 19984 3052
rect 20036 3040 20042 3052
rect 20073 3043 20131 3049
rect 20073 3040 20085 3043
rect 20036 3012 20085 3040
rect 20036 3000 20042 3012
rect 20073 3009 20085 3012
rect 20119 3009 20131 3043
rect 20073 3003 20131 3009
rect 22281 3043 22339 3049
rect 22281 3009 22293 3043
rect 22327 3040 22339 3043
rect 23566 3040 23572 3052
rect 22327 3012 23572 3040
rect 22327 3009 22339 3012
rect 22281 3003 22339 3009
rect 23566 3000 23572 3012
rect 23624 3000 23630 3052
rect 24121 3043 24179 3049
rect 24121 3009 24133 3043
rect 24167 3040 24179 3043
rect 24210 3040 24216 3052
rect 24167 3012 24216 3040
rect 24167 3009 24179 3012
rect 24121 3003 24179 3009
rect 24210 3000 24216 3012
rect 24268 3000 24274 3052
rect 19334 2932 19340 2984
rect 19392 2932 19398 2984
rect 21269 2975 21327 2981
rect 21269 2941 21281 2975
rect 21315 2972 21327 2975
rect 25038 2972 25044 2984
rect 21315 2944 25044 2972
rect 21315 2941 21327 2944
rect 21269 2935 21327 2941
rect 25038 2932 25044 2944
rect 25096 2932 25102 2984
rect 19794 2796 19800 2848
rect 19852 2836 19858 2848
rect 25866 2836 25872 2848
rect 19852 2808 25872 2836
rect 19852 2796 19858 2808
rect 25866 2796 25872 2808
rect 25924 2796 25930 2848
rect 1104 2746 25852 2768
rect 1104 2694 2950 2746
rect 3002 2694 3014 2746
rect 3066 2694 3078 2746
rect 3130 2694 3142 2746
rect 3194 2694 3206 2746
rect 3258 2694 12950 2746
rect 13002 2694 13014 2746
rect 13066 2694 13078 2746
rect 13130 2694 13142 2746
rect 13194 2694 13206 2746
rect 13258 2694 22950 2746
rect 23002 2694 23014 2746
rect 23066 2694 23078 2746
rect 23130 2694 23142 2746
rect 23194 2694 23206 2746
rect 23258 2694 25852 2746
rect 1104 2672 25852 2694
rect 7006 2592 7012 2644
rect 7064 2632 7070 2644
rect 7469 2635 7527 2641
rect 7469 2632 7481 2635
rect 7064 2604 7481 2632
rect 7064 2592 7070 2604
rect 7469 2601 7481 2604
rect 7515 2601 7527 2635
rect 7469 2595 7527 2601
rect 19334 2592 19340 2644
rect 19392 2632 19398 2644
rect 22186 2632 22192 2644
rect 19392 2604 22192 2632
rect 19392 2592 19398 2604
rect 22186 2592 22192 2604
rect 22244 2592 22250 2644
rect 19794 2524 19800 2576
rect 19852 2524 19858 2576
rect 6825 2431 6883 2437
rect 6825 2428 6837 2431
rect 6748 2400 6837 2428
rect 6748 2304 6776 2400
rect 6825 2397 6837 2400
rect 6871 2397 6883 2431
rect 6825 2391 6883 2397
rect 20257 2431 20315 2437
rect 20257 2397 20269 2431
rect 20303 2428 20315 2431
rect 20622 2428 20628 2440
rect 20303 2400 20628 2428
rect 20303 2397 20315 2400
rect 20257 2391 20315 2397
rect 20622 2388 20628 2400
rect 20680 2388 20686 2440
rect 22833 2431 22891 2437
rect 22833 2397 22845 2431
rect 22879 2428 22891 2431
rect 24578 2428 24584 2440
rect 22879 2400 24584 2428
rect 22879 2397 22891 2400
rect 22833 2391 22891 2397
rect 24578 2388 24584 2400
rect 24636 2388 24642 2440
rect 21269 2363 21327 2369
rect 21269 2329 21281 2363
rect 21315 2360 21327 2363
rect 23382 2360 23388 2372
rect 21315 2332 23388 2360
rect 21315 2329 21327 2332
rect 21269 2323 21327 2329
rect 23382 2320 23388 2332
rect 23440 2320 23446 2372
rect 23845 2363 23903 2369
rect 23845 2329 23857 2363
rect 23891 2360 23903 2363
rect 24946 2360 24952 2372
rect 23891 2332 24952 2360
rect 23891 2329 23903 2332
rect 23845 2323 23903 2329
rect 24946 2320 24952 2332
rect 25004 2320 25010 2372
rect 6549 2295 6607 2301
rect 6549 2261 6561 2295
rect 6595 2292 6607 2295
rect 6730 2292 6736 2304
rect 6595 2264 6736 2292
rect 6595 2261 6607 2264
rect 6549 2255 6607 2261
rect 6730 2252 6736 2264
rect 6788 2252 6794 2304
rect 1104 2202 25852 2224
rect 1104 2150 7950 2202
rect 8002 2150 8014 2202
rect 8066 2150 8078 2202
rect 8130 2150 8142 2202
rect 8194 2150 8206 2202
rect 8258 2150 17950 2202
rect 18002 2150 18014 2202
rect 18066 2150 18078 2202
rect 18130 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 25852 2202
rect 1104 2128 25852 2150
<< via1 >>
rect 3056 26392 3108 26444
rect 3332 26392 3384 26444
rect 2136 26324 2188 26376
rect 22192 26324 22244 26376
rect 9588 26256 9640 26308
rect 21824 26256 21876 26308
rect 7564 25236 7616 25288
rect 26148 25236 26200 25288
rect 3608 25168 3660 25220
rect 25596 25168 25648 25220
rect 5172 25100 5224 25152
rect 15844 25100 15896 25152
rect 1952 25032 2004 25084
rect 14004 25032 14056 25084
rect 6644 24964 6696 25016
rect 9864 24896 9916 24948
rect 17316 24896 17368 24948
rect 8484 24828 8536 24880
rect 18144 24828 18196 24880
rect 20628 24828 20680 24880
rect 23204 24828 23256 24880
rect 5816 24760 5868 24812
rect 8392 24760 8444 24812
rect 9772 24760 9824 24812
rect 16028 24760 16080 24812
rect 25136 24760 25188 24812
rect 6000 24692 6052 24744
rect 14096 24692 14148 24744
rect 7748 24624 7800 24676
rect 5264 24556 5316 24608
rect 8576 24556 8628 24608
rect 16856 24624 16908 24676
rect 20628 24624 20680 24676
rect 19708 24556 19760 24608
rect 2950 24454 3002 24506
rect 3014 24454 3066 24506
rect 3078 24454 3130 24506
rect 3142 24454 3194 24506
rect 3206 24454 3258 24506
rect 12950 24454 13002 24506
rect 13014 24454 13066 24506
rect 13078 24454 13130 24506
rect 13142 24454 13194 24506
rect 13206 24454 13258 24506
rect 22950 24454 23002 24506
rect 23014 24454 23066 24506
rect 23078 24454 23130 24506
rect 23142 24454 23194 24506
rect 23206 24454 23258 24506
rect 14004 24352 14056 24404
rect 6368 24284 6420 24336
rect 6552 24327 6604 24336
rect 6552 24293 6561 24327
rect 6561 24293 6595 24327
rect 6595 24293 6604 24327
rect 6552 24284 6604 24293
rect 6460 24216 6512 24268
rect 8484 24284 8536 24336
rect 8852 24284 8904 24336
rect 12348 24284 12400 24336
rect 1768 24191 1820 24200
rect 1768 24157 1777 24191
rect 1777 24157 1811 24191
rect 1811 24157 1820 24191
rect 1768 24148 1820 24157
rect 3884 24148 3936 24200
rect 4804 24191 4856 24200
rect 4804 24157 4813 24191
rect 4813 24157 4847 24191
rect 4847 24157 4856 24191
rect 4804 24148 4856 24157
rect 9680 24216 9732 24268
rect 10968 24259 11020 24268
rect 10968 24225 10977 24259
rect 10977 24225 11011 24259
rect 11011 24225 11020 24259
rect 10968 24216 11020 24225
rect 11796 24216 11848 24268
rect 6736 24191 6788 24200
rect 6736 24157 6745 24191
rect 6745 24157 6779 24191
rect 6779 24157 6788 24191
rect 6736 24148 6788 24157
rect 5816 24123 5868 24132
rect 5816 24089 5825 24123
rect 5825 24089 5859 24123
rect 5859 24089 5868 24123
rect 5816 24080 5868 24089
rect 3976 24012 4028 24064
rect 9312 24191 9364 24200
rect 9312 24157 9321 24191
rect 9321 24157 9355 24191
rect 9355 24157 9364 24191
rect 9312 24148 9364 24157
rect 18144 24395 18196 24404
rect 18144 24361 18153 24395
rect 18153 24361 18187 24395
rect 18187 24361 18196 24395
rect 18144 24352 18196 24361
rect 16396 24284 16448 24336
rect 18788 24352 18840 24404
rect 19984 24352 20036 24404
rect 20076 24352 20128 24404
rect 22376 24352 22428 24404
rect 16120 24259 16172 24268
rect 16120 24225 16129 24259
rect 16129 24225 16163 24259
rect 16163 24225 16172 24259
rect 16120 24216 16172 24225
rect 15660 24148 15712 24200
rect 16948 24148 17000 24200
rect 17776 24216 17828 24268
rect 18696 24216 18748 24268
rect 18788 24259 18840 24268
rect 18788 24225 18797 24259
rect 18797 24225 18831 24259
rect 18831 24225 18840 24259
rect 18788 24216 18840 24225
rect 19984 24216 20036 24268
rect 22560 24216 22612 24268
rect 25044 24259 25096 24268
rect 25044 24225 25053 24259
rect 25053 24225 25087 24259
rect 25087 24225 25096 24259
rect 25044 24216 25096 24225
rect 20076 24148 20128 24200
rect 7472 24012 7524 24064
rect 14648 24080 14700 24132
rect 22284 24191 22336 24200
rect 22284 24157 22293 24191
rect 22293 24157 22327 24191
rect 22327 24157 22336 24191
rect 22284 24148 22336 24157
rect 23848 24148 23900 24200
rect 20260 24080 20312 24132
rect 9128 24055 9180 24064
rect 9128 24021 9137 24055
rect 9137 24021 9171 24055
rect 9171 24021 9180 24055
rect 9128 24012 9180 24021
rect 11336 24012 11388 24064
rect 16856 24012 16908 24064
rect 17040 24012 17092 24064
rect 17776 24012 17828 24064
rect 17960 24055 18012 24064
rect 17960 24021 17969 24055
rect 17969 24021 18003 24055
rect 18003 24021 18012 24055
rect 17960 24012 18012 24021
rect 19248 24012 19300 24064
rect 19340 24012 19392 24064
rect 20996 24012 21048 24064
rect 21364 24012 21416 24064
rect 21824 24012 21876 24064
rect 23572 24012 23624 24064
rect 23940 24012 23992 24064
rect 24124 24012 24176 24064
rect 25044 24080 25096 24132
rect 7950 23910 8002 23962
rect 8014 23910 8066 23962
rect 8078 23910 8130 23962
rect 8142 23910 8194 23962
rect 8206 23910 8258 23962
rect 17950 23910 18002 23962
rect 18014 23910 18066 23962
rect 18078 23910 18130 23962
rect 18142 23910 18194 23962
rect 18206 23910 18258 23962
rect 4896 23808 4948 23860
rect 5356 23740 5408 23792
rect 7380 23740 7432 23792
rect 1124 23672 1176 23724
rect 1492 23672 1544 23724
rect 3792 23672 3844 23724
rect 9312 23808 9364 23860
rect 11520 23851 11572 23860
rect 11520 23817 11529 23851
rect 11529 23817 11563 23851
rect 11563 23817 11572 23851
rect 11520 23808 11572 23817
rect 10140 23740 10192 23792
rect 10876 23783 10928 23792
rect 10876 23749 10885 23783
rect 10885 23749 10919 23783
rect 10919 23749 10928 23783
rect 10876 23740 10928 23749
rect 14004 23808 14056 23860
rect 14096 23851 14148 23860
rect 14096 23817 14105 23851
rect 14105 23817 14139 23851
rect 14139 23817 14148 23851
rect 14096 23808 14148 23817
rect 15568 23808 15620 23860
rect 15752 23808 15804 23860
rect 16580 23808 16632 23860
rect 19340 23808 19392 23860
rect 20076 23808 20128 23860
rect 22284 23808 22336 23860
rect 23296 23808 23348 23860
rect 6460 23536 6512 23588
rect 7564 23604 7616 23656
rect 8576 23672 8628 23724
rect 9956 23672 10008 23724
rect 11888 23740 11940 23792
rect 18420 23740 18472 23792
rect 18972 23740 19024 23792
rect 19616 23740 19668 23792
rect 22100 23740 22152 23792
rect 11060 23604 11112 23656
rect 7380 23536 7432 23588
rect 7104 23468 7156 23520
rect 9496 23468 9548 23520
rect 15200 23672 15252 23724
rect 11980 23604 12032 23656
rect 14740 23647 14792 23656
rect 14740 23613 14749 23647
rect 14749 23613 14783 23647
rect 14783 23613 14792 23647
rect 14740 23604 14792 23613
rect 15476 23604 15528 23656
rect 15752 23604 15804 23656
rect 11520 23536 11572 23588
rect 14556 23536 14608 23588
rect 15660 23536 15712 23588
rect 15844 23536 15896 23588
rect 17776 23672 17828 23724
rect 24032 23740 24084 23792
rect 25136 23783 25188 23792
rect 25136 23749 25145 23783
rect 25145 23749 25179 23783
rect 25179 23749 25188 23783
rect 25136 23740 25188 23749
rect 16304 23604 16356 23656
rect 17316 23647 17368 23656
rect 17316 23613 17325 23647
rect 17325 23613 17359 23647
rect 17359 23613 17368 23647
rect 17316 23604 17368 23613
rect 11704 23468 11756 23520
rect 14924 23468 14976 23520
rect 16764 23468 16816 23520
rect 16856 23511 16908 23520
rect 16856 23477 16865 23511
rect 16865 23477 16899 23511
rect 16899 23477 16908 23511
rect 16856 23468 16908 23477
rect 18052 23647 18104 23656
rect 18052 23613 18061 23647
rect 18061 23613 18095 23647
rect 18095 23613 18104 23647
rect 18052 23604 18104 23613
rect 17960 23536 18012 23588
rect 18420 23604 18472 23656
rect 19340 23604 19392 23656
rect 20628 23647 20680 23656
rect 20628 23613 20637 23647
rect 20637 23613 20671 23647
rect 20671 23613 20680 23647
rect 20628 23604 20680 23613
rect 22560 23647 22612 23656
rect 22560 23613 22569 23647
rect 22569 23613 22603 23647
rect 22603 23613 22612 23647
rect 22560 23604 22612 23613
rect 24308 23604 24360 23656
rect 19800 23511 19852 23520
rect 19800 23477 19809 23511
rect 19809 23477 19843 23511
rect 19843 23477 19852 23511
rect 19800 23468 19852 23477
rect 19892 23468 19944 23520
rect 20444 23468 20496 23520
rect 23572 23536 23624 23588
rect 25412 23536 25464 23588
rect 24124 23468 24176 23520
rect 25136 23468 25188 23520
rect 2950 23366 3002 23418
rect 3014 23366 3066 23418
rect 3078 23366 3130 23418
rect 3142 23366 3194 23418
rect 3206 23366 3258 23418
rect 12950 23366 13002 23418
rect 13014 23366 13066 23418
rect 13078 23366 13130 23418
rect 13142 23366 13194 23418
rect 13206 23366 13258 23418
rect 22950 23366 23002 23418
rect 23014 23366 23066 23418
rect 23078 23366 23130 23418
rect 23142 23366 23194 23418
rect 23206 23366 23258 23418
rect 1492 23307 1544 23316
rect 1492 23273 1501 23307
rect 1501 23273 1535 23307
rect 1535 23273 1544 23307
rect 1492 23264 1544 23273
rect 6736 23264 6788 23316
rect 7380 23264 7432 23316
rect 11980 23264 12032 23316
rect 12348 23264 12400 23316
rect 12440 23264 12492 23316
rect 12900 23264 12952 23316
rect 13820 23264 13872 23316
rect 13912 23264 13964 23316
rect 16488 23264 16540 23316
rect 16580 23264 16632 23316
rect 17684 23264 17736 23316
rect 17960 23264 18012 23316
rect 18788 23264 18840 23316
rect 22560 23264 22612 23316
rect 4620 23128 4672 23180
rect 7656 23128 7708 23180
rect 9404 23196 9456 23248
rect 8576 23128 8628 23180
rect 11704 23196 11756 23248
rect 13544 23239 13596 23248
rect 13544 23205 13553 23239
rect 13553 23205 13587 23239
rect 13587 23205 13596 23239
rect 13544 23196 13596 23205
rect 17132 23196 17184 23248
rect 18880 23196 18932 23248
rect 18972 23196 19024 23248
rect 19432 23196 19484 23248
rect 10508 23171 10560 23180
rect 10508 23137 10517 23171
rect 10517 23137 10551 23171
rect 10551 23137 10560 23171
rect 10508 23128 10560 23137
rect 11612 23128 11664 23180
rect 2228 23103 2280 23112
rect 2228 23069 2237 23103
rect 2237 23069 2271 23103
rect 2271 23069 2280 23103
rect 2228 23060 2280 23069
rect 3424 23060 3476 23112
rect 5448 23103 5500 23112
rect 5448 23069 5457 23103
rect 5457 23069 5491 23103
rect 5491 23069 5500 23103
rect 5448 23060 5500 23069
rect 7012 23060 7064 23112
rect 5632 22992 5684 23044
rect 6368 22992 6420 23044
rect 7564 22992 7616 23044
rect 4712 22967 4764 22976
rect 4712 22933 4721 22967
rect 4721 22933 4755 22967
rect 4755 22933 4764 22967
rect 4712 22924 4764 22933
rect 11980 22992 12032 23044
rect 14188 23128 14240 23180
rect 18604 23128 18656 23180
rect 19064 23128 19116 23180
rect 20720 23128 20772 23180
rect 22284 23128 22336 23180
rect 24768 23128 24820 23180
rect 12716 23060 12768 23112
rect 13636 23060 13688 23112
rect 13728 23103 13780 23112
rect 13728 23069 13737 23103
rect 13737 23069 13771 23103
rect 13771 23069 13780 23103
rect 13728 23060 13780 23069
rect 13820 23060 13872 23112
rect 16764 23060 16816 23112
rect 18052 23060 18104 23112
rect 19340 23060 19392 23112
rect 12992 22992 13044 23044
rect 14556 22992 14608 23044
rect 15568 22992 15620 23044
rect 11888 22924 11940 22976
rect 15016 22924 15068 22976
rect 18512 23035 18564 23044
rect 18512 23001 18519 23035
rect 18519 23001 18564 23035
rect 18512 22992 18564 23001
rect 18696 22992 18748 23044
rect 18972 22992 19024 23044
rect 19156 22992 19208 23044
rect 16764 22924 16816 22976
rect 17316 22924 17368 22976
rect 18052 22924 18104 22976
rect 19064 22967 19116 22976
rect 19064 22933 19073 22967
rect 19073 22933 19107 22967
rect 19107 22933 19116 22967
rect 19064 22924 19116 22933
rect 19984 22992 20036 23044
rect 22192 22992 22244 23044
rect 22376 22992 22428 23044
rect 23940 22924 23992 22976
rect 24584 22967 24636 22976
rect 24584 22933 24593 22967
rect 24593 22933 24627 22967
rect 24627 22933 24636 22967
rect 24584 22924 24636 22933
rect 24952 22967 25004 22976
rect 24952 22933 24961 22967
rect 24961 22933 24995 22967
rect 24995 22933 25004 22967
rect 24952 22924 25004 22933
rect 7950 22822 8002 22874
rect 8014 22822 8066 22874
rect 8078 22822 8130 22874
rect 8142 22822 8194 22874
rect 8206 22822 8258 22874
rect 17950 22822 18002 22874
rect 18014 22822 18066 22874
rect 18078 22822 18130 22874
rect 18142 22822 18194 22874
rect 18206 22822 18258 22874
rect 2228 22720 2280 22772
rect 3424 22652 3476 22704
rect 4252 22652 4304 22704
rect 4712 22720 4764 22772
rect 1216 22584 1268 22636
rect 1676 22627 1728 22636
rect 1676 22593 1685 22627
rect 1685 22593 1719 22627
rect 1719 22593 1728 22627
rect 1676 22584 1728 22593
rect 3240 22516 3292 22568
rect 3424 22516 3476 22568
rect 3700 22516 3752 22568
rect 5724 22695 5776 22704
rect 5724 22661 5733 22695
rect 5733 22661 5767 22695
rect 5767 22661 5776 22695
rect 5724 22652 5776 22661
rect 7380 22652 7432 22704
rect 8760 22695 8812 22704
rect 8760 22661 8769 22695
rect 8769 22661 8803 22695
rect 8803 22661 8812 22695
rect 8760 22652 8812 22661
rect 5816 22584 5868 22636
rect 6736 22584 6788 22636
rect 6184 22516 6236 22568
rect 9680 22652 9732 22704
rect 9772 22652 9824 22704
rect 9956 22652 10008 22704
rect 11060 22652 11112 22704
rect 9036 22516 9088 22568
rect 12716 22584 12768 22636
rect 13820 22652 13872 22704
rect 14004 22652 14056 22704
rect 14556 22720 14608 22772
rect 14740 22720 14792 22772
rect 15568 22720 15620 22772
rect 16856 22720 16908 22772
rect 16580 22652 16632 22704
rect 1768 22423 1820 22432
rect 1768 22389 1777 22423
rect 1777 22389 1811 22423
rect 1811 22389 1820 22423
rect 1768 22380 1820 22389
rect 3792 22380 3844 22432
rect 5540 22380 5592 22432
rect 9404 22380 9456 22432
rect 12072 22448 12124 22500
rect 12440 22448 12492 22500
rect 12624 22448 12676 22500
rect 12992 22448 13044 22500
rect 11152 22423 11204 22432
rect 11152 22389 11161 22423
rect 11161 22389 11195 22423
rect 11195 22389 11204 22423
rect 11152 22380 11204 22389
rect 11244 22380 11296 22432
rect 12532 22380 12584 22432
rect 12900 22380 12952 22432
rect 15936 22627 15988 22636
rect 15936 22593 15945 22627
rect 15945 22593 15979 22627
rect 15979 22593 15988 22627
rect 15936 22584 15988 22593
rect 17132 22652 17184 22704
rect 18604 22763 18656 22772
rect 18604 22729 18613 22763
rect 18613 22729 18647 22763
rect 18647 22729 18656 22763
rect 18604 22720 18656 22729
rect 20904 22720 20956 22772
rect 23848 22720 23900 22772
rect 15660 22516 15712 22568
rect 16304 22516 16356 22568
rect 19800 22652 19852 22704
rect 15292 22448 15344 22500
rect 15844 22380 15896 22432
rect 16028 22423 16080 22432
rect 16028 22389 16037 22423
rect 16037 22389 16071 22423
rect 16071 22389 16080 22423
rect 16028 22380 16080 22389
rect 16304 22380 16356 22432
rect 16488 22380 16540 22432
rect 19432 22584 19484 22636
rect 19892 22584 19944 22636
rect 20260 22627 20312 22636
rect 20260 22593 20269 22627
rect 20269 22593 20303 22627
rect 20303 22593 20312 22627
rect 20260 22584 20312 22593
rect 22284 22652 22336 22704
rect 24032 22652 24084 22704
rect 20812 22516 20864 22568
rect 22376 22584 22428 22636
rect 22560 22516 22612 22568
rect 23296 22559 23348 22568
rect 23296 22525 23305 22559
rect 23305 22525 23339 22559
rect 23339 22525 23348 22559
rect 23296 22516 23348 22525
rect 24124 22516 24176 22568
rect 25872 22516 25924 22568
rect 19432 22448 19484 22500
rect 20260 22380 20312 22432
rect 21088 22380 21140 22432
rect 23664 22380 23716 22432
rect 24768 22380 24820 22432
rect 25504 22380 25556 22432
rect 2950 22278 3002 22330
rect 3014 22278 3066 22330
rect 3078 22278 3130 22330
rect 3142 22278 3194 22330
rect 3206 22278 3258 22330
rect 12950 22278 13002 22330
rect 13014 22278 13066 22330
rect 13078 22278 13130 22330
rect 13142 22278 13194 22330
rect 13206 22278 13258 22330
rect 22950 22278 23002 22330
rect 23014 22278 23066 22330
rect 23078 22278 23130 22330
rect 23142 22278 23194 22330
rect 23206 22278 23258 22330
rect 1676 22219 1728 22228
rect 1676 22185 1685 22219
rect 1685 22185 1719 22219
rect 1719 22185 1728 22219
rect 1676 22176 1728 22185
rect 1768 22108 1820 22160
rect 10600 22176 10652 22228
rect 12808 22176 12860 22228
rect 14740 22176 14792 22228
rect 3608 22108 3660 22160
rect 3792 22108 3844 22160
rect 2872 22083 2924 22092
rect 2872 22049 2881 22083
rect 2881 22049 2915 22083
rect 2915 22049 2924 22083
rect 2872 22040 2924 22049
rect 6092 22083 6144 22092
rect 6092 22049 6101 22083
rect 6101 22049 6135 22083
rect 6135 22049 6144 22083
rect 6092 22040 6144 22049
rect 8300 22083 8352 22092
rect 8300 22049 8309 22083
rect 8309 22049 8343 22083
rect 8343 22049 8352 22083
rect 8300 22040 8352 22049
rect 4528 21972 4580 22024
rect 5448 22015 5500 22024
rect 5448 21981 5457 22015
rect 5457 21981 5491 22015
rect 5491 21981 5500 22015
rect 5448 21972 5500 21981
rect 7840 21972 7892 22024
rect 8300 21904 8352 21956
rect 9404 22108 9456 22160
rect 12256 22108 12308 22160
rect 13452 22108 13504 22160
rect 9036 22040 9088 22092
rect 11060 22040 11112 22092
rect 11704 22040 11756 22092
rect 12440 22083 12492 22092
rect 12440 22049 12449 22083
rect 12449 22049 12483 22083
rect 12483 22049 12492 22083
rect 12440 22040 12492 22049
rect 13176 22040 13228 22092
rect 13820 22040 13872 22092
rect 15844 22108 15896 22160
rect 17132 22176 17184 22228
rect 18972 22176 19024 22228
rect 19064 22176 19116 22228
rect 21824 22176 21876 22228
rect 22284 22176 22336 22228
rect 25780 22176 25832 22228
rect 17684 22108 17736 22160
rect 20260 22108 20312 22160
rect 21640 22108 21692 22160
rect 22744 22108 22796 22160
rect 17224 22040 17276 22092
rect 18144 22083 18196 22092
rect 18144 22049 18153 22083
rect 18153 22049 18187 22083
rect 18187 22049 18196 22083
rect 18144 22040 18196 22049
rect 4988 21836 5040 21888
rect 9312 21879 9364 21888
rect 9312 21845 9321 21879
rect 9321 21845 9355 21879
rect 9355 21845 9364 21879
rect 9312 21836 9364 21845
rect 10048 21879 10100 21888
rect 10048 21845 10057 21879
rect 10057 21845 10091 21879
rect 10091 21845 10100 21879
rect 10048 21836 10100 21845
rect 13360 21972 13412 22024
rect 11704 21904 11756 21956
rect 12440 21904 12492 21956
rect 14188 21972 14240 22024
rect 13544 21947 13596 21956
rect 13544 21913 13553 21947
rect 13553 21913 13587 21947
rect 13587 21913 13596 21947
rect 13544 21904 13596 21913
rect 14004 21904 14056 21956
rect 12256 21836 12308 21888
rect 12900 21879 12952 21888
rect 12900 21845 12909 21879
rect 12909 21845 12943 21879
rect 12943 21845 12952 21879
rect 12900 21836 12952 21845
rect 13176 21836 13228 21888
rect 15292 21836 15344 21888
rect 17316 21904 17368 21956
rect 17500 21904 17552 21956
rect 20168 22040 20220 22092
rect 16764 21836 16816 21888
rect 17132 21836 17184 21888
rect 17684 21879 17736 21888
rect 17684 21845 17693 21879
rect 17693 21845 17727 21879
rect 17727 21845 17736 21879
rect 17684 21836 17736 21845
rect 17776 21836 17828 21888
rect 18144 21836 18196 21888
rect 19064 21972 19116 22024
rect 19340 21972 19392 22024
rect 22192 22040 22244 22092
rect 22836 21972 22888 22024
rect 23204 22015 23256 22024
rect 23204 21981 23213 22015
rect 23213 21981 23247 22015
rect 23247 21981 23256 22015
rect 23204 21972 23256 21981
rect 23480 22015 23532 22024
rect 23480 21981 23489 22015
rect 23489 21981 23523 22015
rect 23523 21981 23532 22015
rect 23480 21972 23532 21981
rect 24860 22040 24912 22092
rect 25136 22040 25188 22092
rect 25320 22108 25372 22160
rect 25964 21972 26016 22024
rect 19524 21947 19576 21956
rect 19524 21913 19533 21947
rect 19533 21913 19567 21947
rect 19567 21913 19576 21947
rect 19524 21904 19576 21913
rect 20904 21904 20956 21956
rect 18696 21879 18748 21888
rect 18696 21845 18705 21879
rect 18705 21845 18739 21879
rect 18739 21845 18748 21879
rect 18696 21836 18748 21845
rect 19616 21879 19668 21888
rect 19616 21845 19625 21879
rect 19625 21845 19659 21879
rect 19659 21845 19668 21879
rect 19616 21836 19668 21845
rect 20812 21836 20864 21888
rect 23848 21904 23900 21956
rect 24032 21904 24084 21956
rect 21272 21836 21324 21888
rect 21456 21836 21508 21888
rect 22192 21836 22244 21888
rect 22284 21836 22336 21888
rect 23572 21836 23624 21888
rect 23756 21836 23808 21888
rect 26240 21836 26292 21888
rect 7950 21734 8002 21786
rect 8014 21734 8066 21786
rect 8078 21734 8130 21786
rect 8142 21734 8194 21786
rect 8206 21734 8258 21786
rect 17950 21734 18002 21786
rect 18014 21734 18066 21786
rect 18078 21734 18130 21786
rect 18142 21734 18194 21786
rect 18206 21734 18258 21786
rect 3424 21632 3476 21684
rect 6460 21632 6512 21684
rect 8208 21632 8260 21684
rect 8484 21632 8536 21684
rect 10048 21632 10100 21684
rect 13452 21675 13504 21684
rect 13452 21641 13461 21675
rect 13461 21641 13495 21675
rect 13495 21641 13504 21675
rect 13452 21632 13504 21641
rect 5540 21564 5592 21616
rect 4804 21539 4856 21548
rect 4804 21505 4813 21539
rect 4813 21505 4847 21539
rect 4847 21505 4856 21539
rect 4804 21496 4856 21505
rect 9404 21564 9456 21616
rect 9772 21564 9824 21616
rect 16212 21632 16264 21684
rect 20168 21632 20220 21684
rect 20444 21675 20496 21684
rect 20444 21641 20453 21675
rect 20453 21641 20487 21675
rect 20487 21641 20496 21675
rect 20444 21632 20496 21641
rect 17684 21564 17736 21616
rect 18512 21564 18564 21616
rect 21548 21632 21600 21684
rect 22100 21632 22152 21684
rect 24676 21632 24728 21684
rect 23664 21607 23716 21616
rect 23664 21573 23673 21607
rect 23673 21573 23707 21607
rect 23707 21573 23716 21607
rect 23664 21564 23716 21573
rect 24124 21564 24176 21616
rect 7380 21539 7432 21548
rect 7380 21505 7389 21539
rect 7389 21505 7423 21539
rect 7423 21505 7432 21539
rect 7380 21496 7432 21505
rect 9036 21539 9088 21548
rect 9036 21505 9045 21539
rect 9045 21505 9079 21539
rect 9079 21505 9088 21539
rect 9036 21496 9088 21505
rect 11152 21496 11204 21548
rect 13268 21496 13320 21548
rect 14096 21496 14148 21548
rect 14188 21539 14240 21548
rect 14188 21505 14197 21539
rect 14197 21505 14231 21539
rect 14231 21505 14240 21539
rect 14188 21496 14240 21505
rect 14832 21496 14884 21548
rect 15568 21496 15620 21548
rect 16212 21539 16264 21548
rect 16212 21505 16221 21539
rect 16221 21505 16255 21539
rect 16255 21505 16264 21539
rect 16212 21496 16264 21505
rect 16304 21496 16356 21548
rect 16856 21496 16908 21548
rect 17224 21496 17276 21548
rect 17408 21539 17460 21548
rect 17408 21505 17417 21539
rect 17417 21505 17451 21539
rect 17451 21505 17460 21539
rect 17408 21496 17460 21505
rect 17868 21496 17920 21548
rect 20812 21539 20864 21548
rect 20812 21505 20821 21539
rect 20821 21505 20855 21539
rect 20855 21505 20864 21539
rect 20812 21496 20864 21505
rect 21456 21539 21508 21548
rect 21456 21505 21465 21539
rect 21465 21505 21499 21539
rect 21499 21505 21508 21539
rect 21456 21496 21508 21505
rect 22192 21496 22244 21548
rect 23296 21496 23348 21548
rect 3516 21471 3568 21480
rect 3516 21437 3525 21471
rect 3525 21437 3559 21471
rect 3559 21437 3568 21471
rect 3516 21428 3568 21437
rect 5080 21471 5132 21480
rect 5080 21437 5089 21471
rect 5089 21437 5123 21471
rect 5123 21437 5132 21471
rect 5080 21428 5132 21437
rect 7288 21428 7340 21480
rect 10692 21360 10744 21412
rect 12532 21428 12584 21480
rect 11428 21360 11480 21412
rect 12900 21471 12952 21480
rect 12900 21437 12909 21471
rect 12909 21437 12943 21471
rect 12943 21437 12952 21471
rect 12900 21428 12952 21437
rect 13636 21428 13688 21480
rect 15660 21471 15712 21480
rect 15660 21437 15669 21471
rect 15669 21437 15703 21471
rect 15703 21437 15712 21471
rect 15660 21428 15712 21437
rect 16120 21428 16172 21480
rect 1768 21335 1820 21344
rect 1768 21301 1777 21335
rect 1777 21301 1811 21335
rect 1811 21301 1820 21335
rect 1768 21292 1820 21301
rect 7840 21292 7892 21344
rect 10508 21292 10560 21344
rect 11152 21335 11204 21344
rect 11152 21301 11161 21335
rect 11161 21301 11195 21335
rect 11195 21301 11204 21335
rect 11152 21292 11204 21301
rect 11704 21292 11756 21344
rect 11980 21292 12032 21344
rect 12900 21292 12952 21344
rect 16580 21360 16632 21412
rect 17500 21471 17552 21480
rect 17500 21437 17509 21471
rect 17509 21437 17543 21471
rect 17543 21437 17552 21471
rect 17500 21428 17552 21437
rect 17684 21471 17736 21480
rect 17684 21437 17693 21471
rect 17693 21437 17727 21471
rect 17727 21437 17736 21471
rect 17684 21428 17736 21437
rect 18420 21428 18472 21480
rect 18972 21428 19024 21480
rect 20996 21428 21048 21480
rect 21088 21471 21140 21480
rect 21088 21437 21097 21471
rect 21097 21437 21131 21471
rect 21131 21437 21140 21471
rect 21088 21428 21140 21437
rect 22468 21471 22520 21480
rect 22468 21437 22477 21471
rect 22477 21437 22511 21471
rect 22511 21437 22520 21471
rect 22468 21428 22520 21437
rect 22652 21471 22704 21480
rect 22652 21437 22661 21471
rect 22661 21437 22695 21471
rect 22695 21437 22704 21471
rect 22652 21428 22704 21437
rect 22744 21428 22796 21480
rect 23204 21428 23256 21480
rect 25688 21428 25740 21480
rect 13912 21292 13964 21344
rect 15016 21335 15068 21344
rect 15016 21301 15025 21335
rect 15025 21301 15059 21335
rect 15059 21301 15068 21335
rect 15016 21292 15068 21301
rect 15844 21292 15896 21344
rect 16212 21292 16264 21344
rect 16672 21335 16724 21344
rect 16672 21301 16681 21335
rect 16681 21301 16715 21335
rect 16715 21301 16724 21335
rect 16672 21292 16724 21301
rect 19064 21292 19116 21344
rect 19340 21292 19392 21344
rect 19984 21360 20036 21412
rect 21548 21360 21600 21412
rect 22284 21360 22336 21412
rect 24860 21360 24912 21412
rect 21824 21292 21876 21344
rect 22836 21292 22888 21344
rect 23848 21292 23900 21344
rect 2950 21190 3002 21242
rect 3014 21190 3066 21242
rect 3078 21190 3130 21242
rect 3142 21190 3194 21242
rect 3206 21190 3258 21242
rect 12950 21190 13002 21242
rect 13014 21190 13066 21242
rect 13078 21190 13130 21242
rect 13142 21190 13194 21242
rect 13206 21190 13258 21242
rect 22950 21190 23002 21242
rect 23014 21190 23066 21242
rect 23078 21190 23130 21242
rect 23142 21190 23194 21242
rect 23206 21190 23258 21242
rect 1768 21088 1820 21140
rect 10324 21088 10376 21140
rect 8300 21020 8352 21072
rect 8484 21020 8536 21072
rect 2780 20995 2832 21004
rect 2780 20961 2789 20995
rect 2789 20961 2823 20995
rect 2823 20961 2832 20995
rect 2780 20952 2832 20961
rect 4160 20952 4212 21004
rect 5632 20952 5684 21004
rect 5724 20884 5776 20936
rect 6920 20952 6972 21004
rect 8208 20952 8260 21004
rect 10508 20995 10560 21004
rect 10508 20961 10517 20995
rect 10517 20961 10551 20995
rect 10551 20961 10560 20995
rect 10508 20952 10560 20961
rect 11060 20952 11112 21004
rect 11428 20995 11480 21004
rect 11428 20961 11437 20995
rect 11437 20961 11471 20995
rect 11471 20961 11480 20995
rect 11428 20952 11480 20961
rect 7104 20927 7156 20936
rect 7104 20893 7113 20927
rect 7113 20893 7147 20927
rect 7147 20893 7156 20927
rect 7104 20884 7156 20893
rect 7748 20884 7800 20936
rect 12808 21088 12860 21140
rect 13452 21088 13504 21140
rect 13728 21020 13780 21072
rect 15384 21020 15436 21072
rect 15844 20952 15896 21004
rect 16580 21088 16632 21140
rect 16948 21020 17000 21072
rect 18236 21020 18288 21072
rect 16212 20952 16264 21004
rect 18604 21020 18656 21072
rect 20720 21020 20772 21072
rect 21180 21063 21232 21072
rect 21180 21029 21189 21063
rect 21189 21029 21223 21063
rect 21223 21029 21232 21063
rect 21180 21020 21232 21029
rect 22284 21020 22336 21072
rect 22652 21020 22704 21072
rect 13360 20884 13412 20936
rect 14464 20884 14516 20936
rect 14556 20884 14608 20936
rect 18696 20952 18748 21004
rect 19340 20884 19392 20936
rect 20720 20884 20772 20936
rect 21548 20952 21600 21004
rect 22008 20952 22060 21004
rect 22836 20952 22888 21004
rect 23664 21020 23716 21072
rect 24124 21063 24176 21072
rect 24124 21029 24133 21063
rect 24133 21029 24167 21063
rect 24167 21029 24176 21063
rect 24124 21020 24176 21029
rect 25136 20995 25188 21004
rect 25136 20961 25145 20995
rect 25145 20961 25179 20995
rect 25179 20961 25188 20995
rect 25136 20952 25188 20961
rect 20996 20884 21048 20936
rect 8300 20816 8352 20868
rect 6184 20748 6236 20800
rect 8760 20816 8812 20868
rect 8944 20791 8996 20800
rect 8944 20757 8953 20791
rect 8953 20757 8987 20791
rect 8987 20757 8996 20791
rect 8944 20748 8996 20757
rect 11888 20816 11940 20868
rect 14004 20816 14056 20868
rect 14096 20816 14148 20868
rect 15292 20816 15344 20868
rect 15384 20816 15436 20868
rect 12440 20748 12492 20800
rect 12808 20748 12860 20800
rect 13728 20748 13780 20800
rect 14832 20791 14884 20800
rect 14832 20757 14841 20791
rect 14841 20757 14875 20791
rect 14875 20757 14884 20791
rect 14832 20748 14884 20757
rect 15844 20791 15896 20800
rect 15844 20757 15853 20791
rect 15853 20757 15887 20791
rect 15887 20757 15896 20791
rect 15844 20748 15896 20757
rect 17040 20791 17092 20800
rect 17040 20757 17049 20791
rect 17049 20757 17083 20791
rect 17083 20757 17092 20791
rect 17040 20748 17092 20757
rect 18972 20816 19024 20868
rect 23204 20927 23256 20936
rect 23204 20893 23213 20927
rect 23213 20893 23247 20927
rect 23247 20893 23256 20927
rect 23204 20884 23256 20893
rect 19248 20748 19300 20800
rect 21180 20748 21232 20800
rect 21916 20748 21968 20800
rect 22100 20791 22152 20800
rect 22100 20757 22109 20791
rect 22109 20757 22143 20791
rect 22143 20757 22152 20791
rect 22100 20748 22152 20757
rect 26056 20748 26108 20800
rect 7950 20646 8002 20698
rect 8014 20646 8066 20698
rect 8078 20646 8130 20698
rect 8142 20646 8194 20698
rect 8206 20646 8258 20698
rect 17950 20646 18002 20698
rect 18014 20646 18066 20698
rect 18078 20646 18130 20698
rect 18142 20646 18194 20698
rect 18206 20646 18258 20698
rect 3976 20544 4028 20596
rect 4712 20544 4764 20596
rect 5172 20587 5224 20596
rect 5172 20553 5181 20587
rect 5181 20553 5215 20587
rect 5215 20553 5224 20587
rect 5172 20544 5224 20553
rect 6552 20587 6604 20596
rect 6552 20553 6561 20587
rect 6561 20553 6595 20587
rect 6595 20553 6604 20587
rect 6552 20544 6604 20553
rect 7196 20544 7248 20596
rect 7748 20587 7800 20596
rect 7748 20553 7757 20587
rect 7757 20553 7791 20587
rect 7791 20553 7800 20587
rect 7748 20544 7800 20553
rect 5356 20476 5408 20528
rect 5540 20408 5592 20460
rect 7196 20408 7248 20460
rect 3332 20383 3384 20392
rect 3332 20349 3341 20383
rect 3341 20349 3375 20383
rect 3375 20349 3384 20383
rect 3332 20340 3384 20349
rect 6552 20340 6604 20392
rect 7012 20340 7064 20392
rect 7748 20340 7800 20392
rect 8392 20340 8444 20392
rect 10140 20544 10192 20596
rect 10324 20544 10376 20596
rect 8944 20476 8996 20528
rect 9772 20476 9824 20528
rect 9036 20451 9088 20460
rect 9036 20417 9045 20451
rect 9045 20417 9079 20451
rect 9079 20417 9088 20451
rect 9036 20408 9088 20417
rect 10784 20544 10836 20596
rect 12348 20544 12400 20596
rect 12440 20587 12492 20596
rect 12440 20553 12449 20587
rect 12449 20553 12483 20587
rect 12483 20553 12492 20587
rect 12440 20544 12492 20553
rect 12532 20544 12584 20596
rect 12808 20544 12860 20596
rect 11152 20519 11204 20528
rect 11152 20485 11161 20519
rect 11161 20485 11195 20519
rect 11195 20485 11204 20519
rect 11152 20476 11204 20485
rect 11888 20476 11940 20528
rect 14832 20544 14884 20596
rect 15384 20544 15436 20596
rect 14096 20476 14148 20528
rect 15292 20476 15344 20528
rect 16764 20476 16816 20528
rect 18604 20544 18656 20596
rect 18696 20587 18748 20596
rect 18696 20553 18705 20587
rect 18705 20553 18739 20587
rect 18739 20553 18748 20587
rect 18696 20544 18748 20553
rect 8944 20340 8996 20392
rect 10508 20340 10560 20392
rect 5172 20272 5224 20324
rect 4160 20204 4212 20256
rect 6828 20204 6880 20256
rect 8392 20247 8444 20256
rect 8392 20213 8401 20247
rect 8401 20213 8435 20247
rect 8435 20213 8444 20247
rect 8392 20204 8444 20213
rect 9404 20204 9456 20256
rect 10784 20247 10836 20256
rect 10784 20213 10793 20247
rect 10793 20213 10827 20247
rect 10827 20213 10836 20247
rect 10784 20204 10836 20213
rect 12164 20340 12216 20392
rect 12808 20340 12860 20392
rect 15844 20451 15896 20460
rect 15844 20417 15853 20451
rect 15853 20417 15887 20451
rect 15887 20417 15896 20451
rect 15844 20408 15896 20417
rect 18328 20408 18380 20460
rect 13452 20272 13504 20324
rect 12256 20204 12308 20256
rect 13820 20340 13872 20392
rect 16488 20340 16540 20392
rect 17224 20383 17276 20392
rect 17224 20349 17233 20383
rect 17233 20349 17267 20383
rect 17267 20349 17276 20383
rect 20904 20544 20956 20596
rect 25136 20544 25188 20596
rect 22468 20519 22520 20528
rect 22468 20485 22477 20519
rect 22477 20485 22511 20519
rect 22511 20485 22520 20519
rect 22468 20476 22520 20485
rect 23664 20476 23716 20528
rect 23848 20476 23900 20528
rect 24216 20476 24268 20528
rect 20628 20408 20680 20460
rect 17224 20340 17276 20349
rect 19248 20383 19300 20392
rect 19248 20349 19257 20383
rect 19257 20349 19291 20383
rect 19291 20349 19300 20383
rect 19248 20340 19300 20349
rect 19892 20340 19944 20392
rect 20812 20340 20864 20392
rect 14832 20272 14884 20324
rect 13636 20204 13688 20256
rect 15936 20247 15988 20256
rect 15936 20213 15945 20247
rect 15945 20213 15979 20247
rect 15979 20213 15988 20247
rect 15936 20204 15988 20213
rect 20904 20272 20956 20324
rect 22652 20383 22704 20392
rect 22652 20349 22661 20383
rect 22661 20349 22695 20383
rect 22695 20349 22704 20383
rect 22652 20340 22704 20349
rect 23296 20408 23348 20460
rect 24124 20340 24176 20392
rect 24768 20340 24820 20392
rect 18604 20204 18656 20256
rect 19616 20204 19668 20256
rect 20536 20204 20588 20256
rect 22836 20204 22888 20256
rect 23940 20204 23992 20256
rect 25228 20247 25280 20256
rect 25228 20213 25237 20247
rect 25237 20213 25271 20247
rect 25271 20213 25280 20247
rect 25228 20204 25280 20213
rect 2950 20102 3002 20154
rect 3014 20102 3066 20154
rect 3078 20102 3130 20154
rect 3142 20102 3194 20154
rect 3206 20102 3258 20154
rect 12950 20102 13002 20154
rect 13014 20102 13066 20154
rect 13078 20102 13130 20154
rect 13142 20102 13194 20154
rect 13206 20102 13258 20154
rect 22950 20102 23002 20154
rect 23014 20102 23066 20154
rect 23078 20102 23130 20154
rect 23142 20102 23194 20154
rect 23206 20102 23258 20154
rect 3976 20000 4028 20052
rect 2044 19864 2096 19916
rect 5264 19864 5316 19916
rect 4712 19839 4764 19848
rect 4712 19805 4721 19839
rect 4721 19805 4755 19839
rect 4755 19805 4764 19839
rect 4712 19796 4764 19805
rect 5816 19796 5868 19848
rect 6644 19839 6696 19848
rect 6644 19805 6653 19839
rect 6653 19805 6687 19839
rect 6687 19805 6696 19839
rect 6644 19796 6696 19805
rect 7196 20000 7248 20052
rect 7472 19864 7524 19916
rect 15200 20000 15252 20052
rect 18328 20000 18380 20052
rect 20628 20000 20680 20052
rect 21088 20000 21140 20052
rect 13360 19975 13412 19984
rect 13360 19941 13369 19975
rect 13369 19941 13403 19975
rect 13403 19941 13412 19975
rect 13360 19932 13412 19941
rect 13452 19932 13504 19984
rect 10968 19907 11020 19916
rect 10968 19873 10977 19907
rect 10977 19873 11011 19907
rect 11011 19873 11020 19907
rect 10968 19864 11020 19873
rect 12256 19864 12308 19916
rect 12348 19864 12400 19916
rect 15660 19864 15712 19916
rect 17960 19864 18012 19916
rect 18604 19932 18656 19984
rect 23388 20000 23440 20052
rect 23940 20000 23992 20052
rect 24216 20000 24268 20052
rect 20904 19864 20956 19916
rect 23296 19864 23348 19916
rect 24492 19864 24544 19916
rect 25044 19907 25096 19916
rect 25044 19873 25053 19907
rect 25053 19873 25087 19907
rect 25087 19873 25096 19907
rect 25044 19864 25096 19873
rect 25964 19864 26016 19916
rect 11060 19796 11112 19848
rect 14096 19796 14148 19848
rect 14188 19796 14240 19848
rect 15108 19796 15160 19848
rect 18420 19796 18472 19848
rect 18880 19839 18932 19848
rect 18880 19805 18889 19839
rect 18889 19805 18923 19839
rect 18923 19805 18932 19839
rect 18880 19796 18932 19805
rect 19708 19796 19760 19848
rect 24032 19796 24084 19848
rect 8300 19728 8352 19780
rect 5540 19660 5592 19712
rect 7012 19660 7064 19712
rect 7472 19660 7524 19712
rect 9128 19703 9180 19712
rect 9128 19669 9137 19703
rect 9137 19669 9171 19703
rect 9171 19669 9180 19703
rect 9128 19660 9180 19669
rect 10876 19660 10928 19712
rect 11520 19660 11572 19712
rect 11796 19660 11848 19712
rect 13728 19728 13780 19780
rect 14556 19728 14608 19780
rect 14648 19728 14700 19780
rect 14832 19728 14884 19780
rect 15016 19728 15068 19780
rect 15384 19771 15436 19780
rect 15384 19737 15393 19771
rect 15393 19737 15427 19771
rect 15427 19737 15436 19771
rect 15384 19728 15436 19737
rect 16212 19771 16264 19780
rect 16212 19737 16221 19771
rect 16221 19737 16255 19771
rect 16255 19737 16264 19771
rect 16212 19728 16264 19737
rect 16764 19728 16816 19780
rect 18236 19728 18288 19780
rect 20536 19728 20588 19780
rect 21364 19771 21416 19780
rect 21364 19737 21373 19771
rect 21373 19737 21407 19771
rect 21407 19737 21416 19771
rect 21364 19728 21416 19737
rect 21640 19728 21692 19780
rect 24308 19728 24360 19780
rect 13912 19660 13964 19712
rect 16304 19703 16356 19712
rect 16304 19669 16313 19703
rect 16313 19669 16347 19703
rect 16347 19669 16356 19703
rect 16304 19660 16356 19669
rect 16580 19660 16632 19712
rect 18420 19660 18472 19712
rect 18604 19660 18656 19712
rect 18788 19660 18840 19712
rect 19524 19660 19576 19712
rect 20720 19660 20772 19712
rect 22008 19660 22060 19712
rect 23572 19660 23624 19712
rect 24584 19703 24636 19712
rect 24584 19669 24593 19703
rect 24593 19669 24627 19703
rect 24627 19669 24636 19703
rect 24584 19660 24636 19669
rect 24860 19660 24912 19712
rect 25964 19660 26016 19712
rect 7950 19558 8002 19610
rect 8014 19558 8066 19610
rect 8078 19558 8130 19610
rect 8142 19558 8194 19610
rect 8206 19558 8258 19610
rect 17950 19558 18002 19610
rect 18014 19558 18066 19610
rect 18078 19558 18130 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 3884 19499 3936 19508
rect 3884 19465 3893 19499
rect 3893 19465 3927 19499
rect 3927 19465 3936 19499
rect 3884 19456 3936 19465
rect 5816 19499 5868 19508
rect 5816 19465 5825 19499
rect 5825 19465 5859 19499
rect 5859 19465 5868 19499
rect 5816 19456 5868 19465
rect 6736 19456 6788 19508
rect 12164 19456 12216 19508
rect 12348 19456 12400 19508
rect 13360 19456 13412 19508
rect 14372 19456 14424 19508
rect 14556 19456 14608 19508
rect 14832 19456 14884 19508
rect 18696 19456 18748 19508
rect 3792 19320 3844 19372
rect 8300 19388 8352 19440
rect 4896 19320 4948 19372
rect 6000 19363 6052 19372
rect 6000 19329 6009 19363
rect 6009 19329 6043 19363
rect 6043 19329 6052 19363
rect 6000 19320 6052 19329
rect 1860 19252 1912 19304
rect 3332 19252 3384 19304
rect 6460 19295 6512 19304
rect 6460 19261 6469 19295
rect 6469 19261 6503 19295
rect 6503 19261 6512 19295
rect 6460 19252 6512 19261
rect 7748 19320 7800 19372
rect 9220 19388 9272 19440
rect 9772 19388 9824 19440
rect 14280 19388 14332 19440
rect 7196 19252 7248 19304
rect 7656 19252 7708 19304
rect 6920 19184 6972 19236
rect 5356 19116 5408 19168
rect 7012 19116 7064 19168
rect 7288 19116 7340 19168
rect 7656 19116 7708 19168
rect 9036 19363 9088 19372
rect 9036 19329 9045 19363
rect 9045 19329 9079 19363
rect 9079 19329 9088 19363
rect 9036 19320 9088 19329
rect 12256 19320 12308 19372
rect 14096 19320 14148 19372
rect 15292 19320 15344 19372
rect 10784 19252 10836 19304
rect 12072 19295 12124 19304
rect 12072 19261 12081 19295
rect 12081 19261 12115 19295
rect 12115 19261 12124 19295
rect 12072 19252 12124 19261
rect 13636 19252 13688 19304
rect 15108 19252 15160 19304
rect 15660 19320 15712 19372
rect 16672 19388 16724 19440
rect 18328 19388 18380 19440
rect 19340 19456 19392 19508
rect 20812 19499 20864 19508
rect 20812 19465 20821 19499
rect 20821 19465 20855 19499
rect 20855 19465 20864 19499
rect 20812 19456 20864 19465
rect 21272 19456 21324 19508
rect 22100 19456 22152 19508
rect 22468 19456 22520 19508
rect 19892 19388 19944 19440
rect 23020 19388 23072 19440
rect 16488 19320 16540 19372
rect 19064 19320 19116 19372
rect 16028 19252 16080 19304
rect 17684 19252 17736 19304
rect 19892 19295 19944 19304
rect 19892 19261 19901 19295
rect 19901 19261 19935 19295
rect 19935 19261 19944 19295
rect 19892 19252 19944 19261
rect 20444 19320 20496 19372
rect 20904 19363 20956 19372
rect 20904 19329 20913 19363
rect 20913 19329 20947 19363
rect 20947 19329 20956 19363
rect 20904 19320 20956 19329
rect 21364 19320 21416 19372
rect 23848 19456 23900 19508
rect 23940 19456 23992 19508
rect 25044 19499 25096 19508
rect 25044 19465 25053 19499
rect 25053 19465 25087 19499
rect 25087 19465 25096 19499
rect 25044 19456 25096 19465
rect 23296 19363 23348 19372
rect 23296 19329 23305 19363
rect 23305 19329 23339 19363
rect 23339 19329 23348 19363
rect 23296 19320 23348 19329
rect 21640 19252 21692 19304
rect 8208 19184 8260 19236
rect 8668 19184 8720 19236
rect 10324 19184 10376 19236
rect 11428 19184 11480 19236
rect 14372 19184 14424 19236
rect 14740 19184 14792 19236
rect 17040 19184 17092 19236
rect 18420 19184 18472 19236
rect 22100 19184 22152 19236
rect 7932 19116 7984 19168
rect 9496 19116 9548 19168
rect 10784 19159 10836 19168
rect 10784 19125 10793 19159
rect 10793 19125 10827 19159
rect 10827 19125 10836 19159
rect 10784 19116 10836 19125
rect 10968 19116 11020 19168
rect 11244 19159 11296 19168
rect 11244 19125 11253 19159
rect 11253 19125 11287 19159
rect 11287 19125 11296 19159
rect 11244 19116 11296 19125
rect 11796 19159 11848 19168
rect 11796 19125 11805 19159
rect 11805 19125 11839 19159
rect 11839 19125 11848 19159
rect 11796 19116 11848 19125
rect 11888 19116 11940 19168
rect 13360 19116 13412 19168
rect 13728 19116 13780 19168
rect 14832 19116 14884 19168
rect 15568 19116 15620 19168
rect 16120 19159 16172 19168
rect 16120 19125 16129 19159
rect 16129 19125 16163 19159
rect 16163 19125 16172 19159
rect 16120 19116 16172 19125
rect 17132 19116 17184 19168
rect 18788 19116 18840 19168
rect 20720 19116 20772 19168
rect 20996 19116 21048 19168
rect 21916 19159 21968 19168
rect 21916 19125 21925 19159
rect 21925 19125 21959 19159
rect 21959 19125 21968 19159
rect 22560 19295 22612 19304
rect 22560 19261 22569 19295
rect 22569 19261 22603 19295
rect 22603 19261 22612 19295
rect 22560 19252 22612 19261
rect 25228 19252 25280 19304
rect 21916 19116 21968 19125
rect 24032 19116 24084 19168
rect 24676 19116 24728 19168
rect 2950 19014 3002 19066
rect 3014 19014 3066 19066
rect 3078 19014 3130 19066
rect 3142 19014 3194 19066
rect 3206 19014 3258 19066
rect 12950 19014 13002 19066
rect 13014 19014 13066 19066
rect 13078 19014 13130 19066
rect 13142 19014 13194 19066
rect 13206 19014 13258 19066
rect 22950 19014 23002 19066
rect 23014 19014 23066 19066
rect 23078 19014 23130 19066
rect 23142 19014 23194 19066
rect 23206 19014 23258 19066
rect 1952 18955 2004 18964
rect 1952 18921 1961 18955
rect 1961 18921 1995 18955
rect 1995 18921 2004 18955
rect 1952 18912 2004 18921
rect 5908 18912 5960 18964
rect 6736 18912 6788 18964
rect 7012 18912 7064 18964
rect 2596 18887 2648 18896
rect 2596 18853 2605 18887
rect 2605 18853 2639 18887
rect 2639 18853 2648 18887
rect 2596 18844 2648 18853
rect 8116 18844 8168 18896
rect 8300 18912 8352 18964
rect 9680 18912 9732 18964
rect 14280 18955 14332 18964
rect 14280 18921 14289 18955
rect 14289 18921 14323 18955
rect 14323 18921 14332 18955
rect 14280 18912 14332 18921
rect 9496 18844 9548 18896
rect 11888 18844 11940 18896
rect 6092 18776 6144 18828
rect 7564 18776 7616 18828
rect 10048 18776 10100 18828
rect 11152 18776 11204 18828
rect 17224 18887 17276 18896
rect 17224 18853 17233 18887
rect 17233 18853 17267 18887
rect 17267 18853 17276 18887
rect 17224 18844 17276 18853
rect 2136 18751 2188 18760
rect 2136 18717 2145 18751
rect 2145 18717 2179 18751
rect 2179 18717 2188 18751
rect 2136 18708 2188 18717
rect 4160 18708 4212 18760
rect 4712 18751 4764 18760
rect 4712 18717 4721 18751
rect 4721 18717 4755 18751
rect 4755 18717 4764 18751
rect 4712 18708 4764 18717
rect 3884 18683 3936 18692
rect 3884 18649 3893 18683
rect 3893 18649 3927 18683
rect 3927 18649 3936 18683
rect 3884 18640 3936 18649
rect 6000 18751 6052 18760
rect 6000 18717 6009 18751
rect 6009 18717 6043 18751
rect 6043 18717 6052 18751
rect 6000 18708 6052 18717
rect 6460 18708 6512 18760
rect 8392 18708 8444 18760
rect 7932 18640 7984 18692
rect 9128 18708 9180 18760
rect 9772 18708 9824 18760
rect 10324 18708 10376 18760
rect 11796 18708 11848 18760
rect 11888 18708 11940 18760
rect 12624 18776 12676 18828
rect 12716 18776 12768 18828
rect 13452 18776 13504 18828
rect 13636 18819 13688 18828
rect 13636 18785 13645 18819
rect 13645 18785 13679 18819
rect 13679 18785 13688 18819
rect 13636 18776 13688 18785
rect 14556 18776 14608 18828
rect 14740 18819 14792 18828
rect 14740 18785 14749 18819
rect 14749 18785 14783 18819
rect 14783 18785 14792 18819
rect 14740 18776 14792 18785
rect 15108 18776 15160 18828
rect 15292 18776 15344 18828
rect 16488 18776 16540 18828
rect 9312 18640 9364 18692
rect 13820 18708 13872 18760
rect 14924 18708 14976 18760
rect 17868 18776 17920 18828
rect 18328 18776 18380 18828
rect 18788 18912 18840 18964
rect 21824 18912 21876 18964
rect 24860 18844 24912 18896
rect 18420 18751 18472 18760
rect 18420 18717 18429 18751
rect 18429 18717 18463 18751
rect 18463 18717 18472 18751
rect 18420 18708 18472 18717
rect 22928 18776 22980 18828
rect 18788 18708 18840 18760
rect 19616 18751 19668 18760
rect 19616 18717 19625 18751
rect 19625 18717 19659 18751
rect 19659 18717 19668 18751
rect 19616 18708 19668 18717
rect 13728 18640 13780 18692
rect 8852 18572 8904 18624
rect 9496 18572 9548 18624
rect 10508 18572 10560 18624
rect 11704 18615 11756 18624
rect 11704 18581 11713 18615
rect 11713 18581 11747 18615
rect 11747 18581 11756 18615
rect 11704 18572 11756 18581
rect 12624 18572 12676 18624
rect 12716 18615 12768 18624
rect 12716 18581 12725 18615
rect 12725 18581 12759 18615
rect 12759 18581 12768 18615
rect 12716 18572 12768 18581
rect 13452 18615 13504 18624
rect 13452 18581 13461 18615
rect 13461 18581 13495 18615
rect 13495 18581 13504 18615
rect 13452 18572 13504 18581
rect 13636 18572 13688 18624
rect 15200 18640 15252 18692
rect 16028 18640 16080 18692
rect 17132 18640 17184 18692
rect 17960 18640 18012 18692
rect 18328 18640 18380 18692
rect 19248 18640 19300 18692
rect 22376 18708 22428 18760
rect 25228 18819 25280 18828
rect 25228 18785 25237 18819
rect 25237 18785 25271 18819
rect 25271 18785 25280 18819
rect 25228 18776 25280 18785
rect 23480 18708 23532 18760
rect 20628 18683 20680 18692
rect 20628 18649 20637 18683
rect 20637 18649 20671 18683
rect 20671 18649 20680 18683
rect 20628 18640 20680 18649
rect 21640 18640 21692 18692
rect 15016 18572 15068 18624
rect 17684 18615 17736 18624
rect 17684 18581 17693 18615
rect 17693 18581 17727 18615
rect 17727 18581 17736 18615
rect 17684 18572 17736 18581
rect 18420 18572 18472 18624
rect 19524 18572 19576 18624
rect 20444 18572 20496 18624
rect 20904 18572 20956 18624
rect 22468 18640 22520 18692
rect 22192 18572 22244 18624
rect 22560 18615 22612 18624
rect 22560 18581 22569 18615
rect 22569 18581 22603 18615
rect 22603 18581 22612 18615
rect 22560 18572 22612 18581
rect 22744 18640 22796 18692
rect 23940 18640 23992 18692
rect 25504 18640 25556 18692
rect 23204 18572 23256 18624
rect 24584 18615 24636 18624
rect 24584 18581 24593 18615
rect 24593 18581 24627 18615
rect 24627 18581 24636 18615
rect 24584 18572 24636 18581
rect 7950 18470 8002 18522
rect 8014 18470 8066 18522
rect 8078 18470 8130 18522
rect 8142 18470 8194 18522
rect 8206 18470 8258 18522
rect 17950 18470 18002 18522
rect 18014 18470 18066 18522
rect 18078 18470 18130 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 3516 18368 3568 18420
rect 3700 18368 3752 18420
rect 4988 18368 5040 18420
rect 5724 18368 5776 18420
rect 6000 18368 6052 18420
rect 2228 18343 2280 18352
rect 2228 18309 2237 18343
rect 2237 18309 2271 18343
rect 2271 18309 2280 18343
rect 2228 18300 2280 18309
rect 4620 18300 4672 18352
rect 6828 18300 6880 18352
rect 5540 18232 5592 18284
rect 6920 18232 6972 18284
rect 7196 18275 7248 18284
rect 7196 18241 7205 18275
rect 7205 18241 7239 18275
rect 7239 18241 7248 18275
rect 7196 18232 7248 18241
rect 8576 18300 8628 18352
rect 10784 18368 10836 18420
rect 10968 18368 11020 18420
rect 11888 18368 11940 18420
rect 12072 18368 12124 18420
rect 13820 18368 13872 18420
rect 14556 18368 14608 18420
rect 15568 18368 15620 18420
rect 9772 18300 9824 18352
rect 10600 18300 10652 18352
rect 11796 18300 11848 18352
rect 18512 18368 18564 18420
rect 19708 18411 19760 18420
rect 19708 18377 19717 18411
rect 19717 18377 19751 18411
rect 19751 18377 19760 18411
rect 19708 18368 19760 18377
rect 20076 18368 20128 18420
rect 21640 18368 21692 18420
rect 23020 18368 23072 18420
rect 23112 18368 23164 18420
rect 23296 18411 23348 18420
rect 23296 18377 23305 18411
rect 23305 18377 23339 18411
rect 23339 18377 23348 18411
rect 23296 18368 23348 18377
rect 24676 18368 24728 18420
rect 24860 18368 24912 18420
rect 16488 18343 16540 18352
rect 16488 18309 16497 18343
rect 16497 18309 16531 18343
rect 16531 18309 16540 18343
rect 16488 18300 16540 18309
rect 17132 18300 17184 18352
rect 20628 18300 20680 18352
rect 21088 18300 21140 18352
rect 21456 18300 21508 18352
rect 25596 18300 25648 18352
rect 6276 18164 6328 18216
rect 8484 18275 8536 18284
rect 8484 18241 8493 18275
rect 8493 18241 8527 18275
rect 8527 18241 8536 18275
rect 8484 18232 8536 18241
rect 8944 18275 8996 18284
rect 8944 18241 8953 18275
rect 8953 18241 8987 18275
rect 8987 18241 8996 18275
rect 8944 18232 8996 18241
rect 10508 18232 10560 18284
rect 9312 18164 9364 18216
rect 3608 18096 3660 18148
rect 4620 18096 4672 18148
rect 6368 18096 6420 18148
rect 7012 18139 7064 18148
rect 7012 18105 7021 18139
rect 7021 18105 7055 18139
rect 7055 18105 7064 18139
rect 7012 18096 7064 18105
rect 4068 18028 4120 18080
rect 7288 18028 7340 18080
rect 7656 18071 7708 18080
rect 7656 18037 7665 18071
rect 7665 18037 7699 18071
rect 7699 18037 7708 18071
rect 7656 18028 7708 18037
rect 9772 18028 9824 18080
rect 11152 18028 11204 18080
rect 12348 18207 12400 18216
rect 12348 18173 12357 18207
rect 12357 18173 12391 18207
rect 12391 18173 12400 18207
rect 12348 18164 12400 18173
rect 12624 18164 12676 18216
rect 15108 18164 15160 18216
rect 16856 18232 16908 18284
rect 17224 18275 17276 18284
rect 17224 18241 17233 18275
rect 17233 18241 17267 18275
rect 17267 18241 17276 18275
rect 17224 18232 17276 18241
rect 17500 18232 17552 18284
rect 19524 18232 19576 18284
rect 20444 18232 20496 18284
rect 20812 18275 20864 18284
rect 20812 18241 20821 18275
rect 20821 18241 20855 18275
rect 20855 18241 20864 18275
rect 20812 18232 20864 18241
rect 21180 18232 21232 18284
rect 22560 18232 22612 18284
rect 25320 18232 25372 18284
rect 17408 18207 17460 18216
rect 17408 18173 17417 18207
rect 17417 18173 17451 18207
rect 17451 18173 17460 18207
rect 17408 18164 17460 18173
rect 18236 18164 18288 18216
rect 18696 18207 18748 18216
rect 18696 18173 18705 18207
rect 18705 18173 18739 18207
rect 18739 18173 18748 18207
rect 18696 18164 18748 18173
rect 19064 18096 19116 18148
rect 19432 18164 19484 18216
rect 19800 18164 19852 18216
rect 20812 18096 20864 18148
rect 21916 18164 21968 18216
rect 22100 18164 22152 18216
rect 22468 18164 22520 18216
rect 23940 18164 23992 18216
rect 25412 18164 25464 18216
rect 21180 18096 21232 18148
rect 17500 18028 17552 18080
rect 19892 18028 19944 18080
rect 20444 18071 20496 18080
rect 20444 18037 20453 18071
rect 20453 18037 20487 18071
rect 20487 18037 20496 18071
rect 20444 18028 20496 18037
rect 22560 18028 22612 18080
rect 23112 18028 23164 18080
rect 2950 17926 3002 17978
rect 3014 17926 3066 17978
rect 3078 17926 3130 17978
rect 3142 17926 3194 17978
rect 3206 17926 3258 17978
rect 12950 17926 13002 17978
rect 13014 17926 13066 17978
rect 13078 17926 13130 17978
rect 13142 17926 13194 17978
rect 13206 17926 13258 17978
rect 22950 17926 23002 17978
rect 23014 17926 23066 17978
rect 23078 17926 23130 17978
rect 23142 17926 23194 17978
rect 23206 17926 23258 17978
rect 3332 17824 3384 17876
rect 5448 17824 5500 17876
rect 7104 17824 7156 17876
rect 6920 17756 6972 17808
rect 7196 17756 7248 17808
rect 3424 17663 3476 17672
rect 3424 17629 3433 17663
rect 3433 17629 3467 17663
rect 3467 17629 3476 17663
rect 3424 17620 3476 17629
rect 5448 17663 5500 17672
rect 5448 17629 5457 17663
rect 5457 17629 5491 17663
rect 5491 17629 5500 17663
rect 5448 17620 5500 17629
rect 6184 17620 6236 17672
rect 7288 17663 7340 17672
rect 7288 17629 7297 17663
rect 7297 17629 7331 17663
rect 7331 17629 7340 17663
rect 7288 17620 7340 17629
rect 7840 17620 7892 17672
rect 9680 17756 9732 17808
rect 11244 17756 11296 17808
rect 11888 17756 11940 17808
rect 13452 17824 13504 17876
rect 13912 17756 13964 17808
rect 20628 17824 20680 17876
rect 22192 17824 22244 17876
rect 22652 17824 22704 17876
rect 24952 17824 25004 17876
rect 8944 17688 8996 17740
rect 11704 17688 11756 17740
rect 12808 17688 12860 17740
rect 13268 17688 13320 17740
rect 13728 17688 13780 17740
rect 14924 17731 14976 17740
rect 14924 17697 14933 17731
rect 14933 17697 14967 17731
rect 14967 17697 14976 17731
rect 14924 17688 14976 17697
rect 15752 17688 15804 17740
rect 17868 17756 17920 17808
rect 19432 17756 19484 17808
rect 20168 17756 20220 17808
rect 8300 17552 8352 17604
rect 16304 17620 16356 17672
rect 16488 17620 16540 17672
rect 16856 17688 16908 17740
rect 19800 17688 19852 17740
rect 22560 17756 22612 17808
rect 23296 17756 23348 17808
rect 23756 17731 23808 17740
rect 23756 17697 23765 17731
rect 23765 17697 23799 17731
rect 23799 17697 23808 17731
rect 23756 17688 23808 17697
rect 23848 17731 23900 17740
rect 23848 17697 23857 17731
rect 23857 17697 23891 17731
rect 23891 17697 23900 17731
rect 23848 17688 23900 17697
rect 25872 17688 25924 17740
rect 17040 17620 17092 17672
rect 18604 17620 18656 17672
rect 18880 17620 18932 17672
rect 20076 17620 20128 17672
rect 22744 17620 22796 17672
rect 9956 17552 10008 17604
rect 10048 17595 10100 17604
rect 10048 17561 10057 17595
rect 10057 17561 10091 17595
rect 10091 17561 10100 17595
rect 10048 17552 10100 17561
rect 10324 17552 10376 17604
rect 10508 17552 10560 17604
rect 4252 17527 4304 17536
rect 4252 17493 4261 17527
rect 4261 17493 4295 17527
rect 4295 17493 4304 17527
rect 4252 17484 4304 17493
rect 6828 17484 6880 17536
rect 7104 17527 7156 17536
rect 7104 17493 7113 17527
rect 7113 17493 7147 17527
rect 7147 17493 7156 17527
rect 7104 17484 7156 17493
rect 8392 17527 8444 17536
rect 8392 17493 8401 17527
rect 8401 17493 8435 17527
rect 8435 17493 8444 17527
rect 8392 17484 8444 17493
rect 9128 17527 9180 17536
rect 9128 17493 9137 17527
rect 9137 17493 9171 17527
rect 9171 17493 9180 17527
rect 9128 17484 9180 17493
rect 9312 17484 9364 17536
rect 12164 17552 12216 17604
rect 12716 17552 12768 17604
rect 14556 17552 14608 17604
rect 15108 17552 15160 17604
rect 15200 17595 15252 17604
rect 15200 17561 15209 17595
rect 15209 17561 15243 17595
rect 15243 17561 15252 17595
rect 15200 17552 15252 17561
rect 11428 17484 11480 17536
rect 12256 17484 12308 17536
rect 17408 17552 17460 17604
rect 16580 17484 16632 17536
rect 17684 17484 17736 17536
rect 19524 17484 19576 17536
rect 20260 17484 20312 17536
rect 22468 17552 22520 17604
rect 23756 17552 23808 17604
rect 24676 17552 24728 17604
rect 21916 17484 21968 17536
rect 23388 17484 23440 17536
rect 23848 17484 23900 17536
rect 7950 17382 8002 17434
rect 8014 17382 8066 17434
rect 8078 17382 8130 17434
rect 8142 17382 8194 17434
rect 8206 17382 8258 17434
rect 17950 17382 18002 17434
rect 18014 17382 18066 17434
rect 18078 17382 18130 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 3976 17280 4028 17332
rect 4252 17280 4304 17332
rect 7012 17280 7064 17332
rect 7196 17323 7248 17332
rect 7196 17289 7205 17323
rect 7205 17289 7239 17323
rect 7239 17289 7248 17323
rect 7196 17280 7248 17289
rect 7380 17280 7432 17332
rect 8392 17280 8444 17332
rect 15936 17280 15988 17332
rect 5172 17212 5224 17264
rect 6920 17144 6972 17196
rect 7288 17144 7340 17196
rect 7748 17144 7800 17196
rect 8760 17187 8812 17196
rect 8760 17153 8769 17187
rect 8769 17153 8803 17187
rect 8803 17153 8812 17187
rect 8760 17144 8812 17153
rect 4804 17119 4856 17128
rect 4804 17085 4813 17119
rect 4813 17085 4847 17119
rect 4847 17085 4856 17119
rect 4804 17076 4856 17085
rect 5448 17076 5500 17128
rect 9404 17212 9456 17264
rect 9772 17212 9824 17264
rect 11428 17212 11480 17264
rect 12716 17212 12768 17264
rect 16212 17212 16264 17264
rect 16856 17212 16908 17264
rect 17868 17212 17920 17264
rect 8944 17144 8996 17196
rect 10600 17144 10652 17196
rect 11704 17187 11756 17196
rect 11704 17153 11713 17187
rect 11713 17153 11747 17187
rect 11747 17153 11756 17187
rect 11704 17144 11756 17153
rect 14556 17144 14608 17196
rect 15016 17187 15068 17196
rect 15016 17153 15025 17187
rect 15025 17153 15059 17187
rect 15059 17153 15068 17187
rect 15016 17144 15068 17153
rect 10048 17076 10100 17128
rect 13268 17076 13320 17128
rect 13820 17076 13872 17128
rect 14096 17076 14148 17128
rect 16948 17144 17000 17196
rect 8668 17008 8720 17060
rect 6552 16983 6604 16992
rect 6552 16949 6561 16983
rect 6561 16949 6595 16983
rect 6595 16949 6604 16983
rect 6552 16940 6604 16949
rect 9496 16940 9548 16992
rect 9956 16940 10008 16992
rect 11060 16940 11112 16992
rect 14832 16983 14884 16992
rect 14832 16949 14841 16983
rect 14841 16949 14875 16983
rect 14875 16949 14884 16983
rect 14832 16940 14884 16949
rect 15016 16940 15068 16992
rect 16856 17051 16908 17060
rect 16856 17017 16865 17051
rect 16865 17017 16899 17051
rect 16899 17017 16908 17051
rect 16856 17008 16908 17017
rect 16488 16940 16540 16992
rect 16580 16940 16632 16992
rect 17684 17076 17736 17128
rect 18972 17280 19024 17332
rect 20168 17280 20220 17332
rect 20536 17323 20588 17332
rect 20536 17289 20545 17323
rect 20545 17289 20579 17323
rect 20579 17289 20588 17323
rect 20536 17280 20588 17289
rect 20628 17280 20680 17332
rect 24768 17280 24820 17332
rect 18328 17187 18380 17196
rect 18328 17153 18337 17187
rect 18337 17153 18371 17187
rect 18371 17153 18380 17187
rect 18328 17144 18380 17153
rect 22008 17212 22060 17264
rect 22468 17212 22520 17264
rect 24676 17212 24728 17264
rect 22560 17187 22612 17196
rect 22560 17153 22569 17187
rect 22569 17153 22603 17187
rect 22603 17153 22612 17187
rect 22560 17144 22612 17153
rect 24860 17187 24912 17196
rect 24860 17153 24869 17187
rect 24869 17153 24903 17187
rect 24903 17153 24912 17187
rect 24860 17144 24912 17153
rect 21088 17076 21140 17128
rect 23480 17076 23532 17128
rect 20168 17008 20220 17060
rect 22468 17008 22520 17060
rect 23940 17008 23992 17060
rect 19616 16940 19668 16992
rect 25044 16940 25096 16992
rect 2950 16838 3002 16890
rect 3014 16838 3066 16890
rect 3078 16838 3130 16890
rect 3142 16838 3194 16890
rect 3206 16838 3258 16890
rect 12950 16838 13002 16890
rect 13014 16838 13066 16890
rect 13078 16838 13130 16890
rect 13142 16838 13194 16890
rect 13206 16838 13258 16890
rect 22950 16838 23002 16890
rect 23014 16838 23066 16890
rect 23078 16838 23130 16890
rect 23142 16838 23194 16890
rect 23206 16838 23258 16890
rect 7288 16779 7340 16788
rect 7288 16745 7297 16779
rect 7297 16745 7331 16779
rect 7331 16745 7340 16779
rect 7288 16736 7340 16745
rect 8392 16779 8444 16788
rect 8392 16745 8401 16779
rect 8401 16745 8435 16779
rect 8435 16745 8444 16779
rect 8392 16736 8444 16745
rect 9312 16736 9364 16788
rect 9588 16736 9640 16788
rect 9772 16736 9824 16788
rect 10692 16736 10744 16788
rect 3424 16668 3476 16720
rect 11152 16668 11204 16720
rect 6920 16643 6972 16652
rect 6920 16609 6929 16643
rect 6929 16609 6963 16643
rect 6963 16609 6972 16643
rect 6920 16600 6972 16609
rect 9128 16600 9180 16652
rect 9956 16600 10008 16652
rect 4160 16575 4212 16584
rect 4160 16541 4169 16575
rect 4169 16541 4203 16575
rect 4203 16541 4212 16575
rect 4160 16532 4212 16541
rect 7380 16532 7432 16584
rect 7932 16575 7984 16584
rect 7932 16541 7941 16575
rect 7941 16541 7975 16575
rect 7975 16541 7984 16575
rect 7932 16532 7984 16541
rect 8576 16575 8628 16584
rect 8576 16541 8585 16575
rect 8585 16541 8619 16575
rect 8619 16541 8628 16575
rect 8576 16532 8628 16541
rect 9588 16532 9640 16584
rect 11060 16600 11112 16652
rect 15016 16736 15068 16788
rect 16028 16779 16080 16788
rect 16028 16745 16037 16779
rect 16037 16745 16071 16779
rect 16071 16745 16080 16779
rect 16028 16736 16080 16745
rect 16120 16736 16172 16788
rect 17868 16736 17920 16788
rect 10876 16532 10928 16584
rect 9404 16396 9456 16448
rect 11060 16464 11112 16516
rect 12256 16643 12308 16652
rect 12256 16609 12265 16643
rect 12265 16609 12299 16643
rect 12299 16609 12308 16643
rect 12256 16600 12308 16609
rect 14924 16600 14976 16652
rect 15016 16600 15068 16652
rect 16856 16600 16908 16652
rect 17132 16643 17184 16652
rect 17132 16609 17141 16643
rect 17141 16609 17175 16643
rect 17175 16609 17184 16643
rect 17132 16600 17184 16609
rect 19432 16736 19484 16788
rect 20720 16736 20772 16788
rect 21088 16736 21140 16788
rect 21364 16736 21416 16788
rect 22560 16779 22612 16788
rect 22560 16745 22590 16779
rect 22590 16745 22612 16779
rect 22560 16736 22612 16745
rect 21548 16668 21600 16720
rect 22560 16600 22612 16652
rect 23756 16600 23808 16652
rect 11704 16532 11756 16584
rect 12256 16464 12308 16516
rect 12716 16464 12768 16516
rect 14556 16507 14608 16516
rect 14556 16473 14565 16507
rect 14565 16473 14599 16507
rect 14599 16473 14608 16507
rect 14556 16464 14608 16473
rect 16304 16464 16356 16516
rect 21088 16532 21140 16584
rect 24400 16532 24452 16584
rect 24768 16532 24820 16584
rect 16856 16464 16908 16516
rect 17684 16464 17736 16516
rect 9680 16396 9732 16448
rect 10048 16396 10100 16448
rect 10140 16439 10192 16448
rect 10140 16405 10149 16439
rect 10149 16405 10183 16439
rect 10183 16405 10192 16439
rect 10140 16396 10192 16405
rect 10784 16439 10836 16448
rect 10784 16405 10793 16439
rect 10793 16405 10827 16439
rect 10827 16405 10836 16439
rect 10784 16396 10836 16405
rect 12348 16396 12400 16448
rect 16488 16439 16540 16448
rect 16488 16405 16497 16439
rect 16497 16405 16531 16439
rect 16531 16405 16540 16439
rect 16488 16396 16540 16405
rect 16672 16396 16724 16448
rect 17592 16396 17644 16448
rect 18328 16396 18380 16448
rect 18880 16439 18932 16448
rect 18880 16405 18889 16439
rect 18889 16405 18923 16439
rect 18923 16405 18932 16439
rect 18880 16396 18932 16405
rect 22008 16464 22060 16516
rect 22192 16464 22244 16516
rect 22652 16464 22704 16516
rect 23848 16396 23900 16448
rect 23940 16396 23992 16448
rect 7950 16294 8002 16346
rect 8014 16294 8066 16346
rect 8078 16294 8130 16346
rect 8142 16294 8194 16346
rect 8206 16294 8258 16346
rect 17950 16294 18002 16346
rect 18014 16294 18066 16346
rect 18078 16294 18130 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 4160 16192 4212 16244
rect 8760 16192 8812 16244
rect 9220 16192 9272 16244
rect 5632 16124 5684 16176
rect 9312 16099 9364 16108
rect 9312 16065 9321 16099
rect 9321 16065 9355 16099
rect 9355 16065 9364 16099
rect 9312 16056 9364 16065
rect 9588 15988 9640 16040
rect 9956 16099 10008 16108
rect 9956 16065 9965 16099
rect 9965 16065 9999 16099
rect 9999 16065 10008 16099
rect 9956 16056 10008 16065
rect 10140 16192 10192 16244
rect 15568 16192 15620 16244
rect 12716 16124 12768 16176
rect 15752 16124 15804 16176
rect 11428 16056 11480 16108
rect 13912 16056 13964 16108
rect 16304 16192 16356 16244
rect 16856 16192 16908 16244
rect 17776 16192 17828 16244
rect 18512 16192 18564 16244
rect 19064 16192 19116 16244
rect 20628 16192 20680 16244
rect 20904 16235 20956 16244
rect 20904 16201 20913 16235
rect 20913 16201 20947 16235
rect 20947 16201 20956 16235
rect 20904 16192 20956 16201
rect 21088 16192 21140 16244
rect 21640 16192 21692 16244
rect 22284 16192 22336 16244
rect 24400 16192 24452 16244
rect 17224 16124 17276 16176
rect 18972 16056 19024 16108
rect 19064 16056 19116 16108
rect 20628 16056 20680 16108
rect 10784 15988 10836 16040
rect 11060 16031 11112 16040
rect 11060 15997 11069 16031
rect 11069 15997 11103 16031
rect 11103 15997 11112 16031
rect 11060 15988 11112 15997
rect 11704 16031 11756 16040
rect 11704 15997 11713 16031
rect 11713 15997 11747 16031
rect 11747 15997 11756 16031
rect 11704 15988 11756 15997
rect 12348 15988 12400 16040
rect 12716 15988 12768 16040
rect 7472 15920 7524 15972
rect 8484 15895 8536 15904
rect 8484 15861 8493 15895
rect 8493 15861 8527 15895
rect 8527 15861 8536 15895
rect 8484 15852 8536 15861
rect 9128 15963 9180 15972
rect 9128 15929 9137 15963
rect 9137 15929 9171 15963
rect 9171 15929 9180 15963
rect 9128 15920 9180 15929
rect 9772 15963 9824 15972
rect 9772 15929 9781 15963
rect 9781 15929 9815 15963
rect 9815 15929 9824 15963
rect 9772 15920 9824 15929
rect 13452 16031 13504 16040
rect 13452 15997 13461 16031
rect 13461 15997 13495 16031
rect 13495 15997 13504 16031
rect 13452 15988 13504 15997
rect 14096 15988 14148 16040
rect 14556 16031 14608 16040
rect 14556 15997 14565 16031
rect 14565 15997 14599 16031
rect 14599 15997 14608 16031
rect 14556 15988 14608 15997
rect 15844 15988 15896 16040
rect 16028 16031 16080 16040
rect 16028 15997 16037 16031
rect 16037 15997 16071 16031
rect 16071 15997 16080 16031
rect 16028 15988 16080 15997
rect 16304 15988 16356 16040
rect 13544 15852 13596 15904
rect 15108 15852 15160 15904
rect 15384 15852 15436 15904
rect 16028 15852 16080 15904
rect 20260 15988 20312 16040
rect 21088 16031 21140 16040
rect 21088 15997 21097 16031
rect 21097 15997 21131 16031
rect 21131 15997 21140 16031
rect 21088 15988 21140 15997
rect 23848 16124 23900 16176
rect 22284 16056 22336 16108
rect 24124 16056 24176 16108
rect 24676 16099 24728 16108
rect 24676 16065 24685 16099
rect 24685 16065 24719 16099
rect 24719 16065 24728 16099
rect 24676 16056 24728 16065
rect 22652 16031 22704 16040
rect 22652 15997 22661 16031
rect 22661 15997 22695 16031
rect 22695 15997 22704 16031
rect 22652 15988 22704 15997
rect 22836 15988 22888 16040
rect 23940 16031 23992 16040
rect 23940 15997 23949 16031
rect 23949 15997 23983 16031
rect 23983 15997 23992 16031
rect 23940 15988 23992 15997
rect 25872 15988 25924 16040
rect 26240 15988 26292 16040
rect 24952 15920 25004 15972
rect 16488 15852 16540 15904
rect 20352 15852 20404 15904
rect 20536 15895 20588 15904
rect 20536 15861 20545 15895
rect 20545 15861 20579 15895
rect 20579 15861 20588 15895
rect 20536 15852 20588 15861
rect 22192 15852 22244 15904
rect 23296 15852 23348 15904
rect 2950 15750 3002 15802
rect 3014 15750 3066 15802
rect 3078 15750 3130 15802
rect 3142 15750 3194 15802
rect 3206 15750 3258 15802
rect 12950 15750 13002 15802
rect 13014 15750 13066 15802
rect 13078 15750 13130 15802
rect 13142 15750 13194 15802
rect 13206 15750 13258 15802
rect 22950 15750 23002 15802
rect 23014 15750 23066 15802
rect 23078 15750 23130 15802
rect 23142 15750 23194 15802
rect 23206 15750 23258 15802
rect 9864 15691 9916 15700
rect 9864 15657 9873 15691
rect 9873 15657 9907 15691
rect 9907 15657 9916 15691
rect 9864 15648 9916 15657
rect 10968 15648 11020 15700
rect 11152 15648 11204 15700
rect 12256 15623 12308 15632
rect 12256 15589 12265 15623
rect 12265 15589 12299 15623
rect 12299 15589 12308 15623
rect 12256 15580 12308 15589
rect 13452 15648 13504 15700
rect 14004 15648 14056 15700
rect 15016 15648 15068 15700
rect 15200 15648 15252 15700
rect 16672 15691 16724 15700
rect 16672 15657 16681 15691
rect 16681 15657 16715 15691
rect 16715 15657 16724 15691
rect 16672 15648 16724 15657
rect 18604 15648 18656 15700
rect 19340 15648 19392 15700
rect 16856 15580 16908 15632
rect 19248 15580 19300 15632
rect 21180 15580 21232 15632
rect 14188 15512 14240 15564
rect 14280 15555 14332 15564
rect 14280 15521 14289 15555
rect 14289 15521 14323 15555
rect 14323 15521 14332 15555
rect 14280 15512 14332 15521
rect 8760 15487 8812 15496
rect 8760 15453 8769 15487
rect 8769 15453 8803 15487
rect 8803 15453 8812 15487
rect 8760 15444 8812 15453
rect 9404 15487 9456 15496
rect 9404 15453 9413 15487
rect 9413 15453 9447 15487
rect 9447 15453 9456 15487
rect 9404 15444 9456 15453
rect 10232 15444 10284 15496
rect 13820 15444 13872 15496
rect 18880 15512 18932 15564
rect 20168 15512 20220 15564
rect 21364 15555 21416 15564
rect 21364 15521 21373 15555
rect 21373 15521 21407 15555
rect 21407 15521 21416 15555
rect 21364 15512 21416 15521
rect 16856 15444 16908 15496
rect 19984 15487 20036 15496
rect 19984 15453 19993 15487
rect 19993 15453 20027 15487
rect 20027 15453 20036 15487
rect 19984 15444 20036 15453
rect 10692 15376 10744 15428
rect 12716 15376 12768 15428
rect 7564 15308 7616 15360
rect 11152 15308 11204 15360
rect 11428 15308 11480 15360
rect 13544 15376 13596 15428
rect 15108 15376 15160 15428
rect 16212 15308 16264 15360
rect 17684 15376 17736 15428
rect 21640 15376 21692 15428
rect 22008 15487 22060 15496
rect 22008 15453 22019 15487
rect 22019 15453 22053 15487
rect 22053 15453 22060 15487
rect 22008 15444 22060 15453
rect 22652 15444 22704 15496
rect 24860 15648 24912 15700
rect 19708 15308 19760 15360
rect 21272 15308 21324 15360
rect 22652 15308 22704 15360
rect 23204 15376 23256 15428
rect 25412 15444 25464 15496
rect 24860 15419 24912 15428
rect 24860 15385 24869 15419
rect 24869 15385 24903 15419
rect 24903 15385 24912 15419
rect 24860 15376 24912 15385
rect 25044 15419 25096 15428
rect 25044 15385 25053 15419
rect 25053 15385 25087 15419
rect 25087 15385 25096 15419
rect 25044 15376 25096 15385
rect 7950 15206 8002 15258
rect 8014 15206 8066 15258
rect 8078 15206 8130 15258
rect 8142 15206 8194 15258
rect 8206 15206 8258 15258
rect 17950 15206 18002 15258
rect 18014 15206 18066 15258
rect 18078 15206 18130 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 9404 15147 9456 15156
rect 9404 15113 9413 15147
rect 9413 15113 9447 15147
rect 9447 15113 9456 15147
rect 9404 15104 9456 15113
rect 10232 15104 10284 15156
rect 10968 15147 11020 15156
rect 10968 15113 10977 15147
rect 10977 15113 11011 15147
rect 11011 15113 11020 15147
rect 10968 15104 11020 15113
rect 11060 15104 11112 15156
rect 12072 15104 12124 15156
rect 13912 15147 13964 15156
rect 13912 15113 13921 15147
rect 13921 15113 13955 15147
rect 13955 15113 13964 15147
rect 13912 15104 13964 15113
rect 15292 15147 15344 15156
rect 15292 15113 15301 15147
rect 15301 15113 15335 15147
rect 15335 15113 15344 15147
rect 15292 15104 15344 15113
rect 12716 15036 12768 15088
rect 10508 15011 10560 15020
rect 10508 14977 10517 15011
rect 10517 14977 10551 15011
rect 10551 14977 10560 15011
rect 10508 14968 10560 14977
rect 11152 15011 11204 15020
rect 11152 14977 11161 15011
rect 11161 14977 11195 15011
rect 11195 14977 11204 15011
rect 11152 14968 11204 14977
rect 17040 15104 17092 15156
rect 18604 15104 18656 15156
rect 18972 15147 19024 15156
rect 18972 15113 18981 15147
rect 18981 15113 19015 15147
rect 19015 15113 19024 15147
rect 18972 15104 19024 15113
rect 20628 15104 20680 15156
rect 21456 15147 21508 15156
rect 21456 15113 21465 15147
rect 21465 15113 21499 15147
rect 21499 15113 21508 15147
rect 21456 15104 21508 15113
rect 17684 15036 17736 15088
rect 20904 15036 20956 15088
rect 22100 15104 22152 15156
rect 23940 15104 23992 15156
rect 24492 15104 24544 15156
rect 23756 15036 23808 15088
rect 10692 14900 10744 14952
rect 11704 14943 11756 14952
rect 11704 14909 11713 14943
rect 11713 14909 11747 14943
rect 11747 14909 11756 14943
rect 11704 14900 11756 14909
rect 12440 14900 12492 14952
rect 15384 14900 15436 14952
rect 16120 14943 16172 14952
rect 16120 14909 16129 14943
rect 16129 14909 16163 14943
rect 16163 14909 16172 14943
rect 16120 14900 16172 14909
rect 10048 14807 10100 14816
rect 10048 14773 10057 14807
rect 10057 14773 10091 14807
rect 10091 14773 10100 14807
rect 10048 14764 10100 14773
rect 14096 14832 14148 14884
rect 14740 14832 14792 14884
rect 16488 14900 16540 14952
rect 16672 14832 16724 14884
rect 16488 14764 16540 14816
rect 17868 14900 17920 14952
rect 18880 14968 18932 15020
rect 19340 14943 19392 14952
rect 17132 14764 17184 14816
rect 19340 14909 19349 14943
rect 19349 14909 19383 14943
rect 19383 14909 19392 14943
rect 19340 14900 19392 14909
rect 21272 14900 21324 14952
rect 18880 14832 18932 14884
rect 22560 14900 22612 14952
rect 18604 14807 18656 14816
rect 18604 14773 18613 14807
rect 18613 14773 18647 14807
rect 18647 14773 18656 14807
rect 18604 14764 18656 14773
rect 22468 14832 22520 14884
rect 22744 14832 22796 14884
rect 2950 14662 3002 14714
rect 3014 14662 3066 14714
rect 3078 14662 3130 14714
rect 3142 14662 3194 14714
rect 3206 14662 3258 14714
rect 12950 14662 13002 14714
rect 13014 14662 13066 14714
rect 13078 14662 13130 14714
rect 13142 14662 13194 14714
rect 13206 14662 13258 14714
rect 22950 14662 23002 14714
rect 23014 14662 23066 14714
rect 23078 14662 23130 14714
rect 23142 14662 23194 14714
rect 23206 14662 23258 14714
rect 10508 14560 10560 14612
rect 11152 14560 11204 14612
rect 12256 14424 12308 14476
rect 10692 14399 10744 14408
rect 10692 14365 10701 14399
rect 10701 14365 10735 14399
rect 10735 14365 10744 14399
rect 10692 14356 10744 14365
rect 12440 14603 12492 14612
rect 12440 14569 12449 14603
rect 12449 14569 12483 14603
rect 12483 14569 12492 14603
rect 12440 14560 12492 14569
rect 13360 14560 13412 14612
rect 15936 14560 15988 14612
rect 16120 14560 16172 14612
rect 16212 14492 16264 14544
rect 18696 14492 18748 14544
rect 19984 14560 20036 14612
rect 20260 14560 20312 14612
rect 20904 14560 20956 14612
rect 22100 14560 22152 14612
rect 22560 14560 22612 14612
rect 23756 14560 23808 14612
rect 25136 14560 25188 14612
rect 26148 14560 26200 14612
rect 14280 14467 14332 14476
rect 14280 14433 14289 14467
rect 14289 14433 14323 14467
rect 14323 14433 14332 14467
rect 14280 14424 14332 14433
rect 14556 14467 14608 14476
rect 14556 14433 14565 14467
rect 14565 14433 14599 14467
rect 14599 14433 14608 14467
rect 14556 14424 14608 14433
rect 18604 14424 18656 14476
rect 14004 14356 14056 14408
rect 16488 14399 16540 14408
rect 16488 14365 16497 14399
rect 16497 14365 16531 14399
rect 16531 14365 16540 14399
rect 16488 14356 16540 14365
rect 19892 14399 19944 14408
rect 19892 14365 19901 14399
rect 19901 14365 19935 14399
rect 19935 14365 19944 14399
rect 19892 14356 19944 14365
rect 10048 14220 10100 14272
rect 14096 14288 14148 14340
rect 15016 14288 15068 14340
rect 16672 14288 16724 14340
rect 20536 14492 20588 14544
rect 25596 14492 25648 14544
rect 23388 14424 23440 14476
rect 23572 14424 23624 14476
rect 24584 14424 24636 14476
rect 25228 14424 25280 14476
rect 20536 14356 20588 14408
rect 21456 14356 21508 14408
rect 12716 14220 12768 14272
rect 13636 14220 13688 14272
rect 16764 14220 16816 14272
rect 18604 14220 18656 14272
rect 19156 14220 19208 14272
rect 20628 14288 20680 14340
rect 22560 14331 22612 14340
rect 22560 14297 22569 14331
rect 22569 14297 22603 14331
rect 22603 14297 22612 14331
rect 22560 14288 22612 14297
rect 22836 14288 22888 14340
rect 23664 14356 23716 14408
rect 25596 14356 25648 14408
rect 25872 14356 25924 14408
rect 23664 14263 23716 14272
rect 23664 14229 23673 14263
rect 23673 14229 23707 14263
rect 23707 14229 23716 14263
rect 23664 14220 23716 14229
rect 24308 14220 24360 14272
rect 7950 14118 8002 14170
rect 8014 14118 8066 14170
rect 8078 14118 8130 14170
rect 8142 14118 8194 14170
rect 8206 14118 8258 14170
rect 17950 14118 18002 14170
rect 18014 14118 18066 14170
rect 18078 14118 18130 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 11796 14059 11848 14068
rect 11796 14025 11805 14059
rect 11805 14025 11839 14059
rect 11839 14025 11848 14059
rect 11796 14016 11848 14025
rect 12532 14016 12584 14068
rect 13636 14016 13688 14068
rect 13728 14016 13780 14068
rect 11980 13923 12032 13932
rect 11980 13889 11989 13923
rect 11989 13889 12023 13923
rect 12023 13889 12032 13923
rect 11980 13880 12032 13889
rect 13544 13948 13596 14000
rect 14280 13948 14332 14000
rect 14648 14016 14700 14068
rect 16396 14016 16448 14068
rect 17500 14059 17552 14068
rect 17500 14025 17509 14059
rect 17509 14025 17543 14059
rect 17543 14025 17552 14059
rect 17500 14016 17552 14025
rect 15016 13880 15068 13932
rect 14004 13812 14056 13864
rect 14372 13812 14424 13864
rect 17408 13923 17460 13932
rect 17408 13889 17417 13923
rect 17417 13889 17451 13923
rect 17451 13889 17460 13923
rect 17408 13880 17460 13889
rect 16672 13855 16724 13864
rect 16672 13821 16681 13855
rect 16681 13821 16715 13855
rect 16715 13821 16724 13855
rect 16672 13812 16724 13821
rect 17592 13855 17644 13864
rect 17592 13821 17601 13855
rect 17601 13821 17635 13855
rect 17635 13821 17644 13855
rect 17592 13812 17644 13821
rect 15568 13744 15620 13796
rect 18512 13948 18564 14000
rect 19340 14016 19392 14068
rect 20260 14059 20312 14068
rect 20260 14025 20269 14059
rect 20269 14025 20303 14059
rect 20303 14025 20312 14059
rect 20260 14016 20312 14025
rect 20444 14016 20496 14068
rect 20076 13948 20128 14000
rect 22744 14016 22796 14068
rect 19432 13880 19484 13932
rect 23388 13948 23440 14000
rect 23756 13948 23808 14000
rect 25136 13991 25188 14000
rect 25136 13957 25145 13991
rect 25145 13957 25179 13991
rect 25179 13957 25188 13991
rect 25136 13948 25188 13957
rect 22560 13880 22612 13932
rect 19248 13812 19300 13864
rect 20260 13812 20312 13864
rect 21272 13855 21324 13864
rect 21272 13821 21281 13855
rect 21281 13821 21315 13855
rect 21315 13821 21324 13855
rect 21272 13812 21324 13821
rect 22284 13855 22336 13864
rect 22284 13821 22293 13855
rect 22293 13821 22327 13855
rect 22327 13821 22336 13855
rect 22284 13812 22336 13821
rect 24492 13812 24544 13864
rect 24584 13855 24636 13864
rect 24584 13821 24593 13855
rect 24593 13821 24627 13855
rect 24627 13821 24636 13855
rect 24584 13812 24636 13821
rect 25872 13812 25924 13864
rect 15200 13676 15252 13728
rect 17040 13719 17092 13728
rect 17040 13685 17049 13719
rect 17049 13685 17083 13719
rect 17083 13685 17092 13719
rect 17040 13676 17092 13685
rect 19892 13676 19944 13728
rect 20076 13676 20128 13728
rect 20720 13719 20772 13728
rect 20720 13685 20729 13719
rect 20729 13685 20763 13719
rect 20763 13685 20772 13719
rect 20720 13676 20772 13685
rect 2950 13574 3002 13626
rect 3014 13574 3066 13626
rect 3078 13574 3130 13626
rect 3142 13574 3194 13626
rect 3206 13574 3258 13626
rect 12950 13574 13002 13626
rect 13014 13574 13066 13626
rect 13078 13574 13130 13626
rect 13142 13574 13194 13626
rect 13206 13574 13258 13626
rect 22950 13574 23002 13626
rect 23014 13574 23066 13626
rect 23078 13574 23130 13626
rect 23142 13574 23194 13626
rect 23206 13574 23258 13626
rect 12716 13472 12768 13524
rect 13728 13472 13780 13524
rect 15200 13472 15252 13524
rect 16304 13472 16356 13524
rect 16580 13472 16632 13524
rect 19064 13472 19116 13524
rect 13360 13404 13412 13456
rect 12072 13379 12124 13388
rect 12072 13345 12081 13379
rect 12081 13345 12115 13379
rect 12115 13345 12124 13379
rect 12072 13336 12124 13345
rect 14280 13379 14332 13388
rect 14280 13345 14289 13379
rect 14289 13345 14323 13379
rect 14323 13345 14332 13379
rect 14280 13336 14332 13345
rect 16488 13379 16540 13388
rect 16488 13345 16497 13379
rect 16497 13345 16531 13379
rect 16531 13345 16540 13379
rect 16488 13336 16540 13345
rect 18696 13336 18748 13388
rect 19616 13472 19668 13524
rect 20536 13472 20588 13524
rect 21272 13472 21324 13524
rect 23204 13472 23256 13524
rect 23480 13472 23532 13524
rect 23756 13404 23808 13456
rect 21916 13379 21968 13388
rect 11520 13200 11572 13252
rect 10048 13132 10100 13184
rect 10692 13132 10744 13184
rect 19432 13268 19484 13320
rect 21916 13345 21925 13379
rect 21925 13345 21959 13379
rect 21959 13345 21968 13379
rect 21916 13336 21968 13345
rect 22652 13336 22704 13388
rect 22836 13336 22888 13388
rect 23204 13336 23256 13388
rect 25320 13268 25372 13320
rect 12716 13200 12768 13252
rect 14188 13200 14240 13252
rect 14556 13243 14608 13252
rect 14556 13209 14565 13243
rect 14565 13209 14599 13243
rect 14599 13209 14608 13243
rect 14556 13200 14608 13209
rect 13728 13132 13780 13184
rect 15016 13200 15068 13252
rect 16488 13200 16540 13252
rect 17224 13200 17276 13252
rect 19892 13200 19944 13252
rect 16304 13132 16356 13184
rect 17592 13132 17644 13184
rect 20260 13200 20312 13252
rect 23756 13200 23808 13252
rect 24032 13200 24084 13252
rect 20812 13132 20864 13184
rect 24492 13132 24544 13184
rect 7950 13030 8002 13082
rect 8014 13030 8066 13082
rect 8078 13030 8130 13082
rect 8142 13030 8194 13082
rect 8206 13030 8258 13082
rect 17950 13030 18002 13082
rect 18014 13030 18066 13082
rect 18078 13030 18130 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 11520 12971 11572 12980
rect 11520 12937 11529 12971
rect 11529 12937 11563 12971
rect 11563 12937 11572 12971
rect 11520 12928 11572 12937
rect 12716 12928 12768 12980
rect 13820 12928 13872 12980
rect 14280 12971 14332 12980
rect 14280 12937 14289 12971
rect 14289 12937 14323 12971
rect 14323 12937 14332 12971
rect 14280 12928 14332 12937
rect 15016 12928 15068 12980
rect 16488 12928 16540 12980
rect 15568 12860 15620 12912
rect 17868 12928 17920 12980
rect 18696 12928 18748 12980
rect 19524 12928 19576 12980
rect 21456 12928 21508 12980
rect 23204 12928 23256 12980
rect 25688 12928 25740 12980
rect 17224 12860 17276 12912
rect 17592 12860 17644 12912
rect 18788 12860 18840 12912
rect 22376 12860 22428 12912
rect 25964 12860 26016 12912
rect 16856 12835 16908 12844
rect 16856 12801 16865 12835
rect 16865 12801 16899 12835
rect 16899 12801 16908 12835
rect 16856 12792 16908 12801
rect 18512 12792 18564 12844
rect 20628 12835 20680 12844
rect 20628 12801 20637 12835
rect 20637 12801 20671 12835
rect 20671 12801 20680 12835
rect 20628 12792 20680 12801
rect 15200 12767 15252 12776
rect 15200 12733 15209 12767
rect 15209 12733 15243 12767
rect 15243 12733 15252 12767
rect 15200 12724 15252 12733
rect 16672 12724 16724 12776
rect 17592 12724 17644 12776
rect 17868 12724 17920 12776
rect 18420 12724 18472 12776
rect 18604 12699 18656 12708
rect 18604 12665 18613 12699
rect 18613 12665 18647 12699
rect 18647 12665 18656 12699
rect 20260 12724 20312 12776
rect 21916 12792 21968 12844
rect 23756 12792 23808 12844
rect 24216 12835 24268 12844
rect 24216 12801 24225 12835
rect 24225 12801 24259 12835
rect 24259 12801 24268 12835
rect 24216 12792 24268 12801
rect 24400 12792 24452 12844
rect 18604 12656 18656 12665
rect 20444 12656 20496 12708
rect 20996 12724 21048 12776
rect 21548 12724 21600 12776
rect 22284 12767 22336 12776
rect 22284 12733 22293 12767
rect 22293 12733 22327 12767
rect 22327 12733 22336 12767
rect 22284 12724 22336 12733
rect 23480 12656 23532 12708
rect 19800 12588 19852 12640
rect 20260 12631 20312 12640
rect 20260 12597 20269 12631
rect 20269 12597 20303 12631
rect 20303 12597 20312 12631
rect 20260 12588 20312 12597
rect 2950 12486 3002 12538
rect 3014 12486 3066 12538
rect 3078 12486 3130 12538
rect 3142 12486 3194 12538
rect 3206 12486 3258 12538
rect 12950 12486 13002 12538
rect 13014 12486 13066 12538
rect 13078 12486 13130 12538
rect 13142 12486 13194 12538
rect 13206 12486 13258 12538
rect 22950 12486 23002 12538
rect 23014 12486 23066 12538
rect 23078 12486 23130 12538
rect 23142 12486 23194 12538
rect 23206 12486 23258 12538
rect 4068 12384 4120 12436
rect 8576 12384 8628 12436
rect 13728 12427 13780 12436
rect 13728 12393 13737 12427
rect 13737 12393 13771 12427
rect 13771 12393 13780 12427
rect 13728 12384 13780 12393
rect 14004 12384 14056 12436
rect 15568 12384 15620 12436
rect 17592 12384 17644 12436
rect 22744 12384 22796 12436
rect 24216 12316 24268 12368
rect 16764 12248 16816 12300
rect 17408 12248 17460 12300
rect 19800 12248 19852 12300
rect 20444 12248 20496 12300
rect 21364 12248 21416 12300
rect 21916 12248 21968 12300
rect 24584 12248 24636 12300
rect 15568 12180 15620 12232
rect 19340 12180 19392 12232
rect 16304 12112 16356 12164
rect 16488 12112 16540 12164
rect 19616 12112 19668 12164
rect 19708 12155 19760 12164
rect 19708 12121 19717 12155
rect 19717 12121 19751 12155
rect 19751 12121 19760 12155
rect 19708 12112 19760 12121
rect 20168 12112 20220 12164
rect 19984 12044 20036 12096
rect 20628 12044 20680 12096
rect 24216 12112 24268 12164
rect 22376 12044 22428 12096
rect 7950 11942 8002 11994
rect 8014 11942 8066 11994
rect 8078 11942 8130 11994
rect 8142 11942 8194 11994
rect 8206 11942 8258 11994
rect 17950 11942 18002 11994
rect 18014 11942 18066 11994
rect 18078 11942 18130 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 13820 11840 13872 11892
rect 14556 11883 14608 11892
rect 14556 11849 14565 11883
rect 14565 11849 14599 11883
rect 14599 11849 14608 11883
rect 14556 11840 14608 11849
rect 13360 11772 13412 11824
rect 13728 11772 13780 11824
rect 15752 11840 15804 11892
rect 16764 11704 16816 11756
rect 16856 11636 16908 11688
rect 19340 11840 19392 11892
rect 17684 11772 17736 11824
rect 19156 11772 19208 11824
rect 19800 11772 19852 11824
rect 20168 11772 20220 11824
rect 24860 11772 24912 11824
rect 25136 11815 25188 11824
rect 25136 11781 25145 11815
rect 25145 11781 25179 11815
rect 25179 11781 25188 11815
rect 25136 11772 25188 11781
rect 19432 11747 19484 11756
rect 19432 11713 19441 11747
rect 19441 11713 19475 11747
rect 19475 11713 19484 11747
rect 19432 11704 19484 11713
rect 22192 11747 22244 11756
rect 22192 11713 22201 11747
rect 22201 11713 22235 11747
rect 22235 11713 22244 11747
rect 22192 11704 22244 11713
rect 18604 11636 18656 11688
rect 14464 11568 14516 11620
rect 18512 11568 18564 11620
rect 20904 11636 20956 11688
rect 20812 11568 20864 11620
rect 21088 11568 21140 11620
rect 21640 11568 21692 11620
rect 14648 11500 14700 11552
rect 16764 11543 16816 11552
rect 16764 11509 16773 11543
rect 16773 11509 16807 11543
rect 16807 11509 16816 11543
rect 16764 11500 16816 11509
rect 18788 11500 18840 11552
rect 19708 11500 19760 11552
rect 21272 11500 21324 11552
rect 21548 11500 21600 11552
rect 24492 11500 24544 11552
rect 2950 11398 3002 11450
rect 3014 11398 3066 11450
rect 3078 11398 3130 11450
rect 3142 11398 3194 11450
rect 3206 11398 3258 11450
rect 12950 11398 13002 11450
rect 13014 11398 13066 11450
rect 13078 11398 13130 11450
rect 13142 11398 13194 11450
rect 13206 11398 13258 11450
rect 22950 11398 23002 11450
rect 23014 11398 23066 11450
rect 23078 11398 23130 11450
rect 23142 11398 23194 11450
rect 23206 11398 23258 11450
rect 12532 11296 12584 11348
rect 13728 11296 13780 11348
rect 14648 11339 14700 11348
rect 14648 11305 14657 11339
rect 14657 11305 14691 11339
rect 14691 11305 14700 11339
rect 14648 11296 14700 11305
rect 15476 11339 15528 11348
rect 15476 11305 15485 11339
rect 15485 11305 15519 11339
rect 15519 11305 15528 11339
rect 15476 11296 15528 11305
rect 16120 11339 16172 11348
rect 16120 11305 16129 11339
rect 16129 11305 16163 11339
rect 16163 11305 16172 11339
rect 16120 11296 16172 11305
rect 16948 11296 17000 11348
rect 17500 11296 17552 11348
rect 19248 11339 19300 11348
rect 19248 11305 19257 11339
rect 19257 11305 19291 11339
rect 19291 11305 19300 11339
rect 19248 11296 19300 11305
rect 19524 11339 19576 11348
rect 19524 11305 19533 11339
rect 19533 11305 19567 11339
rect 19567 11305 19576 11339
rect 19524 11296 19576 11305
rect 19616 11296 19668 11348
rect 20812 11339 20864 11348
rect 20812 11305 20821 11339
rect 20821 11305 20855 11339
rect 20855 11305 20864 11339
rect 20812 11296 20864 11305
rect 23388 11296 23440 11348
rect 24584 11339 24636 11348
rect 24584 11305 24593 11339
rect 24593 11305 24627 11339
rect 24627 11305 24636 11339
rect 24584 11296 24636 11305
rect 24768 11296 24820 11348
rect 25688 11296 25740 11348
rect 19800 11228 19852 11280
rect 20260 11228 20312 11280
rect 22376 11228 22428 11280
rect 22652 11228 22704 11280
rect 25964 11228 26016 11280
rect 18420 11160 18472 11212
rect 15660 11135 15712 11144
rect 15660 11101 15669 11135
rect 15669 11101 15703 11135
rect 15703 11101 15712 11135
rect 15660 11092 15712 11101
rect 16028 11092 16080 11144
rect 17132 11092 17184 11144
rect 18512 11092 18564 11144
rect 21548 11160 21600 11212
rect 24860 11160 24912 11212
rect 19156 11092 19208 11144
rect 20076 11092 20128 11144
rect 22284 11092 22336 11144
rect 22652 11135 22704 11144
rect 22652 11101 22661 11135
rect 22661 11101 22695 11135
rect 22695 11101 22704 11135
rect 22652 11092 22704 11101
rect 24768 11135 24820 11144
rect 24768 11101 24777 11135
rect 24777 11101 24811 11135
rect 24811 11101 24820 11135
rect 24768 11092 24820 11101
rect 15568 11024 15620 11076
rect 23940 11024 23992 11076
rect 20076 10999 20128 11008
rect 20076 10965 20085 10999
rect 20085 10965 20119 10999
rect 20119 10965 20128 10999
rect 20076 10956 20128 10965
rect 20168 10956 20220 11008
rect 21088 10956 21140 11008
rect 21272 10956 21324 11008
rect 21732 10956 21784 11008
rect 7950 10854 8002 10906
rect 8014 10854 8066 10906
rect 8078 10854 8130 10906
rect 8142 10854 8194 10906
rect 8206 10854 8258 10906
rect 17950 10854 18002 10906
rect 18014 10854 18066 10906
rect 18078 10854 18130 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 15660 10752 15712 10804
rect 16028 10752 16080 10804
rect 17132 10795 17184 10804
rect 17132 10761 17141 10795
rect 17141 10761 17175 10795
rect 17175 10761 17184 10795
rect 17132 10752 17184 10761
rect 17868 10752 17920 10804
rect 18328 10752 18380 10804
rect 20996 10752 21048 10804
rect 21088 10752 21140 10804
rect 21916 10752 21968 10804
rect 18696 10616 18748 10668
rect 20536 10684 20588 10736
rect 20168 10659 20220 10668
rect 20168 10625 20177 10659
rect 20177 10625 20211 10659
rect 20211 10625 20220 10659
rect 20168 10616 20220 10625
rect 20444 10616 20496 10668
rect 20720 10616 20772 10668
rect 24860 10684 24912 10736
rect 21272 10548 21324 10600
rect 23940 10659 23992 10668
rect 23940 10625 23949 10659
rect 23949 10625 23983 10659
rect 23983 10625 23992 10659
rect 23940 10616 23992 10625
rect 23296 10548 23348 10600
rect 24676 10591 24728 10600
rect 24676 10557 24685 10591
rect 24685 10557 24719 10591
rect 24719 10557 24728 10591
rect 24676 10548 24728 10557
rect 17316 10480 17368 10532
rect 23940 10480 23992 10532
rect 16672 10412 16724 10464
rect 20444 10412 20496 10464
rect 20812 10412 20864 10464
rect 21272 10455 21324 10464
rect 21272 10421 21281 10455
rect 21281 10421 21315 10455
rect 21315 10421 21324 10455
rect 21272 10412 21324 10421
rect 21548 10412 21600 10464
rect 22100 10412 22152 10464
rect 2950 10310 3002 10362
rect 3014 10310 3066 10362
rect 3078 10310 3130 10362
rect 3142 10310 3194 10362
rect 3206 10310 3258 10362
rect 12950 10310 13002 10362
rect 13014 10310 13066 10362
rect 13078 10310 13130 10362
rect 13142 10310 13194 10362
rect 13206 10310 13258 10362
rect 22950 10310 23002 10362
rect 23014 10310 23066 10362
rect 23078 10310 23130 10362
rect 23142 10310 23194 10362
rect 23206 10310 23258 10362
rect 20168 10208 20220 10260
rect 20720 10251 20772 10260
rect 20720 10217 20729 10251
rect 20729 10217 20763 10251
rect 20763 10217 20772 10251
rect 20720 10208 20772 10217
rect 21732 10208 21784 10260
rect 19432 10183 19484 10192
rect 19432 10149 19441 10183
rect 19441 10149 19475 10183
rect 19475 10149 19484 10183
rect 19432 10140 19484 10149
rect 21272 10072 21324 10124
rect 21364 10115 21416 10124
rect 21364 10081 21373 10115
rect 21373 10081 21407 10115
rect 21407 10081 21416 10115
rect 21364 10072 21416 10081
rect 21640 10115 21692 10124
rect 21640 10081 21649 10115
rect 21649 10081 21683 10115
rect 21683 10081 21692 10115
rect 21640 10072 21692 10081
rect 23664 10072 23716 10124
rect 17592 10047 17644 10056
rect 17592 10013 17601 10047
rect 17601 10013 17635 10047
rect 17635 10013 17644 10047
rect 17592 10004 17644 10013
rect 20720 10004 20772 10056
rect 23112 10004 23164 10056
rect 20444 9868 20496 9920
rect 21548 9936 21600 9988
rect 21640 9936 21692 9988
rect 21916 9936 21968 9988
rect 25228 9936 25280 9988
rect 23112 9911 23164 9920
rect 23112 9877 23121 9911
rect 23121 9877 23155 9911
rect 23155 9877 23164 9911
rect 23112 9868 23164 9877
rect 7950 9766 8002 9818
rect 8014 9766 8066 9818
rect 8078 9766 8130 9818
rect 8142 9766 8194 9818
rect 8206 9766 8258 9818
rect 17950 9766 18002 9818
rect 18014 9766 18066 9818
rect 18078 9766 18130 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 17040 9596 17092 9648
rect 8484 9528 8536 9580
rect 19064 9528 19116 9580
rect 19524 9571 19576 9580
rect 19524 9537 19533 9571
rect 19533 9537 19567 9571
rect 19567 9537 19576 9571
rect 19524 9528 19576 9537
rect 20260 9528 20312 9580
rect 20628 9664 20680 9716
rect 23112 9664 23164 9716
rect 20444 9596 20496 9648
rect 21272 9571 21324 9580
rect 21272 9537 21281 9571
rect 21281 9537 21315 9571
rect 21315 9537 21324 9571
rect 21272 9528 21324 9537
rect 21640 9528 21692 9580
rect 23296 9639 23348 9648
rect 23296 9605 23305 9639
rect 23305 9605 23339 9639
rect 23339 9605 23348 9639
rect 23296 9596 23348 9605
rect 23940 9571 23992 9580
rect 23940 9537 23949 9571
rect 23949 9537 23983 9571
rect 23983 9537 23992 9571
rect 23940 9528 23992 9537
rect 22652 9460 22704 9512
rect 24768 9503 24820 9512
rect 24768 9469 24777 9503
rect 24777 9469 24811 9503
rect 24811 9469 24820 9503
rect 24768 9460 24820 9469
rect 19340 9435 19392 9444
rect 19340 9401 19349 9435
rect 19349 9401 19383 9435
rect 19383 9401 19392 9435
rect 19340 9392 19392 9401
rect 17776 9324 17828 9376
rect 20536 9324 20588 9376
rect 20720 9367 20772 9376
rect 20720 9333 20729 9367
rect 20729 9333 20763 9367
rect 20763 9333 20772 9367
rect 20720 9324 20772 9333
rect 2950 9222 3002 9274
rect 3014 9222 3066 9274
rect 3078 9222 3130 9274
rect 3142 9222 3194 9274
rect 3206 9222 3258 9274
rect 12950 9222 13002 9274
rect 13014 9222 13066 9274
rect 13078 9222 13130 9274
rect 13142 9222 13194 9274
rect 13206 9222 13258 9274
rect 22950 9222 23002 9274
rect 23014 9222 23066 9274
rect 23078 9222 23130 9274
rect 23142 9222 23194 9274
rect 23206 9222 23258 9274
rect 14740 9120 14792 9172
rect 19064 9163 19116 9172
rect 19064 9129 19073 9163
rect 19073 9129 19107 9163
rect 19107 9129 19116 9163
rect 19064 9120 19116 9129
rect 19524 9120 19576 9172
rect 21364 9120 21416 9172
rect 22008 9120 22060 9172
rect 23848 9120 23900 9172
rect 25780 9120 25832 9172
rect 10048 9027 10100 9036
rect 10048 8993 10057 9027
rect 10057 8993 10091 9027
rect 10091 8993 10100 9027
rect 10048 8984 10100 8993
rect 22100 9052 22152 9104
rect 22836 9052 22888 9104
rect 22744 8984 22796 9036
rect 24860 8984 24912 9036
rect 21180 8916 21232 8968
rect 21548 8916 21600 8968
rect 9312 8848 9364 8900
rect 12532 8848 12584 8900
rect 20720 8848 20772 8900
rect 21640 8848 21692 8900
rect 21916 8848 21968 8900
rect 20536 8780 20588 8832
rect 21364 8780 21416 8832
rect 22008 8823 22060 8832
rect 22008 8789 22017 8823
rect 22017 8789 22051 8823
rect 22051 8789 22060 8823
rect 22008 8780 22060 8789
rect 22284 8780 22336 8832
rect 7950 8678 8002 8730
rect 8014 8678 8066 8730
rect 8078 8678 8130 8730
rect 8142 8678 8194 8730
rect 8206 8678 8258 8730
rect 17950 8678 18002 8730
rect 18014 8678 18066 8730
rect 18078 8678 18130 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 22192 8576 22244 8628
rect 14832 8440 14884 8492
rect 21364 8508 21416 8560
rect 19892 8372 19944 8424
rect 22008 8440 22060 8492
rect 24860 8508 24912 8560
rect 21456 8415 21508 8424
rect 21456 8381 21465 8415
rect 21465 8381 21499 8415
rect 21499 8381 21508 8415
rect 21456 8372 21508 8381
rect 24952 8440 25004 8492
rect 24584 8415 24636 8424
rect 24584 8381 24593 8415
rect 24593 8381 24627 8415
rect 24627 8381 24636 8415
rect 24584 8372 24636 8381
rect 19708 8304 19760 8356
rect 24400 8304 24452 8356
rect 2950 8134 3002 8186
rect 3014 8134 3066 8186
rect 3078 8134 3130 8186
rect 3142 8134 3194 8186
rect 3206 8134 3258 8186
rect 12950 8134 13002 8186
rect 13014 8134 13066 8186
rect 13078 8134 13130 8186
rect 13142 8134 13194 8186
rect 13206 8134 13258 8186
rect 22950 8134 23002 8186
rect 23014 8134 23066 8186
rect 23078 8134 23130 8186
rect 23142 8134 23194 8186
rect 23206 8134 23258 8186
rect 20904 8032 20956 8084
rect 21916 8032 21968 8084
rect 24032 7964 24084 8016
rect 19800 7828 19852 7880
rect 23480 7896 23532 7948
rect 24952 7896 25004 7948
rect 22008 7828 22060 7880
rect 23388 7828 23440 7880
rect 25596 7760 25648 7812
rect 20720 7735 20772 7744
rect 20720 7701 20729 7735
rect 20729 7701 20763 7735
rect 20763 7701 20772 7735
rect 20720 7692 20772 7701
rect 23480 7692 23532 7744
rect 7950 7590 8002 7642
rect 8014 7590 8066 7642
rect 8078 7590 8130 7642
rect 8142 7590 8194 7642
rect 8206 7590 8258 7642
rect 17950 7590 18002 7642
rect 18014 7590 18066 7642
rect 18078 7590 18130 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 21272 7531 21324 7540
rect 21272 7497 21281 7531
rect 21281 7497 21315 7531
rect 21315 7497 21324 7531
rect 21272 7488 21324 7497
rect 20720 7420 20772 7472
rect 20352 7352 20404 7404
rect 21824 7352 21876 7404
rect 24860 7420 24912 7472
rect 25044 7352 25096 7404
rect 24676 7327 24728 7336
rect 24676 7293 24685 7327
rect 24685 7293 24719 7327
rect 24719 7293 24728 7327
rect 24676 7284 24728 7293
rect 23388 7148 23440 7200
rect 2950 7046 3002 7098
rect 3014 7046 3066 7098
rect 3078 7046 3130 7098
rect 3142 7046 3194 7098
rect 3206 7046 3258 7098
rect 12950 7046 13002 7098
rect 13014 7046 13066 7098
rect 13078 7046 13130 7098
rect 13142 7046 13194 7098
rect 13206 7046 13258 7098
rect 22950 7046 23002 7098
rect 23014 7046 23066 7098
rect 23078 7046 23130 7098
rect 23142 7046 23194 7098
rect 23206 7046 23258 7098
rect 20812 6783 20864 6792
rect 20812 6749 20821 6783
rect 20821 6749 20855 6783
rect 20855 6749 20864 6783
rect 20812 6740 20864 6749
rect 20996 6740 21048 6792
rect 21640 6740 21692 6792
rect 15200 6672 15252 6724
rect 22192 6783 22244 6792
rect 22192 6749 22201 6783
rect 22201 6749 22235 6783
rect 22235 6749 22244 6783
rect 22192 6740 22244 6749
rect 24860 6808 24912 6860
rect 21548 6604 21600 6656
rect 25044 6672 25096 6724
rect 7950 6502 8002 6554
rect 8014 6502 8066 6554
rect 8078 6502 8130 6554
rect 8142 6502 8194 6554
rect 8206 6502 8258 6554
rect 17950 6502 18002 6554
rect 18014 6502 18066 6554
rect 18078 6502 18130 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 9312 6443 9364 6452
rect 9312 6409 9321 6443
rect 9321 6409 9355 6443
rect 9355 6409 9364 6443
rect 9312 6400 9364 6409
rect 21824 6400 21876 6452
rect 24860 6332 24912 6384
rect 6828 6264 6880 6316
rect 22284 6307 22336 6316
rect 22284 6273 22293 6307
rect 22293 6273 22327 6307
rect 22327 6273 22336 6307
rect 22284 6264 22336 6273
rect 23664 6264 23716 6316
rect 24768 6239 24820 6248
rect 24768 6205 24777 6239
rect 24777 6205 24811 6239
rect 24811 6205 24820 6239
rect 24768 6196 24820 6205
rect 2950 5958 3002 6010
rect 3014 5958 3066 6010
rect 3078 5958 3130 6010
rect 3142 5958 3194 6010
rect 3206 5958 3258 6010
rect 12950 5958 13002 6010
rect 13014 5958 13066 6010
rect 13078 5958 13130 6010
rect 13142 5958 13194 6010
rect 13206 5958 13258 6010
rect 22950 5958 23002 6010
rect 23014 5958 23066 6010
rect 23078 5958 23130 6010
rect 23142 5958 23194 6010
rect 23206 5958 23258 6010
rect 20536 5856 20588 5908
rect 24584 5788 24636 5840
rect 21732 5652 21784 5704
rect 22376 5652 22428 5704
rect 23480 5652 23532 5704
rect 24400 5652 24452 5704
rect 24952 5584 25004 5636
rect 23480 5516 23532 5568
rect 7950 5414 8002 5466
rect 8014 5414 8066 5466
rect 8078 5414 8130 5466
rect 8142 5414 8194 5466
rect 8206 5414 8258 5466
rect 17950 5414 18002 5466
rect 18014 5414 18066 5466
rect 18078 5414 18130 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 24860 5244 24912 5296
rect 22468 5176 22520 5228
rect 22744 5176 22796 5228
rect 24676 5151 24728 5160
rect 24676 5117 24685 5151
rect 24685 5117 24719 5151
rect 24719 5117 24728 5151
rect 24676 5108 24728 5117
rect 2950 4870 3002 4922
rect 3014 4870 3066 4922
rect 3078 4870 3130 4922
rect 3142 4870 3194 4922
rect 3206 4870 3258 4922
rect 12950 4870 13002 4922
rect 13014 4870 13066 4922
rect 13078 4870 13130 4922
rect 13142 4870 13194 4922
rect 13206 4870 13258 4922
rect 22950 4870 23002 4922
rect 23014 4870 23066 4922
rect 23078 4870 23130 4922
rect 23142 4870 23194 4922
rect 23206 4870 23258 4922
rect 22376 4811 22428 4820
rect 22376 4777 22385 4811
rect 22385 4777 22419 4811
rect 22419 4777 22428 4811
rect 22376 4768 22428 4777
rect 22652 4607 22704 4616
rect 22652 4573 22661 4607
rect 22661 4573 22695 4607
rect 22695 4573 22704 4607
rect 22652 4564 22704 4573
rect 23388 4564 23440 4616
rect 24952 4496 25004 4548
rect 23572 4428 23624 4480
rect 7950 4326 8002 4378
rect 8014 4326 8066 4378
rect 8078 4326 8130 4378
rect 8142 4326 8194 4378
rect 8206 4326 8258 4378
rect 17950 4326 18002 4378
rect 18014 4326 18066 4378
rect 18078 4326 18130 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 20260 4131 20312 4140
rect 20260 4097 20269 4131
rect 20269 4097 20303 4131
rect 20303 4097 20312 4131
rect 20260 4088 20312 4097
rect 18972 4020 19024 4072
rect 20168 4020 20220 4072
rect 22100 4020 22152 4072
rect 25136 4088 25188 4140
rect 24768 4063 24820 4072
rect 24768 4029 24777 4063
rect 24777 4029 24811 4063
rect 24811 4029 24820 4063
rect 24768 4020 24820 4029
rect 24952 3952 25004 4004
rect 25044 3884 25096 3936
rect 2950 3782 3002 3834
rect 3014 3782 3066 3834
rect 3078 3782 3130 3834
rect 3142 3782 3194 3834
rect 3206 3782 3258 3834
rect 12950 3782 13002 3834
rect 13014 3782 13066 3834
rect 13078 3782 13130 3834
rect 13142 3782 13194 3834
rect 13206 3782 13258 3834
rect 22950 3782 23002 3834
rect 23014 3782 23066 3834
rect 23078 3782 23130 3834
rect 23142 3782 23194 3834
rect 23206 3782 23258 3834
rect 20076 3476 20128 3528
rect 23480 3476 23532 3528
rect 24584 3476 24636 3528
rect 22008 3451 22060 3460
rect 22008 3417 22017 3451
rect 22017 3417 22051 3451
rect 22051 3417 22060 3451
rect 22008 3408 22060 3417
rect 24952 3408 25004 3460
rect 24584 3383 24636 3392
rect 24584 3349 24593 3383
rect 24593 3349 24627 3383
rect 24627 3349 24636 3383
rect 24584 3340 24636 3349
rect 7950 3238 8002 3290
rect 8014 3238 8066 3290
rect 8078 3238 8130 3290
rect 8142 3238 8194 3290
rect 8206 3238 8258 3290
rect 17950 3238 18002 3290
rect 18014 3238 18066 3290
rect 18078 3238 18130 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 6828 3179 6880 3188
rect 6828 3145 6837 3179
rect 6837 3145 6871 3179
rect 6871 3145 6880 3179
rect 6828 3136 6880 3145
rect 24860 3068 24912 3120
rect 25136 3111 25188 3120
rect 25136 3077 25145 3111
rect 25145 3077 25179 3111
rect 25179 3077 25188 3111
rect 25136 3068 25188 3077
rect 7012 3043 7064 3052
rect 7012 3009 7021 3043
rect 7021 3009 7055 3043
rect 7055 3009 7064 3043
rect 7012 3000 7064 3009
rect 19800 3000 19852 3052
rect 19984 3000 20036 3052
rect 23572 3000 23624 3052
rect 24216 3000 24268 3052
rect 19340 2975 19392 2984
rect 19340 2941 19349 2975
rect 19349 2941 19383 2975
rect 19383 2941 19392 2975
rect 19340 2932 19392 2941
rect 25044 2932 25096 2984
rect 19800 2796 19852 2848
rect 25872 2796 25924 2848
rect 2950 2694 3002 2746
rect 3014 2694 3066 2746
rect 3078 2694 3130 2746
rect 3142 2694 3194 2746
rect 3206 2694 3258 2746
rect 12950 2694 13002 2746
rect 13014 2694 13066 2746
rect 13078 2694 13130 2746
rect 13142 2694 13194 2746
rect 13206 2694 13258 2746
rect 22950 2694 23002 2746
rect 23014 2694 23066 2746
rect 23078 2694 23130 2746
rect 23142 2694 23194 2746
rect 23206 2694 23258 2746
rect 7012 2592 7064 2644
rect 19340 2592 19392 2644
rect 22192 2592 22244 2644
rect 19800 2567 19852 2576
rect 19800 2533 19809 2567
rect 19809 2533 19843 2567
rect 19843 2533 19852 2567
rect 19800 2524 19852 2533
rect 20628 2388 20680 2440
rect 24584 2388 24636 2440
rect 23388 2320 23440 2372
rect 24952 2320 25004 2372
rect 6736 2252 6788 2304
rect 7950 2150 8002 2202
rect 8014 2150 8066 2202
rect 8078 2150 8130 2202
rect 8142 2150 8194 2202
rect 8206 2150 8258 2202
rect 17950 2150 18002 2202
rect 18014 2150 18066 2202
rect 18078 2150 18130 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
<< metal2 >>
rect 1674 26200 1730 27000
rect 2042 26200 2098 27000
rect 2136 26376 2188 26382
rect 2136 26318 2188 26324
rect 2410 26330 2466 27000
rect 2778 26466 2834 27000
rect 2778 26450 3096 26466
rect 2778 26444 3108 26450
rect 2778 26438 3056 26444
rect 1688 24290 1716 26200
rect 1952 25084 2004 25090
rect 1952 25026 2004 25032
rect 1688 24262 1900 24290
rect 1768 24200 1820 24206
rect 1766 24168 1768 24177
rect 1820 24168 1822 24177
rect 1766 24103 1822 24112
rect 1122 23760 1178 23769
rect 1122 23695 1124 23704
rect 1176 23695 1178 23704
rect 1492 23724 1544 23730
rect 1124 23666 1176 23672
rect 1492 23666 1544 23672
rect 1504 23322 1532 23666
rect 1492 23316 1544 23322
rect 1492 23258 1544 23264
rect 1214 22672 1270 22681
rect 1214 22607 1216 22616
rect 1268 22607 1270 22616
rect 1676 22636 1728 22642
rect 1216 22578 1268 22584
rect 1676 22578 1728 22584
rect 1688 22234 1716 22578
rect 1768 22432 1820 22438
rect 1768 22374 1820 22380
rect 1676 22228 1728 22234
rect 1676 22170 1728 22176
rect 1780 22166 1808 22374
rect 1768 22160 1820 22166
rect 1768 22102 1820 22108
rect 1768 21344 1820 21350
rect 1768 21286 1820 21292
rect 1780 21146 1808 21286
rect 1768 21140 1820 21146
rect 1768 21082 1820 21088
rect 1872 19310 1900 24262
rect 1860 19304 1912 19310
rect 1860 19246 1912 19252
rect 1964 18970 1992 25026
rect 2056 19922 2084 26200
rect 2044 19916 2096 19922
rect 2044 19858 2096 19864
rect 1952 18964 2004 18970
rect 1952 18906 2004 18912
rect 2148 18766 2176 26318
rect 2410 26302 2728 26330
rect 2410 26200 2466 26302
rect 2700 23474 2728 26302
rect 2778 26200 2834 26438
rect 3056 26386 3108 26392
rect 3146 26330 3202 27000
rect 3332 26444 3384 26450
rect 3332 26386 3384 26392
rect 2884 26302 3202 26330
rect 2700 23446 2820 23474
rect 2228 23112 2280 23118
rect 2228 23054 2280 23060
rect 2240 22778 2268 23054
rect 2228 22772 2280 22778
rect 2228 22714 2280 22720
rect 2792 21010 2820 23446
rect 2884 22098 2912 26302
rect 3146 26200 3202 26302
rect 2950 24508 3258 24517
rect 2950 24506 2956 24508
rect 3012 24506 3036 24508
rect 3092 24506 3116 24508
rect 3172 24506 3196 24508
rect 3252 24506 3258 24508
rect 3012 24454 3014 24506
rect 3194 24454 3196 24506
rect 2950 24452 2956 24454
rect 3012 24452 3036 24454
rect 3092 24452 3116 24454
rect 3172 24452 3196 24454
rect 3252 24452 3258 24454
rect 2950 24443 3258 24452
rect 2950 23420 3258 23429
rect 2950 23418 2956 23420
rect 3012 23418 3036 23420
rect 3092 23418 3116 23420
rect 3172 23418 3196 23420
rect 3252 23418 3258 23420
rect 3012 23366 3014 23418
rect 3194 23366 3196 23418
rect 2950 23364 2956 23366
rect 3012 23364 3036 23366
rect 3092 23364 3116 23366
rect 3172 23364 3196 23366
rect 3252 23364 3258 23366
rect 2950 23355 3258 23364
rect 3240 22568 3292 22574
rect 3238 22536 3240 22545
rect 3292 22536 3294 22545
rect 3238 22471 3294 22480
rect 2950 22332 3258 22341
rect 2950 22330 2956 22332
rect 3012 22330 3036 22332
rect 3092 22330 3116 22332
rect 3172 22330 3196 22332
rect 3252 22330 3258 22332
rect 3012 22278 3014 22330
rect 3194 22278 3196 22330
rect 2950 22276 2956 22278
rect 3012 22276 3036 22278
rect 3092 22276 3116 22278
rect 3172 22276 3196 22278
rect 3252 22276 3258 22278
rect 2950 22267 3258 22276
rect 2872 22092 2924 22098
rect 2872 22034 2924 22040
rect 2950 21244 3258 21253
rect 2950 21242 2956 21244
rect 3012 21242 3036 21244
rect 3092 21242 3116 21244
rect 3172 21242 3196 21244
rect 3252 21242 3258 21244
rect 3012 21190 3014 21242
rect 3194 21190 3196 21242
rect 2950 21188 2956 21190
rect 3012 21188 3036 21190
rect 3092 21188 3116 21190
rect 3172 21188 3196 21190
rect 3252 21188 3258 21190
rect 2950 21179 3258 21188
rect 2780 21004 2832 21010
rect 2780 20946 2832 20952
rect 3344 20398 3372 26386
rect 3514 26200 3570 27000
rect 3882 26330 3938 27000
rect 3882 26302 4108 26330
rect 3882 26200 3938 26302
rect 3422 24848 3478 24857
rect 3422 24783 3478 24792
rect 3436 23118 3464 24783
rect 3424 23112 3476 23118
rect 3424 23054 3476 23060
rect 3436 22710 3464 23054
rect 3424 22704 3476 22710
rect 3424 22646 3476 22652
rect 3424 22568 3476 22574
rect 3424 22510 3476 22516
rect 3436 21690 3464 22510
rect 3424 21684 3476 21690
rect 3424 21626 3476 21632
rect 3528 21486 3556 26200
rect 3698 25936 3754 25945
rect 3698 25871 3754 25880
rect 3608 25220 3660 25226
rect 3608 25162 3660 25168
rect 3620 22420 3648 25162
rect 3712 22574 3740 25871
rect 3884 24200 3936 24206
rect 3884 24142 3936 24148
rect 3792 23724 3844 23730
rect 3792 23666 3844 23672
rect 3700 22568 3752 22574
rect 3804 22545 3832 23666
rect 3700 22510 3752 22516
rect 3790 22536 3846 22545
rect 3790 22471 3846 22480
rect 3792 22432 3844 22438
rect 3620 22392 3740 22420
rect 3608 22160 3660 22166
rect 3608 22102 3660 22108
rect 3516 21480 3568 21486
rect 3516 21422 3568 21428
rect 3332 20392 3384 20398
rect 3332 20334 3384 20340
rect 3514 20224 3570 20233
rect 2950 20156 3258 20165
rect 3514 20159 3570 20168
rect 2950 20154 2956 20156
rect 3012 20154 3036 20156
rect 3092 20154 3116 20156
rect 3172 20154 3196 20156
rect 3252 20154 3258 20156
rect 3012 20102 3014 20154
rect 3194 20102 3196 20154
rect 2950 20100 2956 20102
rect 3012 20100 3036 20102
rect 3092 20100 3116 20102
rect 3172 20100 3196 20102
rect 3252 20100 3258 20102
rect 2950 20091 3258 20100
rect 3332 19304 3384 19310
rect 3332 19246 3384 19252
rect 2950 19068 3258 19077
rect 2950 19066 2956 19068
rect 3012 19066 3036 19068
rect 3092 19066 3116 19068
rect 3172 19066 3196 19068
rect 3252 19066 3258 19068
rect 3012 19014 3014 19066
rect 3194 19014 3196 19066
rect 2950 19012 2956 19014
rect 3012 19012 3036 19014
rect 3092 19012 3116 19014
rect 3172 19012 3196 19014
rect 3252 19012 3258 19014
rect 2950 19003 3258 19012
rect 2596 18896 2648 18902
rect 2594 18864 2596 18873
rect 2648 18864 2650 18873
rect 2594 18799 2650 18808
rect 2136 18760 2188 18766
rect 2136 18702 2188 18708
rect 2228 18352 2280 18358
rect 2226 18320 2228 18329
rect 2280 18320 2282 18329
rect 2226 18255 2282 18264
rect 2950 17980 3258 17989
rect 2950 17978 2956 17980
rect 3012 17978 3036 17980
rect 3092 17978 3116 17980
rect 3172 17978 3196 17980
rect 3252 17978 3258 17980
rect 3012 17926 3014 17978
rect 3194 17926 3196 17978
rect 2950 17924 2956 17926
rect 3012 17924 3036 17926
rect 3092 17924 3116 17926
rect 3172 17924 3196 17926
rect 3252 17924 3258 17926
rect 2950 17915 3258 17924
rect 3344 17882 3372 19246
rect 3528 18426 3556 20159
rect 3516 18420 3568 18426
rect 3516 18362 3568 18368
rect 3620 18154 3648 22102
rect 3712 18426 3740 22392
rect 3792 22374 3844 22380
rect 3804 22166 3832 22374
rect 3792 22160 3844 22166
rect 3792 22102 3844 22108
rect 3790 21584 3846 21593
rect 3790 21519 3846 21528
rect 3804 19378 3832 21519
rect 3896 19514 3924 24142
rect 3976 24064 4028 24070
rect 3976 24006 4028 24012
rect 3988 20602 4016 24006
rect 4080 22094 4108 26302
rect 4250 26200 4306 27000
rect 4618 26200 4674 27000
rect 4986 26330 5042 27000
rect 4986 26302 5120 26330
rect 4894 26208 4950 26217
rect 4264 22710 4292 26200
rect 4632 23186 4660 26200
rect 4986 26200 5042 26302
rect 4894 26143 4950 26152
rect 4802 24984 4858 24993
rect 4802 24919 4858 24928
rect 4816 24206 4844 24919
rect 4804 24200 4856 24206
rect 4804 24142 4856 24148
rect 4908 24018 4936 26143
rect 4816 23990 4936 24018
rect 4620 23180 4672 23186
rect 4620 23122 4672 23128
rect 4712 22976 4764 22982
rect 4712 22918 4764 22924
rect 4724 22778 4752 22918
rect 4712 22772 4764 22778
rect 4712 22714 4764 22720
rect 4252 22704 4304 22710
rect 4816 22658 4844 23990
rect 4896 23860 4948 23866
rect 4896 23802 4948 23808
rect 4252 22646 4304 22652
rect 4724 22630 4844 22658
rect 4080 22066 4200 22094
rect 4172 21010 4200 22066
rect 4528 22024 4580 22030
rect 4528 21966 4580 21972
rect 4160 21004 4212 21010
rect 4160 20946 4212 20952
rect 3976 20596 4028 20602
rect 3976 20538 4028 20544
rect 4160 20256 4212 20262
rect 4160 20198 4212 20204
rect 3976 20052 4028 20058
rect 3976 19994 4028 20000
rect 3884 19508 3936 19514
rect 3884 19450 3936 19456
rect 3792 19372 3844 19378
rect 3792 19314 3844 19320
rect 3882 18728 3938 18737
rect 3882 18663 3884 18672
rect 3936 18663 3938 18672
rect 3884 18634 3936 18640
rect 3700 18420 3752 18426
rect 3700 18362 3752 18368
rect 3608 18148 3660 18154
rect 3608 18090 3660 18096
rect 3332 17876 3384 17882
rect 3332 17818 3384 17824
rect 3424 17672 3476 17678
rect 3424 17614 3476 17620
rect 2950 16892 3258 16901
rect 2950 16890 2956 16892
rect 3012 16890 3036 16892
rect 3092 16890 3116 16892
rect 3172 16890 3196 16892
rect 3252 16890 3258 16892
rect 3012 16838 3014 16890
rect 3194 16838 3196 16890
rect 2950 16836 2956 16838
rect 3012 16836 3036 16838
rect 3092 16836 3116 16838
rect 3172 16836 3196 16838
rect 3252 16836 3258 16838
rect 2950 16827 3258 16836
rect 3436 16726 3464 17614
rect 3988 17338 4016 19994
rect 4172 18766 4200 20198
rect 4160 18760 4212 18766
rect 4160 18702 4212 18708
rect 4068 18080 4120 18086
rect 4068 18022 4120 18028
rect 3976 17332 4028 17338
rect 3976 17274 4028 17280
rect 3424 16720 3476 16726
rect 3424 16662 3476 16668
rect 2950 15804 3258 15813
rect 2950 15802 2956 15804
rect 3012 15802 3036 15804
rect 3092 15802 3116 15804
rect 3172 15802 3196 15804
rect 3252 15802 3258 15804
rect 3012 15750 3014 15802
rect 3194 15750 3196 15802
rect 2950 15748 2956 15750
rect 3012 15748 3036 15750
rect 3092 15748 3116 15750
rect 3172 15748 3196 15750
rect 3252 15748 3258 15750
rect 2950 15739 3258 15748
rect 2950 14716 3258 14725
rect 2950 14714 2956 14716
rect 3012 14714 3036 14716
rect 3092 14714 3116 14716
rect 3172 14714 3196 14716
rect 3252 14714 3258 14716
rect 3012 14662 3014 14714
rect 3194 14662 3196 14714
rect 2950 14660 2956 14662
rect 3012 14660 3036 14662
rect 3092 14660 3116 14662
rect 3172 14660 3196 14662
rect 3252 14660 3258 14662
rect 2950 14651 3258 14660
rect 2950 13628 3258 13637
rect 2950 13626 2956 13628
rect 3012 13626 3036 13628
rect 3092 13626 3116 13628
rect 3172 13626 3196 13628
rect 3252 13626 3258 13628
rect 3012 13574 3014 13626
rect 3194 13574 3196 13626
rect 2950 13572 2956 13574
rect 3012 13572 3036 13574
rect 3092 13572 3116 13574
rect 3172 13572 3196 13574
rect 3252 13572 3258 13574
rect 2950 13563 3258 13572
rect 2950 12540 3258 12549
rect 2950 12538 2956 12540
rect 3012 12538 3036 12540
rect 3092 12538 3116 12540
rect 3172 12538 3196 12540
rect 3252 12538 3258 12540
rect 3012 12486 3014 12538
rect 3194 12486 3196 12538
rect 2950 12484 2956 12486
rect 3012 12484 3036 12486
rect 3092 12484 3116 12486
rect 3172 12484 3196 12486
rect 3252 12484 3258 12486
rect 2950 12475 3258 12484
rect 4080 12442 4108 18022
rect 4252 17536 4304 17542
rect 4252 17478 4304 17484
rect 4264 17338 4292 17478
rect 4252 17332 4304 17338
rect 4252 17274 4304 17280
rect 4160 16584 4212 16590
rect 4158 16552 4160 16561
rect 4212 16552 4214 16561
rect 4158 16487 4214 16496
rect 4172 16250 4200 16487
rect 4160 16244 4212 16250
rect 4160 16186 4212 16192
rect 4540 14385 4568 21966
rect 4724 20602 4752 22630
rect 4802 22128 4858 22137
rect 4802 22063 4858 22072
rect 4816 21554 4844 22063
rect 4804 21548 4856 21554
rect 4804 21490 4856 21496
rect 4712 20596 4764 20602
rect 4712 20538 4764 20544
rect 4724 19854 4752 20538
rect 4712 19848 4764 19854
rect 4712 19790 4764 19796
rect 4908 19378 4936 23802
rect 4988 21888 5040 21894
rect 4988 21830 5040 21836
rect 4896 19372 4948 19378
rect 4896 19314 4948 19320
rect 4710 19136 4766 19145
rect 4710 19071 4766 19080
rect 4724 18766 4752 19071
rect 4712 18760 4764 18766
rect 4712 18702 4764 18708
rect 5000 18426 5028 21830
rect 5092 21486 5120 26302
rect 5354 26200 5410 27000
rect 5722 26200 5778 27000
rect 6090 26200 6146 27000
rect 6458 26200 6514 27000
rect 6826 26200 6882 27000
rect 7194 26330 7250 27000
rect 7562 26330 7618 27000
rect 7930 26330 7986 27000
rect 7194 26302 7328 26330
rect 7194 26200 7250 26302
rect 5172 25152 5224 25158
rect 5172 25094 5224 25100
rect 5080 21480 5132 21486
rect 5080 21422 5132 21428
rect 5184 20602 5212 25094
rect 5264 24608 5316 24614
rect 5264 24550 5316 24556
rect 5172 20596 5224 20602
rect 5172 20538 5224 20544
rect 5172 20324 5224 20330
rect 5172 20266 5224 20272
rect 4988 18420 5040 18426
rect 4988 18362 5040 18368
rect 4620 18352 4672 18358
rect 4620 18294 4672 18300
rect 4632 18154 4660 18294
rect 4620 18148 4672 18154
rect 4620 18090 4672 18096
rect 5184 17270 5212 20266
rect 5276 19922 5304 24550
rect 5368 23798 5396 26200
rect 5356 23792 5408 23798
rect 5356 23734 5408 23740
rect 5446 23624 5502 23633
rect 5446 23559 5502 23568
rect 5460 23118 5488 23559
rect 5448 23112 5500 23118
rect 5448 23054 5500 23060
rect 5632 23044 5684 23050
rect 5632 22986 5684 22992
rect 5540 22432 5592 22438
rect 5540 22374 5592 22380
rect 5448 22024 5500 22030
rect 5448 21966 5500 21972
rect 5356 20528 5408 20534
rect 5356 20470 5408 20476
rect 5264 19916 5316 19922
rect 5264 19858 5316 19864
rect 5368 19174 5396 20470
rect 5356 19168 5408 19174
rect 5356 19110 5408 19116
rect 5460 17882 5488 21966
rect 5552 21622 5580 22374
rect 5540 21616 5592 21622
rect 5540 21558 5592 21564
rect 5644 21321 5672 22986
rect 5736 22710 5764 26200
rect 5816 24812 5868 24818
rect 5816 24754 5868 24760
rect 5828 24138 5856 24754
rect 6000 24744 6052 24750
rect 6000 24686 6052 24692
rect 5816 24132 5868 24138
rect 5816 24074 5868 24080
rect 5724 22704 5776 22710
rect 5724 22646 5776 22652
rect 5816 22636 5868 22642
rect 5816 22578 5868 22584
rect 5630 21312 5686 21321
rect 5630 21247 5686 21256
rect 5828 21185 5856 22578
rect 5814 21176 5870 21185
rect 5814 21111 5870 21120
rect 5632 21004 5684 21010
rect 5632 20946 5684 20952
rect 5540 20460 5592 20466
rect 5540 20402 5592 20408
rect 5552 20369 5580 20402
rect 5538 20360 5594 20369
rect 5538 20295 5594 20304
rect 5540 19712 5592 19718
rect 5540 19654 5592 19660
rect 5552 18290 5580 19654
rect 5540 18284 5592 18290
rect 5540 18226 5592 18232
rect 5448 17876 5500 17882
rect 5448 17818 5500 17824
rect 5448 17672 5500 17678
rect 5448 17614 5500 17620
rect 5172 17264 5224 17270
rect 5172 17206 5224 17212
rect 5460 17134 5488 17614
rect 4804 17128 4856 17134
rect 4804 17070 4856 17076
rect 5448 17128 5500 17134
rect 5448 17070 5500 17076
rect 4816 16969 4844 17070
rect 4802 16960 4858 16969
rect 4802 16895 4858 16904
rect 5644 16182 5672 20946
rect 5724 20936 5776 20942
rect 5724 20878 5776 20884
rect 5736 18426 5764 20878
rect 5906 20768 5962 20777
rect 5906 20703 5962 20712
rect 5816 19848 5868 19854
rect 5816 19790 5868 19796
rect 5828 19514 5856 19790
rect 5816 19508 5868 19514
rect 5816 19450 5868 19456
rect 5920 18970 5948 20703
rect 6012 19378 6040 24686
rect 6104 22098 6132 26200
rect 6368 24336 6420 24342
rect 6368 24278 6420 24284
rect 6380 23050 6408 24278
rect 6472 24274 6500 26200
rect 6550 25120 6606 25129
rect 6550 25055 6606 25064
rect 6564 24342 6592 25055
rect 6644 25016 6696 25022
rect 6644 24958 6696 24964
rect 6552 24336 6604 24342
rect 6552 24278 6604 24284
rect 6460 24268 6512 24274
rect 6460 24210 6512 24216
rect 6460 23588 6512 23594
rect 6460 23530 6512 23536
rect 6368 23044 6420 23050
rect 6368 22986 6420 22992
rect 6274 22672 6330 22681
rect 6274 22607 6330 22616
rect 6184 22568 6236 22574
rect 6184 22510 6236 22516
rect 6092 22092 6144 22098
rect 6092 22034 6144 22040
rect 6196 20890 6224 22510
rect 6104 20862 6224 20890
rect 6000 19372 6052 19378
rect 6000 19314 6052 19320
rect 5908 18964 5960 18970
rect 5908 18906 5960 18912
rect 6104 18834 6132 20862
rect 6184 20800 6236 20806
rect 6184 20742 6236 20748
rect 6092 18828 6144 18834
rect 6092 18770 6144 18776
rect 6000 18760 6052 18766
rect 6000 18702 6052 18708
rect 6012 18426 6040 18702
rect 5724 18420 5776 18426
rect 5724 18362 5776 18368
rect 6000 18420 6052 18426
rect 6000 18362 6052 18368
rect 6196 17678 6224 20742
rect 6288 18222 6316 22607
rect 6366 22264 6422 22273
rect 6366 22199 6422 22208
rect 6276 18216 6328 18222
rect 6276 18158 6328 18164
rect 6380 18154 6408 22199
rect 6472 21690 6500 23530
rect 6656 22094 6684 24958
rect 6736 24200 6788 24206
rect 6736 24142 6788 24148
rect 6748 23361 6776 24142
rect 6734 23352 6790 23361
rect 6734 23287 6736 23296
rect 6788 23287 6790 23296
rect 6736 23258 6788 23264
rect 6736 22636 6788 22642
rect 6736 22578 6788 22584
rect 6564 22066 6684 22094
rect 6460 21684 6512 21690
rect 6460 21626 6512 21632
rect 6564 20602 6592 22066
rect 6552 20596 6604 20602
rect 6552 20538 6604 20544
rect 6552 20392 6604 20398
rect 6552 20334 6604 20340
rect 6460 19304 6512 19310
rect 6458 19272 6460 19281
rect 6512 19272 6514 19281
rect 6458 19207 6514 19216
rect 6472 18766 6500 19207
rect 6460 18760 6512 18766
rect 6460 18702 6512 18708
rect 6368 18148 6420 18154
rect 6368 18090 6420 18096
rect 6564 17921 6592 20334
rect 6644 19848 6696 19854
rect 6644 19790 6696 19796
rect 6656 19417 6684 19790
rect 6748 19514 6776 22578
rect 6840 22094 6868 26200
rect 7104 23520 7156 23526
rect 7104 23462 7156 23468
rect 7012 23112 7064 23118
rect 7012 23054 7064 23060
rect 6840 22066 6960 22094
rect 6932 21010 6960 22066
rect 6920 21004 6972 21010
rect 6920 20946 6972 20952
rect 7024 20777 7052 23054
rect 7116 21026 7144 23462
rect 7300 21486 7328 26302
rect 7392 26302 7618 26330
rect 7392 23798 7420 26302
rect 7562 26200 7618 26302
rect 7668 26302 7986 26330
rect 7564 25288 7616 25294
rect 7564 25230 7616 25236
rect 7472 24064 7524 24070
rect 7472 24006 7524 24012
rect 7380 23792 7432 23798
rect 7380 23734 7432 23740
rect 7380 23588 7432 23594
rect 7380 23530 7432 23536
rect 7392 23322 7420 23530
rect 7380 23316 7432 23322
rect 7380 23258 7432 23264
rect 7392 22710 7420 23258
rect 7380 22704 7432 22710
rect 7380 22646 7432 22652
rect 7380 21548 7432 21554
rect 7380 21490 7432 21496
rect 7288 21480 7340 21486
rect 7288 21422 7340 21428
rect 7116 20998 7236 21026
rect 7104 20936 7156 20942
rect 7104 20878 7156 20884
rect 7010 20768 7066 20777
rect 7010 20703 7066 20712
rect 7012 20392 7064 20398
rect 7012 20334 7064 20340
rect 6828 20256 6880 20262
rect 6828 20198 6880 20204
rect 6736 19508 6788 19514
rect 6736 19450 6788 19456
rect 6642 19408 6698 19417
rect 6642 19343 6698 19352
rect 6736 18964 6788 18970
rect 6736 18906 6788 18912
rect 6550 17912 6606 17921
rect 6550 17847 6606 17856
rect 6184 17672 6236 17678
rect 6184 17614 6236 17620
rect 6552 16992 6604 16998
rect 6552 16934 6604 16940
rect 5632 16176 5684 16182
rect 5632 16118 5684 16124
rect 6564 14929 6592 16934
rect 6550 14920 6606 14929
rect 6550 14855 6606 14864
rect 4526 14376 4582 14385
rect 4526 14311 4582 14320
rect 6748 12889 6776 18906
rect 6840 18358 6868 20198
rect 7024 19718 7052 20334
rect 7012 19712 7064 19718
rect 7012 19654 7064 19660
rect 6920 19236 6972 19242
rect 6920 19178 6972 19184
rect 6828 18352 6880 18358
rect 6828 18294 6880 18300
rect 6932 18290 6960 19178
rect 7012 19168 7064 19174
rect 7012 19110 7064 19116
rect 7024 18970 7052 19110
rect 7012 18964 7064 18970
rect 7012 18906 7064 18912
rect 6920 18284 6972 18290
rect 6920 18226 6972 18232
rect 7010 18184 7066 18193
rect 7010 18119 7012 18128
rect 7064 18119 7066 18128
rect 7012 18090 7064 18096
rect 7116 17882 7144 20878
rect 7208 20602 7236 20998
rect 7196 20596 7248 20602
rect 7196 20538 7248 20544
rect 7196 20460 7248 20466
rect 7196 20402 7248 20408
rect 7208 20058 7236 20402
rect 7196 20052 7248 20058
rect 7196 19994 7248 20000
rect 7286 19952 7342 19961
rect 7286 19887 7342 19896
rect 7196 19304 7248 19310
rect 7196 19246 7248 19252
rect 7208 18290 7236 19246
rect 7300 19174 7328 19887
rect 7288 19168 7340 19174
rect 7288 19110 7340 19116
rect 7196 18284 7248 18290
rect 7196 18226 7248 18232
rect 7288 18080 7340 18086
rect 7286 18048 7288 18057
rect 7340 18048 7342 18057
rect 7286 17983 7342 17992
rect 7104 17876 7156 17882
rect 7104 17818 7156 17824
rect 6920 17808 6972 17814
rect 6918 17776 6920 17785
rect 7196 17808 7248 17814
rect 6972 17776 6974 17785
rect 7196 17750 7248 17756
rect 6918 17711 6974 17720
rect 7102 17640 7158 17649
rect 7102 17575 7158 17584
rect 7116 17542 7144 17575
rect 6828 17536 6880 17542
rect 6828 17478 6880 17484
rect 7104 17536 7156 17542
rect 7104 17478 7156 17484
rect 6840 16153 6868 17478
rect 7208 17338 7236 17750
rect 7300 17678 7328 17983
rect 7288 17672 7340 17678
rect 7288 17614 7340 17620
rect 7392 17338 7420 21490
rect 7484 19922 7512 24006
rect 7576 23662 7604 25230
rect 7564 23656 7616 23662
rect 7564 23598 7616 23604
rect 7668 23186 7696 26302
rect 7930 26200 7986 26302
rect 8298 26200 8354 27000
rect 8666 26330 8722 27000
rect 9034 26330 9090 27000
rect 8404 26302 8722 26330
rect 7748 24676 7800 24682
rect 7748 24618 7800 24624
rect 7656 23180 7708 23186
rect 7656 23122 7708 23128
rect 7564 23044 7616 23050
rect 7564 22986 7616 22992
rect 7472 19916 7524 19922
rect 7472 19858 7524 19864
rect 7472 19712 7524 19718
rect 7472 19654 7524 19660
rect 7012 17332 7064 17338
rect 7012 17274 7064 17280
rect 7196 17332 7248 17338
rect 7196 17274 7248 17280
rect 7380 17332 7432 17338
rect 7380 17274 7432 17280
rect 6920 17196 6972 17202
rect 6920 17138 6972 17144
rect 6932 16658 6960 17138
rect 7024 16833 7052 17274
rect 7288 17196 7340 17202
rect 7288 17138 7340 17144
rect 7010 16824 7066 16833
rect 7300 16794 7328 17138
rect 7010 16759 7066 16768
rect 7288 16788 7340 16794
rect 7288 16730 7340 16736
rect 6920 16652 6972 16658
rect 6920 16594 6972 16600
rect 7380 16584 7432 16590
rect 7380 16526 7432 16532
rect 6826 16144 6882 16153
rect 6826 16079 6882 16088
rect 7392 13841 7420 16526
rect 7484 15978 7512 19654
rect 7576 18834 7604 22986
rect 7760 22094 7788 24618
rect 7950 23964 8258 23973
rect 7950 23962 7956 23964
rect 8012 23962 8036 23964
rect 8092 23962 8116 23964
rect 8172 23962 8196 23964
rect 8252 23962 8258 23964
rect 8012 23910 8014 23962
rect 8194 23910 8196 23962
rect 7950 23908 7956 23910
rect 8012 23908 8036 23910
rect 8092 23908 8116 23910
rect 8172 23908 8196 23910
rect 8252 23908 8258 23910
rect 7950 23899 8258 23908
rect 7950 22876 8258 22885
rect 7950 22874 7956 22876
rect 8012 22874 8036 22876
rect 8092 22874 8116 22876
rect 8172 22874 8196 22876
rect 8252 22874 8258 22876
rect 8012 22822 8014 22874
rect 8194 22822 8196 22874
rect 7950 22820 7956 22822
rect 8012 22820 8036 22822
rect 8092 22820 8116 22822
rect 8172 22820 8196 22822
rect 8252 22820 8258 22822
rect 7950 22811 8258 22820
rect 8312 22098 8340 26200
rect 8404 24818 8432 26302
rect 8666 26200 8722 26302
rect 8772 26302 9090 26330
rect 8484 24880 8536 24886
rect 8484 24822 8536 24828
rect 8392 24812 8444 24818
rect 8392 24754 8444 24760
rect 8496 24342 8524 24822
rect 8576 24608 8628 24614
rect 8576 24550 8628 24556
rect 8484 24336 8536 24342
rect 8484 24278 8536 24284
rect 8588 23730 8616 24550
rect 8666 23760 8722 23769
rect 8576 23724 8628 23730
rect 8666 23695 8722 23704
rect 8576 23666 8628 23672
rect 8574 23352 8630 23361
rect 8574 23287 8630 23296
rect 8390 23216 8446 23225
rect 8588 23186 8616 23287
rect 8390 23151 8446 23160
rect 8576 23180 8628 23186
rect 7668 22066 7788 22094
rect 8300 22092 8352 22098
rect 7668 19310 7696 22066
rect 8300 22034 8352 22040
rect 7840 22024 7892 22030
rect 7840 21966 7892 21972
rect 7852 21457 7880 21966
rect 8300 21956 8352 21962
rect 8300 21898 8352 21904
rect 7950 21788 8258 21797
rect 7950 21786 7956 21788
rect 8012 21786 8036 21788
rect 8092 21786 8116 21788
rect 8172 21786 8196 21788
rect 8252 21786 8258 21788
rect 8012 21734 8014 21786
rect 8194 21734 8196 21786
rect 7950 21732 7956 21734
rect 8012 21732 8036 21734
rect 8092 21732 8116 21734
rect 8172 21732 8196 21734
rect 8252 21732 8258 21734
rect 7950 21723 8258 21732
rect 8208 21684 8260 21690
rect 8208 21626 8260 21632
rect 7838 21448 7894 21457
rect 7838 21383 7894 21392
rect 7840 21344 7892 21350
rect 7840 21286 7892 21292
rect 7748 20936 7800 20942
rect 7748 20878 7800 20884
rect 7760 20602 7788 20878
rect 7748 20596 7800 20602
rect 7748 20538 7800 20544
rect 7748 20392 7800 20398
rect 7748 20334 7800 20340
rect 7760 19378 7788 20334
rect 7748 19372 7800 19378
rect 7748 19314 7800 19320
rect 7656 19304 7708 19310
rect 7656 19246 7708 19252
rect 7746 19272 7802 19281
rect 7746 19207 7802 19216
rect 7656 19168 7708 19174
rect 7656 19110 7708 19116
rect 7564 18828 7616 18834
rect 7564 18770 7616 18776
rect 7668 18170 7696 19110
rect 7576 18142 7696 18170
rect 7472 15972 7524 15978
rect 7472 15914 7524 15920
rect 7576 15366 7604 18142
rect 7656 18080 7708 18086
rect 7656 18022 7708 18028
rect 7668 17241 7696 18022
rect 7654 17232 7710 17241
rect 7760 17202 7788 19207
rect 7852 17678 7880 21286
rect 8220 21010 8248 21626
rect 8312 21078 8340 21898
rect 8300 21072 8352 21078
rect 8300 21014 8352 21020
rect 8208 21004 8260 21010
rect 8208 20946 8260 20952
rect 8298 20904 8354 20913
rect 8298 20839 8300 20848
rect 8352 20839 8354 20848
rect 8300 20810 8352 20816
rect 7950 20700 8258 20709
rect 7950 20698 7956 20700
rect 8012 20698 8036 20700
rect 8092 20698 8116 20700
rect 8172 20698 8196 20700
rect 8252 20698 8258 20700
rect 8012 20646 8014 20698
rect 8194 20646 8196 20698
rect 7950 20644 7956 20646
rect 8012 20644 8036 20646
rect 8092 20644 8116 20646
rect 8172 20644 8196 20646
rect 8252 20644 8258 20646
rect 7950 20635 8258 20644
rect 8404 20398 8432 23151
rect 8576 23122 8628 23128
rect 8574 23080 8630 23089
rect 8574 23015 8630 23024
rect 8482 21720 8538 21729
rect 8482 21655 8484 21664
rect 8536 21655 8538 21664
rect 8484 21626 8536 21632
rect 8484 21072 8536 21078
rect 8484 21014 8536 21020
rect 8392 20392 8444 20398
rect 8392 20334 8444 20340
rect 8392 20256 8444 20262
rect 8392 20198 8444 20204
rect 8298 19816 8354 19825
rect 8298 19751 8300 19760
rect 8352 19751 8354 19760
rect 8300 19722 8352 19728
rect 7950 19612 8258 19621
rect 7950 19610 7956 19612
rect 8012 19610 8036 19612
rect 8092 19610 8116 19612
rect 8172 19610 8196 19612
rect 8252 19610 8258 19612
rect 8012 19558 8014 19610
rect 8194 19558 8196 19610
rect 7950 19556 7956 19558
rect 8012 19556 8036 19558
rect 8092 19556 8116 19558
rect 8172 19556 8196 19558
rect 8252 19556 8258 19558
rect 7950 19547 8258 19556
rect 8300 19440 8352 19446
rect 8300 19382 8352 19388
rect 8208 19236 8260 19242
rect 8208 19178 8260 19184
rect 7932 19168 7984 19174
rect 7932 19110 7984 19116
rect 7944 18698 7972 19110
rect 8116 18896 8168 18902
rect 8116 18838 8168 18844
rect 8128 18737 8156 18838
rect 8114 18728 8170 18737
rect 7932 18692 7984 18698
rect 8114 18663 8170 18672
rect 7932 18634 7984 18640
rect 8220 18612 8248 19178
rect 8312 18970 8340 19382
rect 8300 18964 8352 18970
rect 8300 18906 8352 18912
rect 8404 18766 8432 20198
rect 8392 18760 8444 18766
rect 8392 18702 8444 18708
rect 8220 18584 8340 18612
rect 7950 18524 8258 18533
rect 7950 18522 7956 18524
rect 8012 18522 8036 18524
rect 8092 18522 8116 18524
rect 8172 18522 8196 18524
rect 8252 18522 8258 18524
rect 8012 18470 8014 18522
rect 8194 18470 8196 18522
rect 7950 18468 7956 18470
rect 8012 18468 8036 18470
rect 8092 18468 8116 18470
rect 8172 18468 8196 18470
rect 8252 18468 8258 18470
rect 7950 18459 8258 18468
rect 7840 17672 7892 17678
rect 7840 17614 7892 17620
rect 8312 17610 8340 18584
rect 8496 18290 8524 21014
rect 8588 18358 8616 23015
rect 8680 19242 8708 23695
rect 8772 22710 8800 26302
rect 9034 26200 9090 26302
rect 9402 26200 9458 27000
rect 9770 26330 9826 27000
rect 9588 26308 9640 26314
rect 9588 26250 9640 26256
rect 9692 26302 9826 26330
rect 8852 24336 8904 24342
rect 8852 24278 8904 24284
rect 8760 22704 8812 22710
rect 8760 22646 8812 22652
rect 8758 21040 8814 21049
rect 8758 20975 8814 20984
rect 8772 20874 8800 20975
rect 8760 20868 8812 20874
rect 8760 20810 8812 20816
rect 8668 19236 8720 19242
rect 8668 19178 8720 19184
rect 8864 18714 8892 24278
rect 9312 24200 9364 24206
rect 9312 24142 9364 24148
rect 9128 24064 9180 24070
rect 9128 24006 9180 24012
rect 9140 23497 9168 24006
rect 9324 23866 9352 24142
rect 9312 23860 9364 23866
rect 9312 23802 9364 23808
rect 9126 23488 9182 23497
rect 9126 23423 9182 23432
rect 9416 23254 9444 26200
rect 9496 23520 9548 23526
rect 9496 23462 9548 23468
rect 9404 23248 9456 23254
rect 9404 23190 9456 23196
rect 9036 22568 9088 22574
rect 9036 22510 9088 22516
rect 9048 22098 9076 22510
rect 9404 22432 9456 22438
rect 9404 22374 9456 22380
rect 9416 22166 9444 22374
rect 9404 22160 9456 22166
rect 9404 22102 9456 22108
rect 9036 22092 9088 22098
rect 9036 22034 9088 22040
rect 9048 21554 9076 22034
rect 9312 21888 9364 21894
rect 9312 21830 9364 21836
rect 9036 21548 9088 21554
rect 9036 21490 9088 21496
rect 8944 20800 8996 20806
rect 8944 20742 8996 20748
rect 8956 20534 8984 20742
rect 8944 20528 8996 20534
rect 8944 20470 8996 20476
rect 8956 20398 8984 20470
rect 9048 20466 9076 21490
rect 9324 20505 9352 21830
rect 9404 21616 9456 21622
rect 9404 21558 9456 21564
rect 9310 20496 9366 20505
rect 9036 20460 9088 20466
rect 9310 20431 9366 20440
rect 9036 20402 9088 20408
rect 8944 20392 8996 20398
rect 8944 20334 8996 20340
rect 9048 19378 9076 20402
rect 9416 20262 9444 21558
rect 9404 20256 9456 20262
rect 9404 20198 9456 20204
rect 9508 19938 9536 23462
rect 9416 19910 9536 19938
rect 9128 19712 9180 19718
rect 9128 19654 9180 19660
rect 9036 19372 9088 19378
rect 8680 18686 8892 18714
rect 8956 19332 9036 19360
rect 8576 18352 8628 18358
rect 8576 18294 8628 18300
rect 8484 18284 8536 18290
rect 8484 18226 8536 18232
rect 8300 17604 8352 17610
rect 8300 17546 8352 17552
rect 8392 17536 8444 17542
rect 8392 17478 8444 17484
rect 7950 17436 8258 17445
rect 7950 17434 7956 17436
rect 8012 17434 8036 17436
rect 8092 17434 8116 17436
rect 8172 17434 8196 17436
rect 8252 17434 8258 17436
rect 8012 17382 8014 17434
rect 8194 17382 8196 17434
rect 7950 17380 7956 17382
rect 8012 17380 8036 17382
rect 8092 17380 8116 17382
rect 8172 17380 8196 17382
rect 8252 17380 8258 17382
rect 7950 17371 8258 17380
rect 8404 17338 8432 17478
rect 8392 17332 8444 17338
rect 8392 17274 8444 17280
rect 7654 17167 7710 17176
rect 7748 17196 7800 17202
rect 7748 17138 7800 17144
rect 7930 17096 7986 17105
rect 8680 17066 8708 18686
rect 8852 18624 8904 18630
rect 8852 18566 8904 18572
rect 8758 17368 8814 17377
rect 8758 17303 8814 17312
rect 8772 17202 8800 17303
rect 8760 17196 8812 17202
rect 8760 17138 8812 17144
rect 7930 17031 7986 17040
rect 8668 17060 8720 17066
rect 7944 16590 7972 17031
rect 8668 17002 8720 17008
rect 8392 16788 8444 16794
rect 8392 16730 8444 16736
rect 7932 16584 7984 16590
rect 7932 16526 7984 16532
rect 8404 16425 8432 16730
rect 8576 16584 8628 16590
rect 8576 16526 8628 16532
rect 8390 16416 8446 16425
rect 7950 16348 8258 16357
rect 8390 16351 8446 16360
rect 7950 16346 7956 16348
rect 8012 16346 8036 16348
rect 8092 16346 8116 16348
rect 8172 16346 8196 16348
rect 8252 16346 8258 16348
rect 8012 16294 8014 16346
rect 8194 16294 8196 16346
rect 7950 16292 7956 16294
rect 8012 16292 8036 16294
rect 8092 16292 8116 16294
rect 8172 16292 8196 16294
rect 8252 16292 8258 16294
rect 7950 16283 8258 16292
rect 8484 15904 8536 15910
rect 8484 15846 8536 15852
rect 8588 15858 8616 16526
rect 8772 16250 8800 17138
rect 8760 16244 8812 16250
rect 8760 16186 8812 16192
rect 7564 15360 7616 15366
rect 7564 15302 7616 15308
rect 7950 15260 8258 15269
rect 7950 15258 7956 15260
rect 8012 15258 8036 15260
rect 8092 15258 8116 15260
rect 8172 15258 8196 15260
rect 8252 15258 8258 15260
rect 8012 15206 8014 15258
rect 8194 15206 8196 15258
rect 7950 15204 7956 15206
rect 8012 15204 8036 15206
rect 8092 15204 8116 15206
rect 8172 15204 8196 15206
rect 8252 15204 8258 15206
rect 7950 15195 8258 15204
rect 7950 14172 8258 14181
rect 7950 14170 7956 14172
rect 8012 14170 8036 14172
rect 8092 14170 8116 14172
rect 8172 14170 8196 14172
rect 8252 14170 8258 14172
rect 8012 14118 8014 14170
rect 8194 14118 8196 14170
rect 7950 14116 7956 14118
rect 8012 14116 8036 14118
rect 8092 14116 8116 14118
rect 8172 14116 8196 14118
rect 8252 14116 8258 14118
rect 7950 14107 8258 14116
rect 7378 13832 7434 13841
rect 7378 13767 7434 13776
rect 7950 13084 8258 13093
rect 7950 13082 7956 13084
rect 8012 13082 8036 13084
rect 8092 13082 8116 13084
rect 8172 13082 8196 13084
rect 8252 13082 8258 13084
rect 8012 13030 8014 13082
rect 8194 13030 8196 13082
rect 7950 13028 7956 13030
rect 8012 13028 8036 13030
rect 8092 13028 8116 13030
rect 8172 13028 8196 13030
rect 8252 13028 8258 13030
rect 7950 13019 8258 13028
rect 6734 12880 6790 12889
rect 6734 12815 6790 12824
rect 4068 12436 4120 12442
rect 4068 12378 4120 12384
rect 7950 11996 8258 12005
rect 7950 11994 7956 11996
rect 8012 11994 8036 11996
rect 8092 11994 8116 11996
rect 8172 11994 8196 11996
rect 8252 11994 8258 11996
rect 8012 11942 8014 11994
rect 8194 11942 8196 11994
rect 7950 11940 7956 11942
rect 8012 11940 8036 11942
rect 8092 11940 8116 11942
rect 8172 11940 8196 11942
rect 8252 11940 8258 11942
rect 7950 11931 8258 11940
rect 2950 11452 3258 11461
rect 2950 11450 2956 11452
rect 3012 11450 3036 11452
rect 3092 11450 3116 11452
rect 3172 11450 3196 11452
rect 3252 11450 3258 11452
rect 3012 11398 3014 11450
rect 3194 11398 3196 11450
rect 2950 11396 2956 11398
rect 3012 11396 3036 11398
rect 3092 11396 3116 11398
rect 3172 11396 3196 11398
rect 3252 11396 3258 11398
rect 2950 11387 3258 11396
rect 7950 10908 8258 10917
rect 7950 10906 7956 10908
rect 8012 10906 8036 10908
rect 8092 10906 8116 10908
rect 8172 10906 8196 10908
rect 8252 10906 8258 10908
rect 8012 10854 8014 10906
rect 8194 10854 8196 10906
rect 7950 10852 7956 10854
rect 8012 10852 8036 10854
rect 8092 10852 8116 10854
rect 8172 10852 8196 10854
rect 8252 10852 8258 10854
rect 7950 10843 8258 10852
rect 2950 10364 3258 10373
rect 2950 10362 2956 10364
rect 3012 10362 3036 10364
rect 3092 10362 3116 10364
rect 3172 10362 3196 10364
rect 3252 10362 3258 10364
rect 3012 10310 3014 10362
rect 3194 10310 3196 10362
rect 2950 10308 2956 10310
rect 3012 10308 3036 10310
rect 3092 10308 3116 10310
rect 3172 10308 3196 10310
rect 3252 10308 3258 10310
rect 2950 10299 3258 10308
rect 7950 9820 8258 9829
rect 7950 9818 7956 9820
rect 8012 9818 8036 9820
rect 8092 9818 8116 9820
rect 8172 9818 8196 9820
rect 8252 9818 8258 9820
rect 8012 9766 8014 9818
rect 8194 9766 8196 9818
rect 7950 9764 7956 9766
rect 8012 9764 8036 9766
rect 8092 9764 8116 9766
rect 8172 9764 8196 9766
rect 8252 9764 8258 9766
rect 7950 9755 8258 9764
rect 8496 9586 8524 15846
rect 8588 15830 8800 15858
rect 8772 15502 8800 15830
rect 8760 15496 8812 15502
rect 8758 15464 8760 15473
rect 8812 15464 8814 15473
rect 8758 15399 8814 15408
rect 8576 12436 8628 12442
rect 8864 12434 8892 18566
rect 8956 18290 8984 19332
rect 9036 19314 9088 19320
rect 9140 18766 9168 19654
rect 9220 19440 9272 19446
rect 9220 19382 9272 19388
rect 9128 18760 9180 18766
rect 9128 18702 9180 18708
rect 8944 18284 8996 18290
rect 8944 18226 8996 18232
rect 8956 17746 8984 18226
rect 9126 17912 9182 17921
rect 9126 17847 9182 17856
rect 8944 17740 8996 17746
rect 8944 17682 8996 17688
rect 8956 17202 8984 17682
rect 9140 17542 9168 17847
rect 9128 17536 9180 17542
rect 9128 17478 9180 17484
rect 8944 17196 8996 17202
rect 8944 17138 8996 17144
rect 9126 16688 9182 16697
rect 9126 16623 9128 16632
rect 9180 16623 9182 16632
rect 9128 16594 9180 16600
rect 9232 16250 9260 19382
rect 9312 18692 9364 18698
rect 9312 18634 9364 18640
rect 9324 18222 9352 18634
rect 9312 18216 9364 18222
rect 9312 18158 9364 18164
rect 9312 17536 9364 17542
rect 9312 17478 9364 17484
rect 9324 17105 9352 17478
rect 9416 17270 9444 19910
rect 9496 19168 9548 19174
rect 9496 19110 9548 19116
rect 9508 18902 9536 19110
rect 9496 18896 9548 18902
rect 9496 18838 9548 18844
rect 9496 18624 9548 18630
rect 9496 18566 9548 18572
rect 9404 17264 9456 17270
rect 9404 17206 9456 17212
rect 9310 17096 9366 17105
rect 9310 17031 9366 17040
rect 9508 16998 9536 18566
rect 9496 16992 9548 16998
rect 9496 16934 9548 16940
rect 9600 16794 9628 26250
rect 9692 24274 9720 26302
rect 9770 26200 9826 26302
rect 10138 26200 10194 27000
rect 10506 26200 10562 27000
rect 10874 26200 10930 27000
rect 11242 26330 11298 27000
rect 11072 26302 11298 26330
rect 9864 24948 9916 24954
rect 9864 24890 9916 24896
rect 9772 24812 9824 24818
rect 9772 24754 9824 24760
rect 9680 24268 9732 24274
rect 9680 24210 9732 24216
rect 9784 24177 9812 24754
rect 9770 24168 9826 24177
rect 9770 24103 9826 24112
rect 9680 22704 9732 22710
rect 9680 22646 9732 22652
rect 9772 22704 9824 22710
rect 9772 22646 9824 22652
rect 9692 21865 9720 22646
rect 9678 21856 9734 21865
rect 9678 21791 9734 21800
rect 9784 21622 9812 22646
rect 9772 21616 9824 21622
rect 9772 21558 9824 21564
rect 9784 20534 9812 21558
rect 9772 20528 9824 20534
rect 9772 20470 9824 20476
rect 9784 19446 9812 20470
rect 9772 19440 9824 19446
rect 9678 19408 9734 19417
rect 9772 19382 9824 19388
rect 9678 19343 9734 19352
rect 9692 18970 9720 19343
rect 9680 18964 9732 18970
rect 9680 18906 9732 18912
rect 9784 18766 9812 19382
rect 9772 18760 9824 18766
rect 9772 18702 9824 18708
rect 9784 18358 9812 18702
rect 9772 18352 9824 18358
rect 9772 18294 9824 18300
rect 9772 18080 9824 18086
rect 9772 18022 9824 18028
rect 9678 17912 9734 17921
rect 9678 17847 9734 17856
rect 9692 17814 9720 17847
rect 9680 17808 9732 17814
rect 9680 17750 9732 17756
rect 9784 17270 9812 18022
rect 9772 17264 9824 17270
rect 9772 17206 9824 17212
rect 9678 17096 9734 17105
rect 9678 17031 9734 17040
rect 9312 16788 9364 16794
rect 9312 16730 9364 16736
rect 9588 16788 9640 16794
rect 9588 16730 9640 16736
rect 9220 16244 9272 16250
rect 9220 16186 9272 16192
rect 9324 16114 9352 16730
rect 9692 16674 9720 17031
rect 9772 16788 9824 16794
rect 9772 16730 9824 16736
rect 9784 16697 9812 16730
rect 9600 16646 9720 16674
rect 9770 16688 9826 16697
rect 9600 16590 9628 16646
rect 9770 16623 9826 16632
rect 9588 16584 9640 16590
rect 9588 16526 9640 16532
rect 9404 16448 9456 16454
rect 9680 16448 9732 16454
rect 9456 16396 9680 16402
rect 9404 16390 9732 16396
rect 9416 16374 9720 16390
rect 9312 16108 9364 16114
rect 9312 16050 9364 16056
rect 9588 16040 9640 16046
rect 9126 16008 9182 16017
rect 9588 15982 9640 15988
rect 9126 15943 9128 15952
rect 9180 15943 9182 15952
rect 9128 15914 9180 15920
rect 9600 15609 9628 15982
rect 9772 15972 9824 15978
rect 9772 15914 9824 15920
rect 9402 15600 9458 15609
rect 9402 15535 9458 15544
rect 9586 15600 9642 15609
rect 9586 15535 9642 15544
rect 9416 15502 9444 15535
rect 9404 15496 9456 15502
rect 9404 15438 9456 15444
rect 9416 15162 9444 15438
rect 9784 15337 9812 15914
rect 9876 15706 9904 24890
rect 10152 23798 10180 26200
rect 10140 23792 10192 23798
rect 10140 23734 10192 23740
rect 9956 23724 10008 23730
rect 9956 23666 10008 23672
rect 9968 22710 9996 23666
rect 10520 23186 10548 26200
rect 10888 23798 10916 26200
rect 11072 24834 11100 26302
rect 11242 26200 11298 26302
rect 11610 26200 11666 27000
rect 11978 26200 12034 27000
rect 12346 26200 12402 27000
rect 12714 26330 12770 27000
rect 13082 26330 13138 27000
rect 12714 26302 12848 26330
rect 12714 26200 12770 26302
rect 10980 24806 11100 24834
rect 10980 24274 11008 24806
rect 10968 24268 11020 24274
rect 10968 24210 11020 24216
rect 11336 24064 11388 24070
rect 11336 24006 11388 24012
rect 10876 23792 10928 23798
rect 10876 23734 10928 23740
rect 11060 23656 11112 23662
rect 11060 23598 11112 23604
rect 10508 23180 10560 23186
rect 10508 23122 10560 23128
rect 11072 22710 11100 23598
rect 9956 22704 10008 22710
rect 9956 22646 10008 22652
rect 11060 22704 11112 22710
rect 11060 22646 11112 22652
rect 11152 22432 11204 22438
rect 11152 22374 11204 22380
rect 11244 22432 11296 22438
rect 11244 22374 11296 22380
rect 10600 22228 10652 22234
rect 10600 22170 10652 22176
rect 10230 21992 10286 22001
rect 10230 21927 10286 21936
rect 10048 21888 10100 21894
rect 10048 21830 10100 21836
rect 10060 21690 10088 21830
rect 10048 21684 10100 21690
rect 10048 21626 10100 21632
rect 10140 20596 10192 20602
rect 10140 20538 10192 20544
rect 10152 19689 10180 20538
rect 10138 19680 10194 19689
rect 10138 19615 10194 19624
rect 10048 18828 10100 18834
rect 10048 18770 10100 18776
rect 10060 17610 10088 18770
rect 10138 18456 10194 18465
rect 10138 18391 10194 18400
rect 9956 17604 10008 17610
rect 9956 17546 10008 17552
rect 10048 17604 10100 17610
rect 10048 17546 10100 17552
rect 9968 16998 9996 17546
rect 10060 17134 10088 17546
rect 10048 17128 10100 17134
rect 10048 17070 10100 17076
rect 9956 16992 10008 16998
rect 9956 16934 10008 16940
rect 9954 16688 10010 16697
rect 9954 16623 9956 16632
rect 10008 16623 10010 16632
rect 9956 16594 10008 16600
rect 9968 16114 9996 16594
rect 10152 16538 10180 18391
rect 10060 16510 10180 16538
rect 10060 16454 10088 16510
rect 10048 16448 10100 16454
rect 10048 16390 10100 16396
rect 10140 16448 10192 16454
rect 10140 16390 10192 16396
rect 10152 16250 10180 16390
rect 10140 16244 10192 16250
rect 10140 16186 10192 16192
rect 9956 16108 10008 16114
rect 9956 16050 10008 16056
rect 9864 15700 9916 15706
rect 9864 15642 9916 15648
rect 10244 15502 10272 21927
rect 10508 21344 10560 21350
rect 10508 21286 10560 21292
rect 10324 21140 10376 21146
rect 10324 21082 10376 21088
rect 10336 20602 10364 21082
rect 10520 21010 10548 21286
rect 10508 21004 10560 21010
rect 10508 20946 10560 20952
rect 10324 20596 10376 20602
rect 10324 20538 10376 20544
rect 10520 20398 10548 20946
rect 10612 20641 10640 22170
rect 11060 22092 11112 22098
rect 11060 22034 11112 22040
rect 10692 21412 10744 21418
rect 10692 21354 10744 21360
rect 10598 20632 10654 20641
rect 10598 20567 10654 20576
rect 10508 20392 10560 20398
rect 10508 20334 10560 20340
rect 10324 19236 10376 19242
rect 10324 19178 10376 19184
rect 10336 18766 10364 19178
rect 10324 18760 10376 18766
rect 10324 18702 10376 18708
rect 10336 17610 10364 18702
rect 10508 18624 10560 18630
rect 10508 18566 10560 18572
rect 10520 18290 10548 18566
rect 10600 18352 10652 18358
rect 10600 18294 10652 18300
rect 10508 18284 10560 18290
rect 10508 18226 10560 18232
rect 10324 17604 10376 17610
rect 10324 17546 10376 17552
rect 10508 17604 10560 17610
rect 10612 17592 10640 18294
rect 10560 17564 10640 17592
rect 10508 17546 10560 17552
rect 10612 17202 10640 17564
rect 10600 17196 10652 17202
rect 10600 17138 10652 17144
rect 10704 16794 10732 21354
rect 11072 21010 11100 22034
rect 11164 21554 11192 22374
rect 11152 21548 11204 21554
rect 11152 21490 11204 21496
rect 11152 21344 11204 21350
rect 11152 21286 11204 21292
rect 11060 21004 11112 21010
rect 11060 20946 11112 20952
rect 11058 20768 11114 20777
rect 11058 20703 11114 20712
rect 10784 20596 10836 20602
rect 10784 20538 10836 20544
rect 10796 20262 10824 20538
rect 10784 20256 10836 20262
rect 10784 20198 10836 20204
rect 10796 19310 10824 20198
rect 10968 19916 11020 19922
rect 10968 19858 11020 19864
rect 10876 19712 10928 19718
rect 10876 19654 10928 19660
rect 10784 19304 10836 19310
rect 10784 19246 10836 19252
rect 10784 19168 10836 19174
rect 10784 19110 10836 19116
rect 10796 18426 10824 19110
rect 10784 18420 10836 18426
rect 10784 18362 10836 18368
rect 10692 16788 10744 16794
rect 10692 16730 10744 16736
rect 10888 16590 10916 19654
rect 10980 19174 11008 19858
rect 11072 19854 11100 20703
rect 11164 20534 11192 21286
rect 11152 20528 11204 20534
rect 11152 20470 11204 20476
rect 11060 19848 11112 19854
rect 11060 19790 11112 19796
rect 11256 19666 11284 22374
rect 11348 21049 11376 24006
rect 11520 23860 11572 23866
rect 11520 23802 11572 23808
rect 11532 23594 11560 23802
rect 11520 23588 11572 23594
rect 11520 23530 11572 23536
rect 11518 23488 11574 23497
rect 11518 23423 11574 23432
rect 11532 22094 11560 23423
rect 11624 23186 11652 26200
rect 11796 24268 11848 24274
rect 11796 24210 11848 24216
rect 11704 23520 11756 23526
rect 11704 23462 11756 23468
rect 11716 23254 11744 23462
rect 11704 23248 11756 23254
rect 11704 23190 11756 23196
rect 11612 23180 11664 23186
rect 11612 23122 11664 23128
rect 11532 22066 11652 22094
rect 11428 21412 11480 21418
rect 11428 21354 11480 21360
rect 11334 21040 11390 21049
rect 11440 21010 11468 21354
rect 11334 20975 11390 20984
rect 11428 21004 11480 21010
rect 11428 20946 11480 20952
rect 11334 20496 11390 20505
rect 11334 20431 11390 20440
rect 11518 20496 11574 20505
rect 11518 20431 11574 20440
rect 11072 19638 11284 19666
rect 10968 19168 11020 19174
rect 10968 19110 11020 19116
rect 10968 18420 11020 18426
rect 10968 18362 11020 18368
rect 10876 16584 10928 16590
rect 10876 16526 10928 16532
rect 10784 16448 10836 16454
rect 10784 16390 10836 16396
rect 10796 16046 10824 16390
rect 10784 16040 10836 16046
rect 10784 15982 10836 15988
rect 10980 15706 11008 18362
rect 11072 16998 11100 19638
rect 11244 19168 11296 19174
rect 11244 19110 11296 19116
rect 11152 18828 11204 18834
rect 11152 18770 11204 18776
rect 11164 18086 11192 18770
rect 11152 18080 11204 18086
rect 11152 18022 11204 18028
rect 11060 16992 11112 16998
rect 11060 16934 11112 16940
rect 11164 16810 11192 18022
rect 11256 17921 11284 19110
rect 11242 17912 11298 17921
rect 11242 17847 11298 17856
rect 11244 17808 11296 17814
rect 11244 17750 11296 17756
rect 11072 16782 11192 16810
rect 11072 16658 11100 16782
rect 11152 16720 11204 16726
rect 11256 16674 11284 17750
rect 11204 16668 11284 16674
rect 11152 16662 11284 16668
rect 11060 16652 11112 16658
rect 11164 16646 11284 16662
rect 11060 16594 11112 16600
rect 11058 16552 11114 16561
rect 11058 16487 11060 16496
rect 11112 16487 11114 16496
rect 11060 16458 11112 16464
rect 11060 16040 11112 16046
rect 11060 15982 11112 15988
rect 10968 15700 11020 15706
rect 10968 15642 11020 15648
rect 10232 15496 10284 15502
rect 10232 15438 10284 15444
rect 9770 15328 9826 15337
rect 9770 15263 9826 15272
rect 10244 15162 10272 15438
rect 10692 15428 10744 15434
rect 10692 15370 10744 15376
rect 9404 15156 9456 15162
rect 9404 15098 9456 15104
rect 10232 15156 10284 15162
rect 10232 15098 10284 15104
rect 10506 15056 10562 15065
rect 10506 14991 10508 15000
rect 10560 14991 10562 15000
rect 10508 14962 10560 14968
rect 10048 14816 10100 14822
rect 10048 14758 10100 14764
rect 10060 14278 10088 14758
rect 10520 14618 10548 14962
rect 10704 14958 10732 15370
rect 11072 15162 11100 15982
rect 11152 15700 11204 15706
rect 11152 15642 11204 15648
rect 11164 15366 11192 15642
rect 11152 15360 11204 15366
rect 11152 15302 11204 15308
rect 10968 15156 11020 15162
rect 10968 15098 11020 15104
rect 11060 15156 11112 15162
rect 11060 15098 11112 15104
rect 10980 15065 11008 15098
rect 10966 15056 11022 15065
rect 10966 14991 11022 15000
rect 11152 15020 11204 15026
rect 11152 14962 11204 14968
rect 10692 14952 10744 14958
rect 10692 14894 10744 14900
rect 10508 14612 10560 14618
rect 10508 14554 10560 14560
rect 10704 14414 10732 14894
rect 11164 14618 11192 14962
rect 11152 14612 11204 14618
rect 11152 14554 11204 14560
rect 10692 14408 10744 14414
rect 10692 14350 10744 14356
rect 10048 14272 10100 14278
rect 10048 14214 10100 14220
rect 10704 13190 10732 14350
rect 10048 13184 10100 13190
rect 10048 13126 10100 13132
rect 10692 13184 10744 13190
rect 10692 13126 10744 13132
rect 8628 12406 8892 12434
rect 8576 12378 8628 12384
rect 8484 9580 8536 9586
rect 8484 9522 8536 9528
rect 2950 9276 3258 9285
rect 2950 9274 2956 9276
rect 3012 9274 3036 9276
rect 3092 9274 3116 9276
rect 3172 9274 3196 9276
rect 3252 9274 3258 9276
rect 3012 9222 3014 9274
rect 3194 9222 3196 9274
rect 2950 9220 2956 9222
rect 3012 9220 3036 9222
rect 3092 9220 3116 9222
rect 3172 9220 3196 9222
rect 3252 9220 3258 9222
rect 2950 9211 3258 9220
rect 10060 9042 10088 13126
rect 11348 12345 11376 20431
rect 11532 20233 11560 20431
rect 11518 20224 11574 20233
rect 11518 20159 11574 20168
rect 11520 19712 11572 19718
rect 11520 19654 11572 19660
rect 11426 19408 11482 19417
rect 11426 19343 11482 19352
rect 11440 19242 11468 19343
rect 11428 19236 11480 19242
rect 11428 19178 11480 19184
rect 11426 18592 11482 18601
rect 11426 18527 11482 18536
rect 11440 17542 11468 18527
rect 11428 17536 11480 17542
rect 11428 17478 11480 17484
rect 11440 17270 11468 17478
rect 11428 17264 11480 17270
rect 11428 17206 11480 17212
rect 11532 16969 11560 19654
rect 11518 16960 11574 16969
rect 11518 16895 11574 16904
rect 11428 16108 11480 16114
rect 11428 16050 11480 16056
rect 11440 15366 11468 16050
rect 11428 15360 11480 15366
rect 11428 15302 11480 15308
rect 11624 14521 11652 22066
rect 11704 22092 11756 22098
rect 11704 22034 11756 22040
rect 11716 21962 11744 22034
rect 11704 21956 11756 21962
rect 11704 21898 11756 21904
rect 11716 21350 11744 21898
rect 11704 21344 11756 21350
rect 11704 21286 11756 21292
rect 11808 19718 11836 24210
rect 11888 23792 11940 23798
rect 11888 23734 11940 23740
rect 11900 23361 11928 23734
rect 11992 23662 12020 26200
rect 12360 24342 12388 26200
rect 12348 24336 12400 24342
rect 12348 24278 12400 24284
rect 11980 23656 12032 23662
rect 11980 23598 12032 23604
rect 12452 23446 12756 23474
rect 11886 23352 11942 23361
rect 12452 23322 12480 23446
rect 11886 23287 11942 23296
rect 11980 23316 12032 23322
rect 12348 23316 12400 23322
rect 11980 23258 12032 23264
rect 12084 23276 12348 23304
rect 11992 23050 12020 23258
rect 11980 23044 12032 23050
rect 11980 22986 12032 22992
rect 11888 22976 11940 22982
rect 11888 22918 11940 22924
rect 11900 21593 11928 22918
rect 12084 22506 12112 23276
rect 12348 23258 12400 23264
rect 12440 23316 12492 23322
rect 12440 23258 12492 23264
rect 12728 23118 12756 23446
rect 12716 23112 12768 23118
rect 12716 23054 12768 23060
rect 12162 22944 12218 22953
rect 12162 22879 12218 22888
rect 12072 22500 12124 22506
rect 12072 22442 12124 22448
rect 12176 21672 12204 22879
rect 12716 22636 12768 22642
rect 12716 22578 12768 22584
rect 12440 22500 12492 22506
rect 12440 22442 12492 22448
rect 12624 22500 12676 22506
rect 12624 22442 12676 22448
rect 12256 22160 12308 22166
rect 12256 22102 12308 22108
rect 12268 21894 12296 22102
rect 12452 22098 12480 22442
rect 12532 22432 12584 22438
rect 12532 22374 12584 22380
rect 12440 22092 12492 22098
rect 12440 22034 12492 22040
rect 12440 21956 12492 21962
rect 12440 21898 12492 21904
rect 12256 21888 12308 21894
rect 12256 21830 12308 21836
rect 12346 21856 12402 21865
rect 12346 21791 12402 21800
rect 12084 21644 12204 21672
rect 11886 21584 11942 21593
rect 11886 21519 11942 21528
rect 11980 21344 12032 21350
rect 11980 21286 12032 21292
rect 11888 20868 11940 20874
rect 11888 20810 11940 20816
rect 11900 20534 11928 20810
rect 11888 20528 11940 20534
rect 11888 20470 11940 20476
rect 11796 19712 11848 19718
rect 11796 19654 11848 19660
rect 11900 19417 11928 20470
rect 11886 19408 11942 19417
rect 11886 19343 11942 19352
rect 11796 19168 11848 19174
rect 11796 19110 11848 19116
rect 11888 19168 11940 19174
rect 11888 19110 11940 19116
rect 11808 18766 11836 19110
rect 11900 18902 11928 19110
rect 11888 18896 11940 18902
rect 11888 18838 11940 18844
rect 11796 18760 11848 18766
rect 11796 18702 11848 18708
rect 11888 18760 11940 18766
rect 11888 18702 11940 18708
rect 11704 18624 11756 18630
rect 11704 18566 11756 18572
rect 11716 17746 11744 18566
rect 11808 18358 11836 18702
rect 11900 18426 11928 18702
rect 11888 18420 11940 18426
rect 11888 18362 11940 18368
rect 11796 18352 11848 18358
rect 11796 18294 11848 18300
rect 11992 17898 12020 21286
rect 12084 19394 12112 21644
rect 12162 21584 12218 21593
rect 12162 21519 12218 21528
rect 12176 20398 12204 21519
rect 12360 20924 12388 21791
rect 12452 21729 12480 21898
rect 12438 21720 12494 21729
rect 12438 21655 12494 21664
rect 12438 21584 12494 21593
rect 12438 21519 12494 21528
rect 12452 21332 12480 21519
rect 12544 21486 12572 22374
rect 12532 21480 12584 21486
rect 12532 21422 12584 21428
rect 12452 21304 12572 21332
rect 12544 21049 12572 21304
rect 12530 21040 12586 21049
rect 12530 20975 12586 20984
rect 12360 20896 12572 20924
rect 12440 20800 12492 20806
rect 12440 20742 12492 20748
rect 12452 20602 12480 20742
rect 12544 20602 12572 20896
rect 12348 20596 12400 20602
rect 12348 20538 12400 20544
rect 12440 20596 12492 20602
rect 12440 20538 12492 20544
rect 12532 20596 12584 20602
rect 12532 20538 12584 20544
rect 12164 20392 12216 20398
rect 12164 20334 12216 20340
rect 12176 19514 12204 20334
rect 12256 20256 12308 20262
rect 12256 20198 12308 20204
rect 12268 19922 12296 20198
rect 12360 19922 12388 20538
rect 12256 19916 12308 19922
rect 12256 19858 12308 19864
rect 12348 19916 12400 19922
rect 12348 19858 12400 19864
rect 12164 19508 12216 19514
rect 12164 19450 12216 19456
rect 12084 19366 12204 19394
rect 12268 19378 12296 19858
rect 12348 19508 12400 19514
rect 12348 19450 12400 19456
rect 12072 19304 12124 19310
rect 12072 19246 12124 19252
rect 12084 18426 12112 19246
rect 12072 18420 12124 18426
rect 12072 18362 12124 18368
rect 11900 17870 12020 17898
rect 11900 17814 11928 17870
rect 11888 17808 11940 17814
rect 11888 17750 11940 17756
rect 11704 17740 11756 17746
rect 12176 17728 12204 19366
rect 12256 19372 12308 19378
rect 12360 19360 12388 19450
rect 12360 19332 12572 19360
rect 12256 19314 12308 19320
rect 12348 18216 12400 18222
rect 12348 18158 12400 18164
rect 11704 17682 11756 17688
rect 12084 17700 12204 17728
rect 11716 17202 11744 17682
rect 11704 17196 11756 17202
rect 11704 17138 11756 17144
rect 12084 16833 12112 17700
rect 12164 17604 12216 17610
rect 12164 17546 12216 17552
rect 12176 17513 12204 17546
rect 12256 17536 12308 17542
rect 12162 17504 12218 17513
rect 12256 17478 12308 17484
rect 12162 17439 12218 17448
rect 12070 16824 12126 16833
rect 12070 16759 12126 16768
rect 12268 16658 12296 17478
rect 12256 16652 12308 16658
rect 12256 16594 12308 16600
rect 11704 16584 11756 16590
rect 11704 16526 11756 16532
rect 11716 16046 11744 16526
rect 12256 16516 12308 16522
rect 12256 16458 12308 16464
rect 11704 16040 11756 16046
rect 11704 15982 11756 15988
rect 11716 14958 11744 15982
rect 12268 15638 12296 16458
rect 12360 16454 12388 18158
rect 12348 16448 12400 16454
rect 12348 16390 12400 16396
rect 12360 16046 12388 16390
rect 12348 16040 12400 16046
rect 12348 15982 12400 15988
rect 12256 15632 12308 15638
rect 12256 15574 12308 15580
rect 12072 15156 12124 15162
rect 12072 15098 12124 15104
rect 11704 14952 11756 14958
rect 11704 14894 11756 14900
rect 11610 14512 11666 14521
rect 11610 14447 11666 14456
rect 11794 14240 11850 14249
rect 11794 14175 11850 14184
rect 11808 14074 11836 14175
rect 11796 14068 11848 14074
rect 11796 14010 11848 14016
rect 11978 13968 12034 13977
rect 11978 13903 11980 13912
rect 12032 13903 12034 13912
rect 11980 13874 12032 13880
rect 12084 13394 12112 15098
rect 12268 14482 12296 15574
rect 12440 14952 12492 14958
rect 12440 14894 12492 14900
rect 12452 14618 12480 14894
rect 12440 14612 12492 14618
rect 12440 14554 12492 14560
rect 12256 14476 12308 14482
rect 12256 14418 12308 14424
rect 12544 14074 12572 19332
rect 12636 18834 12664 22442
rect 12728 19009 12756 22578
rect 12820 22409 12848 26302
rect 13082 26302 13400 26330
rect 13082 26200 13138 26302
rect 12950 24508 13258 24517
rect 12950 24506 12956 24508
rect 13012 24506 13036 24508
rect 13092 24506 13116 24508
rect 13172 24506 13196 24508
rect 13252 24506 13258 24508
rect 13012 24454 13014 24506
rect 13194 24454 13196 24506
rect 12950 24452 12956 24454
rect 13012 24452 13036 24454
rect 13092 24452 13116 24454
rect 13172 24452 13196 24454
rect 13252 24452 13258 24454
rect 12950 24443 13258 24452
rect 12950 23420 13258 23429
rect 12950 23418 12956 23420
rect 13012 23418 13036 23420
rect 13092 23418 13116 23420
rect 13172 23418 13196 23420
rect 13252 23418 13258 23420
rect 13012 23366 13014 23418
rect 13194 23366 13196 23418
rect 12950 23364 12956 23366
rect 13012 23364 13036 23366
rect 13092 23364 13116 23366
rect 13172 23364 13196 23366
rect 13252 23364 13258 23366
rect 12950 23355 13258 23364
rect 12900 23316 12952 23322
rect 12900 23258 12952 23264
rect 12912 22438 12940 23258
rect 12992 23044 13044 23050
rect 12992 22986 13044 22992
rect 13004 22506 13032 22986
rect 13372 22817 13400 26302
rect 13450 26200 13506 27000
rect 13818 26200 13874 27000
rect 14186 26200 14242 27000
rect 14554 26200 14610 27000
rect 14922 26200 14978 27000
rect 15290 26200 15346 27000
rect 15658 26330 15714 27000
rect 15396 26302 15714 26330
rect 13358 22808 13414 22817
rect 13358 22743 13414 22752
rect 12992 22500 13044 22506
rect 12992 22442 13044 22448
rect 12900 22432 12952 22438
rect 12806 22400 12862 22409
rect 12900 22374 12952 22380
rect 12806 22335 12862 22344
rect 12950 22332 13258 22341
rect 12950 22330 12956 22332
rect 13012 22330 13036 22332
rect 13092 22330 13116 22332
rect 13172 22330 13196 22332
rect 13252 22330 13258 22332
rect 13012 22278 13014 22330
rect 13194 22278 13196 22330
rect 12950 22276 12956 22278
rect 13012 22276 13036 22278
rect 13092 22276 13116 22278
rect 13172 22276 13196 22278
rect 13252 22276 13258 22278
rect 12950 22267 13258 22276
rect 12808 22228 12860 22234
rect 12808 22170 12860 22176
rect 12820 22012 12848 22170
rect 13464 22166 13492 26200
rect 13832 23322 13860 26200
rect 14004 25084 14056 25090
rect 14004 25026 14056 25032
rect 14016 24410 14044 25026
rect 14096 24744 14148 24750
rect 14096 24686 14148 24692
rect 14004 24404 14056 24410
rect 14004 24346 14056 24352
rect 14108 23866 14136 24686
rect 14004 23860 14056 23866
rect 14004 23802 14056 23808
rect 14096 23860 14148 23866
rect 14096 23802 14148 23808
rect 13820 23316 13872 23322
rect 13820 23258 13872 23264
rect 13912 23316 13964 23322
rect 13912 23258 13964 23264
rect 13544 23248 13596 23254
rect 13924 23202 13952 23258
rect 13544 23190 13596 23196
rect 13556 22681 13584 23190
rect 13648 23174 13952 23202
rect 13648 23118 13676 23174
rect 13636 23112 13688 23118
rect 13636 23054 13688 23060
rect 13728 23112 13780 23118
rect 13728 23054 13780 23060
rect 13820 23112 13872 23118
rect 13820 23054 13872 23060
rect 13542 22672 13598 22681
rect 13542 22607 13598 22616
rect 13634 22400 13690 22409
rect 13634 22335 13690 22344
rect 13452 22160 13504 22166
rect 13452 22102 13504 22108
rect 13176 22094 13228 22098
rect 13004 22092 13228 22094
rect 13004 22066 13176 22092
rect 13004 22012 13032 22066
rect 13176 22034 13228 22040
rect 12820 21984 13032 22012
rect 13360 22024 13412 22030
rect 12820 21146 12848 21984
rect 13412 21984 13492 22012
rect 13360 21966 13412 21972
rect 12900 21888 12952 21894
rect 12898 21856 12900 21865
rect 13176 21888 13228 21894
rect 12952 21856 12954 21865
rect 13176 21830 13228 21836
rect 12898 21791 12954 21800
rect 12900 21480 12952 21486
rect 12900 21422 12952 21428
rect 12990 21448 13046 21457
rect 12912 21350 12940 21422
rect 13188 21434 13216 21830
rect 13464 21690 13492 21984
rect 13544 21956 13596 21962
rect 13544 21898 13596 21904
rect 13556 21865 13584 21898
rect 13542 21856 13598 21865
rect 13542 21791 13598 21800
rect 13452 21684 13504 21690
rect 13452 21626 13504 21632
rect 13648 21570 13676 22335
rect 13268 21548 13320 21554
rect 13556 21542 13676 21570
rect 13320 21508 13492 21536
rect 13268 21490 13320 21496
rect 13046 21406 13216 21434
rect 12990 21383 13046 21392
rect 12900 21344 12952 21350
rect 12900 21286 12952 21292
rect 12950 21244 13258 21253
rect 12950 21242 12956 21244
rect 13012 21242 13036 21244
rect 13092 21242 13116 21244
rect 13172 21242 13196 21244
rect 13252 21242 13258 21244
rect 13012 21190 13014 21242
rect 13194 21190 13196 21242
rect 12950 21188 12956 21190
rect 13012 21188 13036 21190
rect 13092 21188 13116 21190
rect 13172 21188 13196 21190
rect 13252 21188 13258 21190
rect 12950 21179 13258 21188
rect 13464 21146 13492 21508
rect 12808 21140 12860 21146
rect 12808 21082 12860 21088
rect 13452 21140 13504 21146
rect 13452 21082 13504 21088
rect 13360 20936 13412 20942
rect 13360 20878 13412 20884
rect 12808 20800 12860 20806
rect 12808 20742 12860 20748
rect 12820 20602 12848 20742
rect 12808 20596 12860 20602
rect 12808 20538 12860 20544
rect 12808 20392 12860 20398
rect 12808 20334 12860 20340
rect 12714 19000 12770 19009
rect 12714 18935 12770 18944
rect 12624 18828 12676 18834
rect 12624 18770 12676 18776
rect 12716 18828 12768 18834
rect 12716 18770 12768 18776
rect 12728 18630 12756 18770
rect 12624 18624 12676 18630
rect 12624 18566 12676 18572
rect 12716 18624 12768 18630
rect 12716 18566 12768 18572
rect 12636 18222 12664 18566
rect 12624 18216 12676 18222
rect 12624 18158 12676 18164
rect 12728 17610 12756 18566
rect 12820 17746 12848 20334
rect 12950 20156 13258 20165
rect 12950 20154 12956 20156
rect 13012 20154 13036 20156
rect 13092 20154 13116 20156
rect 13172 20154 13196 20156
rect 13252 20154 13258 20156
rect 13012 20102 13014 20154
rect 13194 20102 13196 20154
rect 12950 20100 12956 20102
rect 13012 20100 13036 20102
rect 13092 20100 13116 20102
rect 13172 20100 13196 20102
rect 13252 20100 13258 20102
rect 12950 20091 13258 20100
rect 13372 19990 13400 20878
rect 13452 20324 13504 20330
rect 13452 20266 13504 20272
rect 13464 19990 13492 20266
rect 13360 19984 13412 19990
rect 13360 19926 13412 19932
rect 13452 19984 13504 19990
rect 13452 19926 13504 19932
rect 13360 19508 13412 19514
rect 13360 19450 13412 19456
rect 13372 19174 13400 19450
rect 13450 19408 13506 19417
rect 13450 19343 13506 19352
rect 13360 19168 13412 19174
rect 13360 19110 13412 19116
rect 12950 19068 13258 19077
rect 12950 19066 12956 19068
rect 13012 19066 13036 19068
rect 13092 19066 13116 19068
rect 13172 19066 13196 19068
rect 13252 19066 13258 19068
rect 13012 19014 13014 19066
rect 13194 19014 13196 19066
rect 12950 19012 12956 19014
rect 13012 19012 13036 19014
rect 13092 19012 13116 19014
rect 13172 19012 13196 19014
rect 13252 19012 13258 19014
rect 12950 19003 13258 19012
rect 13464 18834 13492 19343
rect 13452 18828 13504 18834
rect 13452 18770 13504 18776
rect 13452 18624 13504 18630
rect 13452 18566 13504 18572
rect 12950 17980 13258 17989
rect 12950 17978 12956 17980
rect 13012 17978 13036 17980
rect 13092 17978 13116 17980
rect 13172 17978 13196 17980
rect 13252 17978 13258 17980
rect 13012 17926 13014 17978
rect 13194 17926 13196 17978
rect 12950 17924 12956 17926
rect 13012 17924 13036 17926
rect 13092 17924 13116 17926
rect 13172 17924 13196 17926
rect 13252 17924 13258 17926
rect 12950 17915 13258 17924
rect 13464 17882 13492 18566
rect 13452 17876 13504 17882
rect 13452 17818 13504 17824
rect 12808 17740 12860 17746
rect 12808 17682 12860 17688
rect 13268 17740 13320 17746
rect 13268 17682 13320 17688
rect 12716 17604 12768 17610
rect 12716 17546 12768 17552
rect 12728 17270 12756 17546
rect 12716 17264 12768 17270
rect 12716 17206 12768 17212
rect 12728 16522 12756 17206
rect 13280 17134 13308 17682
rect 13268 17128 13320 17134
rect 13268 17070 13320 17076
rect 12950 16892 13258 16901
rect 12950 16890 12956 16892
rect 13012 16890 13036 16892
rect 13092 16890 13116 16892
rect 13172 16890 13196 16892
rect 13252 16890 13258 16892
rect 13012 16838 13014 16890
rect 13194 16838 13196 16890
rect 12950 16836 12956 16838
rect 13012 16836 13036 16838
rect 13092 16836 13116 16838
rect 13172 16836 13196 16838
rect 13252 16836 13258 16838
rect 12950 16827 13258 16836
rect 12716 16516 12768 16522
rect 12716 16458 12768 16464
rect 12728 16182 12756 16458
rect 13358 16280 13414 16289
rect 13358 16215 13414 16224
rect 12716 16176 12768 16182
rect 12716 16118 12768 16124
rect 12728 16046 12756 16118
rect 12716 16040 12768 16046
rect 12716 15982 12768 15988
rect 12728 15434 12756 15982
rect 12950 15804 13258 15813
rect 12950 15802 12956 15804
rect 13012 15802 13036 15804
rect 13092 15802 13116 15804
rect 13172 15802 13196 15804
rect 13252 15802 13258 15804
rect 13012 15750 13014 15802
rect 13194 15750 13196 15802
rect 12950 15748 12956 15750
rect 13012 15748 13036 15750
rect 13092 15748 13116 15750
rect 13172 15748 13196 15750
rect 13252 15748 13258 15750
rect 12950 15739 13258 15748
rect 12716 15428 12768 15434
rect 12716 15370 12768 15376
rect 12728 15094 12756 15370
rect 12716 15088 12768 15094
rect 12716 15030 12768 15036
rect 12728 14278 12756 15030
rect 12950 14716 13258 14725
rect 12950 14714 12956 14716
rect 13012 14714 13036 14716
rect 13092 14714 13116 14716
rect 13172 14714 13196 14716
rect 13252 14714 13258 14716
rect 13012 14662 13014 14714
rect 13194 14662 13196 14714
rect 12950 14660 12956 14662
rect 13012 14660 13036 14662
rect 13092 14660 13116 14662
rect 13172 14660 13196 14662
rect 13252 14660 13258 14662
rect 12950 14651 13258 14660
rect 13372 14618 13400 16215
rect 13452 16040 13504 16046
rect 13452 15982 13504 15988
rect 13556 15994 13584 21542
rect 13636 21480 13688 21486
rect 13636 21422 13688 21428
rect 13648 20262 13676 21422
rect 13740 21078 13768 23054
rect 13832 22710 13860 23054
rect 14016 22710 14044 23802
rect 14200 23186 14228 26200
rect 14568 23594 14596 26200
rect 14648 24132 14700 24138
rect 14648 24074 14700 24080
rect 14556 23588 14608 23594
rect 14556 23530 14608 23536
rect 14278 23488 14334 23497
rect 14278 23423 14334 23432
rect 14188 23180 14240 23186
rect 14188 23122 14240 23128
rect 13820 22704 13872 22710
rect 13820 22646 13872 22652
rect 14004 22704 14056 22710
rect 14004 22646 14056 22652
rect 13832 22098 13860 22646
rect 13820 22092 13872 22098
rect 13820 22034 13872 22040
rect 13728 21072 13780 21078
rect 13728 21014 13780 21020
rect 13726 20904 13782 20913
rect 13726 20839 13782 20848
rect 13740 20806 13768 20839
rect 13728 20800 13780 20806
rect 13728 20742 13780 20748
rect 13726 20632 13782 20641
rect 13726 20567 13782 20576
rect 13636 20256 13688 20262
rect 13636 20198 13688 20204
rect 13648 19310 13676 20198
rect 13740 19786 13768 20567
rect 13832 20398 13860 22034
rect 14016 21962 14044 22646
rect 14188 22024 14240 22030
rect 14188 21966 14240 21972
rect 14004 21956 14056 21962
rect 14004 21898 14056 21904
rect 14200 21865 14228 21966
rect 14186 21856 14242 21865
rect 14186 21791 14242 21800
rect 14096 21548 14148 21554
rect 14096 21490 14148 21496
rect 14188 21548 14240 21554
rect 14188 21490 14240 21496
rect 13912 21344 13964 21350
rect 13912 21286 13964 21292
rect 13820 20392 13872 20398
rect 13820 20334 13872 20340
rect 13728 19780 13780 19786
rect 13728 19722 13780 19728
rect 13636 19304 13688 19310
rect 13636 19246 13688 19252
rect 13740 19174 13768 19722
rect 13728 19168 13780 19174
rect 13728 19110 13780 19116
rect 13636 18828 13688 18834
rect 13636 18770 13688 18776
rect 13648 18630 13676 18770
rect 13832 18766 13860 20334
rect 13924 19802 13952 21286
rect 14108 21060 14136 21490
rect 14016 21032 14136 21060
rect 14016 20874 14044 21032
rect 14004 20868 14056 20874
rect 14004 20810 14056 20816
rect 14096 20868 14148 20874
rect 14096 20810 14148 20816
rect 14016 20233 14044 20810
rect 14108 20534 14136 20810
rect 14096 20528 14148 20534
rect 14096 20470 14148 20476
rect 14002 20224 14058 20233
rect 14002 20159 14058 20168
rect 14200 19854 14228 21490
rect 14096 19848 14148 19854
rect 13924 19774 14044 19802
rect 14096 19790 14148 19796
rect 14188 19848 14240 19854
rect 14188 19790 14240 19796
rect 13912 19712 13964 19718
rect 14016 19689 14044 19774
rect 13912 19654 13964 19660
rect 14002 19680 14058 19689
rect 13820 18760 13872 18766
rect 13820 18702 13872 18708
rect 13728 18692 13780 18698
rect 13728 18634 13780 18640
rect 13636 18624 13688 18630
rect 13636 18566 13688 18572
rect 13740 17746 13768 18634
rect 13832 18426 13860 18702
rect 13820 18420 13872 18426
rect 13820 18362 13872 18368
rect 13924 17814 13952 19654
rect 14002 19615 14058 19624
rect 14108 19417 14136 19790
rect 14292 19530 14320 23423
rect 14556 23044 14608 23050
rect 14556 22986 14608 22992
rect 14568 22778 14596 22986
rect 14556 22772 14608 22778
rect 14556 22714 14608 22720
rect 14370 21176 14426 21185
rect 14370 21111 14426 21120
rect 14200 19502 14320 19530
rect 14384 19514 14412 21111
rect 14464 20936 14516 20942
rect 14464 20878 14516 20884
rect 14556 20936 14608 20942
rect 14556 20878 14608 20884
rect 14372 19508 14424 19514
rect 14094 19408 14150 19417
rect 14094 19343 14096 19352
rect 14148 19343 14150 19352
rect 14096 19314 14148 19320
rect 13912 17808 13964 17814
rect 13912 17750 13964 17756
rect 13728 17740 13780 17746
rect 13728 17682 13780 17688
rect 14200 17513 14228 19502
rect 14372 19450 14424 19456
rect 14280 19440 14332 19446
rect 14280 19382 14332 19388
rect 14292 18970 14320 19382
rect 14372 19236 14424 19242
rect 14372 19178 14424 19184
rect 14280 18964 14332 18970
rect 14280 18906 14332 18912
rect 14186 17504 14242 17513
rect 14186 17439 14242 17448
rect 13820 17128 13872 17134
rect 13820 17070 13872 17076
rect 14096 17128 14148 17134
rect 14096 17070 14148 17076
rect 13464 15706 13492 15982
rect 13556 15966 13676 15994
rect 13544 15904 13596 15910
rect 13544 15846 13596 15852
rect 13452 15700 13504 15706
rect 13452 15642 13504 15648
rect 13556 15434 13584 15846
rect 13544 15428 13596 15434
rect 13544 15370 13596 15376
rect 13360 14612 13412 14618
rect 13360 14554 13412 14560
rect 13648 14362 13676 15966
rect 13832 15502 13860 17070
rect 14002 16688 14058 16697
rect 14002 16623 14058 16632
rect 13912 16108 13964 16114
rect 13912 16050 13964 16056
rect 13820 15496 13872 15502
rect 13820 15438 13872 15444
rect 13924 15162 13952 16050
rect 14016 15706 14044 16623
rect 14108 16046 14136 17070
rect 14096 16040 14148 16046
rect 14096 15982 14148 15988
rect 14004 15700 14056 15706
rect 14004 15642 14056 15648
rect 13912 15156 13964 15162
rect 13912 15098 13964 15104
rect 14016 14414 14044 15642
rect 14188 15564 14240 15570
rect 14188 15506 14240 15512
rect 14280 15564 14332 15570
rect 14280 15506 14332 15512
rect 14096 14884 14148 14890
rect 14096 14826 14148 14832
rect 13556 14334 13676 14362
rect 14004 14408 14056 14414
rect 14004 14350 14056 14356
rect 14108 14346 14136 14826
rect 14096 14340 14148 14346
rect 12716 14272 12768 14278
rect 12716 14214 12768 14220
rect 12532 14068 12584 14074
rect 12532 14010 12584 14016
rect 12728 13530 12756 14214
rect 13556 14006 13584 14334
rect 14096 14282 14148 14288
rect 13636 14272 13688 14278
rect 13636 14214 13688 14220
rect 13648 14074 13676 14214
rect 13636 14068 13688 14074
rect 13636 14010 13688 14016
rect 13728 14068 13780 14074
rect 13728 14010 13780 14016
rect 13544 14000 13596 14006
rect 13544 13942 13596 13948
rect 12950 13628 13258 13637
rect 12950 13626 12956 13628
rect 13012 13626 13036 13628
rect 13092 13626 13116 13628
rect 13172 13626 13196 13628
rect 13252 13626 13258 13628
rect 13012 13574 13014 13626
rect 13194 13574 13196 13626
rect 12950 13572 12956 13574
rect 13012 13572 13036 13574
rect 13092 13572 13116 13574
rect 13172 13572 13196 13574
rect 13252 13572 13258 13574
rect 12950 13563 13258 13572
rect 13740 13530 13768 14010
rect 14004 13864 14056 13870
rect 14004 13806 14056 13812
rect 12716 13524 12768 13530
rect 12716 13466 12768 13472
rect 13728 13524 13780 13530
rect 13728 13466 13780 13472
rect 12072 13388 12124 13394
rect 12072 13330 12124 13336
rect 12728 13258 12756 13466
rect 13360 13456 13412 13462
rect 13360 13398 13412 13404
rect 11520 13252 11572 13258
rect 11520 13194 11572 13200
rect 12716 13252 12768 13258
rect 12716 13194 12768 13200
rect 11532 12986 11560 13194
rect 12728 12986 12756 13194
rect 11520 12980 11572 12986
rect 11520 12922 11572 12928
rect 12716 12980 12768 12986
rect 12716 12922 12768 12928
rect 12950 12540 13258 12549
rect 12950 12538 12956 12540
rect 13012 12538 13036 12540
rect 13092 12538 13116 12540
rect 13172 12538 13196 12540
rect 13252 12538 13258 12540
rect 13012 12486 13014 12538
rect 13194 12486 13196 12538
rect 12950 12484 12956 12486
rect 13012 12484 13036 12486
rect 13092 12484 13116 12486
rect 13172 12484 13196 12486
rect 13252 12484 13258 12486
rect 12950 12475 13258 12484
rect 11334 12336 11390 12345
rect 11334 12271 11390 12280
rect 13372 11830 13400 13398
rect 13740 13190 13768 13466
rect 13728 13184 13780 13190
rect 13728 13126 13780 13132
rect 13740 12442 13768 13126
rect 13820 12980 13872 12986
rect 13820 12922 13872 12928
rect 13728 12436 13780 12442
rect 13728 12378 13780 12384
rect 13740 11830 13768 12378
rect 13832 11898 13860 12922
rect 14016 12442 14044 13806
rect 14200 13258 14228 15506
rect 14292 14482 14320 15506
rect 14280 14476 14332 14482
rect 14280 14418 14332 14424
rect 14292 14006 14320 14418
rect 14280 14000 14332 14006
rect 14280 13942 14332 13948
rect 14292 13394 14320 13942
rect 14384 13870 14412 19178
rect 14372 13864 14424 13870
rect 14372 13806 14424 13812
rect 14280 13388 14332 13394
rect 14280 13330 14332 13336
rect 14188 13252 14240 13258
rect 14188 13194 14240 13200
rect 14292 12986 14320 13330
rect 14280 12980 14332 12986
rect 14280 12922 14332 12928
rect 14004 12436 14056 12442
rect 14004 12378 14056 12384
rect 13820 11892 13872 11898
rect 13820 11834 13872 11840
rect 13360 11824 13412 11830
rect 13360 11766 13412 11772
rect 13728 11824 13780 11830
rect 13728 11766 13780 11772
rect 12950 11452 13258 11461
rect 12950 11450 12956 11452
rect 13012 11450 13036 11452
rect 13092 11450 13116 11452
rect 13172 11450 13196 11452
rect 13252 11450 13258 11452
rect 13012 11398 13014 11450
rect 13194 11398 13196 11450
rect 12950 11396 12956 11398
rect 13012 11396 13036 11398
rect 13092 11396 13116 11398
rect 13172 11396 13196 11398
rect 13252 11396 13258 11398
rect 12950 11387 13258 11396
rect 13740 11354 13768 11766
rect 14476 11626 14504 20878
rect 14568 19786 14596 20878
rect 14660 19786 14688 24074
rect 14740 23656 14792 23662
rect 14740 23598 14792 23604
rect 14752 22778 14780 23598
rect 14936 23526 14964 26200
rect 15200 23724 15252 23730
rect 15200 23666 15252 23672
rect 14924 23520 14976 23526
rect 14924 23462 14976 23468
rect 15016 22976 15068 22982
rect 15016 22918 15068 22924
rect 14740 22772 14792 22778
rect 14740 22714 14792 22720
rect 14752 22234 14780 22714
rect 14740 22228 14792 22234
rect 14740 22170 14792 22176
rect 14832 21548 14884 21554
rect 14832 21490 14884 21496
rect 14844 20806 14872 21490
rect 15028 21350 15056 22918
rect 15212 21729 15240 23666
rect 15304 22506 15332 26200
rect 15396 23497 15424 26302
rect 15658 26200 15714 26302
rect 16026 26330 16082 27000
rect 16394 26330 16450 27000
rect 16762 26330 16818 27000
rect 16026 26302 16252 26330
rect 16026 26200 16082 26302
rect 15844 25152 15896 25158
rect 15844 25094 15896 25100
rect 15660 24200 15712 24206
rect 15660 24142 15712 24148
rect 15568 23860 15620 23866
rect 15568 23802 15620 23808
rect 15476 23656 15528 23662
rect 15580 23633 15608 23802
rect 15476 23598 15528 23604
rect 15566 23624 15622 23633
rect 15382 23488 15438 23497
rect 15382 23423 15438 23432
rect 15292 22500 15344 22506
rect 15292 22442 15344 22448
rect 15292 21888 15344 21894
rect 15292 21830 15344 21836
rect 15198 21720 15254 21729
rect 15198 21655 15254 21664
rect 15016 21344 15068 21350
rect 15016 21286 15068 21292
rect 15198 20904 15254 20913
rect 15304 20874 15332 21830
rect 15384 21072 15436 21078
rect 15384 21014 15436 21020
rect 15396 20874 15424 21014
rect 15198 20839 15254 20848
rect 15292 20868 15344 20874
rect 14832 20800 14884 20806
rect 14832 20742 14884 20748
rect 14844 20602 14872 20742
rect 14832 20596 14884 20602
rect 14832 20538 14884 20544
rect 14752 20330 14872 20346
rect 14752 20324 14884 20330
rect 14752 20318 14832 20324
rect 14556 19780 14608 19786
rect 14556 19722 14608 19728
rect 14648 19780 14700 19786
rect 14648 19722 14700 19728
rect 14568 19514 14596 19722
rect 14646 19680 14702 19689
rect 14646 19615 14702 19624
rect 14556 19508 14608 19514
rect 14556 19450 14608 19456
rect 14556 18828 14608 18834
rect 14556 18770 14608 18776
rect 14568 18426 14596 18770
rect 14556 18420 14608 18426
rect 14556 18362 14608 18368
rect 14556 17604 14608 17610
rect 14556 17546 14608 17552
rect 14568 17202 14596 17546
rect 14556 17196 14608 17202
rect 14556 17138 14608 17144
rect 14568 16522 14596 17138
rect 14660 16561 14688 19615
rect 14752 19242 14780 20318
rect 14832 20266 14884 20272
rect 14922 20088 14978 20097
rect 15212 20058 15240 20839
rect 15292 20810 15344 20816
rect 15384 20868 15436 20874
rect 15384 20810 15436 20816
rect 15384 20596 15436 20602
rect 15384 20538 15436 20544
rect 15292 20528 15344 20534
rect 15292 20470 15344 20476
rect 14922 20023 14978 20032
rect 15200 20052 15252 20058
rect 14832 19780 14884 19786
rect 14832 19722 14884 19728
rect 14844 19514 14872 19722
rect 14832 19508 14884 19514
rect 14832 19450 14884 19456
rect 14740 19236 14792 19242
rect 14740 19178 14792 19184
rect 14832 19168 14884 19174
rect 14832 19110 14884 19116
rect 14844 18952 14872 19110
rect 14752 18924 14872 18952
rect 14752 18834 14780 18924
rect 14936 18850 14964 20023
rect 15200 19994 15252 20000
rect 15108 19848 15160 19854
rect 15108 19790 15160 19796
rect 15016 19780 15068 19786
rect 15016 19722 15068 19728
rect 14740 18828 14792 18834
rect 14740 18770 14792 18776
rect 14844 18822 14964 18850
rect 14844 17082 14872 18822
rect 14924 18760 14976 18766
rect 14924 18702 14976 18708
rect 14936 17746 14964 18702
rect 15028 18630 15056 19722
rect 15120 19553 15148 19790
rect 15106 19544 15162 19553
rect 15106 19479 15162 19488
rect 15304 19378 15332 20470
rect 15396 19786 15424 20538
rect 15384 19780 15436 19786
rect 15384 19722 15436 19728
rect 15292 19372 15344 19378
rect 15292 19314 15344 19320
rect 15108 19304 15160 19310
rect 15108 19246 15160 19252
rect 15120 18834 15148 19246
rect 15304 18834 15332 19314
rect 15382 19000 15438 19009
rect 15382 18935 15438 18944
rect 15108 18828 15160 18834
rect 15108 18770 15160 18776
rect 15292 18828 15344 18834
rect 15292 18770 15344 18776
rect 15016 18624 15068 18630
rect 15016 18566 15068 18572
rect 15120 18222 15148 18770
rect 15200 18692 15252 18698
rect 15200 18634 15252 18640
rect 15108 18216 15160 18222
rect 15108 18158 15160 18164
rect 15014 18048 15070 18057
rect 15014 17983 15070 17992
rect 14924 17740 14976 17746
rect 14924 17682 14976 17688
rect 14752 17054 14872 17082
rect 14646 16552 14702 16561
rect 14556 16516 14608 16522
rect 14646 16487 14702 16496
rect 14556 16458 14608 16464
rect 14568 16402 14596 16458
rect 14568 16374 14688 16402
rect 14556 16040 14608 16046
rect 14556 15982 14608 15988
rect 14568 14482 14596 15982
rect 14660 14600 14688 16374
rect 14752 14890 14780 17054
rect 14832 16992 14884 16998
rect 14832 16934 14884 16940
rect 14740 14884 14792 14890
rect 14740 14826 14792 14832
rect 14660 14572 14780 14600
rect 14556 14476 14608 14482
rect 14608 14436 14688 14464
rect 14556 14418 14608 14424
rect 14660 14074 14688 14436
rect 14648 14068 14700 14074
rect 14648 14010 14700 14016
rect 14556 13252 14608 13258
rect 14556 13194 14608 13200
rect 14568 11898 14596 13194
rect 14556 11892 14608 11898
rect 14556 11834 14608 11840
rect 14464 11620 14516 11626
rect 14464 11562 14516 11568
rect 14648 11552 14700 11558
rect 14648 11494 14700 11500
rect 14660 11354 14688 11494
rect 12532 11348 12584 11354
rect 12532 11290 12584 11296
rect 13728 11348 13780 11354
rect 13728 11290 13780 11296
rect 14648 11348 14700 11354
rect 14648 11290 14700 11296
rect 10048 9036 10100 9042
rect 10048 8978 10100 8984
rect 12544 8906 12572 11290
rect 12950 10364 13258 10373
rect 12950 10362 12956 10364
rect 13012 10362 13036 10364
rect 13092 10362 13116 10364
rect 13172 10362 13196 10364
rect 13252 10362 13258 10364
rect 13012 10310 13014 10362
rect 13194 10310 13196 10362
rect 12950 10308 12956 10310
rect 13012 10308 13036 10310
rect 13092 10308 13116 10310
rect 13172 10308 13196 10310
rect 13252 10308 13258 10310
rect 12950 10299 13258 10308
rect 12950 9276 13258 9285
rect 12950 9274 12956 9276
rect 13012 9274 13036 9276
rect 13092 9274 13116 9276
rect 13172 9274 13196 9276
rect 13252 9274 13258 9276
rect 13012 9222 13014 9274
rect 13194 9222 13196 9274
rect 12950 9220 12956 9222
rect 13012 9220 13036 9222
rect 13092 9220 13116 9222
rect 13172 9220 13196 9222
rect 13252 9220 13258 9222
rect 12950 9211 13258 9220
rect 14752 9178 14780 14572
rect 14740 9172 14792 9178
rect 14740 9114 14792 9120
rect 9312 8900 9364 8906
rect 9312 8842 9364 8848
rect 12532 8900 12584 8906
rect 12532 8842 12584 8848
rect 7950 8732 8258 8741
rect 7950 8730 7956 8732
rect 8012 8730 8036 8732
rect 8092 8730 8116 8732
rect 8172 8730 8196 8732
rect 8252 8730 8258 8732
rect 8012 8678 8014 8730
rect 8194 8678 8196 8730
rect 7950 8676 7956 8678
rect 8012 8676 8036 8678
rect 8092 8676 8116 8678
rect 8172 8676 8196 8678
rect 8252 8676 8258 8678
rect 7950 8667 8258 8676
rect 2950 8188 3258 8197
rect 2950 8186 2956 8188
rect 3012 8186 3036 8188
rect 3092 8186 3116 8188
rect 3172 8186 3196 8188
rect 3252 8186 3258 8188
rect 3012 8134 3014 8186
rect 3194 8134 3196 8186
rect 2950 8132 2956 8134
rect 3012 8132 3036 8134
rect 3092 8132 3116 8134
rect 3172 8132 3196 8134
rect 3252 8132 3258 8134
rect 2950 8123 3258 8132
rect 7950 7644 8258 7653
rect 7950 7642 7956 7644
rect 8012 7642 8036 7644
rect 8092 7642 8116 7644
rect 8172 7642 8196 7644
rect 8252 7642 8258 7644
rect 8012 7590 8014 7642
rect 8194 7590 8196 7642
rect 7950 7588 7956 7590
rect 8012 7588 8036 7590
rect 8092 7588 8116 7590
rect 8172 7588 8196 7590
rect 8252 7588 8258 7590
rect 7950 7579 8258 7588
rect 2950 7100 3258 7109
rect 2950 7098 2956 7100
rect 3012 7098 3036 7100
rect 3092 7098 3116 7100
rect 3172 7098 3196 7100
rect 3252 7098 3258 7100
rect 3012 7046 3014 7098
rect 3194 7046 3196 7098
rect 2950 7044 2956 7046
rect 3012 7044 3036 7046
rect 3092 7044 3116 7046
rect 3172 7044 3196 7046
rect 3252 7044 3258 7046
rect 2950 7035 3258 7044
rect 7950 6556 8258 6565
rect 7950 6554 7956 6556
rect 8012 6554 8036 6556
rect 8092 6554 8116 6556
rect 8172 6554 8196 6556
rect 8252 6554 8258 6556
rect 8012 6502 8014 6554
rect 8194 6502 8196 6554
rect 7950 6500 7956 6502
rect 8012 6500 8036 6502
rect 8092 6500 8116 6502
rect 8172 6500 8196 6502
rect 8252 6500 8258 6502
rect 7950 6491 8258 6500
rect 9324 6458 9352 8842
rect 14844 8498 14872 16934
rect 14936 16658 14964 17682
rect 15028 17202 15056 17983
rect 15120 17610 15148 18158
rect 15212 17610 15240 18634
rect 15396 18329 15424 18935
rect 15382 18320 15438 18329
rect 15382 18255 15438 18264
rect 15108 17604 15160 17610
rect 15108 17546 15160 17552
rect 15200 17604 15252 17610
rect 15200 17546 15252 17552
rect 15016 17196 15068 17202
rect 15016 17138 15068 17144
rect 15016 16992 15068 16998
rect 15016 16934 15068 16940
rect 15028 16794 15056 16934
rect 15016 16788 15068 16794
rect 15016 16730 15068 16736
rect 14924 16652 14976 16658
rect 14924 16594 14976 16600
rect 15016 16652 15068 16658
rect 15016 16594 15068 16600
rect 15028 15706 15056 16594
rect 15108 15904 15160 15910
rect 15108 15846 15160 15852
rect 15016 15700 15068 15706
rect 15016 15642 15068 15648
rect 15120 15434 15148 15846
rect 15212 15706 15240 17546
rect 15384 15904 15436 15910
rect 15384 15846 15436 15852
rect 15200 15700 15252 15706
rect 15200 15642 15252 15648
rect 15108 15428 15160 15434
rect 15108 15370 15160 15376
rect 15290 15192 15346 15201
rect 15290 15127 15292 15136
rect 15344 15127 15346 15136
rect 15292 15098 15344 15104
rect 15396 14958 15424 15846
rect 15384 14952 15436 14958
rect 15384 14894 15436 14900
rect 15016 14340 15068 14346
rect 15016 14282 15068 14288
rect 15028 13938 15056 14282
rect 15016 13932 15068 13938
rect 15016 13874 15068 13880
rect 15028 13258 15056 13874
rect 15200 13728 15252 13734
rect 15200 13670 15252 13676
rect 15212 13530 15240 13670
rect 15200 13524 15252 13530
rect 15200 13466 15252 13472
rect 15016 13252 15068 13258
rect 15016 13194 15068 13200
rect 15028 12986 15056 13194
rect 15016 12980 15068 12986
rect 15016 12922 15068 12928
rect 15200 12776 15252 12782
rect 15200 12718 15252 12724
rect 14832 8492 14884 8498
rect 14832 8434 14884 8440
rect 12950 8188 13258 8197
rect 12950 8186 12956 8188
rect 13012 8186 13036 8188
rect 13092 8186 13116 8188
rect 13172 8186 13196 8188
rect 13252 8186 13258 8188
rect 13012 8134 13014 8186
rect 13194 8134 13196 8186
rect 12950 8132 12956 8134
rect 13012 8132 13036 8134
rect 13092 8132 13116 8134
rect 13172 8132 13196 8134
rect 13252 8132 13258 8134
rect 12950 8123 13258 8132
rect 12950 7100 13258 7109
rect 12950 7098 12956 7100
rect 13012 7098 13036 7100
rect 13092 7098 13116 7100
rect 13172 7098 13196 7100
rect 13252 7098 13258 7100
rect 13012 7046 13014 7098
rect 13194 7046 13196 7098
rect 12950 7044 12956 7046
rect 13012 7044 13036 7046
rect 13092 7044 13116 7046
rect 13172 7044 13196 7046
rect 13252 7044 13258 7046
rect 12950 7035 13258 7044
rect 15212 6730 15240 12718
rect 15488 11354 15516 23598
rect 15672 23594 15700 24142
rect 15752 23860 15804 23866
rect 15752 23802 15804 23808
rect 15764 23662 15792 23802
rect 15752 23656 15804 23662
rect 15752 23598 15804 23604
rect 15856 23594 15884 25094
rect 16028 24812 16080 24818
rect 16028 24754 16080 24760
rect 16040 24449 16068 24754
rect 16026 24440 16082 24449
rect 16026 24375 16082 24384
rect 16040 23905 16068 24375
rect 16120 24268 16172 24274
rect 16120 24210 16172 24216
rect 16026 23896 16082 23905
rect 16026 23831 16082 23840
rect 15566 23559 15622 23568
rect 15660 23588 15712 23594
rect 15660 23530 15712 23536
rect 15844 23588 15896 23594
rect 15844 23530 15896 23536
rect 15568 23044 15620 23050
rect 15568 22986 15620 22992
rect 15580 22778 15608 22986
rect 15672 22930 15700 23530
rect 15672 22902 15792 22930
rect 15568 22772 15620 22778
rect 15568 22714 15620 22720
rect 15660 22568 15712 22574
rect 15660 22510 15712 22516
rect 15568 21548 15620 21554
rect 15568 21490 15620 21496
rect 15580 19174 15608 21490
rect 15672 21486 15700 22510
rect 15660 21480 15712 21486
rect 15660 21422 15712 21428
rect 15658 21176 15714 21185
rect 15658 21111 15714 21120
rect 15672 20777 15700 21111
rect 15658 20768 15714 20777
rect 15658 20703 15714 20712
rect 15660 19916 15712 19922
rect 15660 19858 15712 19864
rect 15672 19378 15700 19858
rect 15660 19372 15712 19378
rect 15660 19314 15712 19320
rect 15568 19168 15620 19174
rect 15568 19110 15620 19116
rect 15580 18426 15608 19110
rect 15568 18420 15620 18426
rect 15568 18362 15620 18368
rect 15580 16250 15608 18362
rect 15764 17746 15792 22902
rect 15936 22636 15988 22642
rect 15936 22578 15988 22584
rect 15844 22432 15896 22438
rect 15844 22374 15896 22380
rect 15856 22166 15884 22374
rect 15844 22160 15896 22166
rect 15844 22102 15896 22108
rect 15842 21584 15898 21593
rect 15842 21519 15898 21528
rect 15856 21350 15884 21519
rect 15844 21344 15896 21350
rect 15844 21286 15896 21292
rect 15856 21010 15884 21286
rect 15844 21004 15896 21010
rect 15844 20946 15896 20952
rect 15844 20800 15896 20806
rect 15842 20768 15844 20777
rect 15896 20768 15898 20777
rect 15842 20703 15898 20712
rect 15844 20460 15896 20466
rect 15948 20448 15976 22578
rect 16028 22432 16080 22438
rect 16028 22374 16080 22380
rect 16040 22137 16068 22374
rect 16026 22128 16082 22137
rect 16026 22063 16082 22072
rect 16132 21486 16160 24210
rect 16224 21690 16252 26302
rect 16394 26302 16528 26330
rect 16394 26200 16450 26302
rect 16396 24336 16448 24342
rect 16396 24278 16448 24284
rect 16304 23656 16356 23662
rect 16304 23598 16356 23604
rect 16316 22574 16344 23598
rect 16304 22568 16356 22574
rect 16304 22510 16356 22516
rect 16304 22432 16356 22438
rect 16304 22374 16356 22380
rect 16316 22137 16344 22374
rect 16302 22128 16358 22137
rect 16302 22063 16358 22072
rect 16212 21684 16264 21690
rect 16212 21626 16264 21632
rect 16302 21584 16358 21593
rect 16212 21548 16264 21554
rect 16302 21519 16304 21528
rect 16212 21490 16264 21496
rect 16356 21519 16358 21528
rect 16304 21490 16356 21496
rect 16120 21480 16172 21486
rect 16120 21422 16172 21428
rect 16224 21350 16252 21490
rect 16212 21344 16264 21350
rect 16212 21286 16264 21292
rect 16224 21010 16252 21286
rect 16212 21004 16264 21010
rect 16212 20946 16264 20952
rect 16408 20641 16436 24278
rect 16500 23322 16528 26302
rect 16684 26302 16818 26330
rect 16580 23860 16632 23866
rect 16580 23802 16632 23808
rect 16592 23633 16620 23802
rect 16578 23624 16634 23633
rect 16578 23559 16634 23568
rect 16488 23316 16540 23322
rect 16488 23258 16540 23264
rect 16580 23316 16632 23322
rect 16580 23258 16632 23264
rect 16592 22710 16620 23258
rect 16580 22704 16632 22710
rect 16580 22646 16632 22652
rect 16488 22432 16540 22438
rect 16488 22374 16540 22380
rect 16394 20632 16450 20641
rect 16394 20567 16450 20576
rect 16500 20482 16528 22374
rect 16580 21412 16632 21418
rect 16580 21354 16632 21360
rect 16592 21146 16620 21354
rect 16684 21350 16712 26302
rect 16762 26200 16818 26302
rect 17130 26200 17186 27000
rect 17498 26200 17554 27000
rect 17866 26330 17922 27000
rect 17604 26302 17922 26330
rect 16856 24676 16908 24682
rect 16856 24618 16908 24624
rect 16868 24070 16896 24618
rect 16948 24200 17000 24206
rect 16948 24142 17000 24148
rect 16856 24064 16908 24070
rect 16856 24006 16908 24012
rect 16764 23520 16816 23526
rect 16856 23520 16908 23526
rect 16764 23462 16816 23468
rect 16854 23488 16856 23497
rect 16908 23488 16910 23497
rect 16776 23118 16804 23462
rect 16854 23423 16910 23432
rect 16764 23112 16816 23118
rect 16764 23054 16816 23060
rect 16764 22976 16816 22982
rect 16762 22944 16764 22953
rect 16816 22944 16818 22953
rect 16762 22879 16818 22888
rect 16856 22772 16908 22778
rect 16856 22714 16908 22720
rect 16764 21888 16816 21894
rect 16762 21856 16764 21865
rect 16816 21856 16818 21865
rect 16762 21791 16818 21800
rect 16868 21672 16896 22714
rect 16776 21644 16896 21672
rect 16672 21344 16724 21350
rect 16672 21286 16724 21292
rect 16580 21140 16632 21146
rect 16580 21082 16632 21088
rect 16408 20454 16528 20482
rect 15948 20420 16068 20448
rect 15844 20402 15896 20408
rect 15856 19417 15884 20402
rect 15934 20360 15990 20369
rect 15934 20295 15990 20304
rect 15948 20262 15976 20295
rect 15936 20256 15988 20262
rect 15936 20198 15988 20204
rect 16040 20074 16068 20420
rect 15948 20046 16068 20074
rect 15842 19408 15898 19417
rect 15842 19343 15898 19352
rect 15948 18850 15976 20046
rect 16302 19816 16358 19825
rect 16212 19780 16264 19786
rect 16302 19751 16358 19760
rect 16212 19722 16264 19728
rect 16224 19417 16252 19722
rect 16316 19718 16344 19751
rect 16304 19712 16356 19718
rect 16304 19654 16356 19660
rect 16210 19408 16266 19417
rect 16210 19343 16266 19352
rect 16028 19304 16080 19310
rect 16028 19246 16080 19252
rect 15856 18822 15976 18850
rect 15752 17740 15804 17746
rect 15752 17682 15804 17688
rect 15856 16561 15884 18822
rect 16040 18698 16068 19246
rect 16120 19168 16172 19174
rect 16120 19110 16172 19116
rect 16028 18692 16080 18698
rect 16028 18634 16080 18640
rect 15936 17332 15988 17338
rect 15936 17274 15988 17280
rect 15842 16552 15898 16561
rect 15842 16487 15898 16496
rect 15568 16244 15620 16250
rect 15568 16186 15620 16192
rect 15752 16176 15804 16182
rect 15752 16118 15804 16124
rect 15764 16028 15792 16118
rect 15844 16040 15896 16046
rect 15764 16000 15844 16028
rect 15844 15982 15896 15988
rect 15842 15872 15898 15881
rect 15842 15807 15898 15816
rect 15856 15473 15884 15807
rect 15842 15464 15898 15473
rect 15842 15399 15898 15408
rect 15948 14618 15976 17274
rect 16040 16794 16068 18634
rect 16132 16794 16160 19110
rect 16304 17672 16356 17678
rect 16304 17614 16356 17620
rect 16212 17264 16264 17270
rect 16212 17206 16264 17212
rect 16028 16788 16080 16794
rect 16028 16730 16080 16736
rect 16120 16788 16172 16794
rect 16120 16730 16172 16736
rect 16028 16040 16080 16046
rect 16028 15982 16080 15988
rect 16040 15910 16068 15982
rect 16028 15904 16080 15910
rect 16028 15846 16080 15852
rect 16224 15366 16252 17206
rect 16316 16522 16344 17614
rect 16304 16516 16356 16522
rect 16304 16458 16356 16464
rect 16316 16250 16344 16458
rect 16304 16244 16356 16250
rect 16304 16186 16356 16192
rect 16304 16040 16356 16046
rect 16304 15982 16356 15988
rect 16212 15360 16264 15366
rect 16212 15302 16264 15308
rect 16120 14952 16172 14958
rect 16120 14894 16172 14900
rect 16132 14618 16160 14894
rect 15936 14612 15988 14618
rect 15936 14554 15988 14560
rect 16120 14612 16172 14618
rect 16120 14554 16172 14560
rect 16224 14550 16252 15302
rect 16212 14544 16264 14550
rect 16212 14486 16264 14492
rect 16026 14104 16082 14113
rect 16026 14039 16082 14048
rect 15568 13796 15620 13802
rect 15568 13738 15620 13744
rect 15580 12918 15608 13738
rect 15658 13696 15714 13705
rect 15658 13631 15714 13640
rect 15568 12912 15620 12918
rect 15568 12854 15620 12860
rect 15580 12442 15608 12854
rect 15568 12436 15620 12442
rect 15568 12378 15620 12384
rect 15568 12232 15620 12238
rect 15568 12174 15620 12180
rect 15476 11348 15528 11354
rect 15476 11290 15528 11296
rect 15580 11082 15608 12174
rect 15672 11150 15700 13631
rect 15750 13288 15806 13297
rect 15750 13223 15806 13232
rect 15764 11898 15792 13223
rect 15752 11892 15804 11898
rect 15752 11834 15804 11840
rect 16040 11150 16068 14039
rect 16316 13530 16344 15982
rect 16408 14074 16436 20454
rect 16488 20392 16540 20398
rect 16488 20334 16540 20340
rect 16500 19378 16528 20334
rect 16580 19712 16632 19718
rect 16578 19680 16580 19689
rect 16632 19680 16634 19689
rect 16578 19615 16634 19624
rect 16684 19446 16712 21286
rect 16776 20534 16804 21644
rect 16856 21548 16908 21554
rect 16856 21490 16908 21496
rect 16764 20528 16816 20534
rect 16764 20470 16816 20476
rect 16764 19780 16816 19786
rect 16764 19722 16816 19728
rect 16672 19440 16724 19446
rect 16672 19382 16724 19388
rect 16488 19372 16540 19378
rect 16488 19314 16540 19320
rect 16488 18828 16540 18834
rect 16488 18770 16540 18776
rect 16500 18358 16528 18770
rect 16488 18352 16540 18358
rect 16488 18294 16540 18300
rect 16500 17678 16528 18294
rect 16488 17672 16540 17678
rect 16488 17614 16540 17620
rect 16580 17536 16632 17542
rect 16580 17478 16632 17484
rect 16592 17082 16620 17478
rect 16500 17054 16620 17082
rect 16500 16998 16528 17054
rect 16488 16992 16540 16998
rect 16488 16934 16540 16940
rect 16580 16992 16632 16998
rect 16580 16934 16632 16940
rect 16488 16448 16540 16454
rect 16488 16390 16540 16396
rect 16500 15910 16528 16390
rect 16488 15904 16540 15910
rect 16488 15846 16540 15852
rect 16486 15736 16542 15745
rect 16486 15671 16542 15680
rect 16500 14958 16528 15671
rect 16488 14952 16540 14958
rect 16488 14894 16540 14900
rect 16488 14816 16540 14822
rect 16488 14758 16540 14764
rect 16500 14414 16528 14758
rect 16488 14408 16540 14414
rect 16488 14350 16540 14356
rect 16396 14068 16448 14074
rect 16396 14010 16448 14016
rect 16304 13524 16356 13530
rect 16304 13466 16356 13472
rect 16500 13394 16528 14350
rect 16592 13530 16620 16934
rect 16672 16448 16724 16454
rect 16672 16390 16724 16396
rect 16684 15706 16712 16390
rect 16672 15700 16724 15706
rect 16672 15642 16724 15648
rect 16670 15464 16726 15473
rect 16670 15399 16726 15408
rect 16684 14890 16712 15399
rect 16672 14884 16724 14890
rect 16672 14826 16724 14832
rect 16672 14340 16724 14346
rect 16672 14282 16724 14288
rect 16684 13870 16712 14282
rect 16776 14278 16804 19722
rect 16868 18290 16896 21490
rect 16960 21321 16988 24142
rect 17040 24064 17092 24070
rect 17040 24006 17092 24012
rect 16946 21312 17002 21321
rect 16946 21247 17002 21256
rect 16948 21072 17000 21078
rect 16948 21014 17000 21020
rect 16856 18284 16908 18290
rect 16856 18226 16908 18232
rect 16856 17740 16908 17746
rect 16856 17682 16908 17688
rect 16868 17270 16896 17682
rect 16960 17354 16988 21014
rect 17052 20890 17080 24006
rect 17144 23254 17172 26200
rect 17316 24948 17368 24954
rect 17316 24890 17368 24896
rect 17328 23662 17356 24890
rect 17512 24721 17540 26200
rect 17498 24712 17554 24721
rect 17498 24647 17554 24656
rect 17316 23656 17368 23662
rect 17316 23598 17368 23604
rect 17132 23248 17184 23254
rect 17132 23190 17184 23196
rect 17316 22976 17368 22982
rect 17316 22918 17368 22924
rect 17132 22704 17184 22710
rect 17328 22692 17356 22918
rect 17184 22664 17356 22692
rect 17132 22646 17184 22652
rect 17132 22228 17184 22234
rect 17132 22170 17184 22176
rect 17144 21894 17172 22170
rect 17224 22092 17276 22098
rect 17224 22034 17276 22040
rect 17132 21888 17184 21894
rect 17132 21830 17184 21836
rect 17236 21554 17264 22034
rect 17316 21956 17368 21962
rect 17316 21898 17368 21904
rect 17500 21956 17552 21962
rect 17500 21898 17552 21904
rect 17224 21548 17276 21554
rect 17224 21490 17276 21496
rect 17052 20862 17172 20890
rect 17040 20800 17092 20806
rect 17040 20742 17092 20748
rect 17052 19825 17080 20742
rect 17038 19816 17094 19825
rect 17038 19751 17094 19760
rect 17040 19236 17092 19242
rect 17040 19178 17092 19184
rect 17052 17678 17080 19178
rect 17144 19174 17172 20862
rect 17224 20392 17276 20398
rect 17224 20334 17276 20340
rect 17132 19168 17184 19174
rect 17132 19110 17184 19116
rect 17236 18902 17264 20334
rect 17224 18896 17276 18902
rect 17224 18838 17276 18844
rect 17132 18692 17184 18698
rect 17132 18634 17184 18640
rect 17144 18601 17172 18634
rect 17130 18592 17186 18601
rect 17130 18527 17186 18536
rect 17132 18352 17184 18358
rect 17132 18294 17184 18300
rect 17040 17672 17092 17678
rect 17040 17614 17092 17620
rect 17144 17377 17172 18294
rect 17224 18284 17276 18290
rect 17224 18226 17276 18232
rect 17130 17368 17186 17377
rect 16960 17326 17080 17354
rect 16856 17264 16908 17270
rect 16856 17206 16908 17212
rect 16948 17196 17000 17202
rect 16948 17138 17000 17144
rect 16856 17060 16908 17066
rect 16856 17002 16908 17008
rect 16868 16658 16896 17002
rect 16856 16652 16908 16658
rect 16856 16594 16908 16600
rect 16856 16516 16908 16522
rect 16856 16458 16908 16464
rect 16868 16250 16896 16458
rect 16856 16244 16908 16250
rect 16856 16186 16908 16192
rect 16868 15638 16896 16186
rect 16856 15632 16908 15638
rect 16856 15574 16908 15580
rect 16856 15496 16908 15502
rect 16856 15438 16908 15444
rect 16764 14272 16816 14278
rect 16764 14214 16816 14220
rect 16672 13864 16724 13870
rect 16672 13806 16724 13812
rect 16580 13524 16632 13530
rect 16580 13466 16632 13472
rect 16488 13388 16540 13394
rect 16488 13330 16540 13336
rect 16488 13252 16540 13258
rect 16488 13194 16540 13200
rect 16304 13184 16356 13190
rect 16304 13126 16356 13132
rect 16316 12170 16344 13126
rect 16500 12986 16528 13194
rect 16488 12980 16540 12986
rect 16488 12922 16540 12928
rect 16500 12170 16528 12922
rect 16868 12850 16896 15438
rect 16856 12844 16908 12850
rect 16856 12786 16908 12792
rect 16672 12776 16724 12782
rect 16868 12730 16896 12786
rect 16672 12718 16724 12724
rect 16304 12164 16356 12170
rect 16304 12106 16356 12112
rect 16488 12164 16540 12170
rect 16488 12106 16540 12112
rect 16118 11384 16174 11393
rect 16118 11319 16120 11328
rect 16172 11319 16174 11328
rect 16120 11290 16172 11296
rect 15660 11144 15712 11150
rect 15660 11086 15712 11092
rect 16028 11144 16080 11150
rect 16028 11086 16080 11092
rect 15568 11076 15620 11082
rect 15568 11018 15620 11024
rect 15672 10810 15700 11086
rect 16040 10810 16068 11086
rect 15660 10804 15712 10810
rect 15660 10746 15712 10752
rect 16028 10804 16080 10810
rect 16028 10746 16080 10752
rect 16684 10470 16712 12718
rect 16776 12702 16896 12730
rect 16776 12306 16804 12702
rect 16854 12472 16910 12481
rect 16854 12407 16910 12416
rect 16764 12300 16816 12306
rect 16764 12242 16816 12248
rect 16764 11756 16816 11762
rect 16764 11698 16816 11704
rect 16776 11558 16804 11698
rect 16868 11694 16896 12407
rect 16856 11688 16908 11694
rect 16856 11630 16908 11636
rect 16764 11552 16816 11558
rect 16764 11494 16816 11500
rect 16960 11354 16988 17138
rect 17052 15162 17080 17326
rect 17130 17303 17186 17312
rect 17132 16652 17184 16658
rect 17132 16594 17184 16600
rect 17040 15156 17092 15162
rect 17040 15098 17092 15104
rect 17144 14822 17172 16594
rect 17236 16289 17264 18226
rect 17222 16280 17278 16289
rect 17222 16215 17278 16224
rect 17224 16176 17276 16182
rect 17224 16118 17276 16124
rect 17236 15337 17264 16118
rect 17222 15328 17278 15337
rect 17222 15263 17278 15272
rect 17222 15056 17278 15065
rect 17222 14991 17278 15000
rect 17132 14816 17184 14822
rect 17132 14758 17184 14764
rect 17040 13728 17092 13734
rect 17236 13682 17264 14991
rect 17040 13670 17092 13676
rect 16948 11348 17000 11354
rect 16948 11290 17000 11296
rect 16672 10464 16724 10470
rect 16672 10406 16724 10412
rect 17052 9654 17080 13670
rect 17144 13654 17264 13682
rect 17144 11150 17172 13654
rect 17224 13252 17276 13258
rect 17224 13194 17276 13200
rect 17236 12918 17264 13194
rect 17224 12912 17276 12918
rect 17224 12854 17276 12860
rect 17132 11144 17184 11150
rect 17132 11086 17184 11092
rect 17144 10810 17172 11086
rect 17132 10804 17184 10810
rect 17132 10746 17184 10752
rect 17328 10538 17356 21898
rect 17408 21548 17460 21554
rect 17408 21490 17460 21496
rect 17420 18442 17448 21490
rect 17512 21486 17540 21898
rect 17500 21480 17552 21486
rect 17500 21422 17552 21428
rect 17512 20505 17540 21422
rect 17498 20496 17554 20505
rect 17498 20431 17554 20440
rect 17420 18414 17540 18442
rect 17512 18290 17540 18414
rect 17500 18284 17552 18290
rect 17500 18226 17552 18232
rect 17408 18216 17460 18222
rect 17408 18158 17460 18164
rect 17420 17610 17448 18158
rect 17500 18080 17552 18086
rect 17500 18022 17552 18028
rect 17408 17604 17460 17610
rect 17408 17546 17460 17552
rect 17512 14074 17540 18022
rect 17604 16454 17632 26302
rect 17866 26200 17922 26302
rect 18234 26330 18290 27000
rect 18234 26302 18368 26330
rect 18234 26200 18290 26302
rect 18144 24880 18196 24886
rect 18144 24822 18196 24828
rect 17682 24712 17738 24721
rect 17682 24647 17738 24656
rect 17696 24041 17724 24647
rect 18156 24410 18184 24822
rect 18144 24404 18196 24410
rect 18144 24346 18196 24352
rect 17776 24268 17828 24274
rect 17776 24210 17828 24216
rect 17788 24070 17816 24210
rect 17958 24168 18014 24177
rect 17958 24103 18014 24112
rect 17972 24070 18000 24103
rect 17776 24064 17828 24070
rect 17682 24032 17738 24041
rect 17776 24006 17828 24012
rect 17960 24064 18012 24070
rect 17960 24006 18012 24012
rect 17682 23967 17738 23976
rect 17950 23964 18258 23973
rect 17950 23962 17956 23964
rect 18012 23962 18036 23964
rect 18092 23962 18116 23964
rect 18172 23962 18196 23964
rect 18252 23962 18258 23964
rect 18012 23910 18014 23962
rect 18194 23910 18196 23962
rect 17950 23908 17956 23910
rect 18012 23908 18036 23910
rect 18092 23908 18116 23910
rect 18172 23908 18196 23910
rect 18252 23908 18258 23910
rect 17950 23899 18258 23908
rect 17776 23724 17828 23730
rect 17776 23666 17828 23672
rect 17684 23316 17736 23322
rect 17684 23258 17736 23264
rect 17696 22166 17724 23258
rect 17684 22160 17736 22166
rect 17684 22102 17736 22108
rect 17788 22094 17816 23666
rect 18052 23656 18104 23662
rect 18052 23598 18104 23604
rect 17960 23588 18012 23594
rect 17960 23530 18012 23536
rect 17972 23322 18000 23530
rect 17960 23316 18012 23322
rect 17960 23258 18012 23264
rect 18064 23118 18092 23598
rect 18052 23112 18104 23118
rect 18052 23054 18104 23060
rect 18064 22982 18092 23054
rect 18052 22976 18104 22982
rect 18052 22918 18104 22924
rect 17950 22876 18258 22885
rect 17950 22874 17956 22876
rect 18012 22874 18036 22876
rect 18092 22874 18116 22876
rect 18172 22874 18196 22876
rect 18252 22874 18258 22876
rect 18012 22822 18014 22874
rect 18194 22822 18196 22874
rect 17950 22820 17956 22822
rect 18012 22820 18036 22822
rect 18092 22820 18116 22822
rect 18172 22820 18196 22822
rect 18252 22820 18258 22822
rect 17950 22811 18258 22820
rect 17788 22066 17908 22094
rect 17684 21888 17736 21894
rect 17684 21830 17736 21836
rect 17776 21888 17828 21894
rect 17776 21830 17828 21836
rect 17696 21622 17724 21830
rect 17684 21616 17736 21622
rect 17684 21558 17736 21564
rect 17684 21480 17736 21486
rect 17684 21422 17736 21428
rect 17696 19310 17724 21422
rect 17684 19304 17736 19310
rect 17684 19246 17736 19252
rect 17684 18624 17736 18630
rect 17684 18566 17736 18572
rect 17696 17542 17724 18566
rect 17788 18057 17816 21830
rect 17880 21554 17908 22066
rect 18144 22092 18196 22098
rect 18144 22034 18196 22040
rect 18156 21894 18184 22034
rect 18144 21888 18196 21894
rect 18144 21830 18196 21836
rect 17950 21788 18258 21797
rect 17950 21786 17956 21788
rect 18012 21786 18036 21788
rect 18092 21786 18116 21788
rect 18172 21786 18196 21788
rect 18252 21786 18258 21788
rect 18012 21734 18014 21786
rect 18194 21734 18196 21786
rect 17950 21732 17956 21734
rect 18012 21732 18036 21734
rect 18092 21732 18116 21734
rect 18172 21732 18196 21734
rect 18252 21732 18258 21734
rect 17950 21723 18258 21732
rect 17868 21548 17920 21554
rect 17868 21490 17920 21496
rect 18236 21072 18288 21078
rect 18340 21060 18368 26302
rect 18602 26200 18658 27000
rect 18970 26200 19026 27000
rect 19338 26330 19394 27000
rect 19338 26302 19564 26330
rect 19338 26200 19394 26302
rect 18420 23792 18472 23798
rect 18420 23734 18472 23740
rect 18432 23662 18460 23734
rect 18420 23656 18472 23662
rect 18420 23598 18472 23604
rect 18616 23361 18644 26200
rect 18984 26081 19012 26200
rect 18970 26072 19026 26081
rect 18970 26007 19026 26016
rect 19062 24984 19118 24993
rect 19062 24919 19118 24928
rect 19430 24984 19486 24993
rect 19430 24919 19486 24928
rect 18788 24404 18840 24410
rect 18708 24364 18788 24392
rect 18708 24274 18736 24364
rect 18788 24346 18840 24352
rect 18696 24268 18748 24274
rect 18696 24210 18748 24216
rect 18788 24268 18840 24274
rect 18788 24210 18840 24216
rect 18602 23352 18658 23361
rect 18800 23322 18828 24210
rect 18972 23792 19024 23798
rect 18972 23734 19024 23740
rect 18602 23287 18658 23296
rect 18788 23316 18840 23322
rect 18788 23258 18840 23264
rect 18984 23254 19012 23734
rect 18880 23248 18932 23254
rect 18880 23190 18932 23196
rect 18972 23248 19024 23254
rect 18972 23190 19024 23196
rect 18604 23180 18656 23186
rect 18604 23122 18656 23128
rect 18510 23080 18566 23089
rect 18510 23015 18512 23024
rect 18564 23015 18566 23024
rect 18512 22986 18564 22992
rect 18616 22778 18644 23122
rect 18696 23044 18748 23050
rect 18696 22986 18748 22992
rect 18604 22772 18656 22778
rect 18604 22714 18656 22720
rect 18708 21894 18736 22986
rect 18696 21888 18748 21894
rect 18616 21848 18696 21876
rect 18512 21616 18564 21622
rect 18512 21558 18564 21564
rect 18420 21480 18472 21486
rect 18420 21422 18472 21428
rect 18288 21032 18368 21060
rect 18236 21014 18288 21020
rect 18432 20754 18460 21422
rect 18340 20726 18460 20754
rect 17950 20700 18258 20709
rect 17950 20698 17956 20700
rect 18012 20698 18036 20700
rect 18092 20698 18116 20700
rect 18172 20698 18196 20700
rect 18252 20698 18258 20700
rect 18012 20646 18014 20698
rect 18194 20646 18196 20698
rect 17950 20644 17956 20646
rect 18012 20644 18036 20646
rect 18092 20644 18116 20646
rect 18172 20644 18196 20646
rect 18252 20644 18258 20646
rect 17950 20635 18258 20644
rect 18340 20584 18368 20726
rect 18248 20556 18368 20584
rect 18418 20632 18474 20641
rect 18418 20567 18474 20576
rect 17960 19916 18012 19922
rect 17960 19858 18012 19864
rect 17972 19768 18000 19858
rect 18248 19786 18276 20556
rect 18328 20460 18380 20466
rect 18328 20402 18380 20408
rect 18340 20058 18368 20402
rect 18328 20052 18380 20058
rect 18328 19994 18380 20000
rect 17880 19740 18000 19768
rect 18236 19780 18288 19786
rect 17880 19496 17908 19740
rect 18236 19722 18288 19728
rect 17950 19612 18258 19621
rect 17950 19610 17956 19612
rect 18012 19610 18036 19612
rect 18092 19610 18116 19612
rect 18172 19610 18196 19612
rect 18252 19610 18258 19612
rect 18012 19558 18014 19610
rect 18194 19558 18196 19610
rect 17950 19556 17956 19558
rect 18012 19556 18036 19558
rect 18092 19556 18116 19558
rect 18172 19556 18196 19558
rect 18252 19556 18258 19558
rect 17950 19547 18258 19556
rect 17880 19468 18000 19496
rect 17868 18828 17920 18834
rect 17868 18770 17920 18776
rect 17774 18048 17830 18057
rect 17774 17983 17830 17992
rect 17880 17814 17908 18770
rect 17972 18698 18000 19468
rect 18340 19446 18368 19994
rect 18432 19854 18460 20567
rect 18420 19848 18472 19854
rect 18420 19790 18472 19796
rect 18420 19712 18472 19718
rect 18420 19654 18472 19660
rect 18328 19440 18380 19446
rect 18328 19382 18380 19388
rect 18432 19334 18460 19654
rect 18340 19306 18460 19334
rect 18340 18834 18368 19306
rect 18420 19236 18472 19242
rect 18420 19178 18472 19184
rect 18328 18828 18380 18834
rect 18328 18770 18380 18776
rect 18432 18766 18460 19178
rect 18420 18760 18472 18766
rect 18420 18702 18472 18708
rect 17960 18692 18012 18698
rect 17960 18634 18012 18640
rect 18328 18692 18380 18698
rect 18328 18634 18380 18640
rect 17950 18524 18258 18533
rect 17950 18522 17956 18524
rect 18012 18522 18036 18524
rect 18092 18522 18116 18524
rect 18172 18522 18196 18524
rect 18252 18522 18258 18524
rect 18012 18470 18014 18522
rect 18194 18470 18196 18522
rect 17950 18468 17956 18470
rect 18012 18468 18036 18470
rect 18092 18468 18116 18470
rect 18172 18468 18196 18470
rect 18252 18468 18258 18470
rect 17950 18459 18258 18468
rect 18234 18320 18290 18329
rect 18234 18255 18290 18264
rect 18248 18222 18276 18255
rect 18236 18216 18288 18222
rect 18236 18158 18288 18164
rect 17868 17808 17920 17814
rect 17868 17750 17920 17756
rect 17684 17536 17736 17542
rect 17684 17478 17736 17484
rect 17696 17134 17724 17478
rect 17880 17270 17908 17750
rect 17950 17436 18258 17445
rect 17950 17434 17956 17436
rect 18012 17434 18036 17436
rect 18092 17434 18116 17436
rect 18172 17434 18196 17436
rect 18252 17434 18258 17436
rect 18012 17382 18014 17434
rect 18194 17382 18196 17434
rect 17950 17380 17956 17382
rect 18012 17380 18036 17382
rect 18092 17380 18116 17382
rect 18172 17380 18196 17382
rect 18252 17380 18258 17382
rect 17950 17371 18258 17380
rect 17868 17264 17920 17270
rect 17868 17206 17920 17212
rect 18340 17202 18368 18634
rect 18420 18624 18472 18630
rect 18420 18566 18472 18572
rect 18328 17196 18380 17202
rect 18328 17138 18380 17144
rect 17684 17128 17736 17134
rect 17684 17070 17736 17076
rect 17868 16788 17920 16794
rect 17868 16730 17920 16736
rect 17684 16516 17736 16522
rect 17684 16458 17736 16464
rect 17592 16448 17644 16454
rect 17592 16390 17644 16396
rect 17696 15434 17724 16458
rect 17776 16244 17828 16250
rect 17776 16186 17828 16192
rect 17684 15428 17736 15434
rect 17684 15370 17736 15376
rect 17696 15094 17724 15370
rect 17684 15088 17736 15094
rect 17684 15030 17736 15036
rect 17500 14068 17552 14074
rect 17500 14010 17552 14016
rect 17498 13968 17554 13977
rect 17408 13932 17460 13938
rect 17498 13903 17554 13912
rect 17408 13874 17460 13880
rect 17420 12306 17448 13874
rect 17408 12300 17460 12306
rect 17408 12242 17460 12248
rect 17512 11354 17540 13903
rect 17592 13864 17644 13870
rect 17592 13806 17644 13812
rect 17604 13190 17632 13806
rect 17592 13184 17644 13190
rect 17592 13126 17644 13132
rect 17592 12912 17644 12918
rect 17644 12872 17724 12900
rect 17592 12854 17644 12860
rect 17592 12776 17644 12782
rect 17592 12718 17644 12724
rect 17604 12442 17632 12718
rect 17592 12436 17644 12442
rect 17592 12378 17644 12384
rect 17696 11830 17724 12872
rect 17684 11824 17736 11830
rect 17684 11766 17736 11772
rect 17500 11348 17552 11354
rect 17500 11290 17552 11296
rect 17590 10704 17646 10713
rect 17590 10639 17646 10648
rect 17316 10532 17368 10538
rect 17316 10474 17368 10480
rect 17604 10062 17632 10639
rect 17592 10056 17644 10062
rect 17592 9998 17644 10004
rect 17040 9648 17092 9654
rect 17040 9590 17092 9596
rect 17788 9382 17816 16186
rect 17880 14958 17908 16730
rect 18328 16448 18380 16454
rect 18328 16390 18380 16396
rect 17950 16348 18258 16357
rect 17950 16346 17956 16348
rect 18012 16346 18036 16348
rect 18092 16346 18116 16348
rect 18172 16346 18196 16348
rect 18252 16346 18258 16348
rect 18012 16294 18014 16346
rect 18194 16294 18196 16346
rect 17950 16292 17956 16294
rect 18012 16292 18036 16294
rect 18092 16292 18116 16294
rect 18172 16292 18196 16294
rect 18252 16292 18258 16294
rect 17950 16283 18258 16292
rect 17950 15260 18258 15269
rect 17950 15258 17956 15260
rect 18012 15258 18036 15260
rect 18092 15258 18116 15260
rect 18172 15258 18196 15260
rect 18252 15258 18258 15260
rect 18012 15206 18014 15258
rect 18194 15206 18196 15258
rect 17950 15204 17956 15206
rect 18012 15204 18036 15206
rect 18092 15204 18116 15206
rect 18172 15204 18196 15206
rect 18252 15204 18258 15206
rect 17950 15195 18258 15204
rect 17868 14952 17920 14958
rect 17868 14894 17920 14900
rect 17950 14172 18258 14181
rect 17950 14170 17956 14172
rect 18012 14170 18036 14172
rect 18092 14170 18116 14172
rect 18172 14170 18196 14172
rect 18252 14170 18258 14172
rect 18012 14118 18014 14170
rect 18194 14118 18196 14170
rect 17950 14116 17956 14118
rect 18012 14116 18036 14118
rect 18092 14116 18116 14118
rect 18172 14116 18196 14118
rect 18252 14116 18258 14118
rect 17950 14107 18258 14116
rect 17950 13084 18258 13093
rect 17950 13082 17956 13084
rect 18012 13082 18036 13084
rect 18092 13082 18116 13084
rect 18172 13082 18196 13084
rect 18252 13082 18258 13084
rect 18012 13030 18014 13082
rect 18194 13030 18196 13082
rect 17950 13028 17956 13030
rect 18012 13028 18036 13030
rect 18092 13028 18116 13030
rect 18172 13028 18196 13030
rect 18252 13028 18258 13030
rect 17950 13019 18258 13028
rect 17868 12980 17920 12986
rect 17868 12922 17920 12928
rect 17880 12782 17908 12922
rect 17868 12776 17920 12782
rect 17868 12718 17920 12724
rect 17950 11996 18258 12005
rect 17950 11994 17956 11996
rect 18012 11994 18036 11996
rect 18092 11994 18116 11996
rect 18172 11994 18196 11996
rect 18252 11994 18258 11996
rect 18012 11942 18014 11994
rect 18194 11942 18196 11994
rect 17950 11940 17956 11942
rect 18012 11940 18036 11942
rect 18092 11940 18116 11942
rect 18172 11940 18196 11942
rect 18252 11940 18258 11942
rect 17950 11931 18258 11940
rect 18340 11234 18368 16390
rect 18432 12782 18460 18566
rect 18524 18426 18552 21558
rect 18616 21078 18644 21848
rect 18696 21830 18748 21836
rect 18604 21072 18656 21078
rect 18604 21014 18656 21020
rect 18616 20602 18644 21014
rect 18696 21004 18748 21010
rect 18696 20946 18748 20952
rect 18708 20602 18736 20946
rect 18604 20596 18656 20602
rect 18604 20538 18656 20544
rect 18696 20596 18748 20602
rect 18696 20538 18748 20544
rect 18604 20256 18656 20262
rect 18604 20198 18656 20204
rect 18616 19990 18644 20198
rect 18604 19984 18656 19990
rect 18604 19926 18656 19932
rect 18892 19854 18920 23190
rect 18984 23050 19012 23190
rect 19076 23186 19104 24919
rect 19248 24064 19300 24070
rect 19248 24006 19300 24012
rect 19340 24064 19392 24070
rect 19340 24006 19392 24012
rect 19154 23488 19210 23497
rect 19154 23423 19210 23432
rect 19064 23180 19116 23186
rect 19064 23122 19116 23128
rect 19168 23050 19196 23423
rect 18972 23044 19024 23050
rect 18972 22986 19024 22992
rect 19156 23044 19208 23050
rect 19156 22986 19208 22992
rect 19064 22976 19116 22982
rect 19064 22918 19116 22924
rect 19076 22234 19104 22918
rect 18972 22228 19024 22234
rect 18972 22170 19024 22176
rect 19064 22228 19116 22234
rect 19064 22170 19116 22176
rect 18984 21486 19012 22170
rect 19076 22030 19104 22170
rect 19064 22024 19116 22030
rect 19064 21966 19116 21972
rect 18972 21480 19024 21486
rect 18972 21422 19024 21428
rect 19064 21344 19116 21350
rect 19064 21286 19116 21292
rect 18972 20868 19024 20874
rect 18972 20810 19024 20816
rect 18880 19848 18932 19854
rect 18880 19790 18932 19796
rect 18604 19712 18656 19718
rect 18604 19654 18656 19660
rect 18788 19712 18840 19718
rect 18788 19654 18840 19660
rect 18512 18420 18564 18426
rect 18512 18362 18564 18368
rect 18524 16250 18552 18362
rect 18616 17678 18644 19654
rect 18696 19508 18748 19514
rect 18800 19496 18828 19654
rect 18748 19468 18828 19496
rect 18696 19450 18748 19456
rect 18788 19168 18840 19174
rect 18788 19110 18840 19116
rect 18800 18970 18828 19110
rect 18788 18964 18840 18970
rect 18788 18906 18840 18912
rect 18788 18760 18840 18766
rect 18788 18702 18840 18708
rect 18696 18216 18748 18222
rect 18696 18158 18748 18164
rect 18604 17672 18656 17678
rect 18604 17614 18656 17620
rect 18616 17377 18644 17614
rect 18602 17368 18658 17377
rect 18602 17303 18658 17312
rect 18512 16244 18564 16250
rect 18512 16186 18564 16192
rect 18524 14006 18552 16186
rect 18604 15700 18656 15706
rect 18604 15642 18656 15648
rect 18616 15162 18644 15642
rect 18604 15156 18656 15162
rect 18604 15098 18656 15104
rect 18604 14816 18656 14822
rect 18604 14758 18656 14764
rect 18616 14482 18644 14758
rect 18708 14550 18736 18158
rect 18696 14544 18748 14550
rect 18696 14486 18748 14492
rect 18604 14476 18656 14482
rect 18604 14418 18656 14424
rect 18604 14272 18656 14278
rect 18604 14214 18656 14220
rect 18512 14000 18564 14006
rect 18512 13942 18564 13948
rect 18616 12866 18644 14214
rect 18708 13394 18736 14486
rect 18696 13388 18748 13394
rect 18696 13330 18748 13336
rect 18800 13002 18828 18702
rect 18892 17678 18920 19790
rect 18880 17672 18932 17678
rect 18880 17614 18932 17620
rect 18984 17338 19012 20810
rect 19076 19378 19104 21286
rect 19260 20806 19288 24006
rect 19352 23866 19380 24006
rect 19340 23860 19392 23866
rect 19340 23802 19392 23808
rect 19340 23656 19392 23662
rect 19444 23644 19472 24919
rect 19392 23616 19472 23644
rect 19340 23598 19392 23604
rect 19432 23248 19484 23254
rect 19432 23190 19484 23196
rect 19340 23112 19392 23118
rect 19340 23054 19392 23060
rect 19352 22030 19380 23054
rect 19444 22642 19472 23190
rect 19536 22681 19564 26302
rect 19706 26200 19762 27000
rect 20074 26330 20130 27000
rect 20442 26330 20498 27000
rect 19812 26302 20130 26330
rect 19720 24614 19748 26200
rect 19708 24608 19760 24614
rect 19708 24550 19760 24556
rect 19616 23792 19668 23798
rect 19812 23769 19840 26302
rect 20074 26200 20130 26302
rect 20364 26302 20498 26330
rect 20166 25120 20222 25129
rect 20166 25055 20222 25064
rect 19984 24404 20036 24410
rect 19984 24346 20036 24352
rect 20076 24404 20128 24410
rect 20076 24346 20128 24352
rect 19996 24274 20024 24346
rect 19984 24268 20036 24274
rect 19984 24210 20036 24216
rect 19616 23734 19668 23740
rect 19798 23760 19854 23769
rect 19522 22672 19578 22681
rect 19432 22636 19484 22642
rect 19522 22607 19578 22616
rect 19432 22578 19484 22584
rect 19430 22536 19486 22545
rect 19430 22471 19432 22480
rect 19484 22471 19486 22480
rect 19432 22442 19484 22448
rect 19628 22409 19656 23734
rect 19798 23695 19854 23704
rect 19800 23520 19852 23526
rect 19800 23462 19852 23468
rect 19892 23520 19944 23526
rect 19996 23497 20024 24210
rect 20088 24206 20116 24346
rect 20076 24200 20128 24206
rect 20076 24142 20128 24148
rect 20088 23866 20116 24142
rect 20076 23860 20128 23866
rect 20076 23802 20128 23808
rect 20180 23746 20208 25055
rect 20260 24132 20312 24138
rect 20260 24074 20312 24080
rect 20088 23718 20208 23746
rect 19892 23462 19944 23468
rect 19982 23488 20038 23497
rect 19812 22710 19840 23462
rect 19904 23032 19932 23462
rect 19982 23423 20038 23432
rect 19984 23044 20036 23050
rect 19904 23004 19984 23032
rect 19800 22704 19852 22710
rect 19800 22646 19852 22652
rect 19904 22642 19932 23004
rect 19984 22986 20036 22992
rect 19892 22636 19944 22642
rect 19892 22578 19944 22584
rect 19614 22400 19670 22409
rect 19614 22335 19670 22344
rect 19340 22024 19392 22030
rect 19340 21966 19392 21972
rect 19352 21350 19380 21966
rect 19524 21956 19576 21962
rect 19524 21898 19576 21904
rect 19430 21720 19486 21729
rect 19430 21655 19486 21664
rect 19340 21344 19392 21350
rect 19340 21286 19392 21292
rect 19352 20942 19380 21286
rect 19444 21049 19472 21655
rect 19430 21040 19486 21049
rect 19430 20975 19486 20984
rect 19340 20936 19392 20942
rect 19340 20878 19392 20884
rect 19248 20800 19300 20806
rect 19248 20742 19300 20748
rect 19352 20584 19380 20878
rect 19536 20777 19564 21898
rect 19616 21888 19668 21894
rect 19616 21830 19668 21836
rect 19628 21457 19656 21830
rect 19614 21448 19670 21457
rect 19614 21383 19670 21392
rect 19984 21412 20036 21418
rect 19984 21354 20036 21360
rect 19522 20768 19578 20777
rect 19522 20703 19578 20712
rect 19260 20556 19380 20584
rect 19260 20398 19288 20556
rect 19248 20392 19300 20398
rect 19248 20334 19300 20340
rect 19892 20392 19944 20398
rect 19892 20334 19944 20340
rect 19064 19372 19116 19378
rect 19064 19314 19116 19320
rect 19154 19272 19210 19281
rect 19154 19207 19210 19216
rect 19064 18148 19116 18154
rect 19064 18090 19116 18096
rect 18972 17332 19024 17338
rect 18972 17274 19024 17280
rect 18880 16448 18932 16454
rect 18880 16390 18932 16396
rect 18892 15570 18920 16390
rect 19076 16250 19104 18090
rect 19064 16244 19116 16250
rect 19064 16186 19116 16192
rect 18972 16108 19024 16114
rect 18972 16050 19024 16056
rect 19064 16108 19116 16114
rect 19064 16050 19116 16056
rect 18880 15564 18932 15570
rect 18880 15506 18932 15512
rect 18984 15162 19012 16050
rect 18972 15156 19024 15162
rect 18972 15098 19024 15104
rect 18880 15020 18932 15026
rect 18880 14962 18932 14968
rect 18892 14890 18920 14962
rect 18880 14884 18932 14890
rect 18880 14826 18932 14832
rect 18878 14104 18934 14113
rect 18878 14039 18934 14048
rect 18892 13841 18920 14039
rect 18878 13832 18934 13841
rect 18878 13767 18934 13776
rect 18708 12986 18828 13002
rect 18696 12980 18828 12986
rect 18748 12974 18828 12980
rect 18696 12922 18748 12928
rect 18788 12912 18840 12918
rect 18512 12844 18564 12850
rect 18616 12838 18736 12866
rect 18788 12854 18840 12860
rect 18512 12786 18564 12792
rect 18420 12776 18472 12782
rect 18420 12718 18472 12724
rect 18524 12434 18552 12786
rect 18604 12708 18656 12714
rect 18604 12650 18656 12656
rect 17972 11206 18368 11234
rect 18432 12406 18552 12434
rect 18432 11218 18460 12406
rect 18616 11694 18644 12650
rect 18604 11688 18656 11694
rect 18604 11630 18656 11636
rect 18512 11620 18564 11626
rect 18512 11562 18564 11568
rect 18420 11212 18472 11218
rect 17972 11098 18000 11206
rect 18420 11154 18472 11160
rect 18524 11150 18552 11562
rect 18512 11144 18564 11150
rect 17880 11070 18000 11098
rect 18326 11112 18382 11121
rect 17880 10810 17908 11070
rect 18512 11086 18564 11092
rect 18326 11047 18382 11056
rect 17950 10908 18258 10917
rect 17950 10906 17956 10908
rect 18012 10906 18036 10908
rect 18092 10906 18116 10908
rect 18172 10906 18196 10908
rect 18252 10906 18258 10908
rect 18012 10854 18014 10906
rect 18194 10854 18196 10906
rect 17950 10852 17956 10854
rect 18012 10852 18036 10854
rect 18092 10852 18116 10854
rect 18172 10852 18196 10854
rect 18252 10852 18258 10854
rect 17950 10843 18258 10852
rect 18340 10810 18368 11047
rect 17868 10804 17920 10810
rect 17868 10746 17920 10752
rect 18328 10804 18380 10810
rect 18328 10746 18380 10752
rect 18708 10674 18736 12838
rect 18800 11558 18828 12854
rect 18788 11552 18840 11558
rect 18788 11494 18840 11500
rect 18696 10668 18748 10674
rect 18696 10610 18748 10616
rect 17950 9820 18258 9829
rect 17950 9818 17956 9820
rect 18012 9818 18036 9820
rect 18092 9818 18116 9820
rect 18172 9818 18196 9820
rect 18252 9818 18258 9820
rect 18012 9766 18014 9818
rect 18194 9766 18196 9818
rect 17950 9764 17956 9766
rect 18012 9764 18036 9766
rect 18092 9764 18116 9766
rect 18172 9764 18196 9766
rect 18252 9764 18258 9766
rect 17950 9755 18258 9764
rect 17776 9376 17828 9382
rect 17776 9318 17828 9324
rect 17950 8732 18258 8741
rect 17950 8730 17956 8732
rect 18012 8730 18036 8732
rect 18092 8730 18116 8732
rect 18172 8730 18196 8732
rect 18252 8730 18258 8732
rect 18012 8678 18014 8730
rect 18194 8678 18196 8730
rect 17950 8676 17956 8678
rect 18012 8676 18036 8678
rect 18092 8676 18116 8678
rect 18172 8676 18196 8678
rect 18252 8676 18258 8678
rect 17950 8667 18258 8676
rect 17950 7644 18258 7653
rect 17950 7642 17956 7644
rect 18012 7642 18036 7644
rect 18092 7642 18116 7644
rect 18172 7642 18196 7644
rect 18252 7642 18258 7644
rect 18012 7590 18014 7642
rect 18194 7590 18196 7642
rect 17950 7588 17956 7590
rect 18012 7588 18036 7590
rect 18092 7588 18116 7590
rect 18172 7588 18196 7590
rect 18252 7588 18258 7590
rect 17950 7579 18258 7588
rect 15200 6724 15252 6730
rect 15200 6666 15252 6672
rect 17950 6556 18258 6565
rect 17950 6554 17956 6556
rect 18012 6554 18036 6556
rect 18092 6554 18116 6556
rect 18172 6554 18196 6556
rect 18252 6554 18258 6556
rect 18012 6502 18014 6554
rect 18194 6502 18196 6554
rect 17950 6500 17956 6502
rect 18012 6500 18036 6502
rect 18092 6500 18116 6502
rect 18172 6500 18196 6502
rect 18252 6500 18258 6502
rect 17950 6491 18258 6500
rect 9312 6452 9364 6458
rect 9312 6394 9364 6400
rect 6828 6316 6880 6322
rect 6828 6258 6880 6264
rect 2950 6012 3258 6021
rect 2950 6010 2956 6012
rect 3012 6010 3036 6012
rect 3092 6010 3116 6012
rect 3172 6010 3196 6012
rect 3252 6010 3258 6012
rect 3012 5958 3014 6010
rect 3194 5958 3196 6010
rect 2950 5956 2956 5958
rect 3012 5956 3036 5958
rect 3092 5956 3116 5958
rect 3172 5956 3196 5958
rect 3252 5956 3258 5958
rect 2950 5947 3258 5956
rect 2950 4924 3258 4933
rect 2950 4922 2956 4924
rect 3012 4922 3036 4924
rect 3092 4922 3116 4924
rect 3172 4922 3196 4924
rect 3252 4922 3258 4924
rect 3012 4870 3014 4922
rect 3194 4870 3196 4922
rect 2950 4868 2956 4870
rect 3012 4868 3036 4870
rect 3092 4868 3116 4870
rect 3172 4868 3196 4870
rect 3252 4868 3258 4870
rect 2950 4859 3258 4868
rect 2950 3836 3258 3845
rect 2950 3834 2956 3836
rect 3012 3834 3036 3836
rect 3092 3834 3116 3836
rect 3172 3834 3196 3836
rect 3252 3834 3258 3836
rect 3012 3782 3014 3834
rect 3194 3782 3196 3834
rect 2950 3780 2956 3782
rect 3012 3780 3036 3782
rect 3092 3780 3116 3782
rect 3172 3780 3196 3782
rect 3252 3780 3258 3782
rect 2950 3771 3258 3780
rect 6840 3194 6868 6258
rect 12950 6012 13258 6021
rect 12950 6010 12956 6012
rect 13012 6010 13036 6012
rect 13092 6010 13116 6012
rect 13172 6010 13196 6012
rect 13252 6010 13258 6012
rect 13012 5958 13014 6010
rect 13194 5958 13196 6010
rect 12950 5956 12956 5958
rect 13012 5956 13036 5958
rect 13092 5956 13116 5958
rect 13172 5956 13196 5958
rect 13252 5956 13258 5958
rect 12950 5947 13258 5956
rect 7950 5468 8258 5477
rect 7950 5466 7956 5468
rect 8012 5466 8036 5468
rect 8092 5466 8116 5468
rect 8172 5466 8196 5468
rect 8252 5466 8258 5468
rect 8012 5414 8014 5466
rect 8194 5414 8196 5466
rect 7950 5412 7956 5414
rect 8012 5412 8036 5414
rect 8092 5412 8116 5414
rect 8172 5412 8196 5414
rect 8252 5412 8258 5414
rect 7950 5403 8258 5412
rect 17950 5468 18258 5477
rect 17950 5466 17956 5468
rect 18012 5466 18036 5468
rect 18092 5466 18116 5468
rect 18172 5466 18196 5468
rect 18252 5466 18258 5468
rect 18012 5414 18014 5466
rect 18194 5414 18196 5466
rect 17950 5412 17956 5414
rect 18012 5412 18036 5414
rect 18092 5412 18116 5414
rect 18172 5412 18196 5414
rect 18252 5412 18258 5414
rect 17950 5403 18258 5412
rect 12950 4924 13258 4933
rect 12950 4922 12956 4924
rect 13012 4922 13036 4924
rect 13092 4922 13116 4924
rect 13172 4922 13196 4924
rect 13252 4922 13258 4924
rect 13012 4870 13014 4922
rect 13194 4870 13196 4922
rect 12950 4868 12956 4870
rect 13012 4868 13036 4870
rect 13092 4868 13116 4870
rect 13172 4868 13196 4870
rect 13252 4868 13258 4870
rect 12950 4859 13258 4868
rect 7950 4380 8258 4389
rect 7950 4378 7956 4380
rect 8012 4378 8036 4380
rect 8092 4378 8116 4380
rect 8172 4378 8196 4380
rect 8252 4378 8258 4380
rect 8012 4326 8014 4378
rect 8194 4326 8196 4378
rect 7950 4324 7956 4326
rect 8012 4324 8036 4326
rect 8092 4324 8116 4326
rect 8172 4324 8196 4326
rect 8252 4324 8258 4326
rect 7950 4315 8258 4324
rect 17950 4380 18258 4389
rect 17950 4378 17956 4380
rect 18012 4378 18036 4380
rect 18092 4378 18116 4380
rect 18172 4378 18196 4380
rect 18252 4378 18258 4380
rect 18012 4326 18014 4378
rect 18194 4326 18196 4378
rect 17950 4324 17956 4326
rect 18012 4324 18036 4326
rect 18092 4324 18116 4326
rect 18172 4324 18196 4326
rect 18252 4324 18258 4326
rect 17950 4315 18258 4324
rect 18984 4078 19012 15098
rect 19076 13530 19104 16050
rect 19168 14278 19196 19207
rect 19260 18698 19288 20334
rect 19616 20256 19668 20262
rect 19616 20198 19668 20204
rect 19338 19816 19394 19825
rect 19338 19751 19394 19760
rect 19352 19514 19380 19751
rect 19524 19712 19576 19718
rect 19524 19654 19576 19660
rect 19340 19508 19392 19514
rect 19340 19450 19392 19456
rect 19536 19417 19564 19654
rect 19522 19408 19578 19417
rect 19522 19343 19578 19352
rect 19628 18766 19656 20198
rect 19708 19848 19760 19854
rect 19708 19790 19760 19796
rect 19616 18760 19668 18766
rect 19616 18702 19668 18708
rect 19248 18692 19300 18698
rect 19248 18634 19300 18640
rect 19524 18624 19576 18630
rect 19444 18584 19524 18612
rect 19338 18320 19394 18329
rect 19338 18255 19394 18264
rect 19246 16552 19302 16561
rect 19246 16487 19302 16496
rect 19260 15638 19288 16487
rect 19352 15706 19380 18255
rect 19444 18222 19472 18584
rect 19524 18566 19576 18572
rect 19522 18456 19578 18465
rect 19720 18426 19748 19790
rect 19904 19446 19932 20334
rect 19892 19440 19944 19446
rect 19892 19382 19944 19388
rect 19904 19310 19932 19382
rect 19892 19304 19944 19310
rect 19892 19246 19944 19252
rect 19522 18391 19578 18400
rect 19708 18420 19760 18426
rect 19536 18290 19564 18391
rect 19708 18362 19760 18368
rect 19524 18284 19576 18290
rect 19524 18226 19576 18232
rect 19432 18216 19484 18222
rect 19432 18158 19484 18164
rect 19614 17912 19670 17921
rect 19614 17847 19670 17856
rect 19432 17808 19484 17814
rect 19432 17750 19484 17756
rect 19444 16794 19472 17750
rect 19524 17536 19576 17542
rect 19524 17478 19576 17484
rect 19432 16788 19484 16794
rect 19432 16730 19484 16736
rect 19340 15700 19392 15706
rect 19340 15642 19392 15648
rect 19248 15632 19300 15638
rect 19248 15574 19300 15580
rect 19340 14952 19392 14958
rect 19340 14894 19392 14900
rect 19430 14920 19486 14929
rect 19156 14272 19208 14278
rect 19156 14214 19208 14220
rect 19352 14074 19380 14894
rect 19430 14855 19486 14864
rect 19340 14068 19392 14074
rect 19340 14010 19392 14016
rect 19248 13864 19300 13870
rect 19248 13806 19300 13812
rect 19064 13524 19116 13530
rect 19064 13466 19116 13472
rect 19062 13424 19118 13433
rect 19062 13359 19118 13368
rect 19076 9586 19104 13359
rect 19154 12336 19210 12345
rect 19154 12271 19210 12280
rect 19168 11830 19196 12271
rect 19156 11824 19208 11830
rect 19156 11766 19208 11772
rect 19168 11150 19196 11766
rect 19260 11354 19288 13806
rect 19352 12238 19380 14010
rect 19444 13938 19472 14855
rect 19432 13932 19484 13938
rect 19432 13874 19484 13880
rect 19432 13320 19484 13326
rect 19432 13262 19484 13268
rect 19340 12232 19392 12238
rect 19340 12174 19392 12180
rect 19352 11898 19380 12174
rect 19340 11892 19392 11898
rect 19340 11834 19392 11840
rect 19444 11762 19472 13262
rect 19536 12986 19564 17478
rect 19628 16998 19656 17847
rect 19720 17105 19748 18362
rect 19798 18320 19854 18329
rect 19798 18255 19854 18264
rect 19812 18222 19840 18255
rect 19800 18216 19852 18222
rect 19800 18158 19852 18164
rect 19892 18080 19944 18086
rect 19892 18022 19944 18028
rect 19800 17740 19852 17746
rect 19800 17682 19852 17688
rect 19706 17096 19762 17105
rect 19706 17031 19762 17040
rect 19616 16992 19668 16998
rect 19616 16934 19668 16940
rect 19708 15360 19760 15366
rect 19708 15302 19760 15308
rect 19720 14521 19748 15302
rect 19706 14512 19762 14521
rect 19706 14447 19762 14456
rect 19812 14226 19840 17682
rect 19904 14414 19932 18022
rect 19996 15502 20024 21354
rect 20088 18426 20116 23718
rect 20272 22642 20300 24074
rect 20260 22636 20312 22642
rect 20260 22578 20312 22584
rect 20260 22432 20312 22438
rect 20260 22374 20312 22380
rect 20272 22166 20300 22374
rect 20260 22160 20312 22166
rect 20260 22102 20312 22108
rect 20168 22092 20220 22098
rect 20168 22034 20220 22040
rect 20180 21690 20208 22034
rect 20258 21856 20314 21865
rect 20258 21791 20314 21800
rect 20168 21684 20220 21690
rect 20168 21626 20220 21632
rect 20272 21400 20300 21791
rect 20364 21729 20392 26302
rect 20442 26200 20498 26302
rect 20810 26200 20866 27000
rect 21178 26200 21234 27000
rect 21270 26344 21326 26353
rect 21546 26330 21602 27000
rect 21326 26302 21602 26330
rect 21270 26279 21326 26288
rect 21546 26200 21602 26302
rect 21824 26308 21876 26314
rect 21824 26250 21876 26256
rect 20628 24880 20680 24886
rect 20824 24857 20852 26200
rect 20628 24822 20680 24828
rect 20810 24848 20866 24857
rect 20640 24682 20668 24822
rect 20810 24783 20866 24792
rect 20628 24676 20680 24682
rect 20628 24618 20680 24624
rect 20640 23662 20668 24618
rect 20996 24064 21048 24070
rect 20996 24006 21048 24012
rect 20628 23656 20680 23662
rect 20628 23598 20680 23604
rect 20444 23520 20496 23526
rect 20444 23462 20496 23468
rect 20456 23089 20484 23462
rect 20720 23180 20772 23186
rect 20720 23122 20772 23128
rect 20442 23080 20498 23089
rect 20442 23015 20498 23024
rect 20534 22128 20590 22137
rect 20534 22063 20590 22072
rect 20350 21720 20406 21729
rect 20350 21655 20406 21664
rect 20444 21684 20496 21690
rect 20444 21626 20496 21632
rect 20456 21593 20484 21626
rect 20442 21584 20498 21593
rect 20442 21519 20498 21528
rect 20180 21372 20300 21400
rect 20076 18420 20128 18426
rect 20076 18362 20128 18368
rect 20088 17678 20116 18362
rect 20180 17814 20208 21372
rect 20258 21312 20314 21321
rect 20258 21247 20314 21256
rect 20168 17808 20220 17814
rect 20168 17750 20220 17756
rect 20076 17672 20128 17678
rect 20076 17614 20128 17620
rect 20180 17338 20208 17750
rect 20272 17542 20300 21247
rect 20350 21040 20406 21049
rect 20350 20975 20406 20984
rect 20260 17536 20312 17542
rect 20260 17478 20312 17484
rect 20168 17332 20220 17338
rect 20168 17274 20220 17280
rect 20168 17060 20220 17066
rect 20088 17020 20168 17048
rect 19984 15496 20036 15502
rect 19984 15438 20036 15444
rect 19984 14612 20036 14618
rect 19984 14554 20036 14560
rect 19892 14408 19944 14414
rect 19892 14350 19944 14356
rect 19720 14198 19840 14226
rect 19616 13524 19668 13530
rect 19616 13466 19668 13472
rect 19524 12980 19576 12986
rect 19524 12922 19576 12928
rect 19628 12866 19656 13466
rect 19536 12838 19656 12866
rect 19432 11756 19484 11762
rect 19432 11698 19484 11704
rect 19536 11354 19564 12838
rect 19720 12170 19748 14198
rect 19892 13728 19944 13734
rect 19892 13670 19944 13676
rect 19904 13258 19932 13670
rect 19892 13252 19944 13258
rect 19892 13194 19944 13200
rect 19800 12640 19852 12646
rect 19800 12582 19852 12588
rect 19812 12434 19840 12582
rect 19996 12434 20024 14554
rect 20088 14006 20116 17020
rect 20168 17002 20220 17008
rect 20260 16040 20312 16046
rect 20260 15982 20312 15988
rect 20168 15564 20220 15570
rect 20168 15506 20220 15512
rect 20180 14657 20208 15506
rect 20272 14793 20300 15982
rect 20364 15910 20392 20975
rect 20548 20262 20576 22063
rect 20732 21078 20760 23122
rect 20904 22772 20956 22778
rect 20904 22714 20956 22720
rect 20812 22568 20864 22574
rect 20812 22510 20864 22516
rect 20824 21894 20852 22510
rect 20916 21962 20944 22714
rect 20904 21956 20956 21962
rect 20904 21898 20956 21904
rect 20812 21888 20864 21894
rect 20812 21830 20864 21836
rect 20812 21548 20864 21554
rect 20812 21490 20864 21496
rect 20720 21072 20772 21078
rect 20720 21014 20772 21020
rect 20720 20936 20772 20942
rect 20720 20878 20772 20884
rect 20628 20460 20680 20466
rect 20732 20448 20760 20878
rect 20824 20777 20852 21490
rect 20810 20768 20866 20777
rect 20810 20703 20866 20712
rect 20916 20602 20944 21898
rect 21008 21486 21036 24006
rect 21088 22432 21140 22438
rect 21088 22374 21140 22380
rect 21100 21486 21128 22374
rect 21192 22137 21220 26200
rect 21836 26058 21864 26250
rect 21914 26200 21970 27000
rect 22192 26376 22244 26382
rect 22192 26318 22244 26324
rect 21928 26058 21956 26200
rect 21836 26030 21956 26058
rect 22204 26058 22232 26318
rect 22282 26200 22338 27000
rect 22650 26200 22706 27000
rect 23018 26330 23074 27000
rect 22756 26302 23074 26330
rect 22296 26058 22324 26200
rect 22204 26030 22324 26058
rect 22376 24404 22428 24410
rect 22376 24346 22428 24352
rect 22284 24200 22336 24206
rect 22284 24142 22336 24148
rect 21364 24064 21416 24070
rect 21364 24006 21416 24012
rect 21824 24064 21876 24070
rect 21824 24006 21876 24012
rect 21178 22128 21234 22137
rect 21178 22063 21234 22072
rect 21272 21888 21324 21894
rect 21272 21830 21324 21836
rect 20996 21480 21048 21486
rect 20996 21422 21048 21428
rect 21088 21480 21140 21486
rect 21088 21422 21140 21428
rect 21008 20942 21036 21422
rect 21178 21312 21234 21321
rect 21178 21247 21234 21256
rect 21192 21078 21220 21247
rect 21180 21072 21232 21078
rect 21180 21014 21232 21020
rect 20996 20936 21048 20942
rect 21048 20896 21128 20924
rect 20996 20878 21048 20884
rect 20904 20596 20956 20602
rect 20904 20538 20956 20544
rect 20680 20420 20760 20448
rect 20628 20402 20680 20408
rect 20536 20256 20588 20262
rect 20536 20198 20588 20204
rect 20442 20088 20498 20097
rect 20442 20023 20498 20032
rect 20628 20052 20680 20058
rect 20456 19378 20484 20023
rect 20732 20040 20760 20420
rect 20812 20392 20864 20398
rect 20812 20334 20864 20340
rect 20680 20012 20760 20040
rect 20628 19994 20680 20000
rect 20536 19780 20588 19786
rect 20536 19722 20588 19728
rect 20444 19372 20496 19378
rect 20444 19314 20496 19320
rect 20444 18624 20496 18630
rect 20444 18566 20496 18572
rect 20456 18290 20484 18566
rect 20444 18284 20496 18290
rect 20444 18226 20496 18232
rect 20444 18080 20496 18086
rect 20444 18022 20496 18028
rect 20352 15904 20404 15910
rect 20352 15846 20404 15852
rect 20350 15464 20406 15473
rect 20350 15399 20406 15408
rect 20258 14784 20314 14793
rect 20258 14719 20314 14728
rect 20166 14648 20222 14657
rect 20166 14583 20222 14592
rect 20260 14612 20312 14618
rect 20260 14554 20312 14560
rect 20272 14074 20300 14554
rect 20260 14068 20312 14074
rect 20260 14010 20312 14016
rect 20076 14000 20128 14006
rect 20076 13942 20128 13948
rect 20088 13734 20116 13942
rect 20272 13870 20300 14010
rect 20260 13864 20312 13870
rect 20260 13806 20312 13812
rect 20076 13728 20128 13734
rect 20076 13670 20128 13676
rect 20272 13258 20300 13806
rect 20364 13433 20392 15399
rect 20456 14074 20484 18022
rect 20548 17338 20576 19722
rect 20720 19712 20772 19718
rect 20640 19660 20720 19666
rect 20640 19654 20772 19660
rect 20640 19638 20760 19654
rect 20640 18698 20668 19638
rect 20824 19514 20852 20334
rect 20904 20324 20956 20330
rect 20904 20266 20956 20272
rect 20916 19922 20944 20266
rect 20994 20224 21050 20233
rect 20994 20159 21050 20168
rect 20904 19916 20956 19922
rect 20904 19858 20956 19864
rect 20812 19508 20864 19514
rect 20812 19450 20864 19456
rect 20904 19372 20956 19378
rect 20904 19314 20956 19320
rect 20720 19168 20772 19174
rect 20720 19110 20772 19116
rect 20628 18692 20680 18698
rect 20628 18634 20680 18640
rect 20628 18352 20680 18358
rect 20626 18320 20628 18329
rect 20680 18320 20682 18329
rect 20626 18255 20682 18264
rect 20628 17876 20680 17882
rect 20628 17818 20680 17824
rect 20640 17338 20668 17818
rect 20536 17332 20588 17338
rect 20536 17274 20588 17280
rect 20628 17332 20680 17338
rect 20628 17274 20680 17280
rect 20732 16969 20760 19110
rect 20916 18630 20944 19314
rect 21008 19174 21036 20159
rect 21100 20058 21128 20896
rect 21180 20800 21232 20806
rect 21180 20742 21232 20748
rect 21088 20052 21140 20058
rect 21088 19994 21140 20000
rect 21086 19952 21142 19961
rect 21086 19887 21142 19896
rect 20996 19168 21048 19174
rect 20996 19110 21048 19116
rect 20904 18624 20956 18630
rect 20904 18566 20956 18572
rect 20810 18456 20866 18465
rect 20810 18391 20866 18400
rect 20824 18290 20852 18391
rect 20812 18284 20864 18290
rect 20812 18226 20864 18232
rect 20812 18148 20864 18154
rect 20812 18090 20864 18096
rect 20718 16960 20774 16969
rect 20718 16895 20774 16904
rect 20720 16788 20772 16794
rect 20720 16730 20772 16736
rect 20628 16244 20680 16250
rect 20628 16186 20680 16192
rect 20640 16114 20668 16186
rect 20628 16108 20680 16114
rect 20628 16050 20680 16056
rect 20536 15904 20588 15910
rect 20536 15846 20588 15852
rect 20548 14550 20576 15846
rect 20628 15156 20680 15162
rect 20732 15144 20760 16730
rect 20680 15116 20760 15144
rect 20628 15098 20680 15104
rect 20536 14544 20588 14550
rect 20536 14486 20588 14492
rect 20536 14408 20588 14414
rect 20536 14350 20588 14356
rect 20444 14068 20496 14074
rect 20444 14010 20496 14016
rect 20548 13530 20576 14350
rect 20628 14340 20680 14346
rect 20628 14282 20680 14288
rect 20536 13524 20588 13530
rect 20536 13466 20588 13472
rect 20350 13424 20406 13433
rect 20640 13376 20668 14282
rect 20720 13728 20772 13734
rect 20720 13670 20772 13676
rect 20350 13359 20406 13368
rect 20548 13348 20668 13376
rect 20260 13252 20312 13258
rect 20260 13194 20312 13200
rect 20272 12782 20300 13194
rect 20260 12776 20312 12782
rect 20180 12736 20260 12764
rect 19812 12406 19932 12434
rect 19996 12406 20116 12434
rect 19800 12300 19852 12306
rect 19800 12242 19852 12248
rect 19616 12164 19668 12170
rect 19616 12106 19668 12112
rect 19708 12164 19760 12170
rect 19708 12106 19760 12112
rect 19628 11354 19656 12106
rect 19720 11558 19748 12106
rect 19812 11830 19840 12242
rect 19800 11824 19852 11830
rect 19800 11766 19852 11772
rect 19708 11552 19760 11558
rect 19708 11494 19760 11500
rect 19248 11348 19300 11354
rect 19248 11290 19300 11296
rect 19524 11348 19576 11354
rect 19524 11290 19576 11296
rect 19616 11348 19668 11354
rect 19616 11290 19668 11296
rect 19800 11280 19852 11286
rect 19800 11222 19852 11228
rect 19156 11144 19208 11150
rect 19156 11086 19208 11092
rect 19430 11112 19486 11121
rect 19430 11047 19486 11056
rect 19444 10198 19472 11047
rect 19432 10192 19484 10198
rect 19432 10134 19484 10140
rect 19064 9580 19116 9586
rect 19064 9522 19116 9528
rect 19524 9580 19576 9586
rect 19524 9522 19576 9528
rect 19076 9178 19104 9522
rect 19338 9480 19394 9489
rect 19338 9415 19340 9424
rect 19392 9415 19394 9424
rect 19340 9386 19392 9392
rect 19536 9178 19564 9522
rect 19064 9172 19116 9178
rect 19064 9114 19116 9120
rect 19524 9172 19576 9178
rect 19524 9114 19576 9120
rect 19706 8392 19762 8401
rect 19706 8327 19708 8336
rect 19760 8327 19762 8336
rect 19708 8298 19760 8304
rect 19812 7886 19840 11222
rect 19904 8430 19932 12406
rect 19984 12096 20036 12102
rect 19984 12038 20036 12044
rect 19892 8424 19944 8430
rect 19892 8366 19944 8372
rect 19800 7880 19852 7886
rect 19800 7822 19852 7828
rect 18972 4072 19024 4078
rect 18972 4014 19024 4020
rect 12950 3836 13258 3845
rect 12950 3834 12956 3836
rect 13012 3834 13036 3836
rect 13092 3834 13116 3836
rect 13172 3834 13196 3836
rect 13252 3834 13258 3836
rect 13012 3782 13014 3834
rect 13194 3782 13196 3834
rect 12950 3780 12956 3782
rect 13012 3780 13036 3782
rect 13092 3780 13116 3782
rect 13172 3780 13196 3782
rect 13252 3780 13258 3782
rect 12950 3771 13258 3780
rect 7950 3292 8258 3301
rect 7950 3290 7956 3292
rect 8012 3290 8036 3292
rect 8092 3290 8116 3292
rect 8172 3290 8196 3292
rect 8252 3290 8258 3292
rect 8012 3238 8014 3290
rect 8194 3238 8196 3290
rect 7950 3236 7956 3238
rect 8012 3236 8036 3238
rect 8092 3236 8116 3238
rect 8172 3236 8196 3238
rect 8252 3236 8258 3238
rect 7950 3227 8258 3236
rect 17950 3292 18258 3301
rect 17950 3290 17956 3292
rect 18012 3290 18036 3292
rect 18092 3290 18116 3292
rect 18172 3290 18196 3292
rect 18252 3290 18258 3292
rect 18012 3238 18014 3290
rect 18194 3238 18196 3290
rect 17950 3236 17956 3238
rect 18012 3236 18036 3238
rect 18092 3236 18116 3238
rect 18172 3236 18196 3238
rect 18252 3236 18258 3238
rect 17950 3227 18258 3236
rect 6828 3188 6880 3194
rect 6828 3130 6880 3136
rect 19996 3058 20024 12038
rect 20088 11150 20116 12406
rect 20180 12170 20208 12736
rect 20260 12718 20312 12724
rect 20444 12708 20496 12714
rect 20444 12650 20496 12656
rect 20260 12640 20312 12646
rect 20260 12582 20312 12588
rect 20272 12434 20300 12582
rect 20272 12406 20392 12434
rect 20168 12164 20220 12170
rect 20168 12106 20220 12112
rect 20180 11830 20208 12106
rect 20168 11824 20220 11830
rect 20168 11766 20220 11772
rect 20076 11144 20128 11150
rect 20076 11086 20128 11092
rect 20180 11014 20208 11766
rect 20260 11280 20312 11286
rect 20260 11222 20312 11228
rect 20076 11008 20128 11014
rect 20076 10950 20128 10956
rect 20168 11008 20220 11014
rect 20168 10950 20220 10956
rect 20088 3534 20116 10950
rect 20168 10668 20220 10674
rect 20168 10610 20220 10616
rect 20180 10266 20208 10610
rect 20168 10260 20220 10266
rect 20168 10202 20220 10208
rect 20272 9586 20300 11222
rect 20260 9580 20312 9586
rect 20260 9522 20312 9528
rect 20364 7410 20392 12406
rect 20456 12306 20484 12650
rect 20444 12300 20496 12306
rect 20444 12242 20496 12248
rect 20548 10742 20576 13348
rect 20628 12844 20680 12850
rect 20628 12786 20680 12792
rect 20640 12102 20668 12786
rect 20628 12096 20680 12102
rect 20628 12038 20680 12044
rect 20536 10736 20588 10742
rect 20536 10678 20588 10684
rect 20732 10674 20760 13670
rect 20824 13190 20852 18090
rect 20916 16250 20944 18566
rect 20994 18456 21050 18465
rect 20994 18391 21050 18400
rect 20904 16244 20956 16250
rect 20904 16186 20956 16192
rect 20904 15088 20956 15094
rect 20904 15030 20956 15036
rect 20916 14618 20944 15030
rect 20904 14612 20956 14618
rect 20904 14554 20956 14560
rect 20812 13184 20864 13190
rect 20812 13126 20864 13132
rect 21008 12782 21036 18391
rect 21100 18358 21128 19887
rect 21088 18352 21140 18358
rect 21088 18294 21140 18300
rect 21192 18290 21220 20742
rect 21284 20097 21312 21830
rect 21376 21185 21404 24006
rect 21454 22808 21510 22817
rect 21454 22743 21510 22752
rect 21468 21894 21496 22743
rect 21836 22234 21864 24006
rect 22296 23866 22324 24142
rect 22284 23860 22336 23866
rect 22284 23802 22336 23808
rect 22100 23792 22152 23798
rect 22100 23734 22152 23740
rect 22112 23633 22140 23734
rect 22098 23624 22154 23633
rect 22098 23559 22154 23568
rect 22296 23186 22324 23802
rect 22388 23474 22416 24346
rect 22560 24268 22612 24274
rect 22560 24210 22612 24216
rect 22572 23662 22600 24210
rect 22560 23656 22612 23662
rect 22560 23598 22612 23604
rect 22388 23446 22508 23474
rect 22284 23180 22336 23186
rect 22284 23122 22336 23128
rect 22192 23044 22244 23050
rect 22192 22986 22244 22992
rect 22376 23044 22428 23050
rect 22376 22986 22428 22992
rect 21824 22228 21876 22234
rect 21824 22170 21876 22176
rect 21640 22160 21692 22166
rect 21640 22102 21692 22108
rect 21730 22128 21786 22137
rect 21456 21888 21508 21894
rect 21456 21830 21508 21836
rect 21548 21684 21600 21690
rect 21548 21626 21600 21632
rect 21456 21548 21508 21554
rect 21456 21490 21508 21496
rect 21362 21176 21418 21185
rect 21362 21111 21418 21120
rect 21270 20088 21326 20097
rect 21270 20023 21326 20032
rect 21364 19780 21416 19786
rect 21364 19722 21416 19728
rect 21272 19508 21324 19514
rect 21272 19450 21324 19456
rect 21180 18284 21232 18290
rect 21180 18226 21232 18232
rect 21180 18148 21232 18154
rect 21180 18090 21232 18096
rect 21192 18057 21220 18090
rect 21178 18048 21234 18057
rect 21178 17983 21234 17992
rect 21086 17776 21142 17785
rect 21086 17711 21142 17720
rect 21100 17513 21128 17711
rect 21086 17504 21142 17513
rect 21086 17439 21142 17448
rect 21088 17128 21140 17134
rect 21088 17070 21140 17076
rect 21100 16794 21128 17070
rect 21088 16788 21140 16794
rect 21088 16730 21140 16736
rect 21088 16584 21140 16590
rect 21088 16526 21140 16532
rect 21100 16250 21128 16526
rect 21088 16244 21140 16250
rect 21088 16186 21140 16192
rect 21088 16040 21140 16046
rect 21088 15982 21140 15988
rect 20996 12776 21048 12782
rect 20996 12718 21048 12724
rect 20904 11688 20956 11694
rect 20904 11630 20956 11636
rect 20812 11620 20864 11626
rect 20812 11562 20864 11568
rect 20824 11354 20852 11562
rect 20812 11348 20864 11354
rect 20812 11290 20864 11296
rect 20444 10668 20496 10674
rect 20444 10610 20496 10616
rect 20720 10668 20772 10674
rect 20720 10610 20772 10616
rect 20456 10470 20484 10610
rect 20444 10464 20496 10470
rect 20444 10406 20496 10412
rect 20812 10464 20864 10470
rect 20812 10406 20864 10412
rect 20718 10296 20774 10305
rect 20718 10231 20720 10240
rect 20772 10231 20774 10240
rect 20720 10202 20772 10208
rect 20720 10056 20772 10062
rect 20720 9998 20772 10004
rect 20444 9920 20496 9926
rect 20444 9862 20496 9868
rect 20456 9654 20484 9862
rect 20732 9761 20760 9998
rect 20718 9752 20774 9761
rect 20628 9716 20680 9722
rect 20718 9687 20774 9696
rect 20628 9658 20680 9664
rect 20444 9648 20496 9654
rect 20444 9590 20496 9596
rect 20536 9376 20588 9382
rect 20536 9318 20588 9324
rect 20548 8838 20576 9318
rect 20536 8832 20588 8838
rect 20536 8774 20588 8780
rect 20534 7984 20590 7993
rect 20534 7919 20590 7928
rect 20352 7404 20404 7410
rect 20352 7346 20404 7352
rect 20548 5914 20576 7919
rect 20536 5908 20588 5914
rect 20536 5850 20588 5856
rect 20258 5672 20314 5681
rect 20258 5607 20314 5616
rect 20272 4146 20300 5607
rect 20260 4140 20312 4146
rect 20260 4082 20312 4088
rect 20168 4072 20220 4078
rect 20168 4014 20220 4020
rect 20076 3528 20128 3534
rect 20076 3470 20128 3476
rect 7012 3052 7064 3058
rect 7012 2994 7064 3000
rect 19800 3052 19852 3058
rect 19800 2994 19852 3000
rect 19984 3052 20036 3058
rect 19984 2994 20036 3000
rect 2950 2748 3258 2757
rect 2950 2746 2956 2748
rect 3012 2746 3036 2748
rect 3092 2746 3116 2748
rect 3172 2746 3196 2748
rect 3252 2746 3258 2748
rect 3012 2694 3014 2746
rect 3194 2694 3196 2746
rect 2950 2692 2956 2694
rect 3012 2692 3036 2694
rect 3092 2692 3116 2694
rect 3172 2692 3196 2694
rect 3252 2692 3258 2694
rect 2950 2683 3258 2692
rect 7024 2650 7052 2994
rect 19340 2984 19392 2990
rect 19340 2926 19392 2932
rect 12950 2748 13258 2757
rect 12950 2746 12956 2748
rect 13012 2746 13036 2748
rect 13092 2746 13116 2748
rect 13172 2746 13196 2748
rect 13252 2746 13258 2748
rect 13012 2694 13014 2746
rect 13194 2694 13196 2746
rect 12950 2692 12956 2694
rect 13012 2692 13036 2694
rect 13092 2692 13116 2694
rect 13172 2692 13196 2694
rect 13252 2692 13258 2694
rect 12950 2683 13258 2692
rect 19352 2650 19380 2926
rect 19812 2854 19840 2994
rect 19800 2848 19852 2854
rect 19800 2790 19852 2796
rect 7012 2644 7064 2650
rect 7012 2586 7064 2592
rect 19340 2644 19392 2650
rect 19340 2586 19392 2592
rect 19812 2582 19840 2790
rect 19800 2576 19852 2582
rect 19800 2518 19852 2524
rect 6736 2304 6788 2310
rect 6736 2246 6788 2252
rect 6748 800 6776 2246
rect 7950 2204 8258 2213
rect 7950 2202 7956 2204
rect 8012 2202 8036 2204
rect 8092 2202 8116 2204
rect 8172 2202 8196 2204
rect 8252 2202 8258 2204
rect 8012 2150 8014 2202
rect 8194 2150 8196 2202
rect 7950 2148 7956 2150
rect 8012 2148 8036 2150
rect 8092 2148 8116 2150
rect 8172 2148 8196 2150
rect 8252 2148 8258 2150
rect 7950 2139 8258 2148
rect 17950 2204 18258 2213
rect 17950 2202 17956 2204
rect 18012 2202 18036 2204
rect 18092 2202 18116 2204
rect 18172 2202 18196 2204
rect 18252 2202 18258 2204
rect 18012 2150 18014 2202
rect 18194 2150 18196 2202
rect 17950 2148 17956 2150
rect 18012 2148 18036 2150
rect 18092 2148 18116 2150
rect 18172 2148 18196 2150
rect 18252 2148 18258 2150
rect 17950 2139 18258 2148
rect 20180 800 20208 4014
rect 20640 2446 20668 9658
rect 20720 9376 20772 9382
rect 20720 9318 20772 9324
rect 20732 8906 20760 9318
rect 20720 8900 20772 8906
rect 20720 8842 20772 8848
rect 20720 7744 20772 7750
rect 20720 7686 20772 7692
rect 20732 7478 20760 7686
rect 20720 7472 20772 7478
rect 20720 7414 20772 7420
rect 20824 6798 20852 10406
rect 20916 8090 20944 11630
rect 21100 11626 21128 15982
rect 21180 15632 21232 15638
rect 21180 15574 21232 15580
rect 21088 11620 21140 11626
rect 21088 11562 21140 11568
rect 21088 11008 21140 11014
rect 21088 10950 21140 10956
rect 21100 10810 21128 10950
rect 20996 10804 21048 10810
rect 20996 10746 21048 10752
rect 21088 10804 21140 10810
rect 21088 10746 21140 10752
rect 20904 8084 20956 8090
rect 20904 8026 20956 8032
rect 21008 6798 21036 10746
rect 21192 8974 21220 15574
rect 21284 15366 21312 19450
rect 21376 19378 21404 19722
rect 21364 19372 21416 19378
rect 21364 19314 21416 19320
rect 21468 18358 21496 21490
rect 21560 21418 21588 21626
rect 21548 21412 21600 21418
rect 21548 21354 21600 21360
rect 21548 21004 21600 21010
rect 21548 20946 21600 20952
rect 21560 19768 21588 20946
rect 21652 20777 21680 22102
rect 21730 22063 21786 22072
rect 21638 20768 21694 20777
rect 21638 20703 21694 20712
rect 21640 19780 21692 19786
rect 21560 19740 21640 19768
rect 21640 19722 21692 19728
rect 21652 19310 21680 19722
rect 21640 19304 21692 19310
rect 21640 19246 21692 19252
rect 21546 19136 21602 19145
rect 21546 19071 21602 19080
rect 21456 18352 21508 18358
rect 21456 18294 21508 18300
rect 21364 16788 21416 16794
rect 21364 16730 21416 16736
rect 21376 15570 21404 16730
rect 21364 15564 21416 15570
rect 21364 15506 21416 15512
rect 21272 15360 21324 15366
rect 21272 15302 21324 15308
rect 21468 15162 21496 18294
rect 21560 16726 21588 19071
rect 21652 18698 21680 19246
rect 21640 18692 21692 18698
rect 21640 18634 21692 18640
rect 21640 18420 21692 18426
rect 21640 18362 21692 18368
rect 21652 18329 21680 18362
rect 21638 18320 21694 18329
rect 21638 18255 21694 18264
rect 21638 17776 21694 17785
rect 21638 17711 21694 17720
rect 21548 16720 21600 16726
rect 21652 16697 21680 17711
rect 21548 16662 21600 16668
rect 21638 16688 21694 16697
rect 21638 16623 21694 16632
rect 21744 16538 21772 22063
rect 21836 21350 21864 22170
rect 22204 22098 22232 22986
rect 22284 22704 22336 22710
rect 22284 22646 22336 22652
rect 22296 22234 22324 22646
rect 22388 22642 22416 22986
rect 22376 22636 22428 22642
rect 22376 22578 22428 22584
rect 22284 22228 22336 22234
rect 22284 22170 22336 22176
rect 22192 22092 22244 22098
rect 22480 22094 22508 23446
rect 22572 23322 22600 23598
rect 22560 23316 22612 23322
rect 22560 23258 22612 23264
rect 22560 22568 22612 22574
rect 22560 22510 22612 22516
rect 22192 22034 22244 22040
rect 22296 22066 22508 22094
rect 22204 21894 22232 22034
rect 22296 21978 22324 22066
rect 22296 21950 22416 21978
rect 22192 21888 22244 21894
rect 22192 21830 22244 21836
rect 22284 21888 22336 21894
rect 22284 21830 22336 21836
rect 22190 21720 22246 21729
rect 22100 21684 22152 21690
rect 21928 21644 22100 21672
rect 21824 21344 21876 21350
rect 21824 21286 21876 21292
rect 21928 20806 21956 21644
rect 22190 21655 22246 21664
rect 22100 21626 22152 21632
rect 22204 21554 22232 21655
rect 22192 21548 22244 21554
rect 22192 21490 22244 21496
rect 22190 21448 22246 21457
rect 22296 21418 22324 21830
rect 22190 21383 22246 21392
rect 22284 21412 22336 21418
rect 22006 21176 22062 21185
rect 22062 21134 22140 21162
rect 22006 21111 22062 21120
rect 22008 21004 22060 21010
rect 22008 20946 22060 20952
rect 21916 20800 21968 20806
rect 21916 20742 21968 20748
rect 21822 20496 21878 20505
rect 21822 20431 21878 20440
rect 21836 18970 21864 20431
rect 22020 19718 22048 20946
rect 22112 20806 22140 21134
rect 22100 20800 22152 20806
rect 22100 20742 22152 20748
rect 22008 19712 22060 19718
rect 22008 19654 22060 19660
rect 22100 19508 22152 19514
rect 22100 19450 22152 19456
rect 22112 19242 22140 19450
rect 22204 19281 22232 21383
rect 22284 21354 22336 21360
rect 22284 21072 22336 21078
rect 22284 21014 22336 21020
rect 22190 19272 22246 19281
rect 22100 19236 22152 19242
rect 22190 19207 22246 19216
rect 22100 19178 22152 19184
rect 21916 19168 21968 19174
rect 21916 19110 21968 19116
rect 21824 18964 21876 18970
rect 21824 18906 21876 18912
rect 21928 18601 21956 19110
rect 22192 18624 22244 18630
rect 21914 18592 21970 18601
rect 21914 18527 21970 18536
rect 22098 18592 22154 18601
rect 22192 18566 22244 18572
rect 22098 18527 22154 18536
rect 22112 18222 22140 18527
rect 21916 18216 21968 18222
rect 21916 18158 21968 18164
rect 22100 18216 22152 18222
rect 22100 18158 22152 18164
rect 21928 17649 21956 18158
rect 22204 17882 22232 18566
rect 22192 17876 22244 17882
rect 22192 17818 22244 17824
rect 21914 17640 21970 17649
rect 21914 17575 21970 17584
rect 21916 17536 21968 17542
rect 21916 17478 21968 17484
rect 21822 17096 21878 17105
rect 21822 17031 21878 17040
rect 21560 16510 21772 16538
rect 21456 15156 21508 15162
rect 21456 15098 21508 15104
rect 21272 14952 21324 14958
rect 21272 14894 21324 14900
rect 21284 13870 21312 14894
rect 21468 14414 21496 15098
rect 21456 14408 21508 14414
rect 21456 14350 21508 14356
rect 21272 13864 21324 13870
rect 21272 13806 21324 13812
rect 21284 13530 21312 13806
rect 21272 13524 21324 13530
rect 21272 13466 21324 13472
rect 21468 12986 21496 14350
rect 21456 12980 21508 12986
rect 21456 12922 21508 12928
rect 21560 12866 21588 16510
rect 21640 16244 21692 16250
rect 21640 16186 21692 16192
rect 21652 15434 21680 16186
rect 21640 15428 21692 15434
rect 21640 15370 21692 15376
rect 21638 15328 21694 15337
rect 21638 15263 21694 15272
rect 21284 12838 21588 12866
rect 21284 11558 21312 12838
rect 21548 12776 21600 12782
rect 21548 12718 21600 12724
rect 21560 12434 21588 12718
rect 21468 12406 21588 12434
rect 21652 12434 21680 15263
rect 21652 12406 21772 12434
rect 21364 12300 21416 12306
rect 21364 12242 21416 12248
rect 21272 11552 21324 11558
rect 21272 11494 21324 11500
rect 21272 11008 21324 11014
rect 21272 10950 21324 10956
rect 21284 10606 21312 10950
rect 21272 10600 21324 10606
rect 21272 10542 21324 10548
rect 21272 10464 21324 10470
rect 21272 10406 21324 10412
rect 21284 10130 21312 10406
rect 21376 10130 21404 12242
rect 21272 10124 21324 10130
rect 21272 10066 21324 10072
rect 21364 10124 21416 10130
rect 21364 10066 21416 10072
rect 21270 9752 21326 9761
rect 21468 9738 21496 12406
rect 21640 11620 21692 11626
rect 21640 11562 21692 11568
rect 21548 11552 21600 11558
rect 21548 11494 21600 11500
rect 21560 11218 21588 11494
rect 21548 11212 21600 11218
rect 21548 11154 21600 11160
rect 21548 10464 21600 10470
rect 21548 10406 21600 10412
rect 21560 9994 21588 10406
rect 21652 10130 21680 11562
rect 21744 11014 21772 12406
rect 21732 11008 21784 11014
rect 21732 10950 21784 10956
rect 21732 10260 21784 10266
rect 21732 10202 21784 10208
rect 21640 10124 21692 10130
rect 21640 10066 21692 10072
rect 21548 9988 21600 9994
rect 21548 9930 21600 9936
rect 21640 9988 21692 9994
rect 21640 9930 21692 9936
rect 21270 9687 21326 9696
rect 21376 9710 21496 9738
rect 21284 9586 21312 9687
rect 21272 9580 21324 9586
rect 21272 9522 21324 9528
rect 21376 9178 21404 9710
rect 21560 9602 21588 9930
rect 21468 9574 21588 9602
rect 21652 9586 21680 9930
rect 21640 9580 21692 9586
rect 21364 9172 21416 9178
rect 21364 9114 21416 9120
rect 21180 8968 21232 8974
rect 21180 8910 21232 8916
rect 21364 8832 21416 8838
rect 21364 8774 21416 8780
rect 21376 8566 21404 8774
rect 21364 8560 21416 8566
rect 21364 8502 21416 8508
rect 21468 8430 21496 9574
rect 21640 9522 21692 9528
rect 21548 8968 21600 8974
rect 21548 8910 21600 8916
rect 21456 8424 21508 8430
rect 21456 8366 21508 8372
rect 21270 7848 21326 7857
rect 21270 7783 21326 7792
rect 21284 7546 21312 7783
rect 21272 7540 21324 7546
rect 21272 7482 21324 7488
rect 20812 6792 20864 6798
rect 20812 6734 20864 6740
rect 20996 6792 21048 6798
rect 20996 6734 21048 6740
rect 21560 6662 21588 8910
rect 21640 8900 21692 8906
rect 21640 8842 21692 8848
rect 21652 6798 21680 8842
rect 21640 6792 21692 6798
rect 21640 6734 21692 6740
rect 21548 6656 21600 6662
rect 21548 6598 21600 6604
rect 21744 5710 21772 10202
rect 21836 7410 21864 17031
rect 21928 15484 21956 17478
rect 22008 17264 22060 17270
rect 22008 17206 22060 17212
rect 22020 16522 22048 17206
rect 22204 16522 22232 17818
rect 22008 16516 22060 16522
rect 22192 16516 22244 16522
rect 22060 16476 22140 16504
rect 22008 16458 22060 16464
rect 22008 15496 22060 15502
rect 21928 15456 22008 15484
rect 22008 15438 22060 15444
rect 22112 15162 22140 16476
rect 22192 16458 22244 16464
rect 22296 16250 22324 21014
rect 22388 20618 22416 21950
rect 22468 21480 22520 21486
rect 22468 21422 22520 21428
rect 22480 21049 22508 21422
rect 22466 21040 22522 21049
rect 22466 20975 22522 20984
rect 22388 20590 22508 20618
rect 22480 20534 22508 20590
rect 22468 20528 22520 20534
rect 22468 20470 22520 20476
rect 22480 19514 22508 20470
rect 22468 19508 22520 19514
rect 22468 19450 22520 19456
rect 22572 19394 22600 22510
rect 22664 22001 22692 26200
rect 22756 22166 22784 26302
rect 23018 26200 23074 26302
rect 23386 26200 23442 27000
rect 24490 26200 24546 27000
rect 24858 26200 24914 27000
rect 25226 26200 25282 27000
rect 25778 26480 25834 26489
rect 25778 26415 25834 26424
rect 22834 26072 22890 26081
rect 22834 26007 22890 26016
rect 22848 23882 22876 26007
rect 23202 25664 23258 25673
rect 23202 25599 23258 25608
rect 23216 24886 23244 25599
rect 23204 24880 23256 24886
rect 23204 24822 23256 24828
rect 22950 24508 23258 24517
rect 22950 24506 22956 24508
rect 23012 24506 23036 24508
rect 23092 24506 23116 24508
rect 23172 24506 23196 24508
rect 23252 24506 23258 24508
rect 23012 24454 23014 24506
rect 23194 24454 23196 24506
rect 22950 24452 22956 24454
rect 23012 24452 23036 24454
rect 23092 24452 23116 24454
rect 23172 24452 23196 24454
rect 23252 24452 23258 24454
rect 22950 24443 23258 24452
rect 22848 23854 22968 23882
rect 22940 23610 22968 23854
rect 23296 23860 23348 23866
rect 23296 23802 23348 23808
rect 22848 23582 22968 23610
rect 22744 22160 22796 22166
rect 22744 22102 22796 22108
rect 22848 22030 22876 23582
rect 22950 23420 23258 23429
rect 22950 23418 22956 23420
rect 23012 23418 23036 23420
rect 23092 23418 23116 23420
rect 23172 23418 23196 23420
rect 23252 23418 23258 23420
rect 23012 23366 23014 23418
rect 23194 23366 23196 23418
rect 22950 23364 22956 23366
rect 23012 23364 23036 23366
rect 23092 23364 23116 23366
rect 23172 23364 23196 23366
rect 23252 23364 23258 23366
rect 22950 23355 23258 23364
rect 23308 22574 23336 23802
rect 23296 22568 23348 22574
rect 23296 22510 23348 22516
rect 22950 22332 23258 22341
rect 22950 22330 22956 22332
rect 23012 22330 23036 22332
rect 23092 22330 23116 22332
rect 23172 22330 23196 22332
rect 23252 22330 23258 22332
rect 23012 22278 23014 22330
rect 23194 22278 23196 22330
rect 22950 22276 22956 22278
rect 23012 22276 23036 22278
rect 23092 22276 23116 22278
rect 23172 22276 23196 22278
rect 23252 22276 23258 22278
rect 22950 22267 23258 22276
rect 22836 22024 22888 22030
rect 22650 21992 22706 22001
rect 22836 21966 22888 21972
rect 23204 22024 23256 22030
rect 23204 21966 23256 21972
rect 22650 21927 22706 21936
rect 22650 21856 22706 21865
rect 22650 21791 22706 21800
rect 22664 21486 22692 21791
rect 23216 21486 23244 21966
rect 23308 21554 23336 22510
rect 23400 21593 23428 26200
rect 23848 24200 23900 24206
rect 23848 24142 23900 24148
rect 23572 24064 23624 24070
rect 23572 24006 23624 24012
rect 23584 23594 23612 24006
rect 23572 23588 23624 23594
rect 23572 23530 23624 23536
rect 23860 22778 23888 24142
rect 23940 24064 23992 24070
rect 24124 24064 24176 24070
rect 23992 24024 24072 24052
rect 23940 24006 23992 24012
rect 24044 23798 24072 24024
rect 24124 24006 24176 24012
rect 24032 23792 24084 23798
rect 24032 23734 24084 23740
rect 23940 22976 23992 22982
rect 23940 22918 23992 22924
rect 23848 22772 23900 22778
rect 23848 22714 23900 22720
rect 23664 22432 23716 22438
rect 23664 22374 23716 22380
rect 23480 22024 23532 22030
rect 23480 21966 23532 21972
rect 23492 21729 23520 21966
rect 23572 21888 23624 21894
rect 23572 21830 23624 21836
rect 23478 21720 23534 21729
rect 23478 21655 23534 21664
rect 23386 21584 23442 21593
rect 23296 21548 23348 21554
rect 23386 21519 23442 21528
rect 23296 21490 23348 21496
rect 22652 21480 22704 21486
rect 22652 21422 22704 21428
rect 22744 21480 22796 21486
rect 22744 21422 22796 21428
rect 23204 21480 23256 21486
rect 23204 21422 23256 21428
rect 22650 21312 22706 21321
rect 22650 21247 22706 21256
rect 22664 21078 22692 21247
rect 22652 21072 22704 21078
rect 22652 21014 22704 21020
rect 22652 20392 22704 20398
rect 22652 20334 22704 20340
rect 22388 19366 22600 19394
rect 22388 18850 22416 19366
rect 22560 19304 22612 19310
rect 22560 19246 22612 19252
rect 22572 19145 22600 19246
rect 22558 19136 22614 19145
rect 22558 19071 22614 19080
rect 22388 18822 22508 18850
rect 22376 18760 22428 18766
rect 22376 18702 22428 18708
rect 22284 16244 22336 16250
rect 22284 16186 22336 16192
rect 22284 16108 22336 16114
rect 22284 16050 22336 16056
rect 22192 15904 22244 15910
rect 22192 15846 22244 15852
rect 22100 15156 22152 15162
rect 22100 15098 22152 15104
rect 22100 14612 22152 14618
rect 21928 14572 22100 14600
rect 21928 13394 21956 14572
rect 22100 14554 22152 14560
rect 22098 13968 22154 13977
rect 22098 13903 22154 13912
rect 22112 13512 22140 13903
rect 22020 13484 22140 13512
rect 21916 13388 21968 13394
rect 21916 13330 21968 13336
rect 21928 12850 21956 13330
rect 22020 12866 22048 13484
rect 22204 13410 22232 15846
rect 22296 15201 22324 16050
rect 22282 15192 22338 15201
rect 22282 15127 22338 15136
rect 22296 14113 22324 15127
rect 22282 14104 22338 14113
rect 22282 14039 22338 14048
rect 22284 13864 22336 13870
rect 22282 13832 22284 13841
rect 22336 13832 22338 13841
rect 22282 13767 22338 13776
rect 22388 13682 22416 18702
rect 22480 18698 22508 18822
rect 22468 18692 22520 18698
rect 22468 18634 22520 18640
rect 22560 18624 22612 18630
rect 22560 18566 22612 18572
rect 22572 18290 22600 18566
rect 22560 18284 22612 18290
rect 22560 18226 22612 18232
rect 22468 18216 22520 18222
rect 22466 18184 22468 18193
rect 22520 18184 22522 18193
rect 22466 18119 22522 18128
rect 22560 18080 22612 18086
rect 22560 18022 22612 18028
rect 22572 17814 22600 18022
rect 22664 17882 22692 20334
rect 22756 18737 22784 21422
rect 22836 21344 22888 21350
rect 22836 21286 22888 21292
rect 22848 21010 22876 21286
rect 22950 21244 23258 21253
rect 22950 21242 22956 21244
rect 23012 21242 23036 21244
rect 23092 21242 23116 21244
rect 23172 21242 23196 21244
rect 23252 21242 23258 21244
rect 23012 21190 23014 21242
rect 23194 21190 23196 21242
rect 22950 21188 22956 21190
rect 23012 21188 23036 21190
rect 23092 21188 23116 21190
rect 23172 21188 23196 21190
rect 23252 21188 23258 21190
rect 22950 21179 23258 21188
rect 22836 21004 22888 21010
rect 22836 20946 22888 20952
rect 23204 20936 23256 20942
rect 23202 20904 23204 20913
rect 23256 20904 23258 20913
rect 23202 20839 23258 20848
rect 23308 20466 23336 21490
rect 23386 21176 23442 21185
rect 23386 21111 23442 21120
rect 23296 20460 23348 20466
rect 23296 20402 23348 20408
rect 22836 20256 22888 20262
rect 22836 20198 22888 20204
rect 22742 18728 22798 18737
rect 22742 18663 22744 18672
rect 22796 18663 22798 18672
rect 22744 18634 22796 18640
rect 22652 17876 22704 17882
rect 22652 17818 22704 17824
rect 22560 17808 22612 17814
rect 22560 17750 22612 17756
rect 22468 17604 22520 17610
rect 22468 17546 22520 17552
rect 22480 17270 22508 17546
rect 22468 17264 22520 17270
rect 22468 17206 22520 17212
rect 22572 17202 22600 17750
rect 22560 17196 22612 17202
rect 22560 17138 22612 17144
rect 22664 17082 22692 17818
rect 22744 17672 22796 17678
rect 22744 17614 22796 17620
rect 22468 17060 22520 17066
rect 22468 17002 22520 17008
rect 22572 17054 22692 17082
rect 22480 16697 22508 17002
rect 22572 16794 22600 17054
rect 22560 16788 22612 16794
rect 22560 16730 22612 16736
rect 22466 16688 22522 16697
rect 22466 16623 22522 16632
rect 22560 16652 22612 16658
rect 22560 16594 22612 16600
rect 22572 14958 22600 16594
rect 22652 16516 22704 16522
rect 22652 16458 22704 16464
rect 22664 16046 22692 16458
rect 22652 16040 22704 16046
rect 22652 15982 22704 15988
rect 22756 15552 22784 17614
rect 22848 16046 22876 20198
rect 22950 20156 23258 20165
rect 22950 20154 22956 20156
rect 23012 20154 23036 20156
rect 23092 20154 23116 20156
rect 23172 20154 23196 20156
rect 23252 20154 23258 20156
rect 23012 20102 23014 20154
rect 23194 20102 23196 20154
rect 22950 20100 22956 20102
rect 23012 20100 23036 20102
rect 23092 20100 23116 20102
rect 23172 20100 23196 20102
rect 23252 20100 23258 20102
rect 22950 20091 23258 20100
rect 23018 19952 23074 19961
rect 23308 19922 23336 20402
rect 23400 20210 23428 21111
rect 23400 20182 23520 20210
rect 23388 20052 23440 20058
rect 23388 19994 23440 20000
rect 23018 19887 23074 19896
rect 23296 19916 23348 19922
rect 23032 19446 23060 19887
rect 23296 19858 23348 19864
rect 23020 19440 23072 19446
rect 23020 19382 23072 19388
rect 23308 19378 23336 19858
rect 23400 19553 23428 19994
rect 23386 19544 23442 19553
rect 23386 19479 23442 19488
rect 23492 19394 23520 20182
rect 23584 20074 23612 21830
rect 23676 21622 23704 22374
rect 23848 21956 23900 21962
rect 23848 21898 23900 21904
rect 23756 21888 23808 21894
rect 23756 21830 23808 21836
rect 23664 21616 23716 21622
rect 23664 21558 23716 21564
rect 23664 21072 23716 21078
rect 23664 21014 23716 21020
rect 23676 20534 23704 21014
rect 23664 20528 23716 20534
rect 23664 20470 23716 20476
rect 23584 20046 23704 20074
rect 23572 19712 23624 19718
rect 23572 19654 23624 19660
rect 23296 19372 23348 19378
rect 23296 19314 23348 19320
rect 23400 19366 23520 19394
rect 22950 19068 23258 19077
rect 22950 19066 22956 19068
rect 23012 19066 23036 19068
rect 23092 19066 23116 19068
rect 23172 19066 23196 19068
rect 23252 19066 23258 19068
rect 23012 19014 23014 19066
rect 23194 19014 23196 19066
rect 22950 19012 22956 19014
rect 23012 19012 23036 19014
rect 23092 19012 23116 19014
rect 23172 19012 23196 19014
rect 23252 19012 23258 19014
rect 22950 19003 23258 19012
rect 22928 18828 22980 18834
rect 22928 18770 22980 18776
rect 22940 18329 22968 18770
rect 23018 18728 23074 18737
rect 23018 18663 23074 18672
rect 23032 18426 23060 18663
rect 23204 18624 23256 18630
rect 23204 18566 23256 18572
rect 23020 18420 23072 18426
rect 23020 18362 23072 18368
rect 23112 18420 23164 18426
rect 23112 18362 23164 18368
rect 22926 18320 22982 18329
rect 22926 18255 22982 18264
rect 23124 18086 23152 18362
rect 23112 18080 23164 18086
rect 23216 18068 23244 18566
rect 23308 18426 23336 19314
rect 23400 18465 23428 19366
rect 23480 18760 23532 18766
rect 23480 18702 23532 18708
rect 23386 18456 23442 18465
rect 23296 18420 23348 18426
rect 23386 18391 23442 18400
rect 23296 18362 23348 18368
rect 23492 18193 23520 18702
rect 23478 18184 23534 18193
rect 23478 18119 23534 18128
rect 23216 18040 23336 18068
rect 23112 18022 23164 18028
rect 22950 17980 23258 17989
rect 22950 17978 22956 17980
rect 23012 17978 23036 17980
rect 23092 17978 23116 17980
rect 23172 17978 23196 17980
rect 23252 17978 23258 17980
rect 23012 17926 23014 17978
rect 23194 17926 23196 17978
rect 22950 17924 22956 17926
rect 23012 17924 23036 17926
rect 23092 17924 23116 17926
rect 23172 17924 23196 17926
rect 23252 17924 23258 17926
rect 22950 17915 23258 17924
rect 23308 17814 23336 18040
rect 23296 17808 23348 17814
rect 23296 17750 23348 17756
rect 23388 17536 23440 17542
rect 23388 17478 23440 17484
rect 22950 16892 23258 16901
rect 22950 16890 22956 16892
rect 23012 16890 23036 16892
rect 23092 16890 23116 16892
rect 23172 16890 23196 16892
rect 23252 16890 23258 16892
rect 23012 16838 23014 16890
rect 23194 16838 23196 16890
rect 22950 16836 22956 16838
rect 23012 16836 23036 16838
rect 23092 16836 23116 16838
rect 23172 16836 23196 16838
rect 23252 16836 23258 16838
rect 22950 16827 23258 16836
rect 22836 16040 22888 16046
rect 22836 15982 22888 15988
rect 23296 15904 23348 15910
rect 23296 15846 23348 15852
rect 22950 15804 23258 15813
rect 22950 15802 22956 15804
rect 23012 15802 23036 15804
rect 23092 15802 23116 15804
rect 23172 15802 23196 15804
rect 23252 15802 23258 15804
rect 23012 15750 23014 15802
rect 23194 15750 23196 15802
rect 22950 15748 22956 15750
rect 23012 15748 23036 15750
rect 23092 15748 23116 15750
rect 23172 15748 23196 15750
rect 23252 15748 23258 15750
rect 22950 15739 23258 15748
rect 22756 15524 22876 15552
rect 22652 15496 22704 15502
rect 22704 15456 22784 15484
rect 22652 15438 22704 15444
rect 22652 15360 22704 15366
rect 22652 15302 22704 15308
rect 22560 14952 22612 14958
rect 22560 14894 22612 14900
rect 22468 14884 22520 14890
rect 22468 14826 22520 14832
rect 22112 13382 22232 13410
rect 22296 13654 22416 13682
rect 22112 12968 22140 13382
rect 22112 12940 22232 12968
rect 21916 12844 21968 12850
rect 22020 12838 22140 12866
rect 21916 12786 21968 12792
rect 21928 12306 21956 12786
rect 21916 12300 21968 12306
rect 21916 12242 21968 12248
rect 21916 10804 21968 10810
rect 21916 10746 21968 10752
rect 21928 9994 21956 10746
rect 22112 10470 22140 12838
rect 22204 12434 22232 12940
rect 22296 12782 22324 13654
rect 22374 13424 22430 13433
rect 22374 13359 22430 13368
rect 22388 12918 22416 13359
rect 22376 12912 22428 12918
rect 22376 12854 22428 12860
rect 22284 12776 22336 12782
rect 22336 12724 22416 12730
rect 22284 12718 22416 12724
rect 22296 12702 22416 12718
rect 22204 12406 22324 12434
rect 22192 11756 22244 11762
rect 22192 11698 22244 11704
rect 22100 10464 22152 10470
rect 22100 10406 22152 10412
rect 21916 9988 21968 9994
rect 21916 9930 21968 9936
rect 22008 9172 22060 9178
rect 22008 9114 22060 9120
rect 21916 8900 21968 8906
rect 21916 8842 21968 8848
rect 21928 8090 21956 8842
rect 22020 8838 22048 9114
rect 22100 9104 22152 9110
rect 22100 9046 22152 9052
rect 22008 8832 22060 8838
rect 22008 8774 22060 8780
rect 22112 8514 22140 9046
rect 22204 8634 22232 11698
rect 22296 11150 22324 12406
rect 22388 12102 22416 12702
rect 22376 12096 22428 12102
rect 22376 12038 22428 12044
rect 22376 11280 22428 11286
rect 22376 11222 22428 11228
rect 22284 11144 22336 11150
rect 22284 11086 22336 11092
rect 22284 8832 22336 8838
rect 22284 8774 22336 8780
rect 22192 8628 22244 8634
rect 22192 8570 22244 8576
rect 22020 8498 22140 8514
rect 22008 8492 22140 8498
rect 22060 8486 22140 8492
rect 22008 8434 22060 8440
rect 22006 8392 22062 8401
rect 22006 8327 22062 8336
rect 21916 8084 21968 8090
rect 21916 8026 21968 8032
rect 22020 7886 22048 8327
rect 22008 7880 22060 7886
rect 22008 7822 22060 7828
rect 21824 7404 21876 7410
rect 21824 7346 21876 7352
rect 21836 6458 21864 7346
rect 22190 6896 22246 6905
rect 22190 6831 22246 6840
rect 22204 6798 22232 6831
rect 22192 6792 22244 6798
rect 22192 6734 22244 6740
rect 21824 6452 21876 6458
rect 21824 6394 21876 6400
rect 22296 6322 22324 8774
rect 22284 6316 22336 6322
rect 22284 6258 22336 6264
rect 22388 5710 22416 11222
rect 21732 5704 21784 5710
rect 21732 5646 21784 5652
rect 22376 5704 22428 5710
rect 22376 5646 22428 5652
rect 22388 4826 22416 5646
rect 22480 5234 22508 14826
rect 22572 14618 22600 14894
rect 22560 14612 22612 14618
rect 22560 14554 22612 14560
rect 22572 14346 22600 14554
rect 22560 14340 22612 14346
rect 22560 14282 22612 14288
rect 22572 13938 22600 14282
rect 22560 13932 22612 13938
rect 22560 13874 22612 13880
rect 22664 13818 22692 15302
rect 22756 14890 22784 15456
rect 22744 14884 22796 14890
rect 22744 14826 22796 14832
rect 22848 14346 22876 15524
rect 23204 15428 23256 15434
rect 23204 15370 23256 15376
rect 23216 15201 23244 15370
rect 23202 15192 23258 15201
rect 23202 15127 23258 15136
rect 22950 14716 23258 14725
rect 22950 14714 22956 14716
rect 23012 14714 23036 14716
rect 23092 14714 23116 14716
rect 23172 14714 23196 14716
rect 23252 14714 23258 14716
rect 23012 14662 23014 14714
rect 23194 14662 23196 14714
rect 22950 14660 22956 14662
rect 23012 14660 23036 14662
rect 23092 14660 23116 14662
rect 23172 14660 23196 14662
rect 23252 14660 23258 14662
rect 22950 14651 23258 14660
rect 22836 14340 22888 14346
rect 22836 14282 22888 14288
rect 22834 14240 22890 14249
rect 22834 14175 22890 14184
rect 22744 14068 22796 14074
rect 22744 14010 22796 14016
rect 22572 13790 22692 13818
rect 22572 6914 22600 13790
rect 22652 13388 22704 13394
rect 22652 13330 22704 13336
rect 22664 11286 22692 13330
rect 22756 12442 22784 14010
rect 22848 13394 22876 14175
rect 22950 13628 23258 13637
rect 22950 13626 22956 13628
rect 23012 13626 23036 13628
rect 23092 13626 23116 13628
rect 23172 13626 23196 13628
rect 23252 13626 23258 13628
rect 23012 13574 23014 13626
rect 23194 13574 23196 13626
rect 22950 13572 22956 13574
rect 23012 13572 23036 13574
rect 23092 13572 23116 13574
rect 23172 13572 23196 13574
rect 23252 13572 23258 13574
rect 22950 13563 23258 13572
rect 23204 13524 23256 13530
rect 23204 13466 23256 13472
rect 23216 13394 23244 13466
rect 22836 13388 22888 13394
rect 22836 13330 22888 13336
rect 23204 13388 23256 13394
rect 23204 13330 23256 13336
rect 22834 13016 22890 13025
rect 23216 12986 23244 13330
rect 22834 12951 22890 12960
rect 23204 12980 23256 12986
rect 22744 12436 22796 12442
rect 22744 12378 22796 12384
rect 22652 11280 22704 11286
rect 22652 11222 22704 11228
rect 22652 11144 22704 11150
rect 22652 11086 22704 11092
rect 22664 9518 22692 11086
rect 22652 9512 22704 9518
rect 22652 9454 22704 9460
rect 22848 9110 22876 12951
rect 23204 12922 23256 12928
rect 22950 12540 23258 12549
rect 22950 12538 22956 12540
rect 23012 12538 23036 12540
rect 23092 12538 23116 12540
rect 23172 12538 23196 12540
rect 23252 12538 23258 12540
rect 23012 12486 23014 12538
rect 23194 12486 23196 12538
rect 22950 12484 22956 12486
rect 23012 12484 23036 12486
rect 23092 12484 23116 12486
rect 23172 12484 23196 12486
rect 23252 12484 23258 12486
rect 22950 12475 23258 12484
rect 22950 11452 23258 11461
rect 22950 11450 22956 11452
rect 23012 11450 23036 11452
rect 23092 11450 23116 11452
rect 23172 11450 23196 11452
rect 23252 11450 23258 11452
rect 23012 11398 23014 11450
rect 23194 11398 23196 11450
rect 22950 11396 22956 11398
rect 23012 11396 23036 11398
rect 23092 11396 23116 11398
rect 23172 11396 23196 11398
rect 23252 11396 23258 11398
rect 22950 11387 23258 11396
rect 23308 10606 23336 15846
rect 23400 14929 23428 17478
rect 23480 17128 23532 17134
rect 23480 17070 23532 17076
rect 23386 14920 23442 14929
rect 23386 14855 23442 14864
rect 23386 14648 23442 14657
rect 23386 14583 23442 14592
rect 23400 14482 23428 14583
rect 23388 14476 23440 14482
rect 23388 14418 23440 14424
rect 23492 14362 23520 17070
rect 23584 14482 23612 19654
rect 23572 14476 23624 14482
rect 23572 14418 23624 14424
rect 23676 14414 23704 20046
rect 23768 17746 23796 21830
rect 23860 21350 23888 21898
rect 23848 21344 23900 21350
rect 23848 21286 23900 21292
rect 23860 20534 23888 21286
rect 23848 20528 23900 20534
rect 23848 20470 23900 20476
rect 23952 20262 23980 22918
rect 24044 22710 24072 23734
rect 24136 23526 24164 24006
rect 24308 23656 24360 23662
rect 24308 23598 24360 23604
rect 24124 23520 24176 23526
rect 24124 23462 24176 23468
rect 24032 22704 24084 22710
rect 24032 22646 24084 22652
rect 24044 22094 24072 22646
rect 24136 22574 24164 23462
rect 24124 22568 24176 22574
rect 24124 22510 24176 22516
rect 24044 22066 24164 22094
rect 24032 21956 24084 21962
rect 24032 21898 24084 21904
rect 24044 21729 24072 21898
rect 24030 21720 24086 21729
rect 24030 21655 24086 21664
rect 23940 20256 23992 20262
rect 23940 20198 23992 20204
rect 23940 20052 23992 20058
rect 23940 19994 23992 20000
rect 23952 19514 23980 19994
rect 24044 19854 24072 21655
rect 24136 21622 24164 22066
rect 24124 21616 24176 21622
rect 24124 21558 24176 21564
rect 24136 21078 24164 21558
rect 24124 21072 24176 21078
rect 24124 21014 24176 21020
rect 24136 20618 24164 21014
rect 24136 20590 24256 20618
rect 24228 20534 24256 20590
rect 24216 20528 24268 20534
rect 24216 20470 24268 20476
rect 24124 20392 24176 20398
rect 24124 20334 24176 20340
rect 24032 19848 24084 19854
rect 24032 19790 24084 19796
rect 23848 19508 23900 19514
rect 23848 19450 23900 19456
rect 23940 19508 23992 19514
rect 23940 19450 23992 19456
rect 23860 17746 23888 19450
rect 23952 19394 23980 19450
rect 23952 19366 24072 19394
rect 23938 19272 23994 19281
rect 23938 19207 23994 19216
rect 23952 18698 23980 19207
rect 24044 19174 24072 19366
rect 24032 19168 24084 19174
rect 24032 19110 24084 19116
rect 23940 18692 23992 18698
rect 23940 18634 23992 18640
rect 23952 18222 23980 18634
rect 23940 18216 23992 18222
rect 23940 18158 23992 18164
rect 23756 17740 23808 17746
rect 23756 17682 23808 17688
rect 23848 17740 23900 17746
rect 23848 17682 23900 17688
rect 23860 17626 23888 17682
rect 23756 17604 23808 17610
rect 23860 17598 23980 17626
rect 23756 17546 23808 17552
rect 23768 16658 23796 17546
rect 23848 17536 23900 17542
rect 23848 17478 23900 17484
rect 23756 16652 23808 16658
rect 23756 16594 23808 16600
rect 23768 15094 23796 16594
rect 23860 16454 23888 17478
rect 23952 17066 23980 17598
rect 23940 17060 23992 17066
rect 23940 17002 23992 17008
rect 23848 16448 23900 16454
rect 23848 16390 23900 16396
rect 23940 16448 23992 16454
rect 23940 16390 23992 16396
rect 23848 16176 23900 16182
rect 23848 16118 23900 16124
rect 23756 15088 23808 15094
rect 23756 15030 23808 15036
rect 23768 14618 23796 15030
rect 23756 14612 23808 14618
rect 23756 14554 23808 14560
rect 23664 14408 23716 14414
rect 23492 14334 23612 14362
rect 23664 14350 23716 14356
rect 23388 14000 23440 14006
rect 23440 13948 23520 13954
rect 23388 13942 23520 13948
rect 23400 13926 23520 13942
rect 23492 13530 23520 13926
rect 23480 13524 23532 13530
rect 23480 13466 23532 13472
rect 23480 12708 23532 12714
rect 23480 12650 23532 12656
rect 23388 11348 23440 11354
rect 23388 11290 23440 11296
rect 23296 10600 23348 10606
rect 23296 10542 23348 10548
rect 22950 10364 23258 10373
rect 22950 10362 22956 10364
rect 23012 10362 23036 10364
rect 23092 10362 23116 10364
rect 23172 10362 23196 10364
rect 23252 10362 23258 10364
rect 23012 10310 23014 10362
rect 23194 10310 23196 10362
rect 22950 10308 22956 10310
rect 23012 10308 23036 10310
rect 23092 10308 23116 10310
rect 23172 10308 23196 10310
rect 23252 10308 23258 10310
rect 22950 10299 23258 10308
rect 23112 10056 23164 10062
rect 23112 9998 23164 10004
rect 23124 9926 23152 9998
rect 23112 9920 23164 9926
rect 23112 9862 23164 9868
rect 23124 9722 23152 9862
rect 23294 9752 23350 9761
rect 23112 9716 23164 9722
rect 23294 9687 23350 9696
rect 23112 9658 23164 9664
rect 23308 9654 23336 9687
rect 23296 9648 23348 9654
rect 23296 9590 23348 9596
rect 22950 9276 23258 9285
rect 22950 9274 22956 9276
rect 23012 9274 23036 9276
rect 23092 9274 23116 9276
rect 23172 9274 23196 9276
rect 23252 9274 23258 9276
rect 23012 9222 23014 9274
rect 23194 9222 23196 9274
rect 22950 9220 22956 9222
rect 23012 9220 23036 9222
rect 23092 9220 23116 9222
rect 23172 9220 23196 9222
rect 23252 9220 23258 9222
rect 22950 9211 23258 9220
rect 22836 9104 22888 9110
rect 22836 9046 22888 9052
rect 22744 9036 22796 9042
rect 22744 8978 22796 8984
rect 22572 6886 22692 6914
rect 22468 5228 22520 5234
rect 22468 5170 22520 5176
rect 22376 4820 22428 4826
rect 22376 4762 22428 4768
rect 22664 4622 22692 6886
rect 22756 5234 22784 8978
rect 22950 8188 23258 8197
rect 22950 8186 22956 8188
rect 23012 8186 23036 8188
rect 23092 8186 23116 8188
rect 23172 8186 23196 8188
rect 23252 8186 23258 8188
rect 23012 8134 23014 8186
rect 23194 8134 23196 8186
rect 22950 8132 22956 8134
rect 23012 8132 23036 8134
rect 23092 8132 23116 8134
rect 23172 8132 23196 8134
rect 23252 8132 23258 8134
rect 22950 8123 23258 8132
rect 23400 7886 23428 11290
rect 23492 7954 23520 12650
rect 23480 7948 23532 7954
rect 23480 7890 23532 7896
rect 23388 7880 23440 7886
rect 23388 7822 23440 7828
rect 23480 7744 23532 7750
rect 23480 7686 23532 7692
rect 23388 7200 23440 7206
rect 23388 7142 23440 7148
rect 22950 7100 23258 7109
rect 22950 7098 22956 7100
rect 23012 7098 23036 7100
rect 23092 7098 23116 7100
rect 23172 7098 23196 7100
rect 23252 7098 23258 7100
rect 23012 7046 23014 7098
rect 23194 7046 23196 7098
rect 22950 7044 22956 7046
rect 23012 7044 23036 7046
rect 23092 7044 23116 7046
rect 23172 7044 23196 7046
rect 23252 7044 23258 7046
rect 22950 7035 23258 7044
rect 22950 6012 23258 6021
rect 22950 6010 22956 6012
rect 23012 6010 23036 6012
rect 23092 6010 23116 6012
rect 23172 6010 23196 6012
rect 23252 6010 23258 6012
rect 23012 5958 23014 6010
rect 23194 5958 23196 6010
rect 22950 5956 22956 5958
rect 23012 5956 23036 5958
rect 23092 5956 23116 5958
rect 23172 5956 23196 5958
rect 23252 5956 23258 5958
rect 22950 5947 23258 5956
rect 22744 5228 22796 5234
rect 22744 5170 22796 5176
rect 22950 4924 23258 4933
rect 22950 4922 22956 4924
rect 23012 4922 23036 4924
rect 23092 4922 23116 4924
rect 23172 4922 23196 4924
rect 23252 4922 23258 4924
rect 23012 4870 23014 4922
rect 23194 4870 23196 4922
rect 22950 4868 22956 4870
rect 23012 4868 23036 4870
rect 23092 4868 23116 4870
rect 23172 4868 23196 4870
rect 23252 4868 23258 4870
rect 22950 4859 23258 4868
rect 23400 4622 23428 7142
rect 23492 5710 23520 7686
rect 23584 6914 23612 14334
rect 23664 14272 23716 14278
rect 23664 14214 23716 14220
rect 23676 10130 23704 14214
rect 23768 14006 23796 14554
rect 23756 14000 23808 14006
rect 23756 13942 23808 13948
rect 23768 13462 23796 13942
rect 23756 13456 23808 13462
rect 23756 13398 23808 13404
rect 23768 13258 23796 13398
rect 23756 13252 23808 13258
rect 23756 13194 23808 13200
rect 23768 12850 23796 13194
rect 23756 12844 23808 12850
rect 23756 12786 23808 12792
rect 23664 10124 23716 10130
rect 23664 10066 23716 10072
rect 23860 9178 23888 16118
rect 23952 16046 23980 16390
rect 24136 16114 24164 20334
rect 24228 20058 24256 20470
rect 24216 20052 24268 20058
rect 24216 19994 24268 20000
rect 24214 19816 24270 19825
rect 24320 19786 24348 23598
rect 24398 21584 24454 21593
rect 24398 21519 24454 21528
rect 24412 21049 24440 21519
rect 24398 21040 24454 21049
rect 24398 20975 24454 20984
rect 24504 20074 24532 26200
rect 25134 25256 25190 25265
rect 25134 25191 25190 25200
rect 25596 25220 25648 25226
rect 25148 24818 25176 25191
rect 25596 25162 25648 25168
rect 25136 24812 25188 24818
rect 25136 24754 25188 24760
rect 25042 24304 25098 24313
rect 25042 24239 25044 24248
rect 25096 24239 25098 24248
rect 25044 24210 25096 24216
rect 25044 24132 25096 24138
rect 25044 24074 25096 24080
rect 24768 23180 24820 23186
rect 24768 23122 24820 23128
rect 24584 22976 24636 22982
rect 24584 22918 24636 22924
rect 24596 22545 24624 22918
rect 24582 22536 24638 22545
rect 24582 22471 24638 22480
rect 24780 22438 24808 23122
rect 24952 22976 25004 22982
rect 24952 22918 25004 22924
rect 24768 22432 24820 22438
rect 24768 22374 24820 22380
rect 24860 22092 24912 22098
rect 24860 22034 24912 22040
rect 24676 21684 24728 21690
rect 24872 21672 24900 22034
rect 24728 21644 24900 21672
rect 24676 21626 24728 21632
rect 24860 21412 24912 21418
rect 24860 21354 24912 21360
rect 24872 20618 24900 21354
rect 24780 20590 24900 20618
rect 24780 20398 24808 20590
rect 24768 20392 24820 20398
rect 24768 20334 24820 20340
rect 24412 20046 24532 20074
rect 24214 19751 24270 19760
rect 24308 19780 24360 19786
rect 24228 16130 24256 19751
rect 24308 19722 24360 19728
rect 24320 18601 24348 19722
rect 24306 18592 24362 18601
rect 24306 18527 24362 18536
rect 24412 16590 24440 20046
rect 24492 19916 24544 19922
rect 24492 19858 24544 19864
rect 24400 16584 24452 16590
rect 24400 16526 24452 16532
rect 24412 16250 24440 16526
rect 24400 16244 24452 16250
rect 24400 16186 24452 16192
rect 24124 16108 24176 16114
rect 24228 16102 24440 16130
rect 24124 16050 24176 16056
rect 23940 16040 23992 16046
rect 23940 15982 23992 15988
rect 23952 15162 23980 15982
rect 23940 15156 23992 15162
rect 23940 15098 23992 15104
rect 24308 14272 24360 14278
rect 24308 14214 24360 14220
rect 24032 13252 24084 13258
rect 24032 13194 24084 13200
rect 23940 11076 23992 11082
rect 23940 11018 23992 11024
rect 23952 10674 23980 11018
rect 23940 10668 23992 10674
rect 23940 10610 23992 10616
rect 23940 10532 23992 10538
rect 23940 10474 23992 10480
rect 23952 9586 23980 10474
rect 23940 9580 23992 9586
rect 23940 9522 23992 9528
rect 23848 9172 23900 9178
rect 23848 9114 23900 9120
rect 24044 8022 24072 13194
rect 24216 12844 24268 12850
rect 24216 12786 24268 12792
rect 24228 12374 24256 12786
rect 24216 12368 24268 12374
rect 24216 12310 24268 12316
rect 24228 12170 24256 12310
rect 24216 12164 24268 12170
rect 24216 12106 24268 12112
rect 24032 8016 24084 8022
rect 24032 7958 24084 7964
rect 24320 6914 24348 14214
rect 24412 12850 24440 16102
rect 24504 15162 24532 19858
rect 24584 19712 24636 19718
rect 24582 19680 24584 19689
rect 24860 19712 24912 19718
rect 24636 19680 24638 19689
rect 24860 19654 24912 19660
rect 24582 19615 24638 19624
rect 24872 19417 24900 19654
rect 24858 19408 24914 19417
rect 24858 19343 24914 19352
rect 24676 19168 24728 19174
rect 24676 19110 24728 19116
rect 24584 18624 24636 18630
rect 24584 18566 24636 18572
rect 24596 18057 24624 18566
rect 24688 18426 24716 19110
rect 24860 18896 24912 18902
rect 24860 18838 24912 18844
rect 24872 18426 24900 18838
rect 24676 18420 24728 18426
rect 24676 18362 24728 18368
rect 24860 18420 24912 18426
rect 24860 18362 24912 18368
rect 24582 18048 24638 18057
rect 24582 17983 24638 17992
rect 24688 17610 24716 18362
rect 24964 17882 24992 22918
rect 25056 19922 25084 24074
rect 25148 23798 25176 24754
rect 25136 23792 25188 23798
rect 25136 23734 25188 23740
rect 25412 23588 25464 23594
rect 25412 23530 25464 23536
rect 25136 23520 25188 23526
rect 25136 23462 25188 23468
rect 25148 22098 25176 23462
rect 25320 22160 25372 22166
rect 25320 22102 25372 22108
rect 25136 22092 25188 22098
rect 25136 22034 25188 22040
rect 25332 21978 25360 22102
rect 25148 21950 25360 21978
rect 25148 21570 25176 21950
rect 25148 21542 25268 21570
rect 25136 21004 25188 21010
rect 25136 20946 25188 20952
rect 25148 20602 25176 20946
rect 25136 20596 25188 20602
rect 25136 20538 25188 20544
rect 25240 20482 25268 21542
rect 25148 20454 25268 20482
rect 25044 19916 25096 19922
rect 25044 19858 25096 19864
rect 25148 19802 25176 20454
rect 25228 20256 25280 20262
rect 25228 20198 25280 20204
rect 25056 19774 25176 19802
rect 25056 19514 25084 19774
rect 25044 19508 25096 19514
rect 25044 19450 25096 19456
rect 24952 17876 25004 17882
rect 24952 17818 25004 17824
rect 24676 17604 24728 17610
rect 24676 17546 24728 17552
rect 24688 17270 24716 17546
rect 24768 17332 24820 17338
rect 24768 17274 24820 17280
rect 24676 17264 24728 17270
rect 24676 17206 24728 17212
rect 24780 16590 24808 17274
rect 24858 17232 24914 17241
rect 24858 17167 24860 17176
rect 24912 17167 24914 17176
rect 24860 17138 24912 17144
rect 25056 16998 25084 19450
rect 25240 19310 25268 20198
rect 25228 19304 25280 19310
rect 25228 19246 25280 19252
rect 25240 18834 25268 19246
rect 25228 18828 25280 18834
rect 25228 18770 25280 18776
rect 25320 18284 25372 18290
rect 25320 18226 25372 18232
rect 25044 16992 25096 16998
rect 25044 16934 25096 16940
rect 24768 16584 24820 16590
rect 24768 16526 24820 16532
rect 24858 16280 24914 16289
rect 24858 16215 24914 16224
rect 24674 16144 24730 16153
rect 24674 16079 24676 16088
rect 24728 16079 24730 16088
rect 24676 16050 24728 16056
rect 24674 15872 24730 15881
rect 24674 15807 24730 15816
rect 24492 15156 24544 15162
rect 24492 15098 24544 15104
rect 24504 13870 24532 15098
rect 24584 14476 24636 14482
rect 24584 14418 24636 14424
rect 24596 13870 24624 14418
rect 24492 13864 24544 13870
rect 24492 13806 24544 13812
rect 24584 13864 24636 13870
rect 24584 13806 24636 13812
rect 24492 13184 24544 13190
rect 24492 13126 24544 13132
rect 24400 12844 24452 12850
rect 24400 12786 24452 12792
rect 24504 11558 24532 13126
rect 24596 12306 24624 13806
rect 24688 12322 24716 15807
rect 24872 15706 24900 16215
rect 24952 15972 25004 15978
rect 24952 15914 25004 15920
rect 24860 15700 24912 15706
rect 24860 15642 24912 15648
rect 24860 15428 24912 15434
rect 24860 15370 24912 15376
rect 24872 12889 24900 15370
rect 24858 12880 24914 12889
rect 24858 12815 24914 12824
rect 24584 12300 24636 12306
rect 24688 12294 24808 12322
rect 24584 12242 24636 12248
rect 24674 12200 24730 12209
rect 24674 12135 24730 12144
rect 24582 11656 24638 11665
rect 24582 11591 24638 11600
rect 24492 11552 24544 11558
rect 24492 11494 24544 11500
rect 24596 11354 24624 11591
rect 24584 11348 24636 11354
rect 24584 11290 24636 11296
rect 24688 10606 24716 12135
rect 24780 11354 24808 12294
rect 24860 11824 24912 11830
rect 24858 11792 24860 11801
rect 24912 11792 24914 11801
rect 24858 11727 24914 11736
rect 24858 11384 24914 11393
rect 24768 11348 24820 11354
rect 24858 11319 24914 11328
rect 24768 11290 24820 11296
rect 24780 11150 24808 11290
rect 24872 11218 24900 11319
rect 24860 11212 24912 11218
rect 24860 11154 24912 11160
rect 24768 11144 24820 11150
rect 24768 11086 24820 11092
rect 24766 10976 24822 10985
rect 24766 10911 24822 10920
rect 24676 10600 24728 10606
rect 24676 10542 24728 10548
rect 24582 10160 24638 10169
rect 24582 10095 24638 10104
rect 24596 8430 24624 10095
rect 24780 9518 24808 10911
rect 24860 10736 24912 10742
rect 24860 10678 24912 10684
rect 24872 10577 24900 10678
rect 24858 10568 24914 10577
rect 24858 10503 24914 10512
rect 24768 9512 24820 9518
rect 24768 9454 24820 9460
rect 24858 9344 24914 9353
rect 24858 9279 24914 9288
rect 24872 9042 24900 9279
rect 24860 9036 24912 9042
rect 24860 8978 24912 8984
rect 24674 8936 24730 8945
rect 24674 8871 24730 8880
rect 24584 8424 24636 8430
rect 24584 8366 24636 8372
rect 24400 8356 24452 8362
rect 24400 8298 24452 8304
rect 23584 6886 23704 6914
rect 23676 6322 23704 6886
rect 24228 6886 24348 6914
rect 23664 6316 23716 6322
rect 23664 6258 23716 6264
rect 23480 5704 23532 5710
rect 23480 5646 23532 5652
rect 23480 5568 23532 5574
rect 23480 5510 23532 5516
rect 22652 4616 22704 4622
rect 22652 4558 22704 4564
rect 23388 4616 23440 4622
rect 23388 4558 23440 4564
rect 22100 4072 22152 4078
rect 22100 4014 22152 4020
rect 22008 3460 22060 3466
rect 22008 3402 22060 3408
rect 20628 2440 20680 2446
rect 20628 2382 20680 2388
rect 22020 1170 22048 3402
rect 22112 1601 22140 4014
rect 22950 3836 23258 3845
rect 22950 3834 22956 3836
rect 23012 3834 23036 3836
rect 23092 3834 23116 3836
rect 23172 3834 23196 3836
rect 23252 3834 23258 3836
rect 23012 3782 23014 3834
rect 23194 3782 23196 3834
rect 22950 3780 22956 3782
rect 23012 3780 23036 3782
rect 23092 3780 23116 3782
rect 23172 3780 23196 3782
rect 23252 3780 23258 3782
rect 22950 3771 23258 3780
rect 23492 3534 23520 5510
rect 23572 4480 23624 4486
rect 23572 4422 23624 4428
rect 23480 3528 23532 3534
rect 23480 3470 23532 3476
rect 23584 3058 23612 4422
rect 24228 3058 24256 6886
rect 24412 5710 24440 8298
rect 24688 7342 24716 8871
rect 24860 8560 24912 8566
rect 24858 8528 24860 8537
rect 24912 8528 24914 8537
rect 24964 8498 24992 15914
rect 25044 15428 25096 15434
rect 25044 15370 25096 15376
rect 24858 8463 24914 8472
rect 24952 8492 25004 8498
rect 24952 8434 25004 8440
rect 24950 8120 25006 8129
rect 24950 8055 25006 8064
rect 24964 7954 24992 8055
rect 24952 7948 25004 7954
rect 24952 7890 25004 7896
rect 24766 7712 24822 7721
rect 24766 7647 24822 7656
rect 24676 7336 24728 7342
rect 24676 7278 24728 7284
rect 24674 6488 24730 6497
rect 24674 6423 24730 6432
rect 24584 5840 24636 5846
rect 24584 5782 24636 5788
rect 24400 5704 24452 5710
rect 24400 5646 24452 5652
rect 24596 3534 24624 5782
rect 24688 5166 24716 6423
rect 24780 6254 24808 7647
rect 24860 7472 24912 7478
rect 24860 7414 24912 7420
rect 24872 7313 24900 7414
rect 25056 7410 25084 15370
rect 25136 14612 25188 14618
rect 25136 14554 25188 14560
rect 25148 14006 25176 14554
rect 25228 14476 25280 14482
rect 25228 14418 25280 14424
rect 25136 14000 25188 14006
rect 25136 13942 25188 13948
rect 25134 12608 25190 12617
rect 25134 12543 25190 12552
rect 25148 11830 25176 12543
rect 25136 11824 25188 11830
rect 25136 11766 25188 11772
rect 25240 9994 25268 14418
rect 25332 13326 25360 18226
rect 25424 18222 25452 23530
rect 25504 22432 25556 22438
rect 25504 22374 25556 22380
rect 25516 19281 25544 22374
rect 25502 19272 25558 19281
rect 25502 19207 25558 19216
rect 25504 18692 25556 18698
rect 25504 18634 25556 18640
rect 25412 18216 25464 18222
rect 25412 18158 25464 18164
rect 25412 15496 25464 15502
rect 25412 15438 25464 15444
rect 25320 13320 25372 13326
rect 25320 13262 25372 13268
rect 25424 12434 25452 15438
rect 25332 12406 25452 12434
rect 25516 12434 25544 18634
rect 25608 18358 25636 25162
rect 25792 22234 25820 26415
rect 26148 25288 26200 25294
rect 26148 25230 26200 25236
rect 25872 22568 25924 22574
rect 25872 22510 25924 22516
rect 25780 22228 25832 22234
rect 25780 22170 25832 22176
rect 25688 21480 25740 21486
rect 25688 21422 25740 21428
rect 25596 18352 25648 18358
rect 25596 18294 25648 18300
rect 25608 14550 25636 18294
rect 25596 14544 25648 14550
rect 25596 14486 25648 14492
rect 25596 14408 25648 14414
rect 25596 14350 25648 14356
rect 25608 12866 25636 14350
rect 25700 12986 25728 21422
rect 25688 12980 25740 12986
rect 25688 12922 25740 12928
rect 25608 12838 25728 12866
rect 25516 12406 25636 12434
rect 25228 9988 25280 9994
rect 25228 9930 25280 9936
rect 25044 7404 25096 7410
rect 25044 7346 25096 7352
rect 24858 7304 24914 7313
rect 24858 7239 24914 7248
rect 25332 6914 25360 12406
rect 25608 7818 25636 12406
rect 25700 11354 25728 12838
rect 25688 11348 25740 11354
rect 25688 11290 25740 11296
rect 25792 9178 25820 22170
rect 25884 17746 25912 22510
rect 25964 22024 26016 22030
rect 25964 21966 26016 21972
rect 25976 19922 26004 21966
rect 26056 20800 26108 20806
rect 26056 20742 26108 20748
rect 25964 19916 26016 19922
rect 25964 19858 26016 19864
rect 25964 19712 26016 19718
rect 25964 19654 26016 19660
rect 25872 17740 25924 17746
rect 25872 17682 25924 17688
rect 25872 16040 25924 16046
rect 25870 16008 25872 16017
rect 25924 16008 25926 16017
rect 25870 15943 25926 15952
rect 25884 14414 25912 15943
rect 25872 14408 25924 14414
rect 25872 14350 25924 14356
rect 25872 13864 25924 13870
rect 25872 13806 25924 13812
rect 25780 9172 25832 9178
rect 25780 9114 25832 9120
rect 25596 7812 25648 7818
rect 25596 7754 25648 7760
rect 24858 6896 24914 6905
rect 24858 6831 24860 6840
rect 24912 6831 24914 6840
rect 25148 6886 25360 6914
rect 24860 6802 24912 6808
rect 25044 6724 25096 6730
rect 25044 6666 25096 6672
rect 24860 6384 24912 6390
rect 24860 6326 24912 6332
rect 24768 6248 24820 6254
rect 24768 6190 24820 6196
rect 24872 6089 24900 6326
rect 24858 6080 24914 6089
rect 24858 6015 24914 6024
rect 24950 5672 25006 5681
rect 24950 5607 24952 5616
rect 25004 5607 25006 5616
rect 24952 5578 25004 5584
rect 24860 5296 24912 5302
rect 24766 5264 24822 5273
rect 24860 5238 24912 5244
rect 24766 5199 24822 5208
rect 24676 5160 24728 5166
rect 24676 5102 24728 5108
rect 24780 4078 24808 5199
rect 24872 4865 24900 5238
rect 24858 4856 24914 4865
rect 24858 4791 24914 4800
rect 24952 4548 25004 4554
rect 24952 4490 25004 4496
rect 24964 4457 24992 4490
rect 24950 4448 25006 4457
rect 24950 4383 25006 4392
rect 24768 4072 24820 4078
rect 24768 4014 24820 4020
rect 24952 4004 25004 4010
rect 24952 3946 25004 3952
rect 24964 3641 24992 3946
rect 25056 3942 25084 6666
rect 25148 4146 25176 6886
rect 25136 4140 25188 4146
rect 25136 4082 25188 4088
rect 25134 4040 25190 4049
rect 25134 3975 25190 3984
rect 25044 3936 25096 3942
rect 25044 3878 25096 3884
rect 24950 3632 25006 3641
rect 24950 3567 25006 3576
rect 24584 3528 24636 3534
rect 24584 3470 24636 3476
rect 24952 3460 25004 3466
rect 24952 3402 25004 3408
rect 24584 3392 24636 3398
rect 24584 3334 24636 3340
rect 23572 3052 23624 3058
rect 23572 2994 23624 3000
rect 24216 3052 24268 3058
rect 24216 2994 24268 3000
rect 22950 2748 23258 2757
rect 22950 2746 22956 2748
rect 23012 2746 23036 2748
rect 23092 2746 23116 2748
rect 23172 2746 23196 2748
rect 23252 2746 23258 2748
rect 23012 2694 23014 2746
rect 23194 2694 23196 2746
rect 22950 2692 22956 2694
rect 23012 2692 23036 2694
rect 23092 2692 23116 2694
rect 23172 2692 23196 2694
rect 23252 2692 23258 2694
rect 22950 2683 23258 2692
rect 22192 2644 22244 2650
rect 22192 2586 22244 2592
rect 22204 2009 22232 2586
rect 24596 2446 24624 3334
rect 24964 3233 24992 3402
rect 24950 3224 25006 3233
rect 24950 3159 25006 3168
rect 25148 3126 25176 3975
rect 24860 3120 24912 3126
rect 24860 3062 24912 3068
rect 25136 3120 25188 3126
rect 25136 3062 25188 3068
rect 24872 2825 24900 3062
rect 25044 2984 25096 2990
rect 25044 2926 25096 2932
rect 24858 2816 24914 2825
rect 24858 2751 24914 2760
rect 24584 2440 24636 2446
rect 24584 2382 24636 2388
rect 24950 2408 25006 2417
rect 23388 2372 23440 2378
rect 24950 2343 24952 2352
rect 23388 2314 23440 2320
rect 25004 2343 25006 2352
rect 24952 2314 25004 2320
rect 22190 2000 22246 2009
rect 22190 1935 22246 1944
rect 22098 1592 22154 1601
rect 22098 1527 22154 1536
rect 22098 1184 22154 1193
rect 22020 1142 22098 1170
rect 22098 1119 22154 1128
rect 6734 0 6790 800
rect 20166 0 20222 800
rect 23400 377 23428 2314
rect 25056 785 25084 2926
rect 25884 2854 25912 13806
rect 25976 12918 26004 19654
rect 26068 14385 26096 20742
rect 26160 14618 26188 25230
rect 26240 21888 26292 21894
rect 26240 21830 26292 21836
rect 26252 16046 26280 21830
rect 26240 16040 26292 16046
rect 26240 15982 26292 15988
rect 26148 14612 26200 14618
rect 26148 14554 26200 14560
rect 26054 14376 26110 14385
rect 26054 14311 26110 14320
rect 25964 12912 26016 12918
rect 25964 12854 26016 12860
rect 26068 12434 26096 14311
rect 25976 12406 26096 12434
rect 25976 11286 26004 12406
rect 25964 11280 26016 11286
rect 25964 11222 26016 11228
rect 25872 2848 25924 2854
rect 25872 2790 25924 2796
rect 25042 776 25098 785
rect 25042 711 25098 720
rect 23386 368 23442 377
rect 23386 303 23442 312
<< via2 >>
rect 1766 24148 1768 24168
rect 1768 24148 1820 24168
rect 1820 24148 1822 24168
rect 1766 24112 1822 24148
rect 1122 23724 1178 23760
rect 1122 23704 1124 23724
rect 1124 23704 1176 23724
rect 1176 23704 1178 23724
rect 1214 22636 1270 22672
rect 1214 22616 1216 22636
rect 1216 22616 1268 22636
rect 1268 22616 1270 22636
rect 2956 24506 3012 24508
rect 3036 24506 3092 24508
rect 3116 24506 3172 24508
rect 3196 24506 3252 24508
rect 2956 24454 3002 24506
rect 3002 24454 3012 24506
rect 3036 24454 3066 24506
rect 3066 24454 3078 24506
rect 3078 24454 3092 24506
rect 3116 24454 3130 24506
rect 3130 24454 3142 24506
rect 3142 24454 3172 24506
rect 3196 24454 3206 24506
rect 3206 24454 3252 24506
rect 2956 24452 3012 24454
rect 3036 24452 3092 24454
rect 3116 24452 3172 24454
rect 3196 24452 3252 24454
rect 2956 23418 3012 23420
rect 3036 23418 3092 23420
rect 3116 23418 3172 23420
rect 3196 23418 3252 23420
rect 2956 23366 3002 23418
rect 3002 23366 3012 23418
rect 3036 23366 3066 23418
rect 3066 23366 3078 23418
rect 3078 23366 3092 23418
rect 3116 23366 3130 23418
rect 3130 23366 3142 23418
rect 3142 23366 3172 23418
rect 3196 23366 3206 23418
rect 3206 23366 3252 23418
rect 2956 23364 3012 23366
rect 3036 23364 3092 23366
rect 3116 23364 3172 23366
rect 3196 23364 3252 23366
rect 3238 22516 3240 22536
rect 3240 22516 3292 22536
rect 3292 22516 3294 22536
rect 3238 22480 3294 22516
rect 2956 22330 3012 22332
rect 3036 22330 3092 22332
rect 3116 22330 3172 22332
rect 3196 22330 3252 22332
rect 2956 22278 3002 22330
rect 3002 22278 3012 22330
rect 3036 22278 3066 22330
rect 3066 22278 3078 22330
rect 3078 22278 3092 22330
rect 3116 22278 3130 22330
rect 3130 22278 3142 22330
rect 3142 22278 3172 22330
rect 3196 22278 3206 22330
rect 3206 22278 3252 22330
rect 2956 22276 3012 22278
rect 3036 22276 3092 22278
rect 3116 22276 3172 22278
rect 3196 22276 3252 22278
rect 2956 21242 3012 21244
rect 3036 21242 3092 21244
rect 3116 21242 3172 21244
rect 3196 21242 3252 21244
rect 2956 21190 3002 21242
rect 3002 21190 3012 21242
rect 3036 21190 3066 21242
rect 3066 21190 3078 21242
rect 3078 21190 3092 21242
rect 3116 21190 3130 21242
rect 3130 21190 3142 21242
rect 3142 21190 3172 21242
rect 3196 21190 3206 21242
rect 3206 21190 3252 21242
rect 2956 21188 3012 21190
rect 3036 21188 3092 21190
rect 3116 21188 3172 21190
rect 3196 21188 3252 21190
rect 3422 24792 3478 24848
rect 3698 25880 3754 25936
rect 3790 22480 3846 22536
rect 3514 20168 3570 20224
rect 2956 20154 3012 20156
rect 3036 20154 3092 20156
rect 3116 20154 3172 20156
rect 3196 20154 3252 20156
rect 2956 20102 3002 20154
rect 3002 20102 3012 20154
rect 3036 20102 3066 20154
rect 3066 20102 3078 20154
rect 3078 20102 3092 20154
rect 3116 20102 3130 20154
rect 3130 20102 3142 20154
rect 3142 20102 3172 20154
rect 3196 20102 3206 20154
rect 3206 20102 3252 20154
rect 2956 20100 3012 20102
rect 3036 20100 3092 20102
rect 3116 20100 3172 20102
rect 3196 20100 3252 20102
rect 2956 19066 3012 19068
rect 3036 19066 3092 19068
rect 3116 19066 3172 19068
rect 3196 19066 3252 19068
rect 2956 19014 3002 19066
rect 3002 19014 3012 19066
rect 3036 19014 3066 19066
rect 3066 19014 3078 19066
rect 3078 19014 3092 19066
rect 3116 19014 3130 19066
rect 3130 19014 3142 19066
rect 3142 19014 3172 19066
rect 3196 19014 3206 19066
rect 3206 19014 3252 19066
rect 2956 19012 3012 19014
rect 3036 19012 3092 19014
rect 3116 19012 3172 19014
rect 3196 19012 3252 19014
rect 2594 18844 2596 18864
rect 2596 18844 2648 18864
rect 2648 18844 2650 18864
rect 2594 18808 2650 18844
rect 2226 18300 2228 18320
rect 2228 18300 2280 18320
rect 2280 18300 2282 18320
rect 2226 18264 2282 18300
rect 2956 17978 3012 17980
rect 3036 17978 3092 17980
rect 3116 17978 3172 17980
rect 3196 17978 3252 17980
rect 2956 17926 3002 17978
rect 3002 17926 3012 17978
rect 3036 17926 3066 17978
rect 3066 17926 3078 17978
rect 3078 17926 3092 17978
rect 3116 17926 3130 17978
rect 3130 17926 3142 17978
rect 3142 17926 3172 17978
rect 3196 17926 3206 17978
rect 3206 17926 3252 17978
rect 2956 17924 3012 17926
rect 3036 17924 3092 17926
rect 3116 17924 3172 17926
rect 3196 17924 3252 17926
rect 3790 21528 3846 21584
rect 4894 26152 4950 26208
rect 4802 24928 4858 24984
rect 3882 18692 3938 18728
rect 3882 18672 3884 18692
rect 3884 18672 3936 18692
rect 3936 18672 3938 18692
rect 2956 16890 3012 16892
rect 3036 16890 3092 16892
rect 3116 16890 3172 16892
rect 3196 16890 3252 16892
rect 2956 16838 3002 16890
rect 3002 16838 3012 16890
rect 3036 16838 3066 16890
rect 3066 16838 3078 16890
rect 3078 16838 3092 16890
rect 3116 16838 3130 16890
rect 3130 16838 3142 16890
rect 3142 16838 3172 16890
rect 3196 16838 3206 16890
rect 3206 16838 3252 16890
rect 2956 16836 3012 16838
rect 3036 16836 3092 16838
rect 3116 16836 3172 16838
rect 3196 16836 3252 16838
rect 2956 15802 3012 15804
rect 3036 15802 3092 15804
rect 3116 15802 3172 15804
rect 3196 15802 3252 15804
rect 2956 15750 3002 15802
rect 3002 15750 3012 15802
rect 3036 15750 3066 15802
rect 3066 15750 3078 15802
rect 3078 15750 3092 15802
rect 3116 15750 3130 15802
rect 3130 15750 3142 15802
rect 3142 15750 3172 15802
rect 3196 15750 3206 15802
rect 3206 15750 3252 15802
rect 2956 15748 3012 15750
rect 3036 15748 3092 15750
rect 3116 15748 3172 15750
rect 3196 15748 3252 15750
rect 2956 14714 3012 14716
rect 3036 14714 3092 14716
rect 3116 14714 3172 14716
rect 3196 14714 3252 14716
rect 2956 14662 3002 14714
rect 3002 14662 3012 14714
rect 3036 14662 3066 14714
rect 3066 14662 3078 14714
rect 3078 14662 3092 14714
rect 3116 14662 3130 14714
rect 3130 14662 3142 14714
rect 3142 14662 3172 14714
rect 3196 14662 3206 14714
rect 3206 14662 3252 14714
rect 2956 14660 3012 14662
rect 3036 14660 3092 14662
rect 3116 14660 3172 14662
rect 3196 14660 3252 14662
rect 2956 13626 3012 13628
rect 3036 13626 3092 13628
rect 3116 13626 3172 13628
rect 3196 13626 3252 13628
rect 2956 13574 3002 13626
rect 3002 13574 3012 13626
rect 3036 13574 3066 13626
rect 3066 13574 3078 13626
rect 3078 13574 3092 13626
rect 3116 13574 3130 13626
rect 3130 13574 3142 13626
rect 3142 13574 3172 13626
rect 3196 13574 3206 13626
rect 3206 13574 3252 13626
rect 2956 13572 3012 13574
rect 3036 13572 3092 13574
rect 3116 13572 3172 13574
rect 3196 13572 3252 13574
rect 2956 12538 3012 12540
rect 3036 12538 3092 12540
rect 3116 12538 3172 12540
rect 3196 12538 3252 12540
rect 2956 12486 3002 12538
rect 3002 12486 3012 12538
rect 3036 12486 3066 12538
rect 3066 12486 3078 12538
rect 3078 12486 3092 12538
rect 3116 12486 3130 12538
rect 3130 12486 3142 12538
rect 3142 12486 3172 12538
rect 3196 12486 3206 12538
rect 3206 12486 3252 12538
rect 2956 12484 3012 12486
rect 3036 12484 3092 12486
rect 3116 12484 3172 12486
rect 3196 12484 3252 12486
rect 4158 16532 4160 16552
rect 4160 16532 4212 16552
rect 4212 16532 4214 16552
rect 4158 16496 4214 16532
rect 4802 22072 4858 22128
rect 4710 19080 4766 19136
rect 5446 23568 5502 23624
rect 5630 21256 5686 21312
rect 5814 21120 5870 21176
rect 5538 20304 5594 20360
rect 4802 16904 4858 16960
rect 5906 20712 5962 20768
rect 6550 25064 6606 25120
rect 6274 22616 6330 22672
rect 6366 22208 6422 22264
rect 6734 23316 6790 23352
rect 6734 23296 6736 23316
rect 6736 23296 6788 23316
rect 6788 23296 6790 23316
rect 6458 19252 6460 19272
rect 6460 19252 6512 19272
rect 6512 19252 6514 19272
rect 6458 19216 6514 19252
rect 7010 20712 7066 20768
rect 6642 19352 6698 19408
rect 6550 17856 6606 17912
rect 6550 14864 6606 14920
rect 4526 14320 4582 14376
rect 7010 18148 7066 18184
rect 7010 18128 7012 18148
rect 7012 18128 7064 18148
rect 7064 18128 7066 18148
rect 7286 19896 7342 19952
rect 7286 18028 7288 18048
rect 7288 18028 7340 18048
rect 7340 18028 7342 18048
rect 7286 17992 7342 18028
rect 6918 17756 6920 17776
rect 6920 17756 6972 17776
rect 6972 17756 6974 17776
rect 6918 17720 6974 17756
rect 7102 17584 7158 17640
rect 7010 16768 7066 16824
rect 6826 16088 6882 16144
rect 7956 23962 8012 23964
rect 8036 23962 8092 23964
rect 8116 23962 8172 23964
rect 8196 23962 8252 23964
rect 7956 23910 8002 23962
rect 8002 23910 8012 23962
rect 8036 23910 8066 23962
rect 8066 23910 8078 23962
rect 8078 23910 8092 23962
rect 8116 23910 8130 23962
rect 8130 23910 8142 23962
rect 8142 23910 8172 23962
rect 8196 23910 8206 23962
rect 8206 23910 8252 23962
rect 7956 23908 8012 23910
rect 8036 23908 8092 23910
rect 8116 23908 8172 23910
rect 8196 23908 8252 23910
rect 7956 22874 8012 22876
rect 8036 22874 8092 22876
rect 8116 22874 8172 22876
rect 8196 22874 8252 22876
rect 7956 22822 8002 22874
rect 8002 22822 8012 22874
rect 8036 22822 8066 22874
rect 8066 22822 8078 22874
rect 8078 22822 8092 22874
rect 8116 22822 8130 22874
rect 8130 22822 8142 22874
rect 8142 22822 8172 22874
rect 8196 22822 8206 22874
rect 8206 22822 8252 22874
rect 7956 22820 8012 22822
rect 8036 22820 8092 22822
rect 8116 22820 8172 22822
rect 8196 22820 8252 22822
rect 8666 23704 8722 23760
rect 8574 23296 8630 23352
rect 8390 23160 8446 23216
rect 7956 21786 8012 21788
rect 8036 21786 8092 21788
rect 8116 21786 8172 21788
rect 8196 21786 8252 21788
rect 7956 21734 8002 21786
rect 8002 21734 8012 21786
rect 8036 21734 8066 21786
rect 8066 21734 8078 21786
rect 8078 21734 8092 21786
rect 8116 21734 8130 21786
rect 8130 21734 8142 21786
rect 8142 21734 8172 21786
rect 8196 21734 8206 21786
rect 8206 21734 8252 21786
rect 7956 21732 8012 21734
rect 8036 21732 8092 21734
rect 8116 21732 8172 21734
rect 8196 21732 8252 21734
rect 7838 21392 7894 21448
rect 7746 19216 7802 19272
rect 7654 17176 7710 17232
rect 8298 20868 8354 20904
rect 8298 20848 8300 20868
rect 8300 20848 8352 20868
rect 8352 20848 8354 20868
rect 7956 20698 8012 20700
rect 8036 20698 8092 20700
rect 8116 20698 8172 20700
rect 8196 20698 8252 20700
rect 7956 20646 8002 20698
rect 8002 20646 8012 20698
rect 8036 20646 8066 20698
rect 8066 20646 8078 20698
rect 8078 20646 8092 20698
rect 8116 20646 8130 20698
rect 8130 20646 8142 20698
rect 8142 20646 8172 20698
rect 8196 20646 8206 20698
rect 8206 20646 8252 20698
rect 7956 20644 8012 20646
rect 8036 20644 8092 20646
rect 8116 20644 8172 20646
rect 8196 20644 8252 20646
rect 8574 23024 8630 23080
rect 8482 21684 8538 21720
rect 8482 21664 8484 21684
rect 8484 21664 8536 21684
rect 8536 21664 8538 21684
rect 8298 19780 8354 19816
rect 8298 19760 8300 19780
rect 8300 19760 8352 19780
rect 8352 19760 8354 19780
rect 7956 19610 8012 19612
rect 8036 19610 8092 19612
rect 8116 19610 8172 19612
rect 8196 19610 8252 19612
rect 7956 19558 8002 19610
rect 8002 19558 8012 19610
rect 8036 19558 8066 19610
rect 8066 19558 8078 19610
rect 8078 19558 8092 19610
rect 8116 19558 8130 19610
rect 8130 19558 8142 19610
rect 8142 19558 8172 19610
rect 8196 19558 8206 19610
rect 8206 19558 8252 19610
rect 7956 19556 8012 19558
rect 8036 19556 8092 19558
rect 8116 19556 8172 19558
rect 8196 19556 8252 19558
rect 8114 18672 8170 18728
rect 7956 18522 8012 18524
rect 8036 18522 8092 18524
rect 8116 18522 8172 18524
rect 8196 18522 8252 18524
rect 7956 18470 8002 18522
rect 8002 18470 8012 18522
rect 8036 18470 8066 18522
rect 8066 18470 8078 18522
rect 8078 18470 8092 18522
rect 8116 18470 8130 18522
rect 8130 18470 8142 18522
rect 8142 18470 8172 18522
rect 8196 18470 8206 18522
rect 8206 18470 8252 18522
rect 7956 18468 8012 18470
rect 8036 18468 8092 18470
rect 8116 18468 8172 18470
rect 8196 18468 8252 18470
rect 8758 20984 8814 21040
rect 9126 23432 9182 23488
rect 9310 20440 9366 20496
rect 7956 17434 8012 17436
rect 8036 17434 8092 17436
rect 8116 17434 8172 17436
rect 8196 17434 8252 17436
rect 7956 17382 8002 17434
rect 8002 17382 8012 17434
rect 8036 17382 8066 17434
rect 8066 17382 8078 17434
rect 8078 17382 8092 17434
rect 8116 17382 8130 17434
rect 8130 17382 8142 17434
rect 8142 17382 8172 17434
rect 8196 17382 8206 17434
rect 8206 17382 8252 17434
rect 7956 17380 8012 17382
rect 8036 17380 8092 17382
rect 8116 17380 8172 17382
rect 8196 17380 8252 17382
rect 7930 17040 7986 17096
rect 8758 17312 8814 17368
rect 8390 16360 8446 16416
rect 7956 16346 8012 16348
rect 8036 16346 8092 16348
rect 8116 16346 8172 16348
rect 8196 16346 8252 16348
rect 7956 16294 8002 16346
rect 8002 16294 8012 16346
rect 8036 16294 8066 16346
rect 8066 16294 8078 16346
rect 8078 16294 8092 16346
rect 8116 16294 8130 16346
rect 8130 16294 8142 16346
rect 8142 16294 8172 16346
rect 8196 16294 8206 16346
rect 8206 16294 8252 16346
rect 7956 16292 8012 16294
rect 8036 16292 8092 16294
rect 8116 16292 8172 16294
rect 8196 16292 8252 16294
rect 7956 15258 8012 15260
rect 8036 15258 8092 15260
rect 8116 15258 8172 15260
rect 8196 15258 8252 15260
rect 7956 15206 8002 15258
rect 8002 15206 8012 15258
rect 8036 15206 8066 15258
rect 8066 15206 8078 15258
rect 8078 15206 8092 15258
rect 8116 15206 8130 15258
rect 8130 15206 8142 15258
rect 8142 15206 8172 15258
rect 8196 15206 8206 15258
rect 8206 15206 8252 15258
rect 7956 15204 8012 15206
rect 8036 15204 8092 15206
rect 8116 15204 8172 15206
rect 8196 15204 8252 15206
rect 7956 14170 8012 14172
rect 8036 14170 8092 14172
rect 8116 14170 8172 14172
rect 8196 14170 8252 14172
rect 7956 14118 8002 14170
rect 8002 14118 8012 14170
rect 8036 14118 8066 14170
rect 8066 14118 8078 14170
rect 8078 14118 8092 14170
rect 8116 14118 8130 14170
rect 8130 14118 8142 14170
rect 8142 14118 8172 14170
rect 8196 14118 8206 14170
rect 8206 14118 8252 14170
rect 7956 14116 8012 14118
rect 8036 14116 8092 14118
rect 8116 14116 8172 14118
rect 8196 14116 8252 14118
rect 7378 13776 7434 13832
rect 7956 13082 8012 13084
rect 8036 13082 8092 13084
rect 8116 13082 8172 13084
rect 8196 13082 8252 13084
rect 7956 13030 8002 13082
rect 8002 13030 8012 13082
rect 8036 13030 8066 13082
rect 8066 13030 8078 13082
rect 8078 13030 8092 13082
rect 8116 13030 8130 13082
rect 8130 13030 8142 13082
rect 8142 13030 8172 13082
rect 8196 13030 8206 13082
rect 8206 13030 8252 13082
rect 7956 13028 8012 13030
rect 8036 13028 8092 13030
rect 8116 13028 8172 13030
rect 8196 13028 8252 13030
rect 6734 12824 6790 12880
rect 7956 11994 8012 11996
rect 8036 11994 8092 11996
rect 8116 11994 8172 11996
rect 8196 11994 8252 11996
rect 7956 11942 8002 11994
rect 8002 11942 8012 11994
rect 8036 11942 8066 11994
rect 8066 11942 8078 11994
rect 8078 11942 8092 11994
rect 8116 11942 8130 11994
rect 8130 11942 8142 11994
rect 8142 11942 8172 11994
rect 8196 11942 8206 11994
rect 8206 11942 8252 11994
rect 7956 11940 8012 11942
rect 8036 11940 8092 11942
rect 8116 11940 8172 11942
rect 8196 11940 8252 11942
rect 2956 11450 3012 11452
rect 3036 11450 3092 11452
rect 3116 11450 3172 11452
rect 3196 11450 3252 11452
rect 2956 11398 3002 11450
rect 3002 11398 3012 11450
rect 3036 11398 3066 11450
rect 3066 11398 3078 11450
rect 3078 11398 3092 11450
rect 3116 11398 3130 11450
rect 3130 11398 3142 11450
rect 3142 11398 3172 11450
rect 3196 11398 3206 11450
rect 3206 11398 3252 11450
rect 2956 11396 3012 11398
rect 3036 11396 3092 11398
rect 3116 11396 3172 11398
rect 3196 11396 3252 11398
rect 7956 10906 8012 10908
rect 8036 10906 8092 10908
rect 8116 10906 8172 10908
rect 8196 10906 8252 10908
rect 7956 10854 8002 10906
rect 8002 10854 8012 10906
rect 8036 10854 8066 10906
rect 8066 10854 8078 10906
rect 8078 10854 8092 10906
rect 8116 10854 8130 10906
rect 8130 10854 8142 10906
rect 8142 10854 8172 10906
rect 8196 10854 8206 10906
rect 8206 10854 8252 10906
rect 7956 10852 8012 10854
rect 8036 10852 8092 10854
rect 8116 10852 8172 10854
rect 8196 10852 8252 10854
rect 2956 10362 3012 10364
rect 3036 10362 3092 10364
rect 3116 10362 3172 10364
rect 3196 10362 3252 10364
rect 2956 10310 3002 10362
rect 3002 10310 3012 10362
rect 3036 10310 3066 10362
rect 3066 10310 3078 10362
rect 3078 10310 3092 10362
rect 3116 10310 3130 10362
rect 3130 10310 3142 10362
rect 3142 10310 3172 10362
rect 3196 10310 3206 10362
rect 3206 10310 3252 10362
rect 2956 10308 3012 10310
rect 3036 10308 3092 10310
rect 3116 10308 3172 10310
rect 3196 10308 3252 10310
rect 7956 9818 8012 9820
rect 8036 9818 8092 9820
rect 8116 9818 8172 9820
rect 8196 9818 8252 9820
rect 7956 9766 8002 9818
rect 8002 9766 8012 9818
rect 8036 9766 8066 9818
rect 8066 9766 8078 9818
rect 8078 9766 8092 9818
rect 8116 9766 8130 9818
rect 8130 9766 8142 9818
rect 8142 9766 8172 9818
rect 8196 9766 8206 9818
rect 8206 9766 8252 9818
rect 7956 9764 8012 9766
rect 8036 9764 8092 9766
rect 8116 9764 8172 9766
rect 8196 9764 8252 9766
rect 8758 15444 8760 15464
rect 8760 15444 8812 15464
rect 8812 15444 8814 15464
rect 8758 15408 8814 15444
rect 9126 17856 9182 17912
rect 9126 16652 9182 16688
rect 9126 16632 9128 16652
rect 9128 16632 9180 16652
rect 9180 16632 9182 16652
rect 9310 17040 9366 17096
rect 9770 24112 9826 24168
rect 9678 21800 9734 21856
rect 9678 19352 9734 19408
rect 9678 17856 9734 17912
rect 9678 17040 9734 17096
rect 9770 16632 9826 16688
rect 9126 15972 9182 16008
rect 9126 15952 9128 15972
rect 9128 15952 9180 15972
rect 9180 15952 9182 15972
rect 9402 15544 9458 15600
rect 9586 15544 9642 15600
rect 10230 21936 10286 21992
rect 10138 19624 10194 19680
rect 10138 18400 10194 18456
rect 9954 16652 10010 16688
rect 9954 16632 9956 16652
rect 9956 16632 10008 16652
rect 10008 16632 10010 16652
rect 10598 20576 10654 20632
rect 11058 20712 11114 20768
rect 11518 23432 11574 23488
rect 11334 20984 11390 21040
rect 11334 20440 11390 20496
rect 11518 20440 11574 20496
rect 11242 17856 11298 17912
rect 11058 16516 11114 16552
rect 11058 16496 11060 16516
rect 11060 16496 11112 16516
rect 11112 16496 11114 16516
rect 9770 15272 9826 15328
rect 10506 15020 10562 15056
rect 10506 15000 10508 15020
rect 10508 15000 10560 15020
rect 10560 15000 10562 15020
rect 10966 15000 11022 15056
rect 2956 9274 3012 9276
rect 3036 9274 3092 9276
rect 3116 9274 3172 9276
rect 3196 9274 3252 9276
rect 2956 9222 3002 9274
rect 3002 9222 3012 9274
rect 3036 9222 3066 9274
rect 3066 9222 3078 9274
rect 3078 9222 3092 9274
rect 3116 9222 3130 9274
rect 3130 9222 3142 9274
rect 3142 9222 3172 9274
rect 3196 9222 3206 9274
rect 3206 9222 3252 9274
rect 2956 9220 3012 9222
rect 3036 9220 3092 9222
rect 3116 9220 3172 9222
rect 3196 9220 3252 9222
rect 11518 20168 11574 20224
rect 11426 19352 11482 19408
rect 11426 18536 11482 18592
rect 11518 16904 11574 16960
rect 11886 23296 11942 23352
rect 12162 22888 12218 22944
rect 12346 21800 12402 21856
rect 11886 21528 11942 21584
rect 11886 19352 11942 19408
rect 12162 21528 12218 21584
rect 12438 21664 12494 21720
rect 12438 21528 12494 21584
rect 12530 20984 12586 21040
rect 12162 17448 12218 17504
rect 12070 16768 12126 16824
rect 11610 14456 11666 14512
rect 11794 14184 11850 14240
rect 11978 13932 12034 13968
rect 11978 13912 11980 13932
rect 11980 13912 12032 13932
rect 12032 13912 12034 13932
rect 12956 24506 13012 24508
rect 13036 24506 13092 24508
rect 13116 24506 13172 24508
rect 13196 24506 13252 24508
rect 12956 24454 13002 24506
rect 13002 24454 13012 24506
rect 13036 24454 13066 24506
rect 13066 24454 13078 24506
rect 13078 24454 13092 24506
rect 13116 24454 13130 24506
rect 13130 24454 13142 24506
rect 13142 24454 13172 24506
rect 13196 24454 13206 24506
rect 13206 24454 13252 24506
rect 12956 24452 13012 24454
rect 13036 24452 13092 24454
rect 13116 24452 13172 24454
rect 13196 24452 13252 24454
rect 12956 23418 13012 23420
rect 13036 23418 13092 23420
rect 13116 23418 13172 23420
rect 13196 23418 13252 23420
rect 12956 23366 13002 23418
rect 13002 23366 13012 23418
rect 13036 23366 13066 23418
rect 13066 23366 13078 23418
rect 13078 23366 13092 23418
rect 13116 23366 13130 23418
rect 13130 23366 13142 23418
rect 13142 23366 13172 23418
rect 13196 23366 13206 23418
rect 13206 23366 13252 23418
rect 12956 23364 13012 23366
rect 13036 23364 13092 23366
rect 13116 23364 13172 23366
rect 13196 23364 13252 23366
rect 13358 22752 13414 22808
rect 12806 22344 12862 22400
rect 12956 22330 13012 22332
rect 13036 22330 13092 22332
rect 13116 22330 13172 22332
rect 13196 22330 13252 22332
rect 12956 22278 13002 22330
rect 13002 22278 13012 22330
rect 13036 22278 13066 22330
rect 13066 22278 13078 22330
rect 13078 22278 13092 22330
rect 13116 22278 13130 22330
rect 13130 22278 13142 22330
rect 13142 22278 13172 22330
rect 13196 22278 13206 22330
rect 13206 22278 13252 22330
rect 12956 22276 13012 22278
rect 13036 22276 13092 22278
rect 13116 22276 13172 22278
rect 13196 22276 13252 22278
rect 13542 22616 13598 22672
rect 13634 22344 13690 22400
rect 12898 21836 12900 21856
rect 12900 21836 12952 21856
rect 12952 21836 12954 21856
rect 12898 21800 12954 21836
rect 12990 21392 13046 21448
rect 13542 21800 13598 21856
rect 12956 21242 13012 21244
rect 13036 21242 13092 21244
rect 13116 21242 13172 21244
rect 13196 21242 13252 21244
rect 12956 21190 13002 21242
rect 13002 21190 13012 21242
rect 13036 21190 13066 21242
rect 13066 21190 13078 21242
rect 13078 21190 13092 21242
rect 13116 21190 13130 21242
rect 13130 21190 13142 21242
rect 13142 21190 13172 21242
rect 13196 21190 13206 21242
rect 13206 21190 13252 21242
rect 12956 21188 13012 21190
rect 13036 21188 13092 21190
rect 13116 21188 13172 21190
rect 13196 21188 13252 21190
rect 12714 18944 12770 19000
rect 12956 20154 13012 20156
rect 13036 20154 13092 20156
rect 13116 20154 13172 20156
rect 13196 20154 13252 20156
rect 12956 20102 13002 20154
rect 13002 20102 13012 20154
rect 13036 20102 13066 20154
rect 13066 20102 13078 20154
rect 13078 20102 13092 20154
rect 13116 20102 13130 20154
rect 13130 20102 13142 20154
rect 13142 20102 13172 20154
rect 13196 20102 13206 20154
rect 13206 20102 13252 20154
rect 12956 20100 13012 20102
rect 13036 20100 13092 20102
rect 13116 20100 13172 20102
rect 13196 20100 13252 20102
rect 13450 19352 13506 19408
rect 12956 19066 13012 19068
rect 13036 19066 13092 19068
rect 13116 19066 13172 19068
rect 13196 19066 13252 19068
rect 12956 19014 13002 19066
rect 13002 19014 13012 19066
rect 13036 19014 13066 19066
rect 13066 19014 13078 19066
rect 13078 19014 13092 19066
rect 13116 19014 13130 19066
rect 13130 19014 13142 19066
rect 13142 19014 13172 19066
rect 13196 19014 13206 19066
rect 13206 19014 13252 19066
rect 12956 19012 13012 19014
rect 13036 19012 13092 19014
rect 13116 19012 13172 19014
rect 13196 19012 13252 19014
rect 12956 17978 13012 17980
rect 13036 17978 13092 17980
rect 13116 17978 13172 17980
rect 13196 17978 13252 17980
rect 12956 17926 13002 17978
rect 13002 17926 13012 17978
rect 13036 17926 13066 17978
rect 13066 17926 13078 17978
rect 13078 17926 13092 17978
rect 13116 17926 13130 17978
rect 13130 17926 13142 17978
rect 13142 17926 13172 17978
rect 13196 17926 13206 17978
rect 13206 17926 13252 17978
rect 12956 17924 13012 17926
rect 13036 17924 13092 17926
rect 13116 17924 13172 17926
rect 13196 17924 13252 17926
rect 12956 16890 13012 16892
rect 13036 16890 13092 16892
rect 13116 16890 13172 16892
rect 13196 16890 13252 16892
rect 12956 16838 13002 16890
rect 13002 16838 13012 16890
rect 13036 16838 13066 16890
rect 13066 16838 13078 16890
rect 13078 16838 13092 16890
rect 13116 16838 13130 16890
rect 13130 16838 13142 16890
rect 13142 16838 13172 16890
rect 13196 16838 13206 16890
rect 13206 16838 13252 16890
rect 12956 16836 13012 16838
rect 13036 16836 13092 16838
rect 13116 16836 13172 16838
rect 13196 16836 13252 16838
rect 13358 16224 13414 16280
rect 12956 15802 13012 15804
rect 13036 15802 13092 15804
rect 13116 15802 13172 15804
rect 13196 15802 13252 15804
rect 12956 15750 13002 15802
rect 13002 15750 13012 15802
rect 13036 15750 13066 15802
rect 13066 15750 13078 15802
rect 13078 15750 13092 15802
rect 13116 15750 13130 15802
rect 13130 15750 13142 15802
rect 13142 15750 13172 15802
rect 13196 15750 13206 15802
rect 13206 15750 13252 15802
rect 12956 15748 13012 15750
rect 13036 15748 13092 15750
rect 13116 15748 13172 15750
rect 13196 15748 13252 15750
rect 12956 14714 13012 14716
rect 13036 14714 13092 14716
rect 13116 14714 13172 14716
rect 13196 14714 13252 14716
rect 12956 14662 13002 14714
rect 13002 14662 13012 14714
rect 13036 14662 13066 14714
rect 13066 14662 13078 14714
rect 13078 14662 13092 14714
rect 13116 14662 13130 14714
rect 13130 14662 13142 14714
rect 13142 14662 13172 14714
rect 13196 14662 13206 14714
rect 13206 14662 13252 14714
rect 12956 14660 13012 14662
rect 13036 14660 13092 14662
rect 13116 14660 13172 14662
rect 13196 14660 13252 14662
rect 14278 23432 14334 23488
rect 13726 20848 13782 20904
rect 13726 20576 13782 20632
rect 14186 21800 14242 21856
rect 14002 20168 14058 20224
rect 14002 19624 14058 19680
rect 14370 21120 14426 21176
rect 14094 19372 14150 19408
rect 14094 19352 14096 19372
rect 14096 19352 14148 19372
rect 14148 19352 14150 19372
rect 14186 17448 14242 17504
rect 14002 16632 14058 16688
rect 12956 13626 13012 13628
rect 13036 13626 13092 13628
rect 13116 13626 13172 13628
rect 13196 13626 13252 13628
rect 12956 13574 13002 13626
rect 13002 13574 13012 13626
rect 13036 13574 13066 13626
rect 13066 13574 13078 13626
rect 13078 13574 13092 13626
rect 13116 13574 13130 13626
rect 13130 13574 13142 13626
rect 13142 13574 13172 13626
rect 13196 13574 13206 13626
rect 13206 13574 13252 13626
rect 12956 13572 13012 13574
rect 13036 13572 13092 13574
rect 13116 13572 13172 13574
rect 13196 13572 13252 13574
rect 12956 12538 13012 12540
rect 13036 12538 13092 12540
rect 13116 12538 13172 12540
rect 13196 12538 13252 12540
rect 12956 12486 13002 12538
rect 13002 12486 13012 12538
rect 13036 12486 13066 12538
rect 13066 12486 13078 12538
rect 13078 12486 13092 12538
rect 13116 12486 13130 12538
rect 13130 12486 13142 12538
rect 13142 12486 13172 12538
rect 13196 12486 13206 12538
rect 13206 12486 13252 12538
rect 12956 12484 13012 12486
rect 13036 12484 13092 12486
rect 13116 12484 13172 12486
rect 13196 12484 13252 12486
rect 11334 12280 11390 12336
rect 12956 11450 13012 11452
rect 13036 11450 13092 11452
rect 13116 11450 13172 11452
rect 13196 11450 13252 11452
rect 12956 11398 13002 11450
rect 13002 11398 13012 11450
rect 13036 11398 13066 11450
rect 13066 11398 13078 11450
rect 13078 11398 13092 11450
rect 13116 11398 13130 11450
rect 13130 11398 13142 11450
rect 13142 11398 13172 11450
rect 13196 11398 13206 11450
rect 13206 11398 13252 11450
rect 12956 11396 13012 11398
rect 13036 11396 13092 11398
rect 13116 11396 13172 11398
rect 13196 11396 13252 11398
rect 15382 23432 15438 23488
rect 15198 21664 15254 21720
rect 15198 20848 15254 20904
rect 14646 19624 14702 19680
rect 14922 20032 14978 20088
rect 15106 19488 15162 19544
rect 15382 18944 15438 19000
rect 15014 17992 15070 18048
rect 14646 16496 14702 16552
rect 12956 10362 13012 10364
rect 13036 10362 13092 10364
rect 13116 10362 13172 10364
rect 13196 10362 13252 10364
rect 12956 10310 13002 10362
rect 13002 10310 13012 10362
rect 13036 10310 13066 10362
rect 13066 10310 13078 10362
rect 13078 10310 13092 10362
rect 13116 10310 13130 10362
rect 13130 10310 13142 10362
rect 13142 10310 13172 10362
rect 13196 10310 13206 10362
rect 13206 10310 13252 10362
rect 12956 10308 13012 10310
rect 13036 10308 13092 10310
rect 13116 10308 13172 10310
rect 13196 10308 13252 10310
rect 12956 9274 13012 9276
rect 13036 9274 13092 9276
rect 13116 9274 13172 9276
rect 13196 9274 13252 9276
rect 12956 9222 13002 9274
rect 13002 9222 13012 9274
rect 13036 9222 13066 9274
rect 13066 9222 13078 9274
rect 13078 9222 13092 9274
rect 13116 9222 13130 9274
rect 13130 9222 13142 9274
rect 13142 9222 13172 9274
rect 13196 9222 13206 9274
rect 13206 9222 13252 9274
rect 12956 9220 13012 9222
rect 13036 9220 13092 9222
rect 13116 9220 13172 9222
rect 13196 9220 13252 9222
rect 7956 8730 8012 8732
rect 8036 8730 8092 8732
rect 8116 8730 8172 8732
rect 8196 8730 8252 8732
rect 7956 8678 8002 8730
rect 8002 8678 8012 8730
rect 8036 8678 8066 8730
rect 8066 8678 8078 8730
rect 8078 8678 8092 8730
rect 8116 8678 8130 8730
rect 8130 8678 8142 8730
rect 8142 8678 8172 8730
rect 8196 8678 8206 8730
rect 8206 8678 8252 8730
rect 7956 8676 8012 8678
rect 8036 8676 8092 8678
rect 8116 8676 8172 8678
rect 8196 8676 8252 8678
rect 2956 8186 3012 8188
rect 3036 8186 3092 8188
rect 3116 8186 3172 8188
rect 3196 8186 3252 8188
rect 2956 8134 3002 8186
rect 3002 8134 3012 8186
rect 3036 8134 3066 8186
rect 3066 8134 3078 8186
rect 3078 8134 3092 8186
rect 3116 8134 3130 8186
rect 3130 8134 3142 8186
rect 3142 8134 3172 8186
rect 3196 8134 3206 8186
rect 3206 8134 3252 8186
rect 2956 8132 3012 8134
rect 3036 8132 3092 8134
rect 3116 8132 3172 8134
rect 3196 8132 3252 8134
rect 7956 7642 8012 7644
rect 8036 7642 8092 7644
rect 8116 7642 8172 7644
rect 8196 7642 8252 7644
rect 7956 7590 8002 7642
rect 8002 7590 8012 7642
rect 8036 7590 8066 7642
rect 8066 7590 8078 7642
rect 8078 7590 8092 7642
rect 8116 7590 8130 7642
rect 8130 7590 8142 7642
rect 8142 7590 8172 7642
rect 8196 7590 8206 7642
rect 8206 7590 8252 7642
rect 7956 7588 8012 7590
rect 8036 7588 8092 7590
rect 8116 7588 8172 7590
rect 8196 7588 8252 7590
rect 2956 7098 3012 7100
rect 3036 7098 3092 7100
rect 3116 7098 3172 7100
rect 3196 7098 3252 7100
rect 2956 7046 3002 7098
rect 3002 7046 3012 7098
rect 3036 7046 3066 7098
rect 3066 7046 3078 7098
rect 3078 7046 3092 7098
rect 3116 7046 3130 7098
rect 3130 7046 3142 7098
rect 3142 7046 3172 7098
rect 3196 7046 3206 7098
rect 3206 7046 3252 7098
rect 2956 7044 3012 7046
rect 3036 7044 3092 7046
rect 3116 7044 3172 7046
rect 3196 7044 3252 7046
rect 7956 6554 8012 6556
rect 8036 6554 8092 6556
rect 8116 6554 8172 6556
rect 8196 6554 8252 6556
rect 7956 6502 8002 6554
rect 8002 6502 8012 6554
rect 8036 6502 8066 6554
rect 8066 6502 8078 6554
rect 8078 6502 8092 6554
rect 8116 6502 8130 6554
rect 8130 6502 8142 6554
rect 8142 6502 8172 6554
rect 8196 6502 8206 6554
rect 8206 6502 8252 6554
rect 7956 6500 8012 6502
rect 8036 6500 8092 6502
rect 8116 6500 8172 6502
rect 8196 6500 8252 6502
rect 15382 18264 15438 18320
rect 15290 15156 15346 15192
rect 15290 15136 15292 15156
rect 15292 15136 15344 15156
rect 15344 15136 15346 15156
rect 12956 8186 13012 8188
rect 13036 8186 13092 8188
rect 13116 8186 13172 8188
rect 13196 8186 13252 8188
rect 12956 8134 13002 8186
rect 13002 8134 13012 8186
rect 13036 8134 13066 8186
rect 13066 8134 13078 8186
rect 13078 8134 13092 8186
rect 13116 8134 13130 8186
rect 13130 8134 13142 8186
rect 13142 8134 13172 8186
rect 13196 8134 13206 8186
rect 13206 8134 13252 8186
rect 12956 8132 13012 8134
rect 13036 8132 13092 8134
rect 13116 8132 13172 8134
rect 13196 8132 13252 8134
rect 12956 7098 13012 7100
rect 13036 7098 13092 7100
rect 13116 7098 13172 7100
rect 13196 7098 13252 7100
rect 12956 7046 13002 7098
rect 13002 7046 13012 7098
rect 13036 7046 13066 7098
rect 13066 7046 13078 7098
rect 13078 7046 13092 7098
rect 13116 7046 13130 7098
rect 13130 7046 13142 7098
rect 13142 7046 13172 7098
rect 13196 7046 13206 7098
rect 13206 7046 13252 7098
rect 12956 7044 13012 7046
rect 13036 7044 13092 7046
rect 13116 7044 13172 7046
rect 13196 7044 13252 7046
rect 15566 23568 15622 23624
rect 16026 24384 16082 24440
rect 16026 23840 16082 23896
rect 15658 21120 15714 21176
rect 15658 20712 15714 20768
rect 15842 21528 15898 21584
rect 15842 20748 15844 20768
rect 15844 20748 15896 20768
rect 15896 20748 15898 20768
rect 15842 20712 15898 20748
rect 16026 22072 16082 22128
rect 16302 22072 16358 22128
rect 16302 21548 16358 21584
rect 16302 21528 16304 21548
rect 16304 21528 16356 21548
rect 16356 21528 16358 21548
rect 16578 23568 16634 23624
rect 16394 20576 16450 20632
rect 16854 23468 16856 23488
rect 16856 23468 16908 23488
rect 16908 23468 16910 23488
rect 16854 23432 16910 23468
rect 16762 22924 16764 22944
rect 16764 22924 16816 22944
rect 16816 22924 16818 22944
rect 16762 22888 16818 22924
rect 16762 21836 16764 21856
rect 16764 21836 16816 21856
rect 16816 21836 16818 21856
rect 16762 21800 16818 21836
rect 15934 20304 15990 20360
rect 15842 19352 15898 19408
rect 16302 19760 16358 19816
rect 16210 19352 16266 19408
rect 15842 16496 15898 16552
rect 15842 15816 15898 15872
rect 15842 15408 15898 15464
rect 16026 14048 16082 14104
rect 15658 13640 15714 13696
rect 15750 13232 15806 13288
rect 16578 19660 16580 19680
rect 16580 19660 16632 19680
rect 16632 19660 16634 19680
rect 16578 19624 16634 19660
rect 16486 15680 16542 15736
rect 16670 15408 16726 15464
rect 16946 21256 17002 21312
rect 17498 24656 17554 24712
rect 17038 19760 17094 19816
rect 17130 18536 17186 18592
rect 16118 11348 16174 11384
rect 16118 11328 16120 11348
rect 16120 11328 16172 11348
rect 16172 11328 16174 11348
rect 16854 12416 16910 12472
rect 17130 17312 17186 17368
rect 17222 16224 17278 16280
rect 17222 15272 17278 15328
rect 17222 15000 17278 15056
rect 17498 20440 17554 20496
rect 17682 24656 17738 24712
rect 17958 24112 18014 24168
rect 17682 23976 17738 24032
rect 17956 23962 18012 23964
rect 18036 23962 18092 23964
rect 18116 23962 18172 23964
rect 18196 23962 18252 23964
rect 17956 23910 18002 23962
rect 18002 23910 18012 23962
rect 18036 23910 18066 23962
rect 18066 23910 18078 23962
rect 18078 23910 18092 23962
rect 18116 23910 18130 23962
rect 18130 23910 18142 23962
rect 18142 23910 18172 23962
rect 18196 23910 18206 23962
rect 18206 23910 18252 23962
rect 17956 23908 18012 23910
rect 18036 23908 18092 23910
rect 18116 23908 18172 23910
rect 18196 23908 18252 23910
rect 17956 22874 18012 22876
rect 18036 22874 18092 22876
rect 18116 22874 18172 22876
rect 18196 22874 18252 22876
rect 17956 22822 18002 22874
rect 18002 22822 18012 22874
rect 18036 22822 18066 22874
rect 18066 22822 18078 22874
rect 18078 22822 18092 22874
rect 18116 22822 18130 22874
rect 18130 22822 18142 22874
rect 18142 22822 18172 22874
rect 18196 22822 18206 22874
rect 18206 22822 18252 22874
rect 17956 22820 18012 22822
rect 18036 22820 18092 22822
rect 18116 22820 18172 22822
rect 18196 22820 18252 22822
rect 17956 21786 18012 21788
rect 18036 21786 18092 21788
rect 18116 21786 18172 21788
rect 18196 21786 18252 21788
rect 17956 21734 18002 21786
rect 18002 21734 18012 21786
rect 18036 21734 18066 21786
rect 18066 21734 18078 21786
rect 18078 21734 18092 21786
rect 18116 21734 18130 21786
rect 18130 21734 18142 21786
rect 18142 21734 18172 21786
rect 18196 21734 18206 21786
rect 18206 21734 18252 21786
rect 17956 21732 18012 21734
rect 18036 21732 18092 21734
rect 18116 21732 18172 21734
rect 18196 21732 18252 21734
rect 18970 26016 19026 26072
rect 19062 24928 19118 24984
rect 19430 24928 19486 24984
rect 18602 23296 18658 23352
rect 18510 23044 18566 23080
rect 18510 23024 18512 23044
rect 18512 23024 18564 23044
rect 18564 23024 18566 23044
rect 17956 20698 18012 20700
rect 18036 20698 18092 20700
rect 18116 20698 18172 20700
rect 18196 20698 18252 20700
rect 17956 20646 18002 20698
rect 18002 20646 18012 20698
rect 18036 20646 18066 20698
rect 18066 20646 18078 20698
rect 18078 20646 18092 20698
rect 18116 20646 18130 20698
rect 18130 20646 18142 20698
rect 18142 20646 18172 20698
rect 18196 20646 18206 20698
rect 18206 20646 18252 20698
rect 17956 20644 18012 20646
rect 18036 20644 18092 20646
rect 18116 20644 18172 20646
rect 18196 20644 18252 20646
rect 18418 20576 18474 20632
rect 17956 19610 18012 19612
rect 18036 19610 18092 19612
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 17956 19558 18002 19610
rect 18002 19558 18012 19610
rect 18036 19558 18066 19610
rect 18066 19558 18078 19610
rect 18078 19558 18092 19610
rect 18116 19558 18130 19610
rect 18130 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 17956 19556 18012 19558
rect 18036 19556 18092 19558
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 17774 17992 17830 18048
rect 17956 18522 18012 18524
rect 18036 18522 18092 18524
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 17956 18470 18002 18522
rect 18002 18470 18012 18522
rect 18036 18470 18066 18522
rect 18066 18470 18078 18522
rect 18078 18470 18092 18522
rect 18116 18470 18130 18522
rect 18130 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 17956 18468 18012 18470
rect 18036 18468 18092 18470
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 18234 18264 18290 18320
rect 17956 17434 18012 17436
rect 18036 17434 18092 17436
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 17956 17382 18002 17434
rect 18002 17382 18012 17434
rect 18036 17382 18066 17434
rect 18066 17382 18078 17434
rect 18078 17382 18092 17434
rect 18116 17382 18130 17434
rect 18130 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 17956 17380 18012 17382
rect 18036 17380 18092 17382
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 17498 13912 17554 13968
rect 17590 10648 17646 10704
rect 17956 16346 18012 16348
rect 18036 16346 18092 16348
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 17956 16294 18002 16346
rect 18002 16294 18012 16346
rect 18036 16294 18066 16346
rect 18066 16294 18078 16346
rect 18078 16294 18092 16346
rect 18116 16294 18130 16346
rect 18130 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 17956 16292 18012 16294
rect 18036 16292 18092 16294
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 17956 15258 18012 15260
rect 18036 15258 18092 15260
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 17956 15206 18002 15258
rect 18002 15206 18012 15258
rect 18036 15206 18066 15258
rect 18066 15206 18078 15258
rect 18078 15206 18092 15258
rect 18116 15206 18130 15258
rect 18130 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 17956 15204 18012 15206
rect 18036 15204 18092 15206
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 17956 14170 18012 14172
rect 18036 14170 18092 14172
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 17956 14118 18002 14170
rect 18002 14118 18012 14170
rect 18036 14118 18066 14170
rect 18066 14118 18078 14170
rect 18078 14118 18092 14170
rect 18116 14118 18130 14170
rect 18130 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 17956 14116 18012 14118
rect 18036 14116 18092 14118
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 17956 13082 18012 13084
rect 18036 13082 18092 13084
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 17956 13030 18002 13082
rect 18002 13030 18012 13082
rect 18036 13030 18066 13082
rect 18066 13030 18078 13082
rect 18078 13030 18092 13082
rect 18116 13030 18130 13082
rect 18130 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 17956 13028 18012 13030
rect 18036 13028 18092 13030
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 17956 11994 18012 11996
rect 18036 11994 18092 11996
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 17956 11942 18002 11994
rect 18002 11942 18012 11994
rect 18036 11942 18066 11994
rect 18066 11942 18078 11994
rect 18078 11942 18092 11994
rect 18116 11942 18130 11994
rect 18130 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 17956 11940 18012 11942
rect 18036 11940 18092 11942
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 19154 23432 19210 23488
rect 18602 17312 18658 17368
rect 20166 25064 20222 25120
rect 19522 22616 19578 22672
rect 19430 22500 19486 22536
rect 19430 22480 19432 22500
rect 19432 22480 19484 22500
rect 19484 22480 19486 22500
rect 19798 23704 19854 23760
rect 19982 23432 20038 23488
rect 19614 22344 19670 22400
rect 19430 21664 19486 21720
rect 19430 20984 19486 21040
rect 19614 21392 19670 21448
rect 19522 20712 19578 20768
rect 19154 19216 19210 19272
rect 18878 14048 18934 14104
rect 18878 13776 18934 13832
rect 18326 11056 18382 11112
rect 17956 10906 18012 10908
rect 18036 10906 18092 10908
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 17956 10854 18002 10906
rect 18002 10854 18012 10906
rect 18036 10854 18066 10906
rect 18066 10854 18078 10906
rect 18078 10854 18092 10906
rect 18116 10854 18130 10906
rect 18130 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 17956 10852 18012 10854
rect 18036 10852 18092 10854
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 17956 9818 18012 9820
rect 18036 9818 18092 9820
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 17956 9766 18002 9818
rect 18002 9766 18012 9818
rect 18036 9766 18066 9818
rect 18066 9766 18078 9818
rect 18078 9766 18092 9818
rect 18116 9766 18130 9818
rect 18130 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 17956 9764 18012 9766
rect 18036 9764 18092 9766
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 17956 8730 18012 8732
rect 18036 8730 18092 8732
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 17956 8678 18002 8730
rect 18002 8678 18012 8730
rect 18036 8678 18066 8730
rect 18066 8678 18078 8730
rect 18078 8678 18092 8730
rect 18116 8678 18130 8730
rect 18130 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 17956 8676 18012 8678
rect 18036 8676 18092 8678
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 17956 7642 18012 7644
rect 18036 7642 18092 7644
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 17956 7590 18002 7642
rect 18002 7590 18012 7642
rect 18036 7590 18066 7642
rect 18066 7590 18078 7642
rect 18078 7590 18092 7642
rect 18116 7590 18130 7642
rect 18130 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 17956 7588 18012 7590
rect 18036 7588 18092 7590
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 17956 6554 18012 6556
rect 18036 6554 18092 6556
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 17956 6502 18002 6554
rect 18002 6502 18012 6554
rect 18036 6502 18066 6554
rect 18066 6502 18078 6554
rect 18078 6502 18092 6554
rect 18116 6502 18130 6554
rect 18130 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 17956 6500 18012 6502
rect 18036 6500 18092 6502
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 2956 6010 3012 6012
rect 3036 6010 3092 6012
rect 3116 6010 3172 6012
rect 3196 6010 3252 6012
rect 2956 5958 3002 6010
rect 3002 5958 3012 6010
rect 3036 5958 3066 6010
rect 3066 5958 3078 6010
rect 3078 5958 3092 6010
rect 3116 5958 3130 6010
rect 3130 5958 3142 6010
rect 3142 5958 3172 6010
rect 3196 5958 3206 6010
rect 3206 5958 3252 6010
rect 2956 5956 3012 5958
rect 3036 5956 3092 5958
rect 3116 5956 3172 5958
rect 3196 5956 3252 5958
rect 2956 4922 3012 4924
rect 3036 4922 3092 4924
rect 3116 4922 3172 4924
rect 3196 4922 3252 4924
rect 2956 4870 3002 4922
rect 3002 4870 3012 4922
rect 3036 4870 3066 4922
rect 3066 4870 3078 4922
rect 3078 4870 3092 4922
rect 3116 4870 3130 4922
rect 3130 4870 3142 4922
rect 3142 4870 3172 4922
rect 3196 4870 3206 4922
rect 3206 4870 3252 4922
rect 2956 4868 3012 4870
rect 3036 4868 3092 4870
rect 3116 4868 3172 4870
rect 3196 4868 3252 4870
rect 2956 3834 3012 3836
rect 3036 3834 3092 3836
rect 3116 3834 3172 3836
rect 3196 3834 3252 3836
rect 2956 3782 3002 3834
rect 3002 3782 3012 3834
rect 3036 3782 3066 3834
rect 3066 3782 3078 3834
rect 3078 3782 3092 3834
rect 3116 3782 3130 3834
rect 3130 3782 3142 3834
rect 3142 3782 3172 3834
rect 3196 3782 3206 3834
rect 3206 3782 3252 3834
rect 2956 3780 3012 3782
rect 3036 3780 3092 3782
rect 3116 3780 3172 3782
rect 3196 3780 3252 3782
rect 12956 6010 13012 6012
rect 13036 6010 13092 6012
rect 13116 6010 13172 6012
rect 13196 6010 13252 6012
rect 12956 5958 13002 6010
rect 13002 5958 13012 6010
rect 13036 5958 13066 6010
rect 13066 5958 13078 6010
rect 13078 5958 13092 6010
rect 13116 5958 13130 6010
rect 13130 5958 13142 6010
rect 13142 5958 13172 6010
rect 13196 5958 13206 6010
rect 13206 5958 13252 6010
rect 12956 5956 13012 5958
rect 13036 5956 13092 5958
rect 13116 5956 13172 5958
rect 13196 5956 13252 5958
rect 7956 5466 8012 5468
rect 8036 5466 8092 5468
rect 8116 5466 8172 5468
rect 8196 5466 8252 5468
rect 7956 5414 8002 5466
rect 8002 5414 8012 5466
rect 8036 5414 8066 5466
rect 8066 5414 8078 5466
rect 8078 5414 8092 5466
rect 8116 5414 8130 5466
rect 8130 5414 8142 5466
rect 8142 5414 8172 5466
rect 8196 5414 8206 5466
rect 8206 5414 8252 5466
rect 7956 5412 8012 5414
rect 8036 5412 8092 5414
rect 8116 5412 8172 5414
rect 8196 5412 8252 5414
rect 17956 5466 18012 5468
rect 18036 5466 18092 5468
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 17956 5414 18002 5466
rect 18002 5414 18012 5466
rect 18036 5414 18066 5466
rect 18066 5414 18078 5466
rect 18078 5414 18092 5466
rect 18116 5414 18130 5466
rect 18130 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 17956 5412 18012 5414
rect 18036 5412 18092 5414
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 12956 4922 13012 4924
rect 13036 4922 13092 4924
rect 13116 4922 13172 4924
rect 13196 4922 13252 4924
rect 12956 4870 13002 4922
rect 13002 4870 13012 4922
rect 13036 4870 13066 4922
rect 13066 4870 13078 4922
rect 13078 4870 13092 4922
rect 13116 4870 13130 4922
rect 13130 4870 13142 4922
rect 13142 4870 13172 4922
rect 13196 4870 13206 4922
rect 13206 4870 13252 4922
rect 12956 4868 13012 4870
rect 13036 4868 13092 4870
rect 13116 4868 13172 4870
rect 13196 4868 13252 4870
rect 7956 4378 8012 4380
rect 8036 4378 8092 4380
rect 8116 4378 8172 4380
rect 8196 4378 8252 4380
rect 7956 4326 8002 4378
rect 8002 4326 8012 4378
rect 8036 4326 8066 4378
rect 8066 4326 8078 4378
rect 8078 4326 8092 4378
rect 8116 4326 8130 4378
rect 8130 4326 8142 4378
rect 8142 4326 8172 4378
rect 8196 4326 8206 4378
rect 8206 4326 8252 4378
rect 7956 4324 8012 4326
rect 8036 4324 8092 4326
rect 8116 4324 8172 4326
rect 8196 4324 8252 4326
rect 17956 4378 18012 4380
rect 18036 4378 18092 4380
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 17956 4326 18002 4378
rect 18002 4326 18012 4378
rect 18036 4326 18066 4378
rect 18066 4326 18078 4378
rect 18078 4326 18092 4378
rect 18116 4326 18130 4378
rect 18130 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 17956 4324 18012 4326
rect 18036 4324 18092 4326
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 19338 19760 19394 19816
rect 19522 19352 19578 19408
rect 19338 18264 19394 18320
rect 19246 16496 19302 16552
rect 19522 18400 19578 18456
rect 19614 17856 19670 17912
rect 19430 14864 19486 14920
rect 19062 13368 19118 13424
rect 19154 12280 19210 12336
rect 19798 18264 19854 18320
rect 19706 17040 19762 17096
rect 19706 14456 19762 14512
rect 20258 21800 20314 21856
rect 21270 26288 21326 26344
rect 20810 24792 20866 24848
rect 20442 23024 20498 23080
rect 20534 22072 20590 22128
rect 20350 21664 20406 21720
rect 20442 21528 20498 21584
rect 20258 21256 20314 21312
rect 20350 20984 20406 21040
rect 20810 20712 20866 20768
rect 21178 22072 21234 22128
rect 21178 21256 21234 21312
rect 20442 20032 20498 20088
rect 20350 15408 20406 15464
rect 20258 14728 20314 14784
rect 20166 14592 20222 14648
rect 20994 20168 21050 20224
rect 20626 18300 20628 18320
rect 20628 18300 20680 18320
rect 20680 18300 20682 18320
rect 20626 18264 20682 18300
rect 21086 19896 21142 19952
rect 20810 18400 20866 18456
rect 20718 16904 20774 16960
rect 20350 13368 20406 13424
rect 19430 11056 19486 11112
rect 19338 9444 19394 9480
rect 19338 9424 19340 9444
rect 19340 9424 19392 9444
rect 19392 9424 19394 9444
rect 19706 8356 19762 8392
rect 19706 8336 19708 8356
rect 19708 8336 19760 8356
rect 19760 8336 19762 8356
rect 12956 3834 13012 3836
rect 13036 3834 13092 3836
rect 13116 3834 13172 3836
rect 13196 3834 13252 3836
rect 12956 3782 13002 3834
rect 13002 3782 13012 3834
rect 13036 3782 13066 3834
rect 13066 3782 13078 3834
rect 13078 3782 13092 3834
rect 13116 3782 13130 3834
rect 13130 3782 13142 3834
rect 13142 3782 13172 3834
rect 13196 3782 13206 3834
rect 13206 3782 13252 3834
rect 12956 3780 13012 3782
rect 13036 3780 13092 3782
rect 13116 3780 13172 3782
rect 13196 3780 13252 3782
rect 7956 3290 8012 3292
rect 8036 3290 8092 3292
rect 8116 3290 8172 3292
rect 8196 3290 8252 3292
rect 7956 3238 8002 3290
rect 8002 3238 8012 3290
rect 8036 3238 8066 3290
rect 8066 3238 8078 3290
rect 8078 3238 8092 3290
rect 8116 3238 8130 3290
rect 8130 3238 8142 3290
rect 8142 3238 8172 3290
rect 8196 3238 8206 3290
rect 8206 3238 8252 3290
rect 7956 3236 8012 3238
rect 8036 3236 8092 3238
rect 8116 3236 8172 3238
rect 8196 3236 8252 3238
rect 17956 3290 18012 3292
rect 18036 3290 18092 3292
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 17956 3238 18002 3290
rect 18002 3238 18012 3290
rect 18036 3238 18066 3290
rect 18066 3238 18078 3290
rect 18078 3238 18092 3290
rect 18116 3238 18130 3290
rect 18130 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 17956 3236 18012 3238
rect 18036 3236 18092 3238
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 20994 18400 21050 18456
rect 21454 22752 21510 22808
rect 22098 23568 22154 23624
rect 21362 21120 21418 21176
rect 21270 20032 21326 20088
rect 21178 17992 21234 18048
rect 21086 17720 21142 17776
rect 21086 17448 21142 17504
rect 20718 10260 20774 10296
rect 20718 10240 20720 10260
rect 20720 10240 20772 10260
rect 20772 10240 20774 10260
rect 20718 9696 20774 9752
rect 20534 7928 20590 7984
rect 20258 5616 20314 5672
rect 2956 2746 3012 2748
rect 3036 2746 3092 2748
rect 3116 2746 3172 2748
rect 3196 2746 3252 2748
rect 2956 2694 3002 2746
rect 3002 2694 3012 2746
rect 3036 2694 3066 2746
rect 3066 2694 3078 2746
rect 3078 2694 3092 2746
rect 3116 2694 3130 2746
rect 3130 2694 3142 2746
rect 3142 2694 3172 2746
rect 3196 2694 3206 2746
rect 3206 2694 3252 2746
rect 2956 2692 3012 2694
rect 3036 2692 3092 2694
rect 3116 2692 3172 2694
rect 3196 2692 3252 2694
rect 12956 2746 13012 2748
rect 13036 2746 13092 2748
rect 13116 2746 13172 2748
rect 13196 2746 13252 2748
rect 12956 2694 13002 2746
rect 13002 2694 13012 2746
rect 13036 2694 13066 2746
rect 13066 2694 13078 2746
rect 13078 2694 13092 2746
rect 13116 2694 13130 2746
rect 13130 2694 13142 2746
rect 13142 2694 13172 2746
rect 13196 2694 13206 2746
rect 13206 2694 13252 2746
rect 12956 2692 13012 2694
rect 13036 2692 13092 2694
rect 13116 2692 13172 2694
rect 13196 2692 13252 2694
rect 7956 2202 8012 2204
rect 8036 2202 8092 2204
rect 8116 2202 8172 2204
rect 8196 2202 8252 2204
rect 7956 2150 8002 2202
rect 8002 2150 8012 2202
rect 8036 2150 8066 2202
rect 8066 2150 8078 2202
rect 8078 2150 8092 2202
rect 8116 2150 8130 2202
rect 8130 2150 8142 2202
rect 8142 2150 8172 2202
rect 8196 2150 8206 2202
rect 8206 2150 8252 2202
rect 7956 2148 8012 2150
rect 8036 2148 8092 2150
rect 8116 2148 8172 2150
rect 8196 2148 8252 2150
rect 17956 2202 18012 2204
rect 18036 2202 18092 2204
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 17956 2150 18002 2202
rect 18002 2150 18012 2202
rect 18036 2150 18066 2202
rect 18066 2150 18078 2202
rect 18078 2150 18092 2202
rect 18116 2150 18130 2202
rect 18130 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 17956 2148 18012 2150
rect 18036 2148 18092 2150
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 21730 22072 21786 22128
rect 21638 20712 21694 20768
rect 21546 19080 21602 19136
rect 21638 18264 21694 18320
rect 21638 17720 21694 17776
rect 21638 16632 21694 16688
rect 22190 21664 22246 21720
rect 22190 21392 22246 21448
rect 22006 21120 22062 21176
rect 21822 20440 21878 20496
rect 22190 19216 22246 19272
rect 21914 18536 21970 18592
rect 22098 18536 22154 18592
rect 21914 17584 21970 17640
rect 21822 17040 21878 17096
rect 21638 15272 21694 15328
rect 21270 9696 21326 9752
rect 21270 7792 21326 7848
rect 22466 20984 22522 21040
rect 25778 26424 25834 26480
rect 22834 26016 22890 26072
rect 23202 25608 23258 25664
rect 22956 24506 23012 24508
rect 23036 24506 23092 24508
rect 23116 24506 23172 24508
rect 23196 24506 23252 24508
rect 22956 24454 23002 24506
rect 23002 24454 23012 24506
rect 23036 24454 23066 24506
rect 23066 24454 23078 24506
rect 23078 24454 23092 24506
rect 23116 24454 23130 24506
rect 23130 24454 23142 24506
rect 23142 24454 23172 24506
rect 23196 24454 23206 24506
rect 23206 24454 23252 24506
rect 22956 24452 23012 24454
rect 23036 24452 23092 24454
rect 23116 24452 23172 24454
rect 23196 24452 23252 24454
rect 22956 23418 23012 23420
rect 23036 23418 23092 23420
rect 23116 23418 23172 23420
rect 23196 23418 23252 23420
rect 22956 23366 23002 23418
rect 23002 23366 23012 23418
rect 23036 23366 23066 23418
rect 23066 23366 23078 23418
rect 23078 23366 23092 23418
rect 23116 23366 23130 23418
rect 23130 23366 23142 23418
rect 23142 23366 23172 23418
rect 23196 23366 23206 23418
rect 23206 23366 23252 23418
rect 22956 23364 23012 23366
rect 23036 23364 23092 23366
rect 23116 23364 23172 23366
rect 23196 23364 23252 23366
rect 22956 22330 23012 22332
rect 23036 22330 23092 22332
rect 23116 22330 23172 22332
rect 23196 22330 23252 22332
rect 22956 22278 23002 22330
rect 23002 22278 23012 22330
rect 23036 22278 23066 22330
rect 23066 22278 23078 22330
rect 23078 22278 23092 22330
rect 23116 22278 23130 22330
rect 23130 22278 23142 22330
rect 23142 22278 23172 22330
rect 23196 22278 23206 22330
rect 23206 22278 23252 22330
rect 22956 22276 23012 22278
rect 23036 22276 23092 22278
rect 23116 22276 23172 22278
rect 23196 22276 23252 22278
rect 22650 21936 22706 21992
rect 22650 21800 22706 21856
rect 23478 21664 23534 21720
rect 23386 21528 23442 21584
rect 22650 21256 22706 21312
rect 22558 19080 22614 19136
rect 22098 13912 22154 13968
rect 22282 15136 22338 15192
rect 22282 14048 22338 14104
rect 22282 13812 22284 13832
rect 22284 13812 22336 13832
rect 22336 13812 22338 13832
rect 22282 13776 22338 13812
rect 22466 18164 22468 18184
rect 22468 18164 22520 18184
rect 22520 18164 22522 18184
rect 22466 18128 22522 18164
rect 22956 21242 23012 21244
rect 23036 21242 23092 21244
rect 23116 21242 23172 21244
rect 23196 21242 23252 21244
rect 22956 21190 23002 21242
rect 23002 21190 23012 21242
rect 23036 21190 23066 21242
rect 23066 21190 23078 21242
rect 23078 21190 23092 21242
rect 23116 21190 23130 21242
rect 23130 21190 23142 21242
rect 23142 21190 23172 21242
rect 23196 21190 23206 21242
rect 23206 21190 23252 21242
rect 22956 21188 23012 21190
rect 23036 21188 23092 21190
rect 23116 21188 23172 21190
rect 23196 21188 23252 21190
rect 23202 20884 23204 20904
rect 23204 20884 23256 20904
rect 23256 20884 23258 20904
rect 23202 20848 23258 20884
rect 23386 21120 23442 21176
rect 22742 18692 22798 18728
rect 22742 18672 22744 18692
rect 22744 18672 22796 18692
rect 22796 18672 22798 18692
rect 22466 16632 22522 16688
rect 22956 20154 23012 20156
rect 23036 20154 23092 20156
rect 23116 20154 23172 20156
rect 23196 20154 23252 20156
rect 22956 20102 23002 20154
rect 23002 20102 23012 20154
rect 23036 20102 23066 20154
rect 23066 20102 23078 20154
rect 23078 20102 23092 20154
rect 23116 20102 23130 20154
rect 23130 20102 23142 20154
rect 23142 20102 23172 20154
rect 23196 20102 23206 20154
rect 23206 20102 23252 20154
rect 22956 20100 23012 20102
rect 23036 20100 23092 20102
rect 23116 20100 23172 20102
rect 23196 20100 23252 20102
rect 23018 19896 23074 19952
rect 23386 19488 23442 19544
rect 22956 19066 23012 19068
rect 23036 19066 23092 19068
rect 23116 19066 23172 19068
rect 23196 19066 23252 19068
rect 22956 19014 23002 19066
rect 23002 19014 23012 19066
rect 23036 19014 23066 19066
rect 23066 19014 23078 19066
rect 23078 19014 23092 19066
rect 23116 19014 23130 19066
rect 23130 19014 23142 19066
rect 23142 19014 23172 19066
rect 23196 19014 23206 19066
rect 23206 19014 23252 19066
rect 22956 19012 23012 19014
rect 23036 19012 23092 19014
rect 23116 19012 23172 19014
rect 23196 19012 23252 19014
rect 23018 18672 23074 18728
rect 22926 18264 22982 18320
rect 23386 18400 23442 18456
rect 23478 18128 23534 18184
rect 22956 17978 23012 17980
rect 23036 17978 23092 17980
rect 23116 17978 23172 17980
rect 23196 17978 23252 17980
rect 22956 17926 23002 17978
rect 23002 17926 23012 17978
rect 23036 17926 23066 17978
rect 23066 17926 23078 17978
rect 23078 17926 23092 17978
rect 23116 17926 23130 17978
rect 23130 17926 23142 17978
rect 23142 17926 23172 17978
rect 23196 17926 23206 17978
rect 23206 17926 23252 17978
rect 22956 17924 23012 17926
rect 23036 17924 23092 17926
rect 23116 17924 23172 17926
rect 23196 17924 23252 17926
rect 22956 16890 23012 16892
rect 23036 16890 23092 16892
rect 23116 16890 23172 16892
rect 23196 16890 23252 16892
rect 22956 16838 23002 16890
rect 23002 16838 23012 16890
rect 23036 16838 23066 16890
rect 23066 16838 23078 16890
rect 23078 16838 23092 16890
rect 23116 16838 23130 16890
rect 23130 16838 23142 16890
rect 23142 16838 23172 16890
rect 23196 16838 23206 16890
rect 23206 16838 23252 16890
rect 22956 16836 23012 16838
rect 23036 16836 23092 16838
rect 23116 16836 23172 16838
rect 23196 16836 23252 16838
rect 22956 15802 23012 15804
rect 23036 15802 23092 15804
rect 23116 15802 23172 15804
rect 23196 15802 23252 15804
rect 22956 15750 23002 15802
rect 23002 15750 23012 15802
rect 23036 15750 23066 15802
rect 23066 15750 23078 15802
rect 23078 15750 23092 15802
rect 23116 15750 23130 15802
rect 23130 15750 23142 15802
rect 23142 15750 23172 15802
rect 23196 15750 23206 15802
rect 23206 15750 23252 15802
rect 22956 15748 23012 15750
rect 23036 15748 23092 15750
rect 23116 15748 23172 15750
rect 23196 15748 23252 15750
rect 22374 13368 22430 13424
rect 22006 8336 22062 8392
rect 22190 6840 22246 6896
rect 23202 15136 23258 15192
rect 22956 14714 23012 14716
rect 23036 14714 23092 14716
rect 23116 14714 23172 14716
rect 23196 14714 23252 14716
rect 22956 14662 23002 14714
rect 23002 14662 23012 14714
rect 23036 14662 23066 14714
rect 23066 14662 23078 14714
rect 23078 14662 23092 14714
rect 23116 14662 23130 14714
rect 23130 14662 23142 14714
rect 23142 14662 23172 14714
rect 23196 14662 23206 14714
rect 23206 14662 23252 14714
rect 22956 14660 23012 14662
rect 23036 14660 23092 14662
rect 23116 14660 23172 14662
rect 23196 14660 23252 14662
rect 22834 14184 22890 14240
rect 22956 13626 23012 13628
rect 23036 13626 23092 13628
rect 23116 13626 23172 13628
rect 23196 13626 23252 13628
rect 22956 13574 23002 13626
rect 23002 13574 23012 13626
rect 23036 13574 23066 13626
rect 23066 13574 23078 13626
rect 23078 13574 23092 13626
rect 23116 13574 23130 13626
rect 23130 13574 23142 13626
rect 23142 13574 23172 13626
rect 23196 13574 23206 13626
rect 23206 13574 23252 13626
rect 22956 13572 23012 13574
rect 23036 13572 23092 13574
rect 23116 13572 23172 13574
rect 23196 13572 23252 13574
rect 22834 12960 22890 13016
rect 22956 12538 23012 12540
rect 23036 12538 23092 12540
rect 23116 12538 23172 12540
rect 23196 12538 23252 12540
rect 22956 12486 23002 12538
rect 23002 12486 23012 12538
rect 23036 12486 23066 12538
rect 23066 12486 23078 12538
rect 23078 12486 23092 12538
rect 23116 12486 23130 12538
rect 23130 12486 23142 12538
rect 23142 12486 23172 12538
rect 23196 12486 23206 12538
rect 23206 12486 23252 12538
rect 22956 12484 23012 12486
rect 23036 12484 23092 12486
rect 23116 12484 23172 12486
rect 23196 12484 23252 12486
rect 22956 11450 23012 11452
rect 23036 11450 23092 11452
rect 23116 11450 23172 11452
rect 23196 11450 23252 11452
rect 22956 11398 23002 11450
rect 23002 11398 23012 11450
rect 23036 11398 23066 11450
rect 23066 11398 23078 11450
rect 23078 11398 23092 11450
rect 23116 11398 23130 11450
rect 23130 11398 23142 11450
rect 23142 11398 23172 11450
rect 23196 11398 23206 11450
rect 23206 11398 23252 11450
rect 22956 11396 23012 11398
rect 23036 11396 23092 11398
rect 23116 11396 23172 11398
rect 23196 11396 23252 11398
rect 23386 14864 23442 14920
rect 23386 14592 23442 14648
rect 24030 21664 24086 21720
rect 23938 19216 23994 19272
rect 22956 10362 23012 10364
rect 23036 10362 23092 10364
rect 23116 10362 23172 10364
rect 23196 10362 23252 10364
rect 22956 10310 23002 10362
rect 23002 10310 23012 10362
rect 23036 10310 23066 10362
rect 23066 10310 23078 10362
rect 23078 10310 23092 10362
rect 23116 10310 23130 10362
rect 23130 10310 23142 10362
rect 23142 10310 23172 10362
rect 23196 10310 23206 10362
rect 23206 10310 23252 10362
rect 22956 10308 23012 10310
rect 23036 10308 23092 10310
rect 23116 10308 23172 10310
rect 23196 10308 23252 10310
rect 23294 9696 23350 9752
rect 22956 9274 23012 9276
rect 23036 9274 23092 9276
rect 23116 9274 23172 9276
rect 23196 9274 23252 9276
rect 22956 9222 23002 9274
rect 23002 9222 23012 9274
rect 23036 9222 23066 9274
rect 23066 9222 23078 9274
rect 23078 9222 23092 9274
rect 23116 9222 23130 9274
rect 23130 9222 23142 9274
rect 23142 9222 23172 9274
rect 23196 9222 23206 9274
rect 23206 9222 23252 9274
rect 22956 9220 23012 9222
rect 23036 9220 23092 9222
rect 23116 9220 23172 9222
rect 23196 9220 23252 9222
rect 22956 8186 23012 8188
rect 23036 8186 23092 8188
rect 23116 8186 23172 8188
rect 23196 8186 23252 8188
rect 22956 8134 23002 8186
rect 23002 8134 23012 8186
rect 23036 8134 23066 8186
rect 23066 8134 23078 8186
rect 23078 8134 23092 8186
rect 23116 8134 23130 8186
rect 23130 8134 23142 8186
rect 23142 8134 23172 8186
rect 23196 8134 23206 8186
rect 23206 8134 23252 8186
rect 22956 8132 23012 8134
rect 23036 8132 23092 8134
rect 23116 8132 23172 8134
rect 23196 8132 23252 8134
rect 22956 7098 23012 7100
rect 23036 7098 23092 7100
rect 23116 7098 23172 7100
rect 23196 7098 23252 7100
rect 22956 7046 23002 7098
rect 23002 7046 23012 7098
rect 23036 7046 23066 7098
rect 23066 7046 23078 7098
rect 23078 7046 23092 7098
rect 23116 7046 23130 7098
rect 23130 7046 23142 7098
rect 23142 7046 23172 7098
rect 23196 7046 23206 7098
rect 23206 7046 23252 7098
rect 22956 7044 23012 7046
rect 23036 7044 23092 7046
rect 23116 7044 23172 7046
rect 23196 7044 23252 7046
rect 22956 6010 23012 6012
rect 23036 6010 23092 6012
rect 23116 6010 23172 6012
rect 23196 6010 23252 6012
rect 22956 5958 23002 6010
rect 23002 5958 23012 6010
rect 23036 5958 23066 6010
rect 23066 5958 23078 6010
rect 23078 5958 23092 6010
rect 23116 5958 23130 6010
rect 23130 5958 23142 6010
rect 23142 5958 23172 6010
rect 23196 5958 23206 6010
rect 23206 5958 23252 6010
rect 22956 5956 23012 5958
rect 23036 5956 23092 5958
rect 23116 5956 23172 5958
rect 23196 5956 23252 5958
rect 22956 4922 23012 4924
rect 23036 4922 23092 4924
rect 23116 4922 23172 4924
rect 23196 4922 23252 4924
rect 22956 4870 23002 4922
rect 23002 4870 23012 4922
rect 23036 4870 23066 4922
rect 23066 4870 23078 4922
rect 23078 4870 23092 4922
rect 23116 4870 23130 4922
rect 23130 4870 23142 4922
rect 23142 4870 23172 4922
rect 23196 4870 23206 4922
rect 23206 4870 23252 4922
rect 22956 4868 23012 4870
rect 23036 4868 23092 4870
rect 23116 4868 23172 4870
rect 23196 4868 23252 4870
rect 24214 19760 24270 19816
rect 24398 21528 24454 21584
rect 24398 20984 24454 21040
rect 25134 25200 25190 25256
rect 25042 24268 25098 24304
rect 25042 24248 25044 24268
rect 25044 24248 25096 24268
rect 25096 24248 25098 24268
rect 24582 22480 24638 22536
rect 24306 18536 24362 18592
rect 24582 19660 24584 19680
rect 24584 19660 24636 19680
rect 24636 19660 24638 19680
rect 24582 19624 24638 19660
rect 24858 19352 24914 19408
rect 24582 17992 24638 18048
rect 24858 17196 24914 17232
rect 24858 17176 24860 17196
rect 24860 17176 24912 17196
rect 24912 17176 24914 17196
rect 24858 16224 24914 16280
rect 24674 16108 24730 16144
rect 24674 16088 24676 16108
rect 24676 16088 24728 16108
rect 24728 16088 24730 16108
rect 24674 15816 24730 15872
rect 24858 12824 24914 12880
rect 24674 12144 24730 12200
rect 24582 11600 24638 11656
rect 24858 11772 24860 11792
rect 24860 11772 24912 11792
rect 24912 11772 24914 11792
rect 24858 11736 24914 11772
rect 24858 11328 24914 11384
rect 24766 10920 24822 10976
rect 24582 10104 24638 10160
rect 24858 10512 24914 10568
rect 24858 9288 24914 9344
rect 24674 8880 24730 8936
rect 22956 3834 23012 3836
rect 23036 3834 23092 3836
rect 23116 3834 23172 3836
rect 23196 3834 23252 3836
rect 22956 3782 23002 3834
rect 23002 3782 23012 3834
rect 23036 3782 23066 3834
rect 23066 3782 23078 3834
rect 23078 3782 23092 3834
rect 23116 3782 23130 3834
rect 23130 3782 23142 3834
rect 23142 3782 23172 3834
rect 23196 3782 23206 3834
rect 23206 3782 23252 3834
rect 22956 3780 23012 3782
rect 23036 3780 23092 3782
rect 23116 3780 23172 3782
rect 23196 3780 23252 3782
rect 24858 8508 24860 8528
rect 24860 8508 24912 8528
rect 24912 8508 24914 8528
rect 24858 8472 24914 8508
rect 24950 8064 25006 8120
rect 24766 7656 24822 7712
rect 24674 6432 24730 6488
rect 25134 12552 25190 12608
rect 25502 19216 25558 19272
rect 24858 7248 24914 7304
rect 25870 15988 25872 16008
rect 25872 15988 25924 16008
rect 25924 15988 25926 16008
rect 25870 15952 25926 15988
rect 24858 6860 24914 6896
rect 24858 6840 24860 6860
rect 24860 6840 24912 6860
rect 24912 6840 24914 6860
rect 24858 6024 24914 6080
rect 24950 5636 25006 5672
rect 24950 5616 24952 5636
rect 24952 5616 25004 5636
rect 25004 5616 25006 5636
rect 24766 5208 24822 5264
rect 24858 4800 24914 4856
rect 24950 4392 25006 4448
rect 25134 3984 25190 4040
rect 24950 3576 25006 3632
rect 22956 2746 23012 2748
rect 23036 2746 23092 2748
rect 23116 2746 23172 2748
rect 23196 2746 23252 2748
rect 22956 2694 23002 2746
rect 23002 2694 23012 2746
rect 23036 2694 23066 2746
rect 23066 2694 23078 2746
rect 23078 2694 23092 2746
rect 23116 2694 23130 2746
rect 23130 2694 23142 2746
rect 23142 2694 23172 2746
rect 23196 2694 23206 2746
rect 23206 2694 23252 2746
rect 22956 2692 23012 2694
rect 23036 2692 23092 2694
rect 23116 2692 23172 2694
rect 23196 2692 23252 2694
rect 24950 3168 25006 3224
rect 24858 2760 24914 2816
rect 24950 2372 25006 2408
rect 24950 2352 24952 2372
rect 24952 2352 25004 2372
rect 25004 2352 25006 2372
rect 22190 1944 22246 2000
rect 22098 1536 22154 1592
rect 22098 1128 22154 1184
rect 26054 14320 26110 14376
rect 25042 720 25098 776
rect 23386 312 23442 368
<< metal3 >>
rect 25773 26482 25839 26485
rect 26200 26482 27000 26512
rect 25773 26480 27000 26482
rect 25773 26424 25778 26480
rect 25834 26424 27000 26480
rect 25773 26422 27000 26424
rect 25773 26419 25839 26422
rect 26200 26392 27000 26422
rect 21265 26346 21331 26349
rect 12390 26344 21331 26346
rect 12390 26288 21270 26344
rect 21326 26288 21331 26344
rect 12390 26286 21331 26288
rect 4889 26210 4955 26213
rect 12390 26210 12450 26286
rect 21265 26283 21331 26286
rect 4889 26208 12450 26210
rect 4889 26152 4894 26208
rect 4950 26152 12450 26208
rect 4889 26150 12450 26152
rect 4889 26147 4955 26150
rect 6494 26012 6500 26076
rect 6564 26074 6570 26076
rect 18965 26074 19031 26077
rect 6564 26072 19031 26074
rect 6564 26016 18970 26072
rect 19026 26016 19031 26072
rect 6564 26014 19031 26016
rect 6564 26012 6570 26014
rect 18965 26011 19031 26014
rect 22829 26074 22895 26077
rect 26200 26074 27000 26104
rect 22829 26072 27000 26074
rect 22829 26016 22834 26072
rect 22890 26016 27000 26072
rect 22829 26014 27000 26016
rect 22829 26011 22895 26014
rect 26200 25984 27000 26014
rect 0 25938 800 25968
rect 3693 25938 3759 25941
rect 0 25936 3759 25938
rect 0 25880 3698 25936
rect 3754 25880 3759 25936
rect 0 25878 3759 25880
rect 0 25848 800 25878
rect 3693 25875 3759 25878
rect 23197 25666 23263 25669
rect 26200 25666 27000 25696
rect 23197 25664 27000 25666
rect 23197 25608 23202 25664
rect 23258 25608 27000 25664
rect 23197 25606 27000 25608
rect 23197 25603 23263 25606
rect 26200 25576 27000 25606
rect 25129 25258 25195 25261
rect 26200 25258 27000 25288
rect 25129 25256 27000 25258
rect 25129 25200 25134 25256
rect 25190 25200 27000 25256
rect 25129 25198 27000 25200
rect 25129 25195 25195 25198
rect 26200 25168 27000 25198
rect 6545 25122 6611 25125
rect 20161 25122 20227 25125
rect 6545 25120 20227 25122
rect 6545 25064 6550 25120
rect 6606 25064 20166 25120
rect 20222 25064 20227 25120
rect 6545 25062 20227 25064
rect 6545 25059 6611 25062
rect 20161 25059 20227 25062
rect 4797 24986 4863 24989
rect 19057 24986 19123 24989
rect 4797 24984 19123 24986
rect 4797 24928 4802 24984
rect 4858 24928 19062 24984
rect 19118 24928 19123 24984
rect 4797 24926 19123 24928
rect 4797 24923 4863 24926
rect 19057 24923 19123 24926
rect 19425 24986 19491 24989
rect 19425 24984 21098 24986
rect 19425 24928 19430 24984
rect 19486 24928 21098 24984
rect 19425 24926 21098 24928
rect 19425 24923 19491 24926
rect 0 24850 800 24880
rect 3417 24850 3483 24853
rect 0 24848 3483 24850
rect 0 24792 3422 24848
rect 3478 24792 3483 24848
rect 0 24790 3483 24792
rect 0 24760 800 24790
rect 3417 24787 3483 24790
rect 9622 24788 9628 24852
rect 9692 24850 9698 24852
rect 20805 24850 20871 24853
rect 9692 24848 20871 24850
rect 9692 24792 20810 24848
rect 20866 24792 20871 24848
rect 9692 24790 20871 24792
rect 21038 24850 21098 24926
rect 26200 24850 27000 24880
rect 21038 24790 27000 24850
rect 9692 24788 9698 24790
rect 20805 24787 20871 24790
rect 26200 24760 27000 24790
rect 8886 24652 8892 24716
rect 8956 24714 8962 24716
rect 17493 24714 17559 24717
rect 8956 24712 17559 24714
rect 8956 24656 17498 24712
rect 17554 24656 17559 24712
rect 8956 24654 17559 24656
rect 8956 24652 8962 24654
rect 17493 24651 17559 24654
rect 17677 24714 17743 24717
rect 17677 24712 24226 24714
rect 17677 24656 17682 24712
rect 17738 24656 24226 24712
rect 17677 24654 24226 24656
rect 17677 24651 17743 24654
rect 2946 24512 3262 24513
rect 2946 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3262 24512
rect 2946 24447 3262 24448
rect 12946 24512 13262 24513
rect 12946 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13262 24512
rect 12946 24447 13262 24448
rect 22946 24512 23262 24513
rect 22946 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23262 24512
rect 22946 24447 23262 24448
rect 16021 24442 16087 24445
rect 24166 24442 24226 24654
rect 26200 24442 27000 24472
rect 16021 24440 22754 24442
rect 16021 24384 16026 24440
rect 16082 24384 22754 24440
rect 16021 24382 22754 24384
rect 24166 24382 27000 24442
rect 16021 24379 16087 24382
rect 12014 24244 12020 24308
rect 12084 24306 12090 24308
rect 22694 24306 22754 24382
rect 26200 24352 27000 24382
rect 25037 24306 25103 24309
rect 12084 24246 22110 24306
rect 22694 24304 25103 24306
rect 22694 24248 25042 24304
rect 25098 24248 25103 24304
rect 22694 24246 25103 24248
rect 12084 24244 12090 24246
rect 1761 24170 1827 24173
rect 9765 24170 9831 24173
rect 1761 24168 9831 24170
rect 1761 24112 1766 24168
rect 1822 24112 9770 24168
rect 9826 24112 9831 24168
rect 1761 24110 9831 24112
rect 1761 24107 1827 24110
rect 9765 24107 9831 24110
rect 14958 24108 14964 24172
rect 15028 24170 15034 24172
rect 17953 24170 18019 24173
rect 15028 24168 18019 24170
rect 15028 24112 17958 24168
rect 18014 24112 18019 24168
rect 15028 24110 18019 24112
rect 15028 24108 15034 24110
rect 17953 24107 18019 24110
rect 10358 23972 10364 24036
rect 10428 24034 10434 24036
rect 17677 24034 17743 24037
rect 10428 24032 17743 24034
rect 10428 23976 17682 24032
rect 17738 23976 17743 24032
rect 10428 23974 17743 23976
rect 22050 24034 22110 24246
rect 25037 24243 25103 24246
rect 26200 24034 27000 24064
rect 22050 23974 27000 24034
rect 10428 23972 10434 23974
rect 17677 23971 17743 23974
rect 7946 23968 8262 23969
rect 7946 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8262 23968
rect 7946 23903 8262 23904
rect 17946 23968 18262 23969
rect 17946 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18262 23968
rect 26200 23944 27000 23974
rect 17946 23903 18262 23904
rect 16021 23898 16087 23901
rect 16246 23898 16252 23900
rect 16021 23896 16252 23898
rect 16021 23840 16026 23896
rect 16082 23840 16252 23896
rect 16021 23838 16252 23840
rect 16021 23835 16087 23838
rect 16246 23836 16252 23838
rect 16316 23836 16322 23900
rect 0 23762 800 23792
rect 1117 23762 1183 23765
rect 0 23760 1183 23762
rect 0 23704 1122 23760
rect 1178 23704 1183 23760
rect 0 23702 1183 23704
rect 0 23672 800 23702
rect 1117 23699 1183 23702
rect 8661 23762 8727 23765
rect 19793 23762 19859 23765
rect 8661 23760 19859 23762
rect 8661 23704 8666 23760
rect 8722 23704 19798 23760
rect 19854 23704 19859 23760
rect 8661 23702 19859 23704
rect 8661 23699 8727 23702
rect 19793 23699 19859 23702
rect 5441 23626 5507 23629
rect 15142 23626 15148 23628
rect 5441 23624 15148 23626
rect 5441 23568 5446 23624
rect 5502 23568 15148 23624
rect 5441 23566 15148 23568
rect 5441 23563 5507 23566
rect 15142 23564 15148 23566
rect 15212 23564 15218 23628
rect 15561 23626 15627 23629
rect 16573 23626 16639 23629
rect 15561 23624 16639 23626
rect 15561 23568 15566 23624
rect 15622 23568 16578 23624
rect 16634 23568 16639 23624
rect 15561 23566 16639 23568
rect 15561 23563 15627 23566
rect 16573 23563 16639 23566
rect 22093 23626 22159 23629
rect 26200 23626 27000 23656
rect 22093 23624 27000 23626
rect 22093 23568 22098 23624
rect 22154 23568 27000 23624
rect 22093 23566 27000 23568
rect 22093 23563 22159 23566
rect 26200 23536 27000 23566
rect 9121 23490 9187 23493
rect 11513 23490 11579 23493
rect 9121 23488 11579 23490
rect 9121 23432 9126 23488
rect 9182 23432 11518 23488
rect 11574 23432 11579 23488
rect 9121 23430 11579 23432
rect 9121 23427 9187 23430
rect 11513 23427 11579 23430
rect 14273 23490 14339 23493
rect 15377 23490 15443 23493
rect 14273 23488 15443 23490
rect 14273 23432 14278 23488
rect 14334 23432 15382 23488
rect 15438 23432 15443 23488
rect 14273 23430 15443 23432
rect 14273 23427 14339 23430
rect 15377 23427 15443 23430
rect 16849 23490 16915 23493
rect 19149 23490 19215 23493
rect 16849 23488 19215 23490
rect 16849 23432 16854 23488
rect 16910 23432 19154 23488
rect 19210 23432 19215 23488
rect 16849 23430 19215 23432
rect 16849 23427 16915 23430
rect 19149 23427 19215 23430
rect 19977 23490 20043 23493
rect 20110 23490 20116 23492
rect 19977 23488 20116 23490
rect 19977 23432 19982 23488
rect 20038 23432 20116 23488
rect 19977 23430 20116 23432
rect 19977 23427 20043 23430
rect 20110 23428 20116 23430
rect 20180 23428 20186 23492
rect 2946 23424 3262 23425
rect 2946 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3262 23424
rect 2946 23359 3262 23360
rect 12946 23424 13262 23425
rect 12946 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13262 23424
rect 12946 23359 13262 23360
rect 22946 23424 23262 23425
rect 22946 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23262 23424
rect 22946 23359 23262 23360
rect 6729 23354 6795 23357
rect 8569 23354 8635 23357
rect 6729 23352 8635 23354
rect 6729 23296 6734 23352
rect 6790 23296 8574 23352
rect 8630 23296 8635 23352
rect 6729 23294 8635 23296
rect 6729 23291 6795 23294
rect 8569 23291 8635 23294
rect 9438 23292 9444 23356
rect 9508 23354 9514 23356
rect 11881 23354 11947 23357
rect 18597 23354 18663 23357
rect 9508 23352 11947 23354
rect 9508 23296 11886 23352
rect 11942 23296 11947 23352
rect 9508 23294 11947 23296
rect 9508 23292 9514 23294
rect 11881 23291 11947 23294
rect 15518 23352 18663 23354
rect 15518 23296 18602 23352
rect 18658 23296 18663 23352
rect 15518 23294 18663 23296
rect 8385 23218 8451 23221
rect 15518 23218 15578 23294
rect 18597 23291 18663 23294
rect 8385 23216 15578 23218
rect 8385 23160 8390 23216
rect 8446 23160 15578 23216
rect 8385 23158 15578 23160
rect 8385 23155 8451 23158
rect 17350 23156 17356 23220
rect 17420 23218 17426 23220
rect 26200 23218 27000 23248
rect 17420 23158 27000 23218
rect 17420 23156 17426 23158
rect 26200 23128 27000 23158
rect 8569 23082 8635 23085
rect 8569 23080 17418 23082
rect 8569 23024 8574 23080
rect 8630 23024 17418 23080
rect 8569 23022 17418 23024
rect 8569 23019 8635 23022
rect 12157 22946 12223 22949
rect 16757 22946 16823 22949
rect 12157 22944 16823 22946
rect 12157 22888 12162 22944
rect 12218 22888 16762 22944
rect 16818 22888 16823 22944
rect 12157 22886 16823 22888
rect 12157 22883 12223 22886
rect 16757 22883 16823 22886
rect 7946 22880 8262 22881
rect 7946 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8262 22880
rect 7946 22815 8262 22816
rect 12382 22810 12388 22812
rect 8756 22750 12388 22810
rect 0 22674 800 22704
rect 1209 22674 1275 22677
rect 0 22672 1275 22674
rect 0 22616 1214 22672
rect 1270 22616 1275 22672
rect 0 22614 1275 22616
rect 0 22584 800 22614
rect 1209 22611 1275 22614
rect 6269 22674 6335 22677
rect 8756 22674 8816 22750
rect 12382 22748 12388 22750
rect 12452 22748 12458 22812
rect 12566 22748 12572 22812
rect 12636 22810 12642 22812
rect 13353 22810 13419 22813
rect 12636 22808 13419 22810
rect 12636 22752 13358 22808
rect 13414 22752 13419 22808
rect 12636 22750 13419 22752
rect 12636 22748 12642 22750
rect 13353 22747 13419 22750
rect 6269 22672 8816 22674
rect 6269 22616 6274 22672
rect 6330 22616 8816 22672
rect 6269 22614 8816 22616
rect 6269 22611 6335 22614
rect 11094 22612 11100 22676
rect 11164 22674 11170 22676
rect 13537 22674 13603 22677
rect 11164 22672 13603 22674
rect 11164 22616 13542 22672
rect 13598 22616 13603 22672
rect 11164 22614 13603 22616
rect 17358 22674 17418 23022
rect 17718 23020 17724 23084
rect 17788 23082 17794 23084
rect 18505 23082 18571 23085
rect 20437 23082 20503 23085
rect 17788 23080 20503 23082
rect 17788 23024 18510 23080
rect 18566 23024 20442 23080
rect 20498 23024 20503 23080
rect 17788 23022 20503 23024
rect 17788 23020 17794 23022
rect 18505 23019 18571 23022
rect 20437 23019 20503 23022
rect 17946 22880 18262 22881
rect 17946 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18262 22880
rect 17946 22815 18262 22816
rect 21449 22810 21515 22813
rect 26200 22810 27000 22840
rect 21449 22808 27000 22810
rect 21449 22752 21454 22808
rect 21510 22752 27000 22808
rect 21449 22750 27000 22752
rect 21449 22747 21515 22750
rect 26200 22720 27000 22750
rect 19517 22674 19583 22677
rect 17358 22672 19583 22674
rect 17358 22616 19522 22672
rect 19578 22616 19583 22672
rect 17358 22614 19583 22616
rect 11164 22612 11170 22614
rect 13537 22611 13603 22614
rect 19517 22611 19583 22614
rect 3233 22538 3299 22541
rect 3785 22538 3851 22541
rect 19425 22538 19491 22541
rect 24577 22540 24643 22541
rect 24526 22538 24532 22540
rect 3233 22536 19491 22538
rect 3233 22480 3238 22536
rect 3294 22480 3790 22536
rect 3846 22480 19430 22536
rect 19486 22480 19491 22536
rect 3233 22478 19491 22480
rect 24486 22478 24532 22538
rect 24596 22536 24643 22540
rect 24638 22480 24643 22536
rect 3233 22475 3299 22478
rect 3785 22475 3851 22478
rect 19425 22475 19491 22478
rect 24526 22476 24532 22478
rect 24596 22476 24643 22480
rect 24577 22475 24643 22476
rect 12801 22402 12867 22405
rect 12574 22400 12867 22402
rect 12574 22344 12806 22400
rect 12862 22344 12867 22400
rect 12574 22342 12867 22344
rect 2946 22336 3262 22337
rect 2946 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3262 22336
rect 2946 22271 3262 22272
rect 6361 22266 6427 22269
rect 12574 22266 12634 22342
rect 12801 22339 12867 22342
rect 13629 22402 13695 22405
rect 19609 22402 19675 22405
rect 26200 22402 27000 22432
rect 13629 22400 19675 22402
rect 13629 22344 13634 22400
rect 13690 22344 19614 22400
rect 19670 22344 19675 22400
rect 13629 22342 19675 22344
rect 13629 22339 13695 22342
rect 19609 22339 19675 22342
rect 24166 22342 27000 22402
rect 12946 22336 13262 22337
rect 12946 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13262 22336
rect 12946 22271 13262 22272
rect 22946 22336 23262 22337
rect 22946 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23262 22336
rect 22946 22271 23262 22272
rect 6361 22264 12634 22266
rect 6361 22208 6366 22264
rect 6422 22208 12634 22264
rect 6361 22206 12634 22208
rect 6361 22203 6427 22206
rect 4797 22130 4863 22133
rect 16021 22130 16087 22133
rect 4797 22128 16087 22130
rect 4797 22072 4802 22128
rect 4858 22072 16026 22128
rect 16082 22072 16087 22128
rect 4797 22070 16087 22072
rect 4797 22067 4863 22070
rect 16021 22067 16087 22070
rect 16297 22130 16363 22133
rect 20529 22130 20595 22133
rect 16297 22128 20595 22130
rect 16297 22072 16302 22128
rect 16358 22072 20534 22128
rect 20590 22072 20595 22128
rect 16297 22070 20595 22072
rect 16297 22067 16363 22070
rect 20529 22067 20595 22070
rect 21030 22068 21036 22132
rect 21100 22130 21106 22132
rect 21173 22130 21239 22133
rect 21100 22128 21239 22130
rect 21100 22072 21178 22128
rect 21234 22072 21239 22128
rect 21100 22070 21239 22072
rect 21100 22068 21106 22070
rect 21173 22067 21239 22070
rect 21725 22130 21791 22133
rect 24166 22130 24226 22342
rect 26200 22312 27000 22342
rect 21725 22128 24226 22130
rect 21725 22072 21730 22128
rect 21786 22072 24226 22128
rect 21725 22070 24226 22072
rect 21725 22067 21791 22070
rect 10225 21994 10291 21997
rect 22645 21994 22711 21997
rect 26200 21994 27000 22024
rect 10225 21992 22711 21994
rect 10225 21936 10230 21992
rect 10286 21936 22650 21992
rect 22706 21936 22711 21992
rect 10225 21934 22711 21936
rect 10225 21931 10291 21934
rect 22645 21931 22711 21934
rect 24166 21934 27000 21994
rect 9673 21858 9739 21861
rect 12341 21858 12407 21861
rect 9673 21856 12407 21858
rect 9673 21800 9678 21856
rect 9734 21800 12346 21856
rect 12402 21800 12407 21856
rect 9673 21798 12407 21800
rect 9673 21795 9739 21798
rect 12341 21795 12407 21798
rect 12893 21858 12959 21861
rect 13537 21860 13603 21861
rect 13486 21858 13492 21860
rect 12893 21856 13492 21858
rect 13556 21858 13603 21860
rect 14181 21858 14247 21861
rect 16757 21858 16823 21861
rect 13556 21856 13648 21858
rect 12893 21800 12898 21856
rect 12954 21800 13492 21856
rect 13598 21800 13648 21856
rect 12893 21798 13492 21800
rect 12893 21795 12959 21798
rect 13486 21796 13492 21798
rect 13556 21798 13648 21800
rect 14181 21856 16823 21858
rect 14181 21800 14186 21856
rect 14242 21800 16762 21856
rect 16818 21800 16823 21856
rect 14181 21798 16823 21800
rect 13556 21796 13603 21798
rect 13537 21795 13603 21796
rect 14181 21795 14247 21798
rect 16757 21795 16823 21798
rect 20253 21858 20319 21861
rect 22645 21858 22711 21861
rect 20253 21856 22711 21858
rect 20253 21800 20258 21856
rect 20314 21800 22650 21856
rect 22706 21800 22711 21856
rect 20253 21798 22711 21800
rect 20253 21795 20319 21798
rect 22645 21795 22711 21798
rect 7946 21792 8262 21793
rect 7946 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8262 21792
rect 7946 21727 8262 21728
rect 17946 21792 18262 21793
rect 17946 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18262 21792
rect 17946 21727 18262 21728
rect 8477 21722 8543 21725
rect 12433 21722 12499 21725
rect 8477 21720 12499 21722
rect 8477 21664 8482 21720
rect 8538 21664 12438 21720
rect 12494 21664 12499 21720
rect 8477 21662 12499 21664
rect 8477 21659 8543 21662
rect 12433 21659 12499 21662
rect 12566 21660 12572 21724
rect 12636 21722 12642 21724
rect 15193 21722 15259 21725
rect 19425 21722 19491 21725
rect 20345 21722 20411 21725
rect 22185 21722 22251 21725
rect 23473 21722 23539 21725
rect 24025 21722 24091 21725
rect 12636 21662 13416 21722
rect 12636 21660 12642 21662
rect 3785 21586 3851 21589
rect 11881 21586 11947 21589
rect 3785 21584 11947 21586
rect 3785 21528 3790 21584
rect 3846 21528 11886 21584
rect 11942 21528 11947 21584
rect 3785 21526 11947 21528
rect 3785 21523 3851 21526
rect 11881 21523 11947 21526
rect 12157 21586 12223 21589
rect 12433 21586 12499 21589
rect 13356 21586 13416 21662
rect 15193 21720 17004 21722
rect 15193 21664 15198 21720
rect 15254 21664 17004 21720
rect 15193 21662 17004 21664
rect 15193 21659 15259 21662
rect 15837 21586 15903 21589
rect 16297 21586 16363 21589
rect 12157 21584 12499 21586
rect 12157 21528 12162 21584
rect 12218 21528 12438 21584
rect 12494 21528 12499 21584
rect 12157 21526 12499 21528
rect 12157 21523 12223 21526
rect 12433 21523 12499 21526
rect 12574 21526 13186 21586
rect 13356 21584 16363 21586
rect 13356 21528 15842 21584
rect 15898 21528 16302 21584
rect 16358 21528 16363 21584
rect 13356 21526 16363 21528
rect 16944 21586 17004 21662
rect 19425 21720 20411 21722
rect 19425 21664 19430 21720
rect 19486 21664 20350 21720
rect 20406 21664 20411 21720
rect 19425 21662 20411 21664
rect 19425 21659 19491 21662
rect 20345 21659 20411 21662
rect 20670 21720 24091 21722
rect 20670 21664 22190 21720
rect 22246 21664 23478 21720
rect 23534 21664 24030 21720
rect 24086 21664 24091 21720
rect 20670 21662 24091 21664
rect 20437 21586 20503 21589
rect 16944 21584 20503 21586
rect 16944 21528 20442 21584
rect 20498 21528 20503 21584
rect 16944 21526 20503 21528
rect 7833 21450 7899 21453
rect 12574 21450 12634 21526
rect 12985 21450 13051 21453
rect 7833 21448 12634 21450
rect 7833 21392 7838 21448
rect 7894 21392 12634 21448
rect 7833 21390 12634 21392
rect 12804 21448 13051 21450
rect 12804 21392 12990 21448
rect 13046 21392 13051 21448
rect 12804 21390 13051 21392
rect 13126 21450 13186 21526
rect 15837 21523 15903 21526
rect 16297 21523 16363 21526
rect 20437 21523 20503 21526
rect 19609 21450 19675 21453
rect 13126 21448 19675 21450
rect 13126 21392 19614 21448
rect 19670 21392 19675 21448
rect 13126 21390 19675 21392
rect 7833 21387 7899 21390
rect 5625 21314 5691 21317
rect 12382 21314 12388 21316
rect 5625 21312 12388 21314
rect 5625 21256 5630 21312
rect 5686 21256 12388 21312
rect 5625 21254 12388 21256
rect 5625 21251 5691 21254
rect 12382 21252 12388 21254
rect 12452 21252 12458 21316
rect 2946 21248 3262 21249
rect 2946 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3262 21248
rect 2946 21183 3262 21184
rect 5809 21178 5875 21181
rect 12804 21178 12864 21390
rect 12985 21387 13051 21390
rect 19609 21387 19675 21390
rect 16941 21314 17007 21317
rect 20253 21314 20319 21317
rect 20670 21314 20730 21662
rect 22185 21659 22251 21662
rect 23473 21659 23539 21662
rect 24025 21659 24091 21662
rect 21398 21524 21404 21588
rect 21468 21586 21474 21588
rect 23381 21586 23447 21589
rect 21468 21584 23447 21586
rect 21468 21528 23386 21584
rect 23442 21528 23447 21584
rect 21468 21526 23447 21528
rect 21468 21524 21474 21526
rect 23381 21523 23447 21526
rect 22185 21450 22251 21453
rect 24166 21450 24226 21934
rect 26200 21904 27000 21934
rect 24393 21586 24459 21589
rect 26200 21586 27000 21616
rect 24393 21584 27000 21586
rect 24393 21528 24398 21584
rect 24454 21528 27000 21584
rect 24393 21526 27000 21528
rect 24393 21523 24459 21526
rect 26200 21496 27000 21526
rect 22185 21448 24226 21450
rect 22185 21392 22190 21448
rect 22246 21392 24226 21448
rect 22185 21390 24226 21392
rect 22185 21387 22251 21390
rect 16941 21312 20730 21314
rect 16941 21256 16946 21312
rect 17002 21256 20258 21312
rect 20314 21256 20730 21312
rect 16941 21254 20730 21256
rect 21173 21314 21239 21317
rect 22645 21314 22711 21317
rect 21173 21312 22711 21314
rect 21173 21256 21178 21312
rect 21234 21256 22650 21312
rect 22706 21256 22711 21312
rect 21173 21254 22711 21256
rect 16941 21251 17007 21254
rect 20253 21251 20319 21254
rect 21173 21251 21239 21254
rect 22645 21251 22711 21254
rect 12946 21248 13262 21249
rect 12946 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13262 21248
rect 12946 21183 13262 21184
rect 22946 21248 23262 21249
rect 22946 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23262 21248
rect 22946 21183 23262 21184
rect 5809 21176 12864 21178
rect 5809 21120 5814 21176
rect 5870 21120 12864 21176
rect 5809 21118 12864 21120
rect 14365 21178 14431 21181
rect 15653 21178 15719 21181
rect 21357 21178 21423 21181
rect 22001 21178 22067 21181
rect 14365 21176 15578 21178
rect 14365 21120 14370 21176
rect 14426 21120 15578 21176
rect 14365 21118 15578 21120
rect 5809 21115 5875 21118
rect 14365 21115 14431 21118
rect 8753 21042 8819 21045
rect 11329 21042 11395 21045
rect 8753 21040 11395 21042
rect 8753 20984 8758 21040
rect 8814 20984 11334 21040
rect 11390 20984 11395 21040
rect 8753 20982 11395 20984
rect 8753 20979 8819 20982
rect 11329 20979 11395 20982
rect 12525 21042 12591 21045
rect 15518 21042 15578 21118
rect 15653 21176 22067 21178
rect 15653 21120 15658 21176
rect 15714 21120 21362 21176
rect 21418 21120 22006 21176
rect 22062 21120 22067 21176
rect 15653 21118 22067 21120
rect 15653 21115 15719 21118
rect 21357 21115 21423 21118
rect 22001 21115 22067 21118
rect 23381 21178 23447 21181
rect 26200 21178 27000 21208
rect 23381 21176 27000 21178
rect 23381 21120 23386 21176
rect 23442 21120 27000 21176
rect 23381 21118 27000 21120
rect 23381 21115 23447 21118
rect 26200 21088 27000 21118
rect 19425 21042 19491 21045
rect 12525 21040 15394 21042
rect 12525 20984 12530 21040
rect 12586 20984 15394 21040
rect 12525 20982 15394 20984
rect 15518 21040 19491 21042
rect 15518 20984 19430 21040
rect 19486 20984 19491 21040
rect 15518 20982 19491 20984
rect 12525 20979 12591 20982
rect 8293 20906 8359 20909
rect 13721 20906 13787 20909
rect 15193 20908 15259 20909
rect 15142 20906 15148 20908
rect 8293 20904 13787 20906
rect 8293 20848 8298 20904
rect 8354 20848 13726 20904
rect 13782 20848 13787 20904
rect 8293 20846 13787 20848
rect 15102 20846 15148 20906
rect 15212 20904 15259 20908
rect 15254 20848 15259 20904
rect 8293 20843 8359 20846
rect 13721 20843 13787 20846
rect 15142 20844 15148 20846
rect 15212 20844 15259 20848
rect 15334 20906 15394 20982
rect 19425 20979 19491 20982
rect 20345 21042 20411 21045
rect 22461 21042 22527 21045
rect 20345 21040 22527 21042
rect 20345 20984 20350 21040
rect 20406 20984 22466 21040
rect 22522 20984 22527 21040
rect 20345 20982 22527 20984
rect 20345 20979 20411 20982
rect 22461 20979 22527 20982
rect 22686 20980 22692 21044
rect 22756 21042 22762 21044
rect 24393 21042 24459 21045
rect 22756 21040 24459 21042
rect 22756 20984 24398 21040
rect 24454 20984 24459 21040
rect 22756 20982 24459 20984
rect 22756 20980 22762 20982
rect 24393 20979 24459 20982
rect 23197 20906 23263 20909
rect 15334 20904 23263 20906
rect 15334 20848 23202 20904
rect 23258 20848 23263 20904
rect 15334 20846 23263 20848
rect 15193 20843 15259 20844
rect 23197 20843 23263 20846
rect 5901 20770 5967 20773
rect 7005 20770 7071 20773
rect 5901 20768 7071 20770
rect 5901 20712 5906 20768
rect 5962 20712 7010 20768
rect 7066 20712 7071 20768
rect 5901 20710 7071 20712
rect 5901 20707 5967 20710
rect 7005 20707 7071 20710
rect 11053 20770 11119 20773
rect 15653 20770 15719 20773
rect 11053 20768 15719 20770
rect 11053 20712 11058 20768
rect 11114 20712 15658 20768
rect 15714 20712 15719 20768
rect 11053 20710 15719 20712
rect 11053 20707 11119 20710
rect 15653 20707 15719 20710
rect 15837 20772 15903 20773
rect 19517 20772 19583 20773
rect 20805 20772 20871 20773
rect 15837 20768 15884 20772
rect 15948 20770 15954 20772
rect 15837 20712 15842 20768
rect 15837 20708 15884 20712
rect 15948 20710 15994 20770
rect 19517 20768 19564 20772
rect 19628 20770 19634 20772
rect 19517 20712 19522 20768
rect 15948 20708 15954 20710
rect 19517 20708 19564 20712
rect 19628 20710 19674 20770
rect 20805 20768 20852 20772
rect 20916 20770 20922 20772
rect 20805 20712 20810 20768
rect 19628 20708 19634 20710
rect 20805 20708 20852 20712
rect 20916 20710 20962 20770
rect 20916 20708 20922 20710
rect 21214 20708 21220 20772
rect 21284 20770 21290 20772
rect 21633 20770 21699 20773
rect 26200 20770 27000 20800
rect 21284 20768 21699 20770
rect 21284 20712 21638 20768
rect 21694 20712 21699 20768
rect 21284 20710 21699 20712
rect 21284 20708 21290 20710
rect 15837 20707 15903 20708
rect 19517 20707 19583 20708
rect 20805 20707 20871 20708
rect 21633 20707 21699 20710
rect 22050 20710 27000 20770
rect 7946 20704 8262 20705
rect 7946 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8262 20704
rect 7946 20639 8262 20640
rect 17946 20704 18262 20705
rect 17946 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18262 20704
rect 17946 20639 18262 20640
rect 10593 20634 10659 20637
rect 13721 20634 13787 20637
rect 10593 20632 13787 20634
rect 10593 20576 10598 20632
rect 10654 20576 13726 20632
rect 13782 20576 13787 20632
rect 10593 20574 13787 20576
rect 10593 20571 10659 20574
rect 13721 20571 13787 20574
rect 16389 20634 16455 20637
rect 18413 20634 18479 20637
rect 22050 20634 22110 20710
rect 26200 20680 27000 20710
rect 16389 20632 17786 20634
rect 16389 20576 16394 20632
rect 16450 20576 17786 20632
rect 16389 20574 17786 20576
rect 16389 20571 16455 20574
rect 9305 20498 9371 20501
rect 11329 20498 11395 20501
rect 9305 20496 11395 20498
rect 9305 20440 9310 20496
rect 9366 20440 11334 20496
rect 11390 20440 11395 20496
rect 9305 20438 11395 20440
rect 9305 20435 9371 20438
rect 11329 20435 11395 20438
rect 11513 20498 11579 20501
rect 17493 20498 17559 20501
rect 11513 20496 17559 20498
rect 11513 20440 11518 20496
rect 11574 20440 17498 20496
rect 17554 20440 17559 20496
rect 11513 20438 17559 20440
rect 17726 20498 17786 20574
rect 18413 20632 22110 20634
rect 18413 20576 18418 20632
rect 18474 20576 22110 20632
rect 18413 20574 22110 20576
rect 18413 20571 18479 20574
rect 21817 20498 21883 20501
rect 17726 20496 21883 20498
rect 17726 20440 21822 20496
rect 21878 20440 21883 20496
rect 17726 20438 21883 20440
rect 11513 20435 11579 20438
rect 17493 20435 17559 20438
rect 21817 20435 21883 20438
rect 5533 20362 5599 20365
rect 15929 20362 15995 20365
rect 5533 20360 15995 20362
rect 5533 20304 5538 20360
rect 5594 20304 15934 20360
rect 15990 20304 15995 20360
rect 5533 20302 15995 20304
rect 5533 20299 5599 20302
rect 15929 20299 15995 20302
rect 19742 20300 19748 20364
rect 19812 20362 19818 20364
rect 26200 20362 27000 20392
rect 19812 20302 27000 20362
rect 19812 20300 19818 20302
rect 26200 20272 27000 20302
rect 3509 20226 3575 20229
rect 11513 20226 11579 20229
rect 3509 20224 11579 20226
rect 3509 20168 3514 20224
rect 3570 20168 11518 20224
rect 11574 20168 11579 20224
rect 3509 20166 11579 20168
rect 3509 20163 3575 20166
rect 11513 20163 11579 20166
rect 13670 20164 13676 20228
rect 13740 20226 13746 20228
rect 13997 20226 14063 20229
rect 20989 20228 21055 20229
rect 20989 20226 21036 20228
rect 13740 20224 14063 20226
rect 13740 20168 14002 20224
rect 14058 20168 14063 20224
rect 13740 20166 14063 20168
rect 20944 20224 21036 20226
rect 20944 20168 20994 20224
rect 20944 20166 21036 20168
rect 13740 20164 13746 20166
rect 13997 20163 14063 20166
rect 20989 20164 21036 20166
rect 21100 20164 21106 20228
rect 20989 20163 21055 20164
rect 2946 20160 3262 20161
rect 2946 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3262 20160
rect 2946 20095 3262 20096
rect 12946 20160 13262 20161
rect 12946 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13262 20160
rect 12946 20095 13262 20096
rect 22946 20160 23262 20161
rect 22946 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23262 20160
rect 22946 20095 23262 20096
rect 14917 20090 14983 20093
rect 20437 20090 20503 20093
rect 14917 20088 20503 20090
rect 14917 20032 14922 20088
rect 14978 20032 20442 20088
rect 20498 20032 20503 20088
rect 14917 20030 20503 20032
rect 14917 20027 14983 20030
rect 20437 20027 20503 20030
rect 21030 20028 21036 20092
rect 21100 20090 21106 20092
rect 21265 20090 21331 20093
rect 21100 20088 21331 20090
rect 21100 20032 21270 20088
rect 21326 20032 21331 20088
rect 21100 20030 21331 20032
rect 21100 20028 21106 20030
rect 21265 20027 21331 20030
rect 7281 19954 7347 19957
rect 21081 19954 21147 19957
rect 7281 19952 21147 19954
rect 7281 19896 7286 19952
rect 7342 19896 21086 19952
rect 21142 19896 21147 19952
rect 7281 19894 21147 19896
rect 7281 19891 7347 19894
rect 21081 19891 21147 19894
rect 23013 19954 23079 19957
rect 26200 19954 27000 19984
rect 23013 19952 27000 19954
rect 23013 19896 23018 19952
rect 23074 19896 27000 19952
rect 23013 19894 27000 19896
rect 23013 19891 23079 19894
rect 26200 19864 27000 19894
rect 8293 19818 8359 19821
rect 16297 19818 16363 19821
rect 8293 19816 16363 19818
rect 8293 19760 8298 19816
rect 8354 19760 16302 19816
rect 16358 19760 16363 19816
rect 8293 19758 16363 19760
rect 8293 19755 8359 19758
rect 16297 19755 16363 19758
rect 17033 19818 17099 19821
rect 18454 19818 18460 19820
rect 17033 19816 18460 19818
rect 17033 19760 17038 19816
rect 17094 19760 18460 19816
rect 17033 19758 18460 19760
rect 17033 19755 17099 19758
rect 18454 19756 18460 19758
rect 18524 19756 18530 19820
rect 19333 19818 19399 19821
rect 24209 19818 24275 19821
rect 19333 19816 24275 19818
rect 19333 19760 19338 19816
rect 19394 19760 24214 19816
rect 24270 19760 24275 19816
rect 19333 19758 24275 19760
rect 19333 19755 19399 19758
rect 24209 19755 24275 19758
rect 10133 19682 10199 19685
rect 13997 19682 14063 19685
rect 10133 19680 14063 19682
rect 10133 19624 10138 19680
rect 10194 19624 14002 19680
rect 14058 19624 14063 19680
rect 10133 19622 14063 19624
rect 10133 19619 10199 19622
rect 13997 19619 14063 19622
rect 14641 19682 14707 19685
rect 16573 19682 16639 19685
rect 24577 19682 24643 19685
rect 14641 19680 16639 19682
rect 14641 19624 14646 19680
rect 14702 19624 16578 19680
rect 16634 19624 16639 19680
rect 14641 19622 16639 19624
rect 14641 19619 14707 19622
rect 16573 19619 16639 19622
rect 18462 19680 24643 19682
rect 18462 19624 24582 19680
rect 24638 19624 24643 19680
rect 18462 19622 24643 19624
rect 7946 19616 8262 19617
rect 7946 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8262 19616
rect 7946 19551 8262 19552
rect 17946 19616 18262 19617
rect 17946 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18262 19616
rect 17946 19551 18262 19552
rect 15101 19546 15167 19549
rect 9814 19544 15167 19546
rect 9814 19488 15106 19544
rect 15162 19488 15167 19544
rect 9814 19486 15167 19488
rect 6637 19410 6703 19413
rect 9673 19410 9739 19413
rect 6637 19408 9739 19410
rect 6637 19352 6642 19408
rect 6698 19352 9678 19408
rect 9734 19352 9739 19408
rect 6637 19350 9739 19352
rect 6637 19347 6703 19350
rect 9673 19347 9739 19350
rect 6453 19276 6519 19277
rect 6453 19274 6500 19276
rect 6408 19272 6500 19274
rect 6408 19216 6458 19272
rect 6408 19214 6500 19216
rect 6453 19212 6500 19214
rect 6564 19212 6570 19276
rect 7741 19274 7807 19277
rect 9814 19274 9874 19486
rect 15101 19483 15167 19486
rect 11421 19410 11487 19413
rect 11881 19410 11947 19413
rect 13445 19410 13511 19413
rect 14089 19410 14155 19413
rect 11421 19408 14155 19410
rect 11421 19352 11426 19408
rect 11482 19352 11886 19408
rect 11942 19352 13450 19408
rect 13506 19352 14094 19408
rect 14150 19352 14155 19408
rect 11421 19350 14155 19352
rect 11421 19347 11487 19350
rect 11881 19347 11947 19350
rect 13445 19347 13511 19350
rect 14089 19347 14155 19350
rect 15837 19410 15903 19413
rect 16062 19410 16068 19412
rect 15837 19408 16068 19410
rect 15837 19352 15842 19408
rect 15898 19352 16068 19408
rect 15837 19350 16068 19352
rect 15837 19347 15903 19350
rect 16062 19348 16068 19350
rect 16132 19348 16138 19412
rect 16205 19410 16271 19413
rect 16430 19410 16436 19412
rect 16205 19408 16436 19410
rect 16205 19352 16210 19408
rect 16266 19352 16436 19408
rect 16205 19350 16436 19352
rect 16205 19347 16271 19350
rect 16430 19348 16436 19350
rect 16500 19348 16506 19412
rect 18462 19274 18522 19622
rect 24577 19619 24643 19622
rect 23381 19546 23447 19549
rect 26200 19546 27000 19576
rect 23381 19544 27000 19546
rect 23381 19488 23386 19544
rect 23442 19488 27000 19544
rect 23381 19486 27000 19488
rect 23381 19483 23447 19486
rect 26200 19456 27000 19486
rect 19374 19348 19380 19412
rect 19444 19410 19450 19412
rect 19517 19410 19583 19413
rect 24853 19410 24919 19413
rect 19444 19408 19583 19410
rect 19444 19352 19522 19408
rect 19578 19352 19583 19408
rect 19444 19350 19583 19352
rect 19444 19348 19450 19350
rect 19517 19347 19583 19350
rect 23798 19408 24919 19410
rect 23798 19352 24858 19408
rect 24914 19352 24919 19408
rect 23798 19350 24919 19352
rect 7741 19272 9874 19274
rect 7741 19216 7746 19272
rect 7802 19216 9874 19272
rect 7741 19214 9874 19216
rect 12390 19214 18522 19274
rect 19149 19274 19215 19277
rect 22185 19274 22251 19277
rect 23798 19274 23858 19350
rect 24853 19347 24919 19350
rect 19149 19272 22251 19274
rect 19149 19216 19154 19272
rect 19210 19216 22190 19272
rect 22246 19216 22251 19272
rect 19149 19214 22251 19216
rect 6453 19211 6519 19212
rect 7741 19211 7807 19214
rect 4705 19138 4771 19141
rect 12390 19138 12450 19214
rect 19149 19211 19215 19214
rect 22185 19211 22251 19214
rect 22694 19214 23858 19274
rect 23933 19274 23999 19277
rect 25497 19274 25563 19277
rect 23933 19272 25563 19274
rect 23933 19216 23938 19272
rect 23994 19216 25502 19272
rect 25558 19216 25563 19272
rect 23933 19214 25563 19216
rect 4705 19136 12450 19138
rect 4705 19080 4710 19136
rect 4766 19080 12450 19136
rect 4705 19078 12450 19080
rect 21541 19138 21607 19141
rect 22553 19138 22619 19141
rect 21541 19136 22619 19138
rect 21541 19080 21546 19136
rect 21602 19080 22558 19136
rect 22614 19080 22619 19136
rect 21541 19078 22619 19080
rect 4705 19075 4771 19078
rect 21541 19075 21607 19078
rect 22553 19075 22619 19078
rect 2946 19072 3262 19073
rect 2946 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3262 19072
rect 2946 19007 3262 19008
rect 12946 19072 13262 19073
rect 12946 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13262 19072
rect 12946 19007 13262 19008
rect 12709 19002 12775 19005
rect 6272 19000 12775 19002
rect 6272 18944 12714 19000
rect 12770 18944 12775 19000
rect 6272 18942 12775 18944
rect 2589 18866 2655 18869
rect 6272 18866 6332 18942
rect 12709 18939 12775 18942
rect 15377 19002 15443 19005
rect 22694 19002 22754 19214
rect 23933 19211 23999 19214
rect 25497 19211 25563 19214
rect 26200 19138 27000 19168
rect 24166 19078 27000 19138
rect 22946 19072 23262 19073
rect 22946 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23262 19072
rect 22946 19007 23262 19008
rect 15377 19000 22754 19002
rect 15377 18944 15382 19000
rect 15438 18944 22754 19000
rect 15377 18942 22754 18944
rect 15377 18939 15443 18942
rect 24166 18866 24226 19078
rect 26200 19048 27000 19078
rect 2589 18864 6332 18866
rect 2589 18808 2594 18864
rect 2650 18808 6332 18864
rect 2589 18806 6332 18808
rect 6456 18806 24226 18866
rect 2589 18803 2655 18806
rect 3877 18730 3943 18733
rect 6456 18730 6516 18806
rect 3877 18728 6516 18730
rect 3877 18672 3882 18728
rect 3938 18672 6516 18728
rect 3877 18670 6516 18672
rect 8109 18730 8175 18733
rect 22737 18730 22803 18733
rect 8109 18728 22803 18730
rect 8109 18672 8114 18728
rect 8170 18672 22742 18728
rect 22798 18672 22803 18728
rect 8109 18670 22803 18672
rect 3877 18667 3943 18670
rect 8109 18667 8175 18670
rect 22737 18667 22803 18670
rect 23013 18730 23079 18733
rect 26200 18730 27000 18760
rect 23013 18728 27000 18730
rect 23013 18672 23018 18728
rect 23074 18672 27000 18728
rect 23013 18670 27000 18672
rect 23013 18667 23079 18670
rect 26200 18640 27000 18670
rect 11421 18594 11487 18597
rect 17125 18594 17191 18597
rect 11421 18592 17191 18594
rect 11421 18536 11426 18592
rect 11482 18536 17130 18592
rect 17186 18536 17191 18592
rect 11421 18534 17191 18536
rect 11421 18531 11487 18534
rect 17125 18531 17191 18534
rect 20662 18532 20668 18596
rect 20732 18594 20738 18596
rect 21909 18594 21975 18597
rect 20732 18592 21975 18594
rect 20732 18536 21914 18592
rect 21970 18536 21975 18592
rect 20732 18534 21975 18536
rect 20732 18532 20738 18534
rect 21909 18531 21975 18534
rect 22093 18594 22159 18597
rect 24301 18594 24367 18597
rect 22093 18592 24367 18594
rect 22093 18536 22098 18592
rect 22154 18536 24306 18592
rect 24362 18536 24367 18592
rect 22093 18534 24367 18536
rect 22093 18531 22159 18534
rect 24301 18531 24367 18534
rect 7946 18528 8262 18529
rect 7946 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8262 18528
rect 7946 18463 8262 18464
rect 17946 18528 18262 18529
rect 17946 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18262 18528
rect 17946 18463 18262 18464
rect 10133 18458 10199 18461
rect 19517 18458 19583 18461
rect 20805 18458 20871 18461
rect 10133 18456 15578 18458
rect 10133 18400 10138 18456
rect 10194 18400 15578 18456
rect 10133 18398 15578 18400
rect 10133 18395 10199 18398
rect 2221 18322 2287 18325
rect 15377 18322 15443 18325
rect 2221 18320 15443 18322
rect 2221 18264 2226 18320
rect 2282 18264 15382 18320
rect 15438 18264 15443 18320
rect 2221 18262 15443 18264
rect 15518 18322 15578 18398
rect 19517 18456 20871 18458
rect 19517 18400 19522 18456
rect 19578 18400 20810 18456
rect 20866 18400 20871 18456
rect 19517 18398 20871 18400
rect 19517 18395 19583 18398
rect 20805 18395 20871 18398
rect 20989 18458 21055 18461
rect 23381 18458 23447 18461
rect 20989 18456 23447 18458
rect 20989 18400 20994 18456
rect 21050 18400 23386 18456
rect 23442 18400 23447 18456
rect 20989 18398 23447 18400
rect 20989 18395 21055 18398
rect 23381 18395 23447 18398
rect 18229 18322 18295 18325
rect 15518 18320 18295 18322
rect 15518 18264 18234 18320
rect 18290 18264 18295 18320
rect 15518 18262 18295 18264
rect 2221 18259 2287 18262
rect 15377 18259 15443 18262
rect 18229 18259 18295 18262
rect 19333 18322 19399 18325
rect 19793 18322 19859 18325
rect 19333 18320 19859 18322
rect 19333 18264 19338 18320
rect 19394 18264 19798 18320
rect 19854 18264 19859 18320
rect 19333 18262 19859 18264
rect 19333 18259 19399 18262
rect 19793 18259 19859 18262
rect 20621 18322 20687 18325
rect 21633 18322 21699 18325
rect 20621 18320 21699 18322
rect 20621 18264 20626 18320
rect 20682 18264 21638 18320
rect 21694 18264 21699 18320
rect 20621 18262 21699 18264
rect 20621 18259 20687 18262
rect 21633 18259 21699 18262
rect 22921 18322 22987 18325
rect 26200 18322 27000 18352
rect 22921 18320 27000 18322
rect 22921 18264 22926 18320
rect 22982 18264 27000 18320
rect 22921 18262 27000 18264
rect 22921 18259 22987 18262
rect 26200 18232 27000 18262
rect 7005 18186 7071 18189
rect 22461 18186 22527 18189
rect 23473 18186 23539 18189
rect 7005 18184 22527 18186
rect 7005 18128 7010 18184
rect 7066 18128 22466 18184
rect 22522 18128 22527 18184
rect 7005 18126 22527 18128
rect 7005 18123 7071 18126
rect 22461 18123 22527 18126
rect 22694 18184 23539 18186
rect 22694 18128 23478 18184
rect 23534 18128 23539 18184
rect 22694 18126 23539 18128
rect 7281 18050 7347 18053
rect 9622 18050 9628 18052
rect 7281 18048 9628 18050
rect 7281 17992 7286 18048
rect 7342 17992 9628 18048
rect 7281 17990 9628 17992
rect 7281 17987 7347 17990
rect 9622 17988 9628 17990
rect 9692 17988 9698 18052
rect 15009 18050 15075 18053
rect 15009 18048 17464 18050
rect 15009 17992 15014 18048
rect 15070 17992 17464 18048
rect 15009 17990 17464 17992
rect 15009 17987 15075 17990
rect 2946 17984 3262 17985
rect 2946 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3262 17984
rect 2946 17919 3262 17920
rect 12946 17984 13262 17985
rect 12946 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13262 17984
rect 12946 17919 13262 17920
rect 6545 17914 6611 17917
rect 9121 17914 9187 17917
rect 6545 17912 9187 17914
rect 6545 17856 6550 17912
rect 6606 17856 9126 17912
rect 9182 17856 9187 17912
rect 6545 17854 9187 17856
rect 6545 17851 6611 17854
rect 9121 17851 9187 17854
rect 9673 17914 9739 17917
rect 11237 17914 11303 17917
rect 17404 17914 17464 17990
rect 17534 17988 17540 18052
rect 17604 18050 17610 18052
rect 17769 18050 17835 18053
rect 21173 18050 21239 18053
rect 17604 18048 17835 18050
rect 17604 17992 17774 18048
rect 17830 17992 17835 18048
rect 17604 17990 17835 17992
rect 17604 17988 17610 17990
rect 17769 17987 17835 17990
rect 17910 18048 21239 18050
rect 17910 17992 21178 18048
rect 21234 17992 21239 18048
rect 17910 17990 21239 17992
rect 17910 17914 17970 17990
rect 21173 17987 21239 17990
rect 9673 17912 12450 17914
rect 9673 17856 9678 17912
rect 9734 17856 11242 17912
rect 11298 17856 12450 17912
rect 9673 17854 12450 17856
rect 17404 17854 17970 17914
rect 19609 17914 19675 17917
rect 22694 17914 22754 18126
rect 23473 18123 23539 18126
rect 23422 17988 23428 18052
rect 23492 18050 23498 18052
rect 24577 18050 24643 18053
rect 23492 18048 24643 18050
rect 23492 17992 24582 18048
rect 24638 17992 24643 18048
rect 23492 17990 24643 17992
rect 23492 17988 23498 17990
rect 24577 17987 24643 17990
rect 22946 17984 23262 17985
rect 22946 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23262 17984
rect 22946 17919 23262 17920
rect 26200 17914 27000 17944
rect 19609 17912 22754 17914
rect 19609 17856 19614 17912
rect 19670 17856 22754 17912
rect 19609 17854 22754 17856
rect 24166 17854 27000 17914
rect 9673 17851 9739 17854
rect 11237 17851 11303 17854
rect 6913 17778 6979 17781
rect 11094 17778 11100 17780
rect 6913 17776 11100 17778
rect 6913 17720 6918 17776
rect 6974 17720 11100 17776
rect 6913 17718 11100 17720
rect 6913 17715 6979 17718
rect 11094 17716 11100 17718
rect 11164 17716 11170 17780
rect 12390 17778 12450 17854
rect 19609 17851 19675 17854
rect 21081 17778 21147 17781
rect 12390 17776 21147 17778
rect 12390 17720 21086 17776
rect 21142 17720 21147 17776
rect 12390 17718 21147 17720
rect 21081 17715 21147 17718
rect 21633 17778 21699 17781
rect 24166 17778 24226 17854
rect 26200 17824 27000 17854
rect 21633 17776 24226 17778
rect 21633 17720 21638 17776
rect 21694 17720 24226 17776
rect 21633 17718 24226 17720
rect 21633 17715 21699 17718
rect 7097 17642 7163 17645
rect 21909 17642 21975 17645
rect 7097 17640 21975 17642
rect 7097 17584 7102 17640
rect 7158 17584 21914 17640
rect 21970 17584 21975 17640
rect 7097 17582 21975 17584
rect 7097 17579 7163 17582
rect 21909 17579 21975 17582
rect 12157 17506 12223 17509
rect 14181 17506 14247 17509
rect 12157 17504 14247 17506
rect 12157 17448 12162 17504
rect 12218 17448 14186 17504
rect 14242 17448 14247 17504
rect 12157 17446 14247 17448
rect 12157 17443 12223 17446
rect 14181 17443 14247 17446
rect 21081 17506 21147 17509
rect 26200 17506 27000 17536
rect 21081 17504 27000 17506
rect 21081 17448 21086 17504
rect 21142 17448 27000 17504
rect 21081 17446 27000 17448
rect 21081 17443 21147 17446
rect 7946 17440 8262 17441
rect 7946 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8262 17440
rect 7946 17375 8262 17376
rect 17946 17440 18262 17441
rect 17946 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18262 17440
rect 26200 17416 27000 17446
rect 17946 17375 18262 17376
rect 8753 17370 8819 17373
rect 17125 17370 17191 17373
rect 8753 17368 17191 17370
rect 8753 17312 8758 17368
rect 8814 17312 17130 17368
rect 17186 17312 17191 17368
rect 8753 17310 17191 17312
rect 8753 17307 8819 17310
rect 17125 17307 17191 17310
rect 18597 17370 18663 17373
rect 19190 17370 19196 17372
rect 18597 17368 19196 17370
rect 18597 17312 18602 17368
rect 18658 17312 19196 17368
rect 18597 17310 19196 17312
rect 18597 17307 18663 17310
rect 19190 17308 19196 17310
rect 19260 17308 19266 17372
rect 7649 17234 7715 17237
rect 24853 17234 24919 17237
rect 7649 17232 24919 17234
rect 7649 17176 7654 17232
rect 7710 17176 24858 17232
rect 24914 17176 24919 17232
rect 7649 17174 24919 17176
rect 7649 17171 7715 17174
rect 24853 17171 24919 17174
rect 7925 17098 7991 17101
rect 9305 17098 9371 17101
rect 7925 17096 9371 17098
rect 7925 17040 7930 17096
rect 7986 17040 9310 17096
rect 9366 17040 9371 17096
rect 7925 17038 9371 17040
rect 7925 17035 7991 17038
rect 9305 17035 9371 17038
rect 9673 17098 9739 17101
rect 19701 17098 19767 17101
rect 9673 17096 19767 17098
rect 9673 17040 9678 17096
rect 9734 17040 19706 17096
rect 19762 17040 19767 17096
rect 9673 17038 19767 17040
rect 9673 17035 9739 17038
rect 19701 17035 19767 17038
rect 21817 17098 21883 17101
rect 26200 17098 27000 17128
rect 21817 17096 27000 17098
rect 21817 17040 21822 17096
rect 21878 17040 27000 17096
rect 21817 17038 27000 17040
rect 21817 17035 21883 17038
rect 26200 17008 27000 17038
rect 4797 16962 4863 16965
rect 11513 16962 11579 16965
rect 20713 16962 20779 16965
rect 4797 16960 11579 16962
rect 4797 16904 4802 16960
rect 4858 16904 11518 16960
rect 11574 16904 11579 16960
rect 4797 16902 11579 16904
rect 4797 16899 4863 16902
rect 11513 16899 11579 16902
rect 13862 16960 20779 16962
rect 13862 16904 20718 16960
rect 20774 16904 20779 16960
rect 13862 16902 20779 16904
rect 2946 16896 3262 16897
rect 2946 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3262 16896
rect 2946 16831 3262 16832
rect 12946 16896 13262 16897
rect 12946 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13262 16896
rect 12946 16831 13262 16832
rect 7005 16826 7071 16829
rect 12065 16826 12131 16829
rect 7005 16824 12131 16826
rect 7005 16768 7010 16824
rect 7066 16768 12070 16824
rect 12126 16768 12131 16824
rect 7005 16766 12131 16768
rect 7005 16763 7071 16766
rect 12065 16763 12131 16766
rect 9121 16690 9187 16693
rect 9765 16690 9831 16693
rect 9121 16688 9831 16690
rect 9121 16632 9126 16688
rect 9182 16632 9770 16688
rect 9826 16632 9831 16688
rect 9121 16630 9831 16632
rect 9121 16627 9187 16630
rect 9765 16627 9831 16630
rect 9949 16690 10015 16693
rect 13862 16690 13922 16902
rect 20713 16899 20779 16902
rect 22946 16896 23262 16897
rect 22946 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23262 16896
rect 22946 16831 23262 16832
rect 16614 16764 16620 16828
rect 16684 16826 16690 16828
rect 19558 16826 19564 16828
rect 16684 16766 19564 16826
rect 16684 16764 16690 16766
rect 19558 16764 19564 16766
rect 19628 16764 19634 16828
rect 9949 16688 13922 16690
rect 9949 16632 9954 16688
rect 10010 16632 13922 16688
rect 9949 16630 13922 16632
rect 13997 16690 14063 16693
rect 21633 16690 21699 16693
rect 13997 16688 21699 16690
rect 13997 16632 14002 16688
rect 14058 16632 21638 16688
rect 21694 16632 21699 16688
rect 13997 16630 21699 16632
rect 9949 16627 10015 16630
rect 13997 16627 14063 16630
rect 21633 16627 21699 16630
rect 22461 16690 22527 16693
rect 26200 16690 27000 16720
rect 22461 16688 27000 16690
rect 22461 16632 22466 16688
rect 22522 16632 27000 16688
rect 22461 16630 27000 16632
rect 22461 16627 22527 16630
rect 26200 16600 27000 16630
rect 4153 16554 4219 16557
rect 8886 16554 8892 16556
rect 4153 16552 8892 16554
rect 4153 16496 4158 16552
rect 4214 16496 8892 16552
rect 4153 16494 8892 16496
rect 4153 16491 4219 16494
rect 8886 16492 8892 16494
rect 8956 16492 8962 16556
rect 11053 16554 11119 16557
rect 14641 16554 14707 16557
rect 11053 16552 14707 16554
rect 11053 16496 11058 16552
rect 11114 16496 14646 16552
rect 14702 16496 14707 16552
rect 11053 16494 14707 16496
rect 11053 16491 11119 16494
rect 14641 16491 14707 16494
rect 15837 16554 15903 16557
rect 19241 16554 19307 16557
rect 15837 16552 19307 16554
rect 15837 16496 15842 16552
rect 15898 16496 19246 16552
rect 19302 16496 19307 16552
rect 15837 16494 19307 16496
rect 15837 16491 15903 16494
rect 19241 16491 19307 16494
rect 8385 16418 8451 16421
rect 17718 16418 17724 16420
rect 8385 16416 17724 16418
rect 8385 16360 8390 16416
rect 8446 16360 17724 16416
rect 8385 16358 17724 16360
rect 8385 16355 8451 16358
rect 17718 16356 17724 16358
rect 17788 16356 17794 16420
rect 7946 16352 8262 16353
rect 7946 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8262 16352
rect 7946 16287 8262 16288
rect 17946 16352 18262 16353
rect 17946 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18262 16352
rect 17946 16287 18262 16288
rect 13353 16282 13419 16285
rect 17217 16282 17283 16285
rect 13353 16280 17283 16282
rect 13353 16224 13358 16280
rect 13414 16224 17222 16280
rect 17278 16224 17283 16280
rect 13353 16222 17283 16224
rect 13353 16219 13419 16222
rect 17217 16219 17283 16222
rect 24853 16282 24919 16285
rect 26200 16282 27000 16312
rect 24853 16280 27000 16282
rect 24853 16224 24858 16280
rect 24914 16224 27000 16280
rect 24853 16222 27000 16224
rect 24853 16219 24919 16222
rect 26200 16192 27000 16222
rect 6821 16146 6887 16149
rect 24669 16146 24735 16149
rect 6821 16144 24735 16146
rect 6821 16088 6826 16144
rect 6882 16088 24674 16144
rect 24730 16088 24735 16144
rect 6821 16086 24735 16088
rect 6821 16083 6887 16086
rect 24669 16083 24735 16086
rect 9121 16010 9187 16013
rect 25865 16010 25931 16013
rect 9121 16008 25931 16010
rect 9121 15952 9126 16008
rect 9182 15952 25870 16008
rect 25926 15952 25931 16008
rect 9121 15950 25931 15952
rect 9121 15947 9187 15950
rect 25865 15947 25931 15950
rect 15837 15874 15903 15877
rect 19742 15874 19748 15876
rect 15837 15872 19748 15874
rect 15837 15816 15842 15872
rect 15898 15816 19748 15872
rect 15837 15814 19748 15816
rect 15837 15811 15903 15814
rect 19742 15812 19748 15814
rect 19812 15812 19818 15876
rect 24669 15874 24735 15877
rect 26200 15874 27000 15904
rect 24669 15872 27000 15874
rect 24669 15816 24674 15872
rect 24730 15816 27000 15872
rect 24669 15814 27000 15816
rect 24669 15811 24735 15814
rect 2946 15808 3262 15809
rect 2946 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3262 15808
rect 2946 15743 3262 15744
rect 12946 15808 13262 15809
rect 12946 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13262 15808
rect 12946 15743 13262 15744
rect 22946 15808 23262 15809
rect 22946 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23262 15808
rect 26200 15784 27000 15814
rect 22946 15743 23262 15744
rect 16481 15738 16547 15741
rect 20662 15738 20668 15740
rect 16481 15736 20668 15738
rect 16481 15680 16486 15736
rect 16542 15680 20668 15736
rect 16481 15678 20668 15680
rect 16481 15675 16547 15678
rect 20662 15676 20668 15678
rect 20732 15676 20738 15740
rect 9397 15604 9463 15605
rect 9397 15602 9444 15604
rect 9352 15600 9444 15602
rect 9352 15544 9402 15600
rect 9352 15542 9444 15544
rect 9397 15540 9444 15542
rect 9508 15540 9514 15604
rect 9581 15602 9647 15605
rect 24526 15602 24532 15604
rect 9581 15600 24532 15602
rect 9581 15544 9586 15600
rect 9642 15544 24532 15600
rect 9581 15542 24532 15544
rect 9397 15539 9463 15540
rect 9581 15539 9647 15542
rect 24526 15540 24532 15542
rect 24596 15540 24602 15604
rect 8753 15466 8819 15469
rect 15837 15466 15903 15469
rect 8753 15464 15903 15466
rect 8753 15408 8758 15464
rect 8814 15408 15842 15464
rect 15898 15408 15903 15464
rect 8753 15406 15903 15408
rect 8753 15403 8819 15406
rect 15837 15403 15903 15406
rect 16665 15466 16731 15469
rect 19374 15466 19380 15468
rect 16665 15464 19380 15466
rect 16665 15408 16670 15464
rect 16726 15408 19380 15464
rect 16665 15406 19380 15408
rect 16665 15403 16731 15406
rect 19374 15404 19380 15406
rect 19444 15404 19450 15468
rect 20345 15466 20411 15469
rect 26200 15466 27000 15496
rect 20345 15464 27000 15466
rect 20345 15408 20350 15464
rect 20406 15408 27000 15464
rect 20345 15406 27000 15408
rect 20345 15403 20411 15406
rect 26200 15376 27000 15406
rect 9765 15330 9831 15333
rect 17217 15330 17283 15333
rect 9765 15328 17283 15330
rect 9765 15272 9770 15328
rect 9826 15272 17222 15328
rect 17278 15272 17283 15328
rect 9765 15270 17283 15272
rect 9765 15267 9831 15270
rect 17217 15267 17283 15270
rect 21633 15330 21699 15333
rect 22686 15330 22692 15332
rect 21633 15328 22692 15330
rect 21633 15272 21638 15328
rect 21694 15272 22692 15328
rect 21633 15270 22692 15272
rect 21633 15267 21699 15270
rect 22686 15268 22692 15270
rect 22756 15268 22762 15332
rect 7946 15264 8262 15265
rect 7946 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8262 15264
rect 7946 15199 8262 15200
rect 17946 15264 18262 15265
rect 17946 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18262 15264
rect 17946 15199 18262 15200
rect 14958 15132 14964 15196
rect 15028 15194 15034 15196
rect 15285 15194 15351 15197
rect 15028 15192 15351 15194
rect 15028 15136 15290 15192
rect 15346 15136 15351 15192
rect 15028 15134 15351 15136
rect 15028 15132 15034 15134
rect 15285 15131 15351 15134
rect 22277 15194 22343 15197
rect 23197 15194 23263 15197
rect 22277 15192 23263 15194
rect 22277 15136 22282 15192
rect 22338 15136 23202 15192
rect 23258 15136 23263 15192
rect 22277 15134 23263 15136
rect 22277 15131 22343 15134
rect 23197 15131 23263 15134
rect 10358 14996 10364 15060
rect 10428 15058 10434 15060
rect 10501 15058 10567 15061
rect 10428 15056 10567 15058
rect 10428 15000 10506 15056
rect 10562 15000 10567 15056
rect 10428 14998 10567 15000
rect 10428 14996 10434 14998
rect 10501 14995 10567 14998
rect 10961 15058 11027 15061
rect 16614 15058 16620 15060
rect 10961 15056 16620 15058
rect 10961 15000 10966 15056
rect 11022 15000 16620 15056
rect 10961 14998 16620 15000
rect 10961 14995 11027 14998
rect 16614 14996 16620 14998
rect 16684 14996 16690 15060
rect 17217 15058 17283 15061
rect 26200 15058 27000 15088
rect 17217 15056 27000 15058
rect 17217 15000 17222 15056
rect 17278 15000 27000 15056
rect 17217 14998 27000 15000
rect 17217 14995 17283 14998
rect 26200 14968 27000 14998
rect 6545 14922 6611 14925
rect 19425 14922 19491 14925
rect 6545 14920 19491 14922
rect 6545 14864 6550 14920
rect 6606 14864 19430 14920
rect 19486 14864 19491 14920
rect 6545 14862 19491 14864
rect 6545 14859 6611 14862
rect 19425 14859 19491 14862
rect 22318 14860 22324 14924
rect 22388 14922 22394 14924
rect 23381 14922 23447 14925
rect 22388 14920 23447 14922
rect 22388 14864 23386 14920
rect 23442 14864 23447 14920
rect 22388 14862 23447 14864
rect 22388 14860 22394 14862
rect 23381 14859 23447 14862
rect 20253 14786 20319 14789
rect 16806 14784 20319 14786
rect 16806 14728 20258 14784
rect 20314 14728 20319 14784
rect 16806 14726 20319 14728
rect 2946 14720 3262 14721
rect 2946 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3262 14720
rect 2946 14655 3262 14656
rect 12946 14720 13262 14721
rect 12946 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13262 14720
rect 12946 14655 13262 14656
rect 11605 14514 11671 14517
rect 16806 14514 16866 14726
rect 20253 14723 20319 14726
rect 22946 14720 23262 14721
rect 22946 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23262 14720
rect 22946 14655 23262 14656
rect 20161 14650 20227 14653
rect 11605 14512 16866 14514
rect 11605 14456 11610 14512
rect 11666 14456 16866 14512
rect 11605 14454 16866 14456
rect 16990 14648 20227 14650
rect 16990 14592 20166 14648
rect 20222 14592 20227 14648
rect 16990 14590 20227 14592
rect 11605 14451 11671 14454
rect 4521 14378 4587 14381
rect 16990 14378 17050 14590
rect 20161 14587 20227 14590
rect 23381 14650 23447 14653
rect 26200 14650 27000 14680
rect 23381 14648 27000 14650
rect 23381 14592 23386 14648
rect 23442 14592 27000 14648
rect 23381 14590 27000 14592
rect 23381 14587 23447 14590
rect 26200 14560 27000 14590
rect 19701 14514 19767 14517
rect 21950 14514 21956 14516
rect 19701 14512 21956 14514
rect 19701 14456 19706 14512
rect 19762 14456 21956 14512
rect 19701 14454 21956 14456
rect 19701 14451 19767 14454
rect 21950 14452 21956 14454
rect 22020 14452 22026 14516
rect 26049 14378 26115 14381
rect 4521 14376 17050 14378
rect 4521 14320 4526 14376
rect 4582 14320 17050 14376
rect 4521 14318 17050 14320
rect 17174 14376 26115 14378
rect 17174 14320 26054 14376
rect 26110 14320 26115 14376
rect 17174 14318 26115 14320
rect 4521 14315 4587 14318
rect 11789 14242 11855 14245
rect 17174 14242 17234 14318
rect 26049 14315 26115 14318
rect 11789 14240 17234 14242
rect 11789 14184 11794 14240
rect 11850 14184 17234 14240
rect 11789 14182 17234 14184
rect 22829 14242 22895 14245
rect 26200 14242 27000 14272
rect 22829 14240 27000 14242
rect 22829 14184 22834 14240
rect 22890 14184 27000 14240
rect 22829 14182 27000 14184
rect 11789 14179 11855 14182
rect 22829 14179 22895 14182
rect 7946 14176 8262 14177
rect 7946 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8262 14176
rect 7946 14111 8262 14112
rect 17946 14176 18262 14177
rect 17946 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18262 14176
rect 26200 14152 27000 14182
rect 17946 14111 18262 14112
rect 16021 14106 16087 14109
rect 18873 14106 18939 14109
rect 22277 14106 22343 14109
rect 16021 14104 17786 14106
rect 16021 14048 16026 14104
rect 16082 14048 17786 14104
rect 16021 14046 17786 14048
rect 16021 14043 16087 14046
rect 11973 13972 12039 13973
rect 17493 13972 17559 13973
rect 11973 13970 12020 13972
rect 11928 13968 12020 13970
rect 11928 13912 11978 13968
rect 11928 13910 12020 13912
rect 11973 13908 12020 13910
rect 12084 13908 12090 13972
rect 17493 13970 17540 13972
rect 17448 13968 17540 13970
rect 17448 13912 17498 13968
rect 17448 13910 17540 13912
rect 17493 13908 17540 13910
rect 17604 13908 17610 13972
rect 17726 13970 17786 14046
rect 18873 14104 22343 14106
rect 18873 14048 18878 14104
rect 18934 14048 22282 14104
rect 22338 14048 22343 14104
rect 18873 14046 22343 14048
rect 18873 14043 18939 14046
rect 22277 14043 22343 14046
rect 21398 13970 21404 13972
rect 17726 13910 21404 13970
rect 21398 13908 21404 13910
rect 21468 13908 21474 13972
rect 22093 13970 22159 13973
rect 22093 13968 22570 13970
rect 22093 13912 22098 13968
rect 22154 13912 22570 13968
rect 22093 13910 22570 13912
rect 11973 13907 12039 13908
rect 17493 13907 17559 13908
rect 22093 13907 22159 13910
rect 7373 13834 7439 13837
rect 18873 13834 18939 13837
rect 7373 13832 18939 13834
rect 7373 13776 7378 13832
rect 7434 13776 18878 13832
rect 18934 13776 18939 13832
rect 7373 13774 18939 13776
rect 7373 13771 7439 13774
rect 18873 13771 18939 13774
rect 20478 13772 20484 13836
rect 20548 13834 20554 13836
rect 22277 13834 22343 13837
rect 20548 13832 22343 13834
rect 20548 13776 22282 13832
rect 22338 13776 22343 13832
rect 20548 13774 22343 13776
rect 22510 13834 22570 13910
rect 26200 13834 27000 13864
rect 22510 13774 27000 13834
rect 20548 13772 20554 13774
rect 22277 13771 22343 13774
rect 26200 13744 27000 13774
rect 15653 13698 15719 13701
rect 17350 13698 17356 13700
rect 15653 13696 17356 13698
rect 15653 13640 15658 13696
rect 15714 13640 17356 13696
rect 15653 13638 17356 13640
rect 15653 13635 15719 13638
rect 17350 13636 17356 13638
rect 17420 13636 17426 13700
rect 2946 13632 3262 13633
rect 2946 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3262 13632
rect 2946 13567 3262 13568
rect 12946 13632 13262 13633
rect 12946 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13262 13632
rect 12946 13567 13262 13568
rect 22946 13632 23262 13633
rect 22946 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23262 13632
rect 22946 13567 23262 13568
rect 13670 13500 13676 13564
rect 13740 13562 13746 13564
rect 17718 13562 17724 13564
rect 13740 13502 17724 13562
rect 13740 13500 13746 13502
rect 17718 13500 17724 13502
rect 17788 13500 17794 13564
rect 19057 13426 19123 13429
rect 20345 13426 20411 13429
rect 19057 13424 20411 13426
rect 19057 13368 19062 13424
rect 19118 13368 20350 13424
rect 20406 13368 20411 13424
rect 19057 13366 20411 13368
rect 19057 13363 19123 13366
rect 20345 13363 20411 13366
rect 22369 13426 22435 13429
rect 26200 13426 27000 13456
rect 22369 13424 27000 13426
rect 22369 13368 22374 13424
rect 22430 13368 27000 13424
rect 22369 13366 27000 13368
rect 22369 13363 22435 13366
rect 26200 13336 27000 13366
rect 15745 13290 15811 13293
rect 21030 13290 21036 13292
rect 15745 13288 21036 13290
rect 15745 13232 15750 13288
rect 15806 13232 21036 13288
rect 15745 13230 21036 13232
rect 15745 13227 15811 13230
rect 21030 13228 21036 13230
rect 21100 13228 21106 13292
rect 7946 13088 8262 13089
rect 7946 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8262 13088
rect 7946 13023 8262 13024
rect 17946 13088 18262 13089
rect 17946 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18262 13088
rect 17946 13023 18262 13024
rect 22829 13018 22895 13021
rect 26200 13018 27000 13048
rect 22829 13016 27000 13018
rect 22829 12960 22834 13016
rect 22890 12960 27000 13016
rect 22829 12958 27000 12960
rect 22829 12955 22895 12958
rect 26200 12928 27000 12958
rect 6729 12882 6795 12885
rect 24853 12882 24919 12885
rect 6729 12880 24919 12882
rect 6729 12824 6734 12880
rect 6790 12824 24858 12880
rect 24914 12824 24919 12880
rect 6729 12822 24919 12824
rect 6729 12819 6795 12822
rect 24853 12819 24919 12822
rect 25129 12610 25195 12613
rect 26200 12610 27000 12640
rect 25129 12608 27000 12610
rect 25129 12552 25134 12608
rect 25190 12552 27000 12608
rect 25129 12550 27000 12552
rect 25129 12547 25195 12550
rect 2946 12544 3262 12545
rect 2946 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3262 12544
rect 2946 12479 3262 12480
rect 12946 12544 13262 12545
rect 12946 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13262 12544
rect 12946 12479 13262 12480
rect 22946 12544 23262 12545
rect 22946 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23262 12544
rect 26200 12520 27000 12550
rect 22946 12479 23262 12480
rect 16849 12474 16915 12477
rect 20846 12474 20852 12476
rect 16849 12472 20852 12474
rect 16849 12416 16854 12472
rect 16910 12416 20852 12472
rect 16849 12414 20852 12416
rect 16849 12411 16915 12414
rect 20846 12412 20852 12414
rect 20916 12412 20922 12476
rect 11329 12338 11395 12341
rect 19149 12338 19215 12341
rect 11329 12336 19215 12338
rect 11329 12280 11334 12336
rect 11390 12280 19154 12336
rect 19210 12280 19215 12336
rect 11329 12278 19215 12280
rect 11329 12275 11395 12278
rect 19149 12275 19215 12278
rect 24669 12202 24735 12205
rect 26200 12202 27000 12232
rect 24669 12200 27000 12202
rect 24669 12144 24674 12200
rect 24730 12144 27000 12200
rect 24669 12142 27000 12144
rect 24669 12139 24735 12142
rect 26200 12112 27000 12142
rect 7946 12000 8262 12001
rect 7946 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8262 12000
rect 7946 11935 8262 11936
rect 17946 12000 18262 12001
rect 17946 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18262 12000
rect 17946 11935 18262 11936
rect 24853 11794 24919 11797
rect 26200 11794 27000 11824
rect 24853 11792 27000 11794
rect 24853 11736 24858 11792
rect 24914 11736 27000 11792
rect 24853 11734 27000 11736
rect 24853 11731 24919 11734
rect 26200 11704 27000 11734
rect 17718 11596 17724 11660
rect 17788 11658 17794 11660
rect 24577 11658 24643 11661
rect 17788 11656 24643 11658
rect 17788 11600 24582 11656
rect 24638 11600 24643 11656
rect 17788 11598 24643 11600
rect 17788 11596 17794 11598
rect 24577 11595 24643 11598
rect 2946 11456 3262 11457
rect 2946 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3262 11456
rect 2946 11391 3262 11392
rect 12946 11456 13262 11457
rect 12946 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13262 11456
rect 12946 11391 13262 11392
rect 22946 11456 23262 11457
rect 22946 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23262 11456
rect 22946 11391 23262 11392
rect 16113 11386 16179 11389
rect 16246 11386 16252 11388
rect 16113 11384 16252 11386
rect 16113 11328 16118 11384
rect 16174 11328 16252 11384
rect 16113 11326 16252 11328
rect 16113 11323 16179 11326
rect 16246 11324 16252 11326
rect 16316 11324 16322 11388
rect 24853 11386 24919 11389
rect 26200 11386 27000 11416
rect 24853 11384 27000 11386
rect 24853 11328 24858 11384
rect 24914 11328 27000 11384
rect 24853 11326 27000 11328
rect 24853 11323 24919 11326
rect 26200 11296 27000 11326
rect 18321 11114 18387 11117
rect 18454 11114 18460 11116
rect 18321 11112 18460 11114
rect 18321 11056 18326 11112
rect 18382 11056 18460 11112
rect 18321 11054 18460 11056
rect 18321 11051 18387 11054
rect 18454 11052 18460 11054
rect 18524 11052 18530 11116
rect 19425 11114 19491 11117
rect 20110 11114 20116 11116
rect 19425 11112 20116 11114
rect 19425 11056 19430 11112
rect 19486 11056 20116 11112
rect 19425 11054 20116 11056
rect 19425 11051 19491 11054
rect 20110 11052 20116 11054
rect 20180 11052 20186 11116
rect 24761 10978 24827 10981
rect 26200 10978 27000 11008
rect 24761 10976 27000 10978
rect 24761 10920 24766 10976
rect 24822 10920 27000 10976
rect 24761 10918 27000 10920
rect 24761 10915 24827 10918
rect 7946 10912 8262 10913
rect 7946 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8262 10912
rect 7946 10847 8262 10848
rect 17946 10912 18262 10913
rect 17946 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18262 10912
rect 26200 10888 27000 10918
rect 17946 10847 18262 10848
rect 17585 10706 17651 10709
rect 23422 10706 23428 10708
rect 17585 10704 23428 10706
rect 17585 10648 17590 10704
rect 17646 10648 23428 10704
rect 17585 10646 23428 10648
rect 17585 10643 17651 10646
rect 23422 10644 23428 10646
rect 23492 10644 23498 10708
rect 24853 10570 24919 10573
rect 26200 10570 27000 10600
rect 24853 10568 27000 10570
rect 24853 10512 24858 10568
rect 24914 10512 27000 10568
rect 24853 10510 27000 10512
rect 24853 10507 24919 10510
rect 26200 10480 27000 10510
rect 2946 10368 3262 10369
rect 2946 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3262 10368
rect 2946 10303 3262 10304
rect 12946 10368 13262 10369
rect 12946 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13262 10368
rect 12946 10303 13262 10304
rect 22946 10368 23262 10369
rect 22946 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23262 10368
rect 22946 10303 23262 10304
rect 16062 10236 16068 10300
rect 16132 10298 16138 10300
rect 20713 10298 20779 10301
rect 16132 10296 20779 10298
rect 16132 10240 20718 10296
rect 20774 10240 20779 10296
rect 16132 10238 20779 10240
rect 16132 10236 16138 10238
rect 20713 10235 20779 10238
rect 24577 10162 24643 10165
rect 26200 10162 27000 10192
rect 24577 10160 27000 10162
rect 24577 10104 24582 10160
rect 24638 10104 27000 10160
rect 24577 10102 27000 10104
rect 24577 10099 24643 10102
rect 26200 10072 27000 10102
rect 7946 9824 8262 9825
rect 7946 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8262 9824
rect 7946 9759 8262 9760
rect 17946 9824 18262 9825
rect 17946 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18262 9824
rect 17946 9759 18262 9760
rect 20713 9754 20779 9757
rect 21265 9756 21331 9757
rect 21214 9754 21220 9756
rect 20713 9752 21220 9754
rect 21284 9754 21331 9756
rect 23289 9754 23355 9757
rect 26200 9754 27000 9784
rect 21284 9752 21376 9754
rect 20713 9696 20718 9752
rect 20774 9696 21220 9752
rect 21326 9696 21376 9752
rect 20713 9694 21220 9696
rect 20713 9691 20779 9694
rect 21214 9692 21220 9694
rect 21284 9694 21376 9696
rect 23289 9752 27000 9754
rect 23289 9696 23294 9752
rect 23350 9696 27000 9752
rect 23289 9694 27000 9696
rect 21284 9692 21331 9694
rect 21265 9691 21331 9692
rect 23289 9691 23355 9694
rect 26200 9664 27000 9694
rect 15878 9420 15884 9484
rect 15948 9482 15954 9484
rect 19333 9482 19399 9485
rect 15948 9480 19399 9482
rect 15948 9424 19338 9480
rect 19394 9424 19399 9480
rect 15948 9422 19399 9424
rect 15948 9420 15954 9422
rect 19333 9419 19399 9422
rect 24853 9346 24919 9349
rect 26200 9346 27000 9376
rect 24853 9344 27000 9346
rect 24853 9288 24858 9344
rect 24914 9288 27000 9344
rect 24853 9286 27000 9288
rect 24853 9283 24919 9286
rect 2946 9280 3262 9281
rect 2946 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3262 9280
rect 2946 9215 3262 9216
rect 12946 9280 13262 9281
rect 12946 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13262 9280
rect 12946 9215 13262 9216
rect 22946 9280 23262 9281
rect 22946 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23262 9280
rect 26200 9256 27000 9286
rect 22946 9215 23262 9216
rect 24669 8938 24735 8941
rect 26200 8938 27000 8968
rect 24669 8936 27000 8938
rect 24669 8880 24674 8936
rect 24730 8880 27000 8936
rect 24669 8878 27000 8880
rect 24669 8875 24735 8878
rect 26200 8848 27000 8878
rect 7946 8736 8262 8737
rect 7946 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8262 8736
rect 7946 8671 8262 8672
rect 17946 8736 18262 8737
rect 17946 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18262 8736
rect 17946 8671 18262 8672
rect 24853 8530 24919 8533
rect 26200 8530 27000 8560
rect 24853 8528 27000 8530
rect 24853 8472 24858 8528
rect 24914 8472 27000 8528
rect 24853 8470 27000 8472
rect 24853 8467 24919 8470
rect 26200 8440 27000 8470
rect 16430 8332 16436 8396
rect 16500 8394 16506 8396
rect 19701 8394 19767 8397
rect 22001 8396 22067 8397
rect 21950 8394 21956 8396
rect 16500 8392 19767 8394
rect 16500 8336 19706 8392
rect 19762 8336 19767 8392
rect 16500 8334 19767 8336
rect 21910 8334 21956 8394
rect 22020 8392 22067 8396
rect 22062 8336 22067 8392
rect 16500 8332 16506 8334
rect 19701 8331 19767 8334
rect 21950 8332 21956 8334
rect 22020 8332 22067 8336
rect 22001 8331 22067 8332
rect 2946 8192 3262 8193
rect 2946 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3262 8192
rect 2946 8127 3262 8128
rect 12946 8192 13262 8193
rect 12946 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13262 8192
rect 12946 8127 13262 8128
rect 22946 8192 23262 8193
rect 22946 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23262 8192
rect 22946 8127 23262 8128
rect 24945 8122 25011 8125
rect 26200 8122 27000 8152
rect 24945 8120 27000 8122
rect 24945 8064 24950 8120
rect 25006 8064 27000 8120
rect 24945 8062 27000 8064
rect 24945 8059 25011 8062
rect 26200 8032 27000 8062
rect 19190 7924 19196 7988
rect 19260 7986 19266 7988
rect 20529 7986 20595 7989
rect 19260 7984 20595 7986
rect 19260 7928 20534 7984
rect 20590 7928 20595 7984
rect 19260 7926 20595 7928
rect 19260 7924 19266 7926
rect 20529 7923 20595 7926
rect 13486 7788 13492 7852
rect 13556 7850 13562 7852
rect 21265 7850 21331 7853
rect 13556 7848 21331 7850
rect 13556 7792 21270 7848
rect 21326 7792 21331 7848
rect 13556 7790 21331 7792
rect 13556 7788 13562 7790
rect 21265 7787 21331 7790
rect 24761 7714 24827 7717
rect 26200 7714 27000 7744
rect 24761 7712 27000 7714
rect 24761 7656 24766 7712
rect 24822 7656 27000 7712
rect 24761 7654 27000 7656
rect 24761 7651 24827 7654
rect 7946 7648 8262 7649
rect 7946 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8262 7648
rect 7946 7583 8262 7584
rect 17946 7648 18262 7649
rect 17946 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18262 7648
rect 26200 7624 27000 7654
rect 17946 7583 18262 7584
rect 24853 7306 24919 7309
rect 26200 7306 27000 7336
rect 24853 7304 27000 7306
rect 24853 7248 24858 7304
rect 24914 7248 27000 7304
rect 24853 7246 27000 7248
rect 24853 7243 24919 7246
rect 26200 7216 27000 7246
rect 2946 7104 3262 7105
rect 2946 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3262 7104
rect 2946 7039 3262 7040
rect 12946 7104 13262 7105
rect 12946 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13262 7104
rect 12946 7039 13262 7040
rect 22946 7104 23262 7105
rect 22946 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23262 7104
rect 22946 7039 23262 7040
rect 22185 6898 22251 6901
rect 22318 6898 22324 6900
rect 22185 6896 22324 6898
rect 22185 6840 22190 6896
rect 22246 6840 22324 6896
rect 22185 6838 22324 6840
rect 22185 6835 22251 6838
rect 22318 6836 22324 6838
rect 22388 6836 22394 6900
rect 24853 6898 24919 6901
rect 26200 6898 27000 6928
rect 24853 6896 27000 6898
rect 24853 6840 24858 6896
rect 24914 6840 27000 6896
rect 24853 6838 27000 6840
rect 24853 6835 24919 6838
rect 26200 6808 27000 6838
rect 7946 6560 8262 6561
rect 7946 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8262 6560
rect 7946 6495 8262 6496
rect 17946 6560 18262 6561
rect 17946 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18262 6560
rect 17946 6495 18262 6496
rect 24669 6490 24735 6493
rect 26200 6490 27000 6520
rect 24669 6488 27000 6490
rect 24669 6432 24674 6488
rect 24730 6432 27000 6488
rect 24669 6430 27000 6432
rect 24669 6427 24735 6430
rect 26200 6400 27000 6430
rect 24853 6082 24919 6085
rect 26200 6082 27000 6112
rect 24853 6080 27000 6082
rect 24853 6024 24858 6080
rect 24914 6024 27000 6080
rect 24853 6022 27000 6024
rect 24853 6019 24919 6022
rect 2946 6016 3262 6017
rect 2946 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3262 6016
rect 2946 5951 3262 5952
rect 12946 6016 13262 6017
rect 12946 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13262 6016
rect 12946 5951 13262 5952
rect 22946 6016 23262 6017
rect 22946 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23262 6016
rect 26200 5992 27000 6022
rect 22946 5951 23262 5952
rect 20253 5674 20319 5677
rect 20478 5674 20484 5676
rect 20253 5672 20484 5674
rect 20253 5616 20258 5672
rect 20314 5616 20484 5672
rect 20253 5614 20484 5616
rect 20253 5611 20319 5614
rect 20478 5612 20484 5614
rect 20548 5612 20554 5676
rect 24945 5674 25011 5677
rect 26200 5674 27000 5704
rect 24945 5672 27000 5674
rect 24945 5616 24950 5672
rect 25006 5616 27000 5672
rect 24945 5614 27000 5616
rect 24945 5611 25011 5614
rect 26200 5584 27000 5614
rect 7946 5472 8262 5473
rect 7946 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8262 5472
rect 7946 5407 8262 5408
rect 17946 5472 18262 5473
rect 17946 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18262 5472
rect 17946 5407 18262 5408
rect 24761 5266 24827 5269
rect 26200 5266 27000 5296
rect 24761 5264 27000 5266
rect 24761 5208 24766 5264
rect 24822 5208 27000 5264
rect 24761 5206 27000 5208
rect 24761 5203 24827 5206
rect 26200 5176 27000 5206
rect 2946 4928 3262 4929
rect 2946 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3262 4928
rect 2946 4863 3262 4864
rect 12946 4928 13262 4929
rect 12946 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13262 4928
rect 12946 4863 13262 4864
rect 22946 4928 23262 4929
rect 22946 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23262 4928
rect 22946 4863 23262 4864
rect 24853 4858 24919 4861
rect 26200 4858 27000 4888
rect 24853 4856 27000 4858
rect 24853 4800 24858 4856
rect 24914 4800 27000 4856
rect 24853 4798 27000 4800
rect 24853 4795 24919 4798
rect 26200 4768 27000 4798
rect 24945 4450 25011 4453
rect 26200 4450 27000 4480
rect 24945 4448 27000 4450
rect 24945 4392 24950 4448
rect 25006 4392 27000 4448
rect 24945 4390 27000 4392
rect 24945 4387 25011 4390
rect 7946 4384 8262 4385
rect 7946 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8262 4384
rect 7946 4319 8262 4320
rect 17946 4384 18262 4385
rect 17946 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18262 4384
rect 26200 4360 27000 4390
rect 17946 4319 18262 4320
rect 25129 4042 25195 4045
rect 26200 4042 27000 4072
rect 25129 4040 27000 4042
rect 25129 3984 25134 4040
rect 25190 3984 27000 4040
rect 25129 3982 27000 3984
rect 25129 3979 25195 3982
rect 26200 3952 27000 3982
rect 2946 3840 3262 3841
rect 2946 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3262 3840
rect 2946 3775 3262 3776
rect 12946 3840 13262 3841
rect 12946 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13262 3840
rect 12946 3775 13262 3776
rect 22946 3840 23262 3841
rect 22946 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23262 3840
rect 22946 3775 23262 3776
rect 24945 3634 25011 3637
rect 26200 3634 27000 3664
rect 24945 3632 27000 3634
rect 24945 3576 24950 3632
rect 25006 3576 27000 3632
rect 24945 3574 27000 3576
rect 24945 3571 25011 3574
rect 26200 3544 27000 3574
rect 7946 3296 8262 3297
rect 7946 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8262 3296
rect 7946 3231 8262 3232
rect 17946 3296 18262 3297
rect 17946 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18262 3296
rect 17946 3231 18262 3232
rect 24945 3226 25011 3229
rect 26200 3226 27000 3256
rect 24945 3224 27000 3226
rect 24945 3168 24950 3224
rect 25006 3168 27000 3224
rect 24945 3166 27000 3168
rect 24945 3163 25011 3166
rect 26200 3136 27000 3166
rect 24853 2818 24919 2821
rect 26200 2818 27000 2848
rect 24853 2816 27000 2818
rect 24853 2760 24858 2816
rect 24914 2760 27000 2816
rect 24853 2758 27000 2760
rect 24853 2755 24919 2758
rect 2946 2752 3262 2753
rect 2946 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3262 2752
rect 2946 2687 3262 2688
rect 12946 2752 13262 2753
rect 12946 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13262 2752
rect 12946 2687 13262 2688
rect 22946 2752 23262 2753
rect 22946 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23262 2752
rect 26200 2728 27000 2758
rect 22946 2687 23262 2688
rect 24945 2410 25011 2413
rect 26200 2410 27000 2440
rect 24945 2408 27000 2410
rect 24945 2352 24950 2408
rect 25006 2352 27000 2408
rect 24945 2350 27000 2352
rect 24945 2347 25011 2350
rect 26200 2320 27000 2350
rect 7946 2208 8262 2209
rect 7946 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8262 2208
rect 7946 2143 8262 2144
rect 17946 2208 18262 2209
rect 17946 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18262 2208
rect 17946 2143 18262 2144
rect 22185 2002 22251 2005
rect 26200 2002 27000 2032
rect 22185 2000 27000 2002
rect 22185 1944 22190 2000
rect 22246 1944 27000 2000
rect 22185 1942 27000 1944
rect 22185 1939 22251 1942
rect 26200 1912 27000 1942
rect 22093 1594 22159 1597
rect 26200 1594 27000 1624
rect 22093 1592 27000 1594
rect 22093 1536 22098 1592
rect 22154 1536 27000 1592
rect 22093 1534 27000 1536
rect 22093 1531 22159 1534
rect 26200 1504 27000 1534
rect 22093 1186 22159 1189
rect 26200 1186 27000 1216
rect 22093 1184 27000 1186
rect 22093 1128 22098 1184
rect 22154 1128 27000 1184
rect 22093 1126 27000 1128
rect 22093 1123 22159 1126
rect 26200 1096 27000 1126
rect 25037 778 25103 781
rect 26200 778 27000 808
rect 25037 776 27000 778
rect 25037 720 25042 776
rect 25098 720 27000 776
rect 25037 718 27000 720
rect 25037 715 25103 718
rect 26200 688 27000 718
rect 23381 370 23447 373
rect 26200 370 27000 400
rect 23381 368 27000 370
rect 23381 312 23386 368
rect 23442 312 27000 368
rect 23381 310 27000 312
rect 23381 307 23447 310
rect 26200 280 27000 310
<< via3 >>
rect 6500 26012 6564 26076
rect 9628 24788 9692 24852
rect 8892 24652 8956 24716
rect 2952 24508 3016 24512
rect 2952 24452 2956 24508
rect 2956 24452 3012 24508
rect 3012 24452 3016 24508
rect 2952 24448 3016 24452
rect 3032 24508 3096 24512
rect 3032 24452 3036 24508
rect 3036 24452 3092 24508
rect 3092 24452 3096 24508
rect 3032 24448 3096 24452
rect 3112 24508 3176 24512
rect 3112 24452 3116 24508
rect 3116 24452 3172 24508
rect 3172 24452 3176 24508
rect 3112 24448 3176 24452
rect 3192 24508 3256 24512
rect 3192 24452 3196 24508
rect 3196 24452 3252 24508
rect 3252 24452 3256 24508
rect 3192 24448 3256 24452
rect 12952 24508 13016 24512
rect 12952 24452 12956 24508
rect 12956 24452 13012 24508
rect 13012 24452 13016 24508
rect 12952 24448 13016 24452
rect 13032 24508 13096 24512
rect 13032 24452 13036 24508
rect 13036 24452 13092 24508
rect 13092 24452 13096 24508
rect 13032 24448 13096 24452
rect 13112 24508 13176 24512
rect 13112 24452 13116 24508
rect 13116 24452 13172 24508
rect 13172 24452 13176 24508
rect 13112 24448 13176 24452
rect 13192 24508 13256 24512
rect 13192 24452 13196 24508
rect 13196 24452 13252 24508
rect 13252 24452 13256 24508
rect 13192 24448 13256 24452
rect 22952 24508 23016 24512
rect 22952 24452 22956 24508
rect 22956 24452 23012 24508
rect 23012 24452 23016 24508
rect 22952 24448 23016 24452
rect 23032 24508 23096 24512
rect 23032 24452 23036 24508
rect 23036 24452 23092 24508
rect 23092 24452 23096 24508
rect 23032 24448 23096 24452
rect 23112 24508 23176 24512
rect 23112 24452 23116 24508
rect 23116 24452 23172 24508
rect 23172 24452 23176 24508
rect 23112 24448 23176 24452
rect 23192 24508 23256 24512
rect 23192 24452 23196 24508
rect 23196 24452 23252 24508
rect 23252 24452 23256 24508
rect 23192 24448 23256 24452
rect 12020 24244 12084 24308
rect 14964 24108 15028 24172
rect 10364 23972 10428 24036
rect 7952 23964 8016 23968
rect 7952 23908 7956 23964
rect 7956 23908 8012 23964
rect 8012 23908 8016 23964
rect 7952 23904 8016 23908
rect 8032 23964 8096 23968
rect 8032 23908 8036 23964
rect 8036 23908 8092 23964
rect 8092 23908 8096 23964
rect 8032 23904 8096 23908
rect 8112 23964 8176 23968
rect 8112 23908 8116 23964
rect 8116 23908 8172 23964
rect 8172 23908 8176 23964
rect 8112 23904 8176 23908
rect 8192 23964 8256 23968
rect 8192 23908 8196 23964
rect 8196 23908 8252 23964
rect 8252 23908 8256 23964
rect 8192 23904 8256 23908
rect 17952 23964 18016 23968
rect 17952 23908 17956 23964
rect 17956 23908 18012 23964
rect 18012 23908 18016 23964
rect 17952 23904 18016 23908
rect 18032 23964 18096 23968
rect 18032 23908 18036 23964
rect 18036 23908 18092 23964
rect 18092 23908 18096 23964
rect 18032 23904 18096 23908
rect 18112 23964 18176 23968
rect 18112 23908 18116 23964
rect 18116 23908 18172 23964
rect 18172 23908 18176 23964
rect 18112 23904 18176 23908
rect 18192 23964 18256 23968
rect 18192 23908 18196 23964
rect 18196 23908 18252 23964
rect 18252 23908 18256 23964
rect 18192 23904 18256 23908
rect 16252 23836 16316 23900
rect 15148 23564 15212 23628
rect 20116 23428 20180 23492
rect 2952 23420 3016 23424
rect 2952 23364 2956 23420
rect 2956 23364 3012 23420
rect 3012 23364 3016 23420
rect 2952 23360 3016 23364
rect 3032 23420 3096 23424
rect 3032 23364 3036 23420
rect 3036 23364 3092 23420
rect 3092 23364 3096 23420
rect 3032 23360 3096 23364
rect 3112 23420 3176 23424
rect 3112 23364 3116 23420
rect 3116 23364 3172 23420
rect 3172 23364 3176 23420
rect 3112 23360 3176 23364
rect 3192 23420 3256 23424
rect 3192 23364 3196 23420
rect 3196 23364 3252 23420
rect 3252 23364 3256 23420
rect 3192 23360 3256 23364
rect 12952 23420 13016 23424
rect 12952 23364 12956 23420
rect 12956 23364 13012 23420
rect 13012 23364 13016 23420
rect 12952 23360 13016 23364
rect 13032 23420 13096 23424
rect 13032 23364 13036 23420
rect 13036 23364 13092 23420
rect 13092 23364 13096 23420
rect 13032 23360 13096 23364
rect 13112 23420 13176 23424
rect 13112 23364 13116 23420
rect 13116 23364 13172 23420
rect 13172 23364 13176 23420
rect 13112 23360 13176 23364
rect 13192 23420 13256 23424
rect 13192 23364 13196 23420
rect 13196 23364 13252 23420
rect 13252 23364 13256 23420
rect 13192 23360 13256 23364
rect 22952 23420 23016 23424
rect 22952 23364 22956 23420
rect 22956 23364 23012 23420
rect 23012 23364 23016 23420
rect 22952 23360 23016 23364
rect 23032 23420 23096 23424
rect 23032 23364 23036 23420
rect 23036 23364 23092 23420
rect 23092 23364 23096 23420
rect 23032 23360 23096 23364
rect 23112 23420 23176 23424
rect 23112 23364 23116 23420
rect 23116 23364 23172 23420
rect 23172 23364 23176 23420
rect 23112 23360 23176 23364
rect 23192 23420 23256 23424
rect 23192 23364 23196 23420
rect 23196 23364 23252 23420
rect 23252 23364 23256 23420
rect 23192 23360 23256 23364
rect 9444 23292 9508 23356
rect 17356 23156 17420 23220
rect 7952 22876 8016 22880
rect 7952 22820 7956 22876
rect 7956 22820 8012 22876
rect 8012 22820 8016 22876
rect 7952 22816 8016 22820
rect 8032 22876 8096 22880
rect 8032 22820 8036 22876
rect 8036 22820 8092 22876
rect 8092 22820 8096 22876
rect 8032 22816 8096 22820
rect 8112 22876 8176 22880
rect 8112 22820 8116 22876
rect 8116 22820 8172 22876
rect 8172 22820 8176 22876
rect 8112 22816 8176 22820
rect 8192 22876 8256 22880
rect 8192 22820 8196 22876
rect 8196 22820 8252 22876
rect 8252 22820 8256 22876
rect 8192 22816 8256 22820
rect 12388 22748 12452 22812
rect 12572 22748 12636 22812
rect 11100 22612 11164 22676
rect 17724 23020 17788 23084
rect 17952 22876 18016 22880
rect 17952 22820 17956 22876
rect 17956 22820 18012 22876
rect 18012 22820 18016 22876
rect 17952 22816 18016 22820
rect 18032 22876 18096 22880
rect 18032 22820 18036 22876
rect 18036 22820 18092 22876
rect 18092 22820 18096 22876
rect 18032 22816 18096 22820
rect 18112 22876 18176 22880
rect 18112 22820 18116 22876
rect 18116 22820 18172 22876
rect 18172 22820 18176 22876
rect 18112 22816 18176 22820
rect 18192 22876 18256 22880
rect 18192 22820 18196 22876
rect 18196 22820 18252 22876
rect 18252 22820 18256 22876
rect 18192 22816 18256 22820
rect 24532 22536 24596 22540
rect 24532 22480 24582 22536
rect 24582 22480 24596 22536
rect 24532 22476 24596 22480
rect 2952 22332 3016 22336
rect 2952 22276 2956 22332
rect 2956 22276 3012 22332
rect 3012 22276 3016 22332
rect 2952 22272 3016 22276
rect 3032 22332 3096 22336
rect 3032 22276 3036 22332
rect 3036 22276 3092 22332
rect 3092 22276 3096 22332
rect 3032 22272 3096 22276
rect 3112 22332 3176 22336
rect 3112 22276 3116 22332
rect 3116 22276 3172 22332
rect 3172 22276 3176 22332
rect 3112 22272 3176 22276
rect 3192 22332 3256 22336
rect 3192 22276 3196 22332
rect 3196 22276 3252 22332
rect 3252 22276 3256 22332
rect 3192 22272 3256 22276
rect 12952 22332 13016 22336
rect 12952 22276 12956 22332
rect 12956 22276 13012 22332
rect 13012 22276 13016 22332
rect 12952 22272 13016 22276
rect 13032 22332 13096 22336
rect 13032 22276 13036 22332
rect 13036 22276 13092 22332
rect 13092 22276 13096 22332
rect 13032 22272 13096 22276
rect 13112 22332 13176 22336
rect 13112 22276 13116 22332
rect 13116 22276 13172 22332
rect 13172 22276 13176 22332
rect 13112 22272 13176 22276
rect 13192 22332 13256 22336
rect 13192 22276 13196 22332
rect 13196 22276 13252 22332
rect 13252 22276 13256 22332
rect 13192 22272 13256 22276
rect 22952 22332 23016 22336
rect 22952 22276 22956 22332
rect 22956 22276 23012 22332
rect 23012 22276 23016 22332
rect 22952 22272 23016 22276
rect 23032 22332 23096 22336
rect 23032 22276 23036 22332
rect 23036 22276 23092 22332
rect 23092 22276 23096 22332
rect 23032 22272 23096 22276
rect 23112 22332 23176 22336
rect 23112 22276 23116 22332
rect 23116 22276 23172 22332
rect 23172 22276 23176 22332
rect 23112 22272 23176 22276
rect 23192 22332 23256 22336
rect 23192 22276 23196 22332
rect 23196 22276 23252 22332
rect 23252 22276 23256 22332
rect 23192 22272 23256 22276
rect 21036 22068 21100 22132
rect 13492 21856 13556 21860
rect 13492 21800 13542 21856
rect 13542 21800 13556 21856
rect 13492 21796 13556 21800
rect 7952 21788 8016 21792
rect 7952 21732 7956 21788
rect 7956 21732 8012 21788
rect 8012 21732 8016 21788
rect 7952 21728 8016 21732
rect 8032 21788 8096 21792
rect 8032 21732 8036 21788
rect 8036 21732 8092 21788
rect 8092 21732 8096 21788
rect 8032 21728 8096 21732
rect 8112 21788 8176 21792
rect 8112 21732 8116 21788
rect 8116 21732 8172 21788
rect 8172 21732 8176 21788
rect 8112 21728 8176 21732
rect 8192 21788 8256 21792
rect 8192 21732 8196 21788
rect 8196 21732 8252 21788
rect 8252 21732 8256 21788
rect 8192 21728 8256 21732
rect 17952 21788 18016 21792
rect 17952 21732 17956 21788
rect 17956 21732 18012 21788
rect 18012 21732 18016 21788
rect 17952 21728 18016 21732
rect 18032 21788 18096 21792
rect 18032 21732 18036 21788
rect 18036 21732 18092 21788
rect 18092 21732 18096 21788
rect 18032 21728 18096 21732
rect 18112 21788 18176 21792
rect 18112 21732 18116 21788
rect 18116 21732 18172 21788
rect 18172 21732 18176 21788
rect 18112 21728 18176 21732
rect 18192 21788 18256 21792
rect 18192 21732 18196 21788
rect 18196 21732 18252 21788
rect 18252 21732 18256 21788
rect 18192 21728 18256 21732
rect 12572 21660 12636 21724
rect 12388 21252 12452 21316
rect 2952 21244 3016 21248
rect 2952 21188 2956 21244
rect 2956 21188 3012 21244
rect 3012 21188 3016 21244
rect 2952 21184 3016 21188
rect 3032 21244 3096 21248
rect 3032 21188 3036 21244
rect 3036 21188 3092 21244
rect 3092 21188 3096 21244
rect 3032 21184 3096 21188
rect 3112 21244 3176 21248
rect 3112 21188 3116 21244
rect 3116 21188 3172 21244
rect 3172 21188 3176 21244
rect 3112 21184 3176 21188
rect 3192 21244 3256 21248
rect 3192 21188 3196 21244
rect 3196 21188 3252 21244
rect 3252 21188 3256 21244
rect 3192 21184 3256 21188
rect 21404 21524 21468 21588
rect 12952 21244 13016 21248
rect 12952 21188 12956 21244
rect 12956 21188 13012 21244
rect 13012 21188 13016 21244
rect 12952 21184 13016 21188
rect 13032 21244 13096 21248
rect 13032 21188 13036 21244
rect 13036 21188 13092 21244
rect 13092 21188 13096 21244
rect 13032 21184 13096 21188
rect 13112 21244 13176 21248
rect 13112 21188 13116 21244
rect 13116 21188 13172 21244
rect 13172 21188 13176 21244
rect 13112 21184 13176 21188
rect 13192 21244 13256 21248
rect 13192 21188 13196 21244
rect 13196 21188 13252 21244
rect 13252 21188 13256 21244
rect 13192 21184 13256 21188
rect 22952 21244 23016 21248
rect 22952 21188 22956 21244
rect 22956 21188 23012 21244
rect 23012 21188 23016 21244
rect 22952 21184 23016 21188
rect 23032 21244 23096 21248
rect 23032 21188 23036 21244
rect 23036 21188 23092 21244
rect 23092 21188 23096 21244
rect 23032 21184 23096 21188
rect 23112 21244 23176 21248
rect 23112 21188 23116 21244
rect 23116 21188 23172 21244
rect 23172 21188 23176 21244
rect 23112 21184 23176 21188
rect 23192 21244 23256 21248
rect 23192 21188 23196 21244
rect 23196 21188 23252 21244
rect 23252 21188 23256 21244
rect 23192 21184 23256 21188
rect 15148 20904 15212 20908
rect 15148 20848 15198 20904
rect 15198 20848 15212 20904
rect 15148 20844 15212 20848
rect 22692 20980 22756 21044
rect 15884 20768 15948 20772
rect 15884 20712 15898 20768
rect 15898 20712 15948 20768
rect 15884 20708 15948 20712
rect 19564 20768 19628 20772
rect 19564 20712 19578 20768
rect 19578 20712 19628 20768
rect 19564 20708 19628 20712
rect 20852 20768 20916 20772
rect 20852 20712 20866 20768
rect 20866 20712 20916 20768
rect 20852 20708 20916 20712
rect 21220 20708 21284 20772
rect 7952 20700 8016 20704
rect 7952 20644 7956 20700
rect 7956 20644 8012 20700
rect 8012 20644 8016 20700
rect 7952 20640 8016 20644
rect 8032 20700 8096 20704
rect 8032 20644 8036 20700
rect 8036 20644 8092 20700
rect 8092 20644 8096 20700
rect 8032 20640 8096 20644
rect 8112 20700 8176 20704
rect 8112 20644 8116 20700
rect 8116 20644 8172 20700
rect 8172 20644 8176 20700
rect 8112 20640 8176 20644
rect 8192 20700 8256 20704
rect 8192 20644 8196 20700
rect 8196 20644 8252 20700
rect 8252 20644 8256 20700
rect 8192 20640 8256 20644
rect 17952 20700 18016 20704
rect 17952 20644 17956 20700
rect 17956 20644 18012 20700
rect 18012 20644 18016 20700
rect 17952 20640 18016 20644
rect 18032 20700 18096 20704
rect 18032 20644 18036 20700
rect 18036 20644 18092 20700
rect 18092 20644 18096 20700
rect 18032 20640 18096 20644
rect 18112 20700 18176 20704
rect 18112 20644 18116 20700
rect 18116 20644 18172 20700
rect 18172 20644 18176 20700
rect 18112 20640 18176 20644
rect 18192 20700 18256 20704
rect 18192 20644 18196 20700
rect 18196 20644 18252 20700
rect 18252 20644 18256 20700
rect 18192 20640 18256 20644
rect 19748 20300 19812 20364
rect 13676 20164 13740 20228
rect 21036 20224 21100 20228
rect 21036 20168 21050 20224
rect 21050 20168 21100 20224
rect 21036 20164 21100 20168
rect 2952 20156 3016 20160
rect 2952 20100 2956 20156
rect 2956 20100 3012 20156
rect 3012 20100 3016 20156
rect 2952 20096 3016 20100
rect 3032 20156 3096 20160
rect 3032 20100 3036 20156
rect 3036 20100 3092 20156
rect 3092 20100 3096 20156
rect 3032 20096 3096 20100
rect 3112 20156 3176 20160
rect 3112 20100 3116 20156
rect 3116 20100 3172 20156
rect 3172 20100 3176 20156
rect 3112 20096 3176 20100
rect 3192 20156 3256 20160
rect 3192 20100 3196 20156
rect 3196 20100 3252 20156
rect 3252 20100 3256 20156
rect 3192 20096 3256 20100
rect 12952 20156 13016 20160
rect 12952 20100 12956 20156
rect 12956 20100 13012 20156
rect 13012 20100 13016 20156
rect 12952 20096 13016 20100
rect 13032 20156 13096 20160
rect 13032 20100 13036 20156
rect 13036 20100 13092 20156
rect 13092 20100 13096 20156
rect 13032 20096 13096 20100
rect 13112 20156 13176 20160
rect 13112 20100 13116 20156
rect 13116 20100 13172 20156
rect 13172 20100 13176 20156
rect 13112 20096 13176 20100
rect 13192 20156 13256 20160
rect 13192 20100 13196 20156
rect 13196 20100 13252 20156
rect 13252 20100 13256 20156
rect 13192 20096 13256 20100
rect 22952 20156 23016 20160
rect 22952 20100 22956 20156
rect 22956 20100 23012 20156
rect 23012 20100 23016 20156
rect 22952 20096 23016 20100
rect 23032 20156 23096 20160
rect 23032 20100 23036 20156
rect 23036 20100 23092 20156
rect 23092 20100 23096 20156
rect 23032 20096 23096 20100
rect 23112 20156 23176 20160
rect 23112 20100 23116 20156
rect 23116 20100 23172 20156
rect 23172 20100 23176 20156
rect 23112 20096 23176 20100
rect 23192 20156 23256 20160
rect 23192 20100 23196 20156
rect 23196 20100 23252 20156
rect 23252 20100 23256 20156
rect 23192 20096 23256 20100
rect 21036 20028 21100 20092
rect 18460 19756 18524 19820
rect 7952 19612 8016 19616
rect 7952 19556 7956 19612
rect 7956 19556 8012 19612
rect 8012 19556 8016 19612
rect 7952 19552 8016 19556
rect 8032 19612 8096 19616
rect 8032 19556 8036 19612
rect 8036 19556 8092 19612
rect 8092 19556 8096 19612
rect 8032 19552 8096 19556
rect 8112 19612 8176 19616
rect 8112 19556 8116 19612
rect 8116 19556 8172 19612
rect 8172 19556 8176 19612
rect 8112 19552 8176 19556
rect 8192 19612 8256 19616
rect 8192 19556 8196 19612
rect 8196 19556 8252 19612
rect 8252 19556 8256 19612
rect 8192 19552 8256 19556
rect 17952 19612 18016 19616
rect 17952 19556 17956 19612
rect 17956 19556 18012 19612
rect 18012 19556 18016 19612
rect 17952 19552 18016 19556
rect 18032 19612 18096 19616
rect 18032 19556 18036 19612
rect 18036 19556 18092 19612
rect 18092 19556 18096 19612
rect 18032 19552 18096 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 6500 19272 6564 19276
rect 6500 19216 6514 19272
rect 6514 19216 6564 19272
rect 6500 19212 6564 19216
rect 16068 19348 16132 19412
rect 16436 19348 16500 19412
rect 19380 19348 19444 19412
rect 2952 19068 3016 19072
rect 2952 19012 2956 19068
rect 2956 19012 3012 19068
rect 3012 19012 3016 19068
rect 2952 19008 3016 19012
rect 3032 19068 3096 19072
rect 3032 19012 3036 19068
rect 3036 19012 3092 19068
rect 3092 19012 3096 19068
rect 3032 19008 3096 19012
rect 3112 19068 3176 19072
rect 3112 19012 3116 19068
rect 3116 19012 3172 19068
rect 3172 19012 3176 19068
rect 3112 19008 3176 19012
rect 3192 19068 3256 19072
rect 3192 19012 3196 19068
rect 3196 19012 3252 19068
rect 3252 19012 3256 19068
rect 3192 19008 3256 19012
rect 12952 19068 13016 19072
rect 12952 19012 12956 19068
rect 12956 19012 13012 19068
rect 13012 19012 13016 19068
rect 12952 19008 13016 19012
rect 13032 19068 13096 19072
rect 13032 19012 13036 19068
rect 13036 19012 13092 19068
rect 13092 19012 13096 19068
rect 13032 19008 13096 19012
rect 13112 19068 13176 19072
rect 13112 19012 13116 19068
rect 13116 19012 13172 19068
rect 13172 19012 13176 19068
rect 13112 19008 13176 19012
rect 13192 19068 13256 19072
rect 13192 19012 13196 19068
rect 13196 19012 13252 19068
rect 13252 19012 13256 19068
rect 13192 19008 13256 19012
rect 22952 19068 23016 19072
rect 22952 19012 22956 19068
rect 22956 19012 23012 19068
rect 23012 19012 23016 19068
rect 22952 19008 23016 19012
rect 23032 19068 23096 19072
rect 23032 19012 23036 19068
rect 23036 19012 23092 19068
rect 23092 19012 23096 19068
rect 23032 19008 23096 19012
rect 23112 19068 23176 19072
rect 23112 19012 23116 19068
rect 23116 19012 23172 19068
rect 23172 19012 23176 19068
rect 23112 19008 23176 19012
rect 23192 19068 23256 19072
rect 23192 19012 23196 19068
rect 23196 19012 23252 19068
rect 23252 19012 23256 19068
rect 23192 19008 23256 19012
rect 20668 18532 20732 18596
rect 7952 18524 8016 18528
rect 7952 18468 7956 18524
rect 7956 18468 8012 18524
rect 8012 18468 8016 18524
rect 7952 18464 8016 18468
rect 8032 18524 8096 18528
rect 8032 18468 8036 18524
rect 8036 18468 8092 18524
rect 8092 18468 8096 18524
rect 8032 18464 8096 18468
rect 8112 18524 8176 18528
rect 8112 18468 8116 18524
rect 8116 18468 8172 18524
rect 8172 18468 8176 18524
rect 8112 18464 8176 18468
rect 8192 18524 8256 18528
rect 8192 18468 8196 18524
rect 8196 18468 8252 18524
rect 8252 18468 8256 18524
rect 8192 18464 8256 18468
rect 17952 18524 18016 18528
rect 17952 18468 17956 18524
rect 17956 18468 18012 18524
rect 18012 18468 18016 18524
rect 17952 18464 18016 18468
rect 18032 18524 18096 18528
rect 18032 18468 18036 18524
rect 18036 18468 18092 18524
rect 18092 18468 18096 18524
rect 18032 18464 18096 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 9628 17988 9692 18052
rect 2952 17980 3016 17984
rect 2952 17924 2956 17980
rect 2956 17924 3012 17980
rect 3012 17924 3016 17980
rect 2952 17920 3016 17924
rect 3032 17980 3096 17984
rect 3032 17924 3036 17980
rect 3036 17924 3092 17980
rect 3092 17924 3096 17980
rect 3032 17920 3096 17924
rect 3112 17980 3176 17984
rect 3112 17924 3116 17980
rect 3116 17924 3172 17980
rect 3172 17924 3176 17980
rect 3112 17920 3176 17924
rect 3192 17980 3256 17984
rect 3192 17924 3196 17980
rect 3196 17924 3252 17980
rect 3252 17924 3256 17980
rect 3192 17920 3256 17924
rect 12952 17980 13016 17984
rect 12952 17924 12956 17980
rect 12956 17924 13012 17980
rect 13012 17924 13016 17980
rect 12952 17920 13016 17924
rect 13032 17980 13096 17984
rect 13032 17924 13036 17980
rect 13036 17924 13092 17980
rect 13092 17924 13096 17980
rect 13032 17920 13096 17924
rect 13112 17980 13176 17984
rect 13112 17924 13116 17980
rect 13116 17924 13172 17980
rect 13172 17924 13176 17980
rect 13112 17920 13176 17924
rect 13192 17980 13256 17984
rect 13192 17924 13196 17980
rect 13196 17924 13252 17980
rect 13252 17924 13256 17980
rect 13192 17920 13256 17924
rect 17540 17988 17604 18052
rect 23428 17988 23492 18052
rect 22952 17980 23016 17984
rect 22952 17924 22956 17980
rect 22956 17924 23012 17980
rect 23012 17924 23016 17980
rect 22952 17920 23016 17924
rect 23032 17980 23096 17984
rect 23032 17924 23036 17980
rect 23036 17924 23092 17980
rect 23092 17924 23096 17980
rect 23032 17920 23096 17924
rect 23112 17980 23176 17984
rect 23112 17924 23116 17980
rect 23116 17924 23172 17980
rect 23172 17924 23176 17980
rect 23112 17920 23176 17924
rect 23192 17980 23256 17984
rect 23192 17924 23196 17980
rect 23196 17924 23252 17980
rect 23252 17924 23256 17980
rect 23192 17920 23256 17924
rect 11100 17716 11164 17780
rect 7952 17436 8016 17440
rect 7952 17380 7956 17436
rect 7956 17380 8012 17436
rect 8012 17380 8016 17436
rect 7952 17376 8016 17380
rect 8032 17436 8096 17440
rect 8032 17380 8036 17436
rect 8036 17380 8092 17436
rect 8092 17380 8096 17436
rect 8032 17376 8096 17380
rect 8112 17436 8176 17440
rect 8112 17380 8116 17436
rect 8116 17380 8172 17436
rect 8172 17380 8176 17436
rect 8112 17376 8176 17380
rect 8192 17436 8256 17440
rect 8192 17380 8196 17436
rect 8196 17380 8252 17436
rect 8252 17380 8256 17436
rect 8192 17376 8256 17380
rect 17952 17436 18016 17440
rect 17952 17380 17956 17436
rect 17956 17380 18012 17436
rect 18012 17380 18016 17436
rect 17952 17376 18016 17380
rect 18032 17436 18096 17440
rect 18032 17380 18036 17436
rect 18036 17380 18092 17436
rect 18092 17380 18096 17436
rect 18032 17376 18096 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 19196 17308 19260 17372
rect 2952 16892 3016 16896
rect 2952 16836 2956 16892
rect 2956 16836 3012 16892
rect 3012 16836 3016 16892
rect 2952 16832 3016 16836
rect 3032 16892 3096 16896
rect 3032 16836 3036 16892
rect 3036 16836 3092 16892
rect 3092 16836 3096 16892
rect 3032 16832 3096 16836
rect 3112 16892 3176 16896
rect 3112 16836 3116 16892
rect 3116 16836 3172 16892
rect 3172 16836 3176 16892
rect 3112 16832 3176 16836
rect 3192 16892 3256 16896
rect 3192 16836 3196 16892
rect 3196 16836 3252 16892
rect 3252 16836 3256 16892
rect 3192 16832 3256 16836
rect 12952 16892 13016 16896
rect 12952 16836 12956 16892
rect 12956 16836 13012 16892
rect 13012 16836 13016 16892
rect 12952 16832 13016 16836
rect 13032 16892 13096 16896
rect 13032 16836 13036 16892
rect 13036 16836 13092 16892
rect 13092 16836 13096 16892
rect 13032 16832 13096 16836
rect 13112 16892 13176 16896
rect 13112 16836 13116 16892
rect 13116 16836 13172 16892
rect 13172 16836 13176 16892
rect 13112 16832 13176 16836
rect 13192 16892 13256 16896
rect 13192 16836 13196 16892
rect 13196 16836 13252 16892
rect 13252 16836 13256 16892
rect 13192 16832 13256 16836
rect 22952 16892 23016 16896
rect 22952 16836 22956 16892
rect 22956 16836 23012 16892
rect 23012 16836 23016 16892
rect 22952 16832 23016 16836
rect 23032 16892 23096 16896
rect 23032 16836 23036 16892
rect 23036 16836 23092 16892
rect 23092 16836 23096 16892
rect 23032 16832 23096 16836
rect 23112 16892 23176 16896
rect 23112 16836 23116 16892
rect 23116 16836 23172 16892
rect 23172 16836 23176 16892
rect 23112 16832 23176 16836
rect 23192 16892 23256 16896
rect 23192 16836 23196 16892
rect 23196 16836 23252 16892
rect 23252 16836 23256 16892
rect 23192 16832 23256 16836
rect 16620 16764 16684 16828
rect 19564 16764 19628 16828
rect 8892 16492 8956 16556
rect 17724 16356 17788 16420
rect 7952 16348 8016 16352
rect 7952 16292 7956 16348
rect 7956 16292 8012 16348
rect 8012 16292 8016 16348
rect 7952 16288 8016 16292
rect 8032 16348 8096 16352
rect 8032 16292 8036 16348
rect 8036 16292 8092 16348
rect 8092 16292 8096 16348
rect 8032 16288 8096 16292
rect 8112 16348 8176 16352
rect 8112 16292 8116 16348
rect 8116 16292 8172 16348
rect 8172 16292 8176 16348
rect 8112 16288 8176 16292
rect 8192 16348 8256 16352
rect 8192 16292 8196 16348
rect 8196 16292 8252 16348
rect 8252 16292 8256 16348
rect 8192 16288 8256 16292
rect 17952 16348 18016 16352
rect 17952 16292 17956 16348
rect 17956 16292 18012 16348
rect 18012 16292 18016 16348
rect 17952 16288 18016 16292
rect 18032 16348 18096 16352
rect 18032 16292 18036 16348
rect 18036 16292 18092 16348
rect 18092 16292 18096 16348
rect 18032 16288 18096 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 19748 15812 19812 15876
rect 2952 15804 3016 15808
rect 2952 15748 2956 15804
rect 2956 15748 3012 15804
rect 3012 15748 3016 15804
rect 2952 15744 3016 15748
rect 3032 15804 3096 15808
rect 3032 15748 3036 15804
rect 3036 15748 3092 15804
rect 3092 15748 3096 15804
rect 3032 15744 3096 15748
rect 3112 15804 3176 15808
rect 3112 15748 3116 15804
rect 3116 15748 3172 15804
rect 3172 15748 3176 15804
rect 3112 15744 3176 15748
rect 3192 15804 3256 15808
rect 3192 15748 3196 15804
rect 3196 15748 3252 15804
rect 3252 15748 3256 15804
rect 3192 15744 3256 15748
rect 12952 15804 13016 15808
rect 12952 15748 12956 15804
rect 12956 15748 13012 15804
rect 13012 15748 13016 15804
rect 12952 15744 13016 15748
rect 13032 15804 13096 15808
rect 13032 15748 13036 15804
rect 13036 15748 13092 15804
rect 13092 15748 13096 15804
rect 13032 15744 13096 15748
rect 13112 15804 13176 15808
rect 13112 15748 13116 15804
rect 13116 15748 13172 15804
rect 13172 15748 13176 15804
rect 13112 15744 13176 15748
rect 13192 15804 13256 15808
rect 13192 15748 13196 15804
rect 13196 15748 13252 15804
rect 13252 15748 13256 15804
rect 13192 15744 13256 15748
rect 22952 15804 23016 15808
rect 22952 15748 22956 15804
rect 22956 15748 23012 15804
rect 23012 15748 23016 15804
rect 22952 15744 23016 15748
rect 23032 15804 23096 15808
rect 23032 15748 23036 15804
rect 23036 15748 23092 15804
rect 23092 15748 23096 15804
rect 23032 15744 23096 15748
rect 23112 15804 23176 15808
rect 23112 15748 23116 15804
rect 23116 15748 23172 15804
rect 23172 15748 23176 15804
rect 23112 15744 23176 15748
rect 23192 15804 23256 15808
rect 23192 15748 23196 15804
rect 23196 15748 23252 15804
rect 23252 15748 23256 15804
rect 23192 15744 23256 15748
rect 20668 15676 20732 15740
rect 9444 15600 9508 15604
rect 9444 15544 9458 15600
rect 9458 15544 9508 15600
rect 9444 15540 9508 15544
rect 24532 15540 24596 15604
rect 19380 15404 19444 15468
rect 22692 15268 22756 15332
rect 7952 15260 8016 15264
rect 7952 15204 7956 15260
rect 7956 15204 8012 15260
rect 8012 15204 8016 15260
rect 7952 15200 8016 15204
rect 8032 15260 8096 15264
rect 8032 15204 8036 15260
rect 8036 15204 8092 15260
rect 8092 15204 8096 15260
rect 8032 15200 8096 15204
rect 8112 15260 8176 15264
rect 8112 15204 8116 15260
rect 8116 15204 8172 15260
rect 8172 15204 8176 15260
rect 8112 15200 8176 15204
rect 8192 15260 8256 15264
rect 8192 15204 8196 15260
rect 8196 15204 8252 15260
rect 8252 15204 8256 15260
rect 8192 15200 8256 15204
rect 17952 15260 18016 15264
rect 17952 15204 17956 15260
rect 17956 15204 18012 15260
rect 18012 15204 18016 15260
rect 17952 15200 18016 15204
rect 18032 15260 18096 15264
rect 18032 15204 18036 15260
rect 18036 15204 18092 15260
rect 18092 15204 18096 15260
rect 18032 15200 18096 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 14964 15132 15028 15196
rect 10364 14996 10428 15060
rect 16620 14996 16684 15060
rect 22324 14860 22388 14924
rect 2952 14716 3016 14720
rect 2952 14660 2956 14716
rect 2956 14660 3012 14716
rect 3012 14660 3016 14716
rect 2952 14656 3016 14660
rect 3032 14716 3096 14720
rect 3032 14660 3036 14716
rect 3036 14660 3092 14716
rect 3092 14660 3096 14716
rect 3032 14656 3096 14660
rect 3112 14716 3176 14720
rect 3112 14660 3116 14716
rect 3116 14660 3172 14716
rect 3172 14660 3176 14716
rect 3112 14656 3176 14660
rect 3192 14716 3256 14720
rect 3192 14660 3196 14716
rect 3196 14660 3252 14716
rect 3252 14660 3256 14716
rect 3192 14656 3256 14660
rect 12952 14716 13016 14720
rect 12952 14660 12956 14716
rect 12956 14660 13012 14716
rect 13012 14660 13016 14716
rect 12952 14656 13016 14660
rect 13032 14716 13096 14720
rect 13032 14660 13036 14716
rect 13036 14660 13092 14716
rect 13092 14660 13096 14716
rect 13032 14656 13096 14660
rect 13112 14716 13176 14720
rect 13112 14660 13116 14716
rect 13116 14660 13172 14716
rect 13172 14660 13176 14716
rect 13112 14656 13176 14660
rect 13192 14716 13256 14720
rect 13192 14660 13196 14716
rect 13196 14660 13252 14716
rect 13252 14660 13256 14716
rect 13192 14656 13256 14660
rect 22952 14716 23016 14720
rect 22952 14660 22956 14716
rect 22956 14660 23012 14716
rect 23012 14660 23016 14716
rect 22952 14656 23016 14660
rect 23032 14716 23096 14720
rect 23032 14660 23036 14716
rect 23036 14660 23092 14716
rect 23092 14660 23096 14716
rect 23032 14656 23096 14660
rect 23112 14716 23176 14720
rect 23112 14660 23116 14716
rect 23116 14660 23172 14716
rect 23172 14660 23176 14716
rect 23112 14656 23176 14660
rect 23192 14716 23256 14720
rect 23192 14660 23196 14716
rect 23196 14660 23252 14716
rect 23252 14660 23256 14716
rect 23192 14656 23256 14660
rect 21956 14452 22020 14516
rect 7952 14172 8016 14176
rect 7952 14116 7956 14172
rect 7956 14116 8012 14172
rect 8012 14116 8016 14172
rect 7952 14112 8016 14116
rect 8032 14172 8096 14176
rect 8032 14116 8036 14172
rect 8036 14116 8092 14172
rect 8092 14116 8096 14172
rect 8032 14112 8096 14116
rect 8112 14172 8176 14176
rect 8112 14116 8116 14172
rect 8116 14116 8172 14172
rect 8172 14116 8176 14172
rect 8112 14112 8176 14116
rect 8192 14172 8256 14176
rect 8192 14116 8196 14172
rect 8196 14116 8252 14172
rect 8252 14116 8256 14172
rect 8192 14112 8256 14116
rect 17952 14172 18016 14176
rect 17952 14116 17956 14172
rect 17956 14116 18012 14172
rect 18012 14116 18016 14172
rect 17952 14112 18016 14116
rect 18032 14172 18096 14176
rect 18032 14116 18036 14172
rect 18036 14116 18092 14172
rect 18092 14116 18096 14172
rect 18032 14112 18096 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 12020 13968 12084 13972
rect 12020 13912 12034 13968
rect 12034 13912 12084 13968
rect 12020 13908 12084 13912
rect 17540 13968 17604 13972
rect 17540 13912 17554 13968
rect 17554 13912 17604 13968
rect 17540 13908 17604 13912
rect 21404 13908 21468 13972
rect 20484 13772 20548 13836
rect 17356 13636 17420 13700
rect 2952 13628 3016 13632
rect 2952 13572 2956 13628
rect 2956 13572 3012 13628
rect 3012 13572 3016 13628
rect 2952 13568 3016 13572
rect 3032 13628 3096 13632
rect 3032 13572 3036 13628
rect 3036 13572 3092 13628
rect 3092 13572 3096 13628
rect 3032 13568 3096 13572
rect 3112 13628 3176 13632
rect 3112 13572 3116 13628
rect 3116 13572 3172 13628
rect 3172 13572 3176 13628
rect 3112 13568 3176 13572
rect 3192 13628 3256 13632
rect 3192 13572 3196 13628
rect 3196 13572 3252 13628
rect 3252 13572 3256 13628
rect 3192 13568 3256 13572
rect 12952 13628 13016 13632
rect 12952 13572 12956 13628
rect 12956 13572 13012 13628
rect 13012 13572 13016 13628
rect 12952 13568 13016 13572
rect 13032 13628 13096 13632
rect 13032 13572 13036 13628
rect 13036 13572 13092 13628
rect 13092 13572 13096 13628
rect 13032 13568 13096 13572
rect 13112 13628 13176 13632
rect 13112 13572 13116 13628
rect 13116 13572 13172 13628
rect 13172 13572 13176 13628
rect 13112 13568 13176 13572
rect 13192 13628 13256 13632
rect 13192 13572 13196 13628
rect 13196 13572 13252 13628
rect 13252 13572 13256 13628
rect 13192 13568 13256 13572
rect 22952 13628 23016 13632
rect 22952 13572 22956 13628
rect 22956 13572 23012 13628
rect 23012 13572 23016 13628
rect 22952 13568 23016 13572
rect 23032 13628 23096 13632
rect 23032 13572 23036 13628
rect 23036 13572 23092 13628
rect 23092 13572 23096 13628
rect 23032 13568 23096 13572
rect 23112 13628 23176 13632
rect 23112 13572 23116 13628
rect 23116 13572 23172 13628
rect 23172 13572 23176 13628
rect 23112 13568 23176 13572
rect 23192 13628 23256 13632
rect 23192 13572 23196 13628
rect 23196 13572 23252 13628
rect 23252 13572 23256 13628
rect 23192 13568 23256 13572
rect 13676 13500 13740 13564
rect 17724 13500 17788 13564
rect 21036 13228 21100 13292
rect 7952 13084 8016 13088
rect 7952 13028 7956 13084
rect 7956 13028 8012 13084
rect 8012 13028 8016 13084
rect 7952 13024 8016 13028
rect 8032 13084 8096 13088
rect 8032 13028 8036 13084
rect 8036 13028 8092 13084
rect 8092 13028 8096 13084
rect 8032 13024 8096 13028
rect 8112 13084 8176 13088
rect 8112 13028 8116 13084
rect 8116 13028 8172 13084
rect 8172 13028 8176 13084
rect 8112 13024 8176 13028
rect 8192 13084 8256 13088
rect 8192 13028 8196 13084
rect 8196 13028 8252 13084
rect 8252 13028 8256 13084
rect 8192 13024 8256 13028
rect 17952 13084 18016 13088
rect 17952 13028 17956 13084
rect 17956 13028 18012 13084
rect 18012 13028 18016 13084
rect 17952 13024 18016 13028
rect 18032 13084 18096 13088
rect 18032 13028 18036 13084
rect 18036 13028 18092 13084
rect 18092 13028 18096 13084
rect 18032 13024 18096 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 2952 12540 3016 12544
rect 2952 12484 2956 12540
rect 2956 12484 3012 12540
rect 3012 12484 3016 12540
rect 2952 12480 3016 12484
rect 3032 12540 3096 12544
rect 3032 12484 3036 12540
rect 3036 12484 3092 12540
rect 3092 12484 3096 12540
rect 3032 12480 3096 12484
rect 3112 12540 3176 12544
rect 3112 12484 3116 12540
rect 3116 12484 3172 12540
rect 3172 12484 3176 12540
rect 3112 12480 3176 12484
rect 3192 12540 3256 12544
rect 3192 12484 3196 12540
rect 3196 12484 3252 12540
rect 3252 12484 3256 12540
rect 3192 12480 3256 12484
rect 12952 12540 13016 12544
rect 12952 12484 12956 12540
rect 12956 12484 13012 12540
rect 13012 12484 13016 12540
rect 12952 12480 13016 12484
rect 13032 12540 13096 12544
rect 13032 12484 13036 12540
rect 13036 12484 13092 12540
rect 13092 12484 13096 12540
rect 13032 12480 13096 12484
rect 13112 12540 13176 12544
rect 13112 12484 13116 12540
rect 13116 12484 13172 12540
rect 13172 12484 13176 12540
rect 13112 12480 13176 12484
rect 13192 12540 13256 12544
rect 13192 12484 13196 12540
rect 13196 12484 13252 12540
rect 13252 12484 13256 12540
rect 13192 12480 13256 12484
rect 22952 12540 23016 12544
rect 22952 12484 22956 12540
rect 22956 12484 23012 12540
rect 23012 12484 23016 12540
rect 22952 12480 23016 12484
rect 23032 12540 23096 12544
rect 23032 12484 23036 12540
rect 23036 12484 23092 12540
rect 23092 12484 23096 12540
rect 23032 12480 23096 12484
rect 23112 12540 23176 12544
rect 23112 12484 23116 12540
rect 23116 12484 23172 12540
rect 23172 12484 23176 12540
rect 23112 12480 23176 12484
rect 23192 12540 23256 12544
rect 23192 12484 23196 12540
rect 23196 12484 23252 12540
rect 23252 12484 23256 12540
rect 23192 12480 23256 12484
rect 20852 12412 20916 12476
rect 7952 11996 8016 12000
rect 7952 11940 7956 11996
rect 7956 11940 8012 11996
rect 8012 11940 8016 11996
rect 7952 11936 8016 11940
rect 8032 11996 8096 12000
rect 8032 11940 8036 11996
rect 8036 11940 8092 11996
rect 8092 11940 8096 11996
rect 8032 11936 8096 11940
rect 8112 11996 8176 12000
rect 8112 11940 8116 11996
rect 8116 11940 8172 11996
rect 8172 11940 8176 11996
rect 8112 11936 8176 11940
rect 8192 11996 8256 12000
rect 8192 11940 8196 11996
rect 8196 11940 8252 11996
rect 8252 11940 8256 11996
rect 8192 11936 8256 11940
rect 17952 11996 18016 12000
rect 17952 11940 17956 11996
rect 17956 11940 18012 11996
rect 18012 11940 18016 11996
rect 17952 11936 18016 11940
rect 18032 11996 18096 12000
rect 18032 11940 18036 11996
rect 18036 11940 18092 11996
rect 18092 11940 18096 11996
rect 18032 11936 18096 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 17724 11596 17788 11660
rect 2952 11452 3016 11456
rect 2952 11396 2956 11452
rect 2956 11396 3012 11452
rect 3012 11396 3016 11452
rect 2952 11392 3016 11396
rect 3032 11452 3096 11456
rect 3032 11396 3036 11452
rect 3036 11396 3092 11452
rect 3092 11396 3096 11452
rect 3032 11392 3096 11396
rect 3112 11452 3176 11456
rect 3112 11396 3116 11452
rect 3116 11396 3172 11452
rect 3172 11396 3176 11452
rect 3112 11392 3176 11396
rect 3192 11452 3256 11456
rect 3192 11396 3196 11452
rect 3196 11396 3252 11452
rect 3252 11396 3256 11452
rect 3192 11392 3256 11396
rect 12952 11452 13016 11456
rect 12952 11396 12956 11452
rect 12956 11396 13012 11452
rect 13012 11396 13016 11452
rect 12952 11392 13016 11396
rect 13032 11452 13096 11456
rect 13032 11396 13036 11452
rect 13036 11396 13092 11452
rect 13092 11396 13096 11452
rect 13032 11392 13096 11396
rect 13112 11452 13176 11456
rect 13112 11396 13116 11452
rect 13116 11396 13172 11452
rect 13172 11396 13176 11452
rect 13112 11392 13176 11396
rect 13192 11452 13256 11456
rect 13192 11396 13196 11452
rect 13196 11396 13252 11452
rect 13252 11396 13256 11452
rect 13192 11392 13256 11396
rect 22952 11452 23016 11456
rect 22952 11396 22956 11452
rect 22956 11396 23012 11452
rect 23012 11396 23016 11452
rect 22952 11392 23016 11396
rect 23032 11452 23096 11456
rect 23032 11396 23036 11452
rect 23036 11396 23092 11452
rect 23092 11396 23096 11452
rect 23032 11392 23096 11396
rect 23112 11452 23176 11456
rect 23112 11396 23116 11452
rect 23116 11396 23172 11452
rect 23172 11396 23176 11452
rect 23112 11392 23176 11396
rect 23192 11452 23256 11456
rect 23192 11396 23196 11452
rect 23196 11396 23252 11452
rect 23252 11396 23256 11452
rect 23192 11392 23256 11396
rect 16252 11324 16316 11388
rect 18460 11052 18524 11116
rect 20116 11052 20180 11116
rect 7952 10908 8016 10912
rect 7952 10852 7956 10908
rect 7956 10852 8012 10908
rect 8012 10852 8016 10908
rect 7952 10848 8016 10852
rect 8032 10908 8096 10912
rect 8032 10852 8036 10908
rect 8036 10852 8092 10908
rect 8092 10852 8096 10908
rect 8032 10848 8096 10852
rect 8112 10908 8176 10912
rect 8112 10852 8116 10908
rect 8116 10852 8172 10908
rect 8172 10852 8176 10908
rect 8112 10848 8176 10852
rect 8192 10908 8256 10912
rect 8192 10852 8196 10908
rect 8196 10852 8252 10908
rect 8252 10852 8256 10908
rect 8192 10848 8256 10852
rect 17952 10908 18016 10912
rect 17952 10852 17956 10908
rect 17956 10852 18012 10908
rect 18012 10852 18016 10908
rect 17952 10848 18016 10852
rect 18032 10908 18096 10912
rect 18032 10852 18036 10908
rect 18036 10852 18092 10908
rect 18092 10852 18096 10908
rect 18032 10848 18096 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 23428 10644 23492 10708
rect 2952 10364 3016 10368
rect 2952 10308 2956 10364
rect 2956 10308 3012 10364
rect 3012 10308 3016 10364
rect 2952 10304 3016 10308
rect 3032 10364 3096 10368
rect 3032 10308 3036 10364
rect 3036 10308 3092 10364
rect 3092 10308 3096 10364
rect 3032 10304 3096 10308
rect 3112 10364 3176 10368
rect 3112 10308 3116 10364
rect 3116 10308 3172 10364
rect 3172 10308 3176 10364
rect 3112 10304 3176 10308
rect 3192 10364 3256 10368
rect 3192 10308 3196 10364
rect 3196 10308 3252 10364
rect 3252 10308 3256 10364
rect 3192 10304 3256 10308
rect 12952 10364 13016 10368
rect 12952 10308 12956 10364
rect 12956 10308 13012 10364
rect 13012 10308 13016 10364
rect 12952 10304 13016 10308
rect 13032 10364 13096 10368
rect 13032 10308 13036 10364
rect 13036 10308 13092 10364
rect 13092 10308 13096 10364
rect 13032 10304 13096 10308
rect 13112 10364 13176 10368
rect 13112 10308 13116 10364
rect 13116 10308 13172 10364
rect 13172 10308 13176 10364
rect 13112 10304 13176 10308
rect 13192 10364 13256 10368
rect 13192 10308 13196 10364
rect 13196 10308 13252 10364
rect 13252 10308 13256 10364
rect 13192 10304 13256 10308
rect 22952 10364 23016 10368
rect 22952 10308 22956 10364
rect 22956 10308 23012 10364
rect 23012 10308 23016 10364
rect 22952 10304 23016 10308
rect 23032 10364 23096 10368
rect 23032 10308 23036 10364
rect 23036 10308 23092 10364
rect 23092 10308 23096 10364
rect 23032 10304 23096 10308
rect 23112 10364 23176 10368
rect 23112 10308 23116 10364
rect 23116 10308 23172 10364
rect 23172 10308 23176 10364
rect 23112 10304 23176 10308
rect 23192 10364 23256 10368
rect 23192 10308 23196 10364
rect 23196 10308 23252 10364
rect 23252 10308 23256 10364
rect 23192 10304 23256 10308
rect 16068 10236 16132 10300
rect 7952 9820 8016 9824
rect 7952 9764 7956 9820
rect 7956 9764 8012 9820
rect 8012 9764 8016 9820
rect 7952 9760 8016 9764
rect 8032 9820 8096 9824
rect 8032 9764 8036 9820
rect 8036 9764 8092 9820
rect 8092 9764 8096 9820
rect 8032 9760 8096 9764
rect 8112 9820 8176 9824
rect 8112 9764 8116 9820
rect 8116 9764 8172 9820
rect 8172 9764 8176 9820
rect 8112 9760 8176 9764
rect 8192 9820 8256 9824
rect 8192 9764 8196 9820
rect 8196 9764 8252 9820
rect 8252 9764 8256 9820
rect 8192 9760 8256 9764
rect 17952 9820 18016 9824
rect 17952 9764 17956 9820
rect 17956 9764 18012 9820
rect 18012 9764 18016 9820
rect 17952 9760 18016 9764
rect 18032 9820 18096 9824
rect 18032 9764 18036 9820
rect 18036 9764 18092 9820
rect 18092 9764 18096 9820
rect 18032 9760 18096 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 21220 9752 21284 9756
rect 21220 9696 21270 9752
rect 21270 9696 21284 9752
rect 21220 9692 21284 9696
rect 15884 9420 15948 9484
rect 2952 9276 3016 9280
rect 2952 9220 2956 9276
rect 2956 9220 3012 9276
rect 3012 9220 3016 9276
rect 2952 9216 3016 9220
rect 3032 9276 3096 9280
rect 3032 9220 3036 9276
rect 3036 9220 3092 9276
rect 3092 9220 3096 9276
rect 3032 9216 3096 9220
rect 3112 9276 3176 9280
rect 3112 9220 3116 9276
rect 3116 9220 3172 9276
rect 3172 9220 3176 9276
rect 3112 9216 3176 9220
rect 3192 9276 3256 9280
rect 3192 9220 3196 9276
rect 3196 9220 3252 9276
rect 3252 9220 3256 9276
rect 3192 9216 3256 9220
rect 12952 9276 13016 9280
rect 12952 9220 12956 9276
rect 12956 9220 13012 9276
rect 13012 9220 13016 9276
rect 12952 9216 13016 9220
rect 13032 9276 13096 9280
rect 13032 9220 13036 9276
rect 13036 9220 13092 9276
rect 13092 9220 13096 9276
rect 13032 9216 13096 9220
rect 13112 9276 13176 9280
rect 13112 9220 13116 9276
rect 13116 9220 13172 9276
rect 13172 9220 13176 9276
rect 13112 9216 13176 9220
rect 13192 9276 13256 9280
rect 13192 9220 13196 9276
rect 13196 9220 13252 9276
rect 13252 9220 13256 9276
rect 13192 9216 13256 9220
rect 22952 9276 23016 9280
rect 22952 9220 22956 9276
rect 22956 9220 23012 9276
rect 23012 9220 23016 9276
rect 22952 9216 23016 9220
rect 23032 9276 23096 9280
rect 23032 9220 23036 9276
rect 23036 9220 23092 9276
rect 23092 9220 23096 9276
rect 23032 9216 23096 9220
rect 23112 9276 23176 9280
rect 23112 9220 23116 9276
rect 23116 9220 23172 9276
rect 23172 9220 23176 9276
rect 23112 9216 23176 9220
rect 23192 9276 23256 9280
rect 23192 9220 23196 9276
rect 23196 9220 23252 9276
rect 23252 9220 23256 9276
rect 23192 9216 23256 9220
rect 7952 8732 8016 8736
rect 7952 8676 7956 8732
rect 7956 8676 8012 8732
rect 8012 8676 8016 8732
rect 7952 8672 8016 8676
rect 8032 8732 8096 8736
rect 8032 8676 8036 8732
rect 8036 8676 8092 8732
rect 8092 8676 8096 8732
rect 8032 8672 8096 8676
rect 8112 8732 8176 8736
rect 8112 8676 8116 8732
rect 8116 8676 8172 8732
rect 8172 8676 8176 8732
rect 8112 8672 8176 8676
rect 8192 8732 8256 8736
rect 8192 8676 8196 8732
rect 8196 8676 8252 8732
rect 8252 8676 8256 8732
rect 8192 8672 8256 8676
rect 17952 8732 18016 8736
rect 17952 8676 17956 8732
rect 17956 8676 18012 8732
rect 18012 8676 18016 8732
rect 17952 8672 18016 8676
rect 18032 8732 18096 8736
rect 18032 8676 18036 8732
rect 18036 8676 18092 8732
rect 18092 8676 18096 8732
rect 18032 8672 18096 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 16436 8332 16500 8396
rect 21956 8392 22020 8396
rect 21956 8336 22006 8392
rect 22006 8336 22020 8392
rect 21956 8332 22020 8336
rect 2952 8188 3016 8192
rect 2952 8132 2956 8188
rect 2956 8132 3012 8188
rect 3012 8132 3016 8188
rect 2952 8128 3016 8132
rect 3032 8188 3096 8192
rect 3032 8132 3036 8188
rect 3036 8132 3092 8188
rect 3092 8132 3096 8188
rect 3032 8128 3096 8132
rect 3112 8188 3176 8192
rect 3112 8132 3116 8188
rect 3116 8132 3172 8188
rect 3172 8132 3176 8188
rect 3112 8128 3176 8132
rect 3192 8188 3256 8192
rect 3192 8132 3196 8188
rect 3196 8132 3252 8188
rect 3252 8132 3256 8188
rect 3192 8128 3256 8132
rect 12952 8188 13016 8192
rect 12952 8132 12956 8188
rect 12956 8132 13012 8188
rect 13012 8132 13016 8188
rect 12952 8128 13016 8132
rect 13032 8188 13096 8192
rect 13032 8132 13036 8188
rect 13036 8132 13092 8188
rect 13092 8132 13096 8188
rect 13032 8128 13096 8132
rect 13112 8188 13176 8192
rect 13112 8132 13116 8188
rect 13116 8132 13172 8188
rect 13172 8132 13176 8188
rect 13112 8128 13176 8132
rect 13192 8188 13256 8192
rect 13192 8132 13196 8188
rect 13196 8132 13252 8188
rect 13252 8132 13256 8188
rect 13192 8128 13256 8132
rect 22952 8188 23016 8192
rect 22952 8132 22956 8188
rect 22956 8132 23012 8188
rect 23012 8132 23016 8188
rect 22952 8128 23016 8132
rect 23032 8188 23096 8192
rect 23032 8132 23036 8188
rect 23036 8132 23092 8188
rect 23092 8132 23096 8188
rect 23032 8128 23096 8132
rect 23112 8188 23176 8192
rect 23112 8132 23116 8188
rect 23116 8132 23172 8188
rect 23172 8132 23176 8188
rect 23112 8128 23176 8132
rect 23192 8188 23256 8192
rect 23192 8132 23196 8188
rect 23196 8132 23252 8188
rect 23252 8132 23256 8188
rect 23192 8128 23256 8132
rect 19196 7924 19260 7988
rect 13492 7788 13556 7852
rect 7952 7644 8016 7648
rect 7952 7588 7956 7644
rect 7956 7588 8012 7644
rect 8012 7588 8016 7644
rect 7952 7584 8016 7588
rect 8032 7644 8096 7648
rect 8032 7588 8036 7644
rect 8036 7588 8092 7644
rect 8092 7588 8096 7644
rect 8032 7584 8096 7588
rect 8112 7644 8176 7648
rect 8112 7588 8116 7644
rect 8116 7588 8172 7644
rect 8172 7588 8176 7644
rect 8112 7584 8176 7588
rect 8192 7644 8256 7648
rect 8192 7588 8196 7644
rect 8196 7588 8252 7644
rect 8252 7588 8256 7644
rect 8192 7584 8256 7588
rect 17952 7644 18016 7648
rect 17952 7588 17956 7644
rect 17956 7588 18012 7644
rect 18012 7588 18016 7644
rect 17952 7584 18016 7588
rect 18032 7644 18096 7648
rect 18032 7588 18036 7644
rect 18036 7588 18092 7644
rect 18092 7588 18096 7644
rect 18032 7584 18096 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 2952 7100 3016 7104
rect 2952 7044 2956 7100
rect 2956 7044 3012 7100
rect 3012 7044 3016 7100
rect 2952 7040 3016 7044
rect 3032 7100 3096 7104
rect 3032 7044 3036 7100
rect 3036 7044 3092 7100
rect 3092 7044 3096 7100
rect 3032 7040 3096 7044
rect 3112 7100 3176 7104
rect 3112 7044 3116 7100
rect 3116 7044 3172 7100
rect 3172 7044 3176 7100
rect 3112 7040 3176 7044
rect 3192 7100 3256 7104
rect 3192 7044 3196 7100
rect 3196 7044 3252 7100
rect 3252 7044 3256 7100
rect 3192 7040 3256 7044
rect 12952 7100 13016 7104
rect 12952 7044 12956 7100
rect 12956 7044 13012 7100
rect 13012 7044 13016 7100
rect 12952 7040 13016 7044
rect 13032 7100 13096 7104
rect 13032 7044 13036 7100
rect 13036 7044 13092 7100
rect 13092 7044 13096 7100
rect 13032 7040 13096 7044
rect 13112 7100 13176 7104
rect 13112 7044 13116 7100
rect 13116 7044 13172 7100
rect 13172 7044 13176 7100
rect 13112 7040 13176 7044
rect 13192 7100 13256 7104
rect 13192 7044 13196 7100
rect 13196 7044 13252 7100
rect 13252 7044 13256 7100
rect 13192 7040 13256 7044
rect 22952 7100 23016 7104
rect 22952 7044 22956 7100
rect 22956 7044 23012 7100
rect 23012 7044 23016 7100
rect 22952 7040 23016 7044
rect 23032 7100 23096 7104
rect 23032 7044 23036 7100
rect 23036 7044 23092 7100
rect 23092 7044 23096 7100
rect 23032 7040 23096 7044
rect 23112 7100 23176 7104
rect 23112 7044 23116 7100
rect 23116 7044 23172 7100
rect 23172 7044 23176 7100
rect 23112 7040 23176 7044
rect 23192 7100 23256 7104
rect 23192 7044 23196 7100
rect 23196 7044 23252 7100
rect 23252 7044 23256 7100
rect 23192 7040 23256 7044
rect 22324 6836 22388 6900
rect 7952 6556 8016 6560
rect 7952 6500 7956 6556
rect 7956 6500 8012 6556
rect 8012 6500 8016 6556
rect 7952 6496 8016 6500
rect 8032 6556 8096 6560
rect 8032 6500 8036 6556
rect 8036 6500 8092 6556
rect 8092 6500 8096 6556
rect 8032 6496 8096 6500
rect 8112 6556 8176 6560
rect 8112 6500 8116 6556
rect 8116 6500 8172 6556
rect 8172 6500 8176 6556
rect 8112 6496 8176 6500
rect 8192 6556 8256 6560
rect 8192 6500 8196 6556
rect 8196 6500 8252 6556
rect 8252 6500 8256 6556
rect 8192 6496 8256 6500
rect 17952 6556 18016 6560
rect 17952 6500 17956 6556
rect 17956 6500 18012 6556
rect 18012 6500 18016 6556
rect 17952 6496 18016 6500
rect 18032 6556 18096 6560
rect 18032 6500 18036 6556
rect 18036 6500 18092 6556
rect 18092 6500 18096 6556
rect 18032 6496 18096 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 2952 6012 3016 6016
rect 2952 5956 2956 6012
rect 2956 5956 3012 6012
rect 3012 5956 3016 6012
rect 2952 5952 3016 5956
rect 3032 6012 3096 6016
rect 3032 5956 3036 6012
rect 3036 5956 3092 6012
rect 3092 5956 3096 6012
rect 3032 5952 3096 5956
rect 3112 6012 3176 6016
rect 3112 5956 3116 6012
rect 3116 5956 3172 6012
rect 3172 5956 3176 6012
rect 3112 5952 3176 5956
rect 3192 6012 3256 6016
rect 3192 5956 3196 6012
rect 3196 5956 3252 6012
rect 3252 5956 3256 6012
rect 3192 5952 3256 5956
rect 12952 6012 13016 6016
rect 12952 5956 12956 6012
rect 12956 5956 13012 6012
rect 13012 5956 13016 6012
rect 12952 5952 13016 5956
rect 13032 6012 13096 6016
rect 13032 5956 13036 6012
rect 13036 5956 13092 6012
rect 13092 5956 13096 6012
rect 13032 5952 13096 5956
rect 13112 6012 13176 6016
rect 13112 5956 13116 6012
rect 13116 5956 13172 6012
rect 13172 5956 13176 6012
rect 13112 5952 13176 5956
rect 13192 6012 13256 6016
rect 13192 5956 13196 6012
rect 13196 5956 13252 6012
rect 13252 5956 13256 6012
rect 13192 5952 13256 5956
rect 22952 6012 23016 6016
rect 22952 5956 22956 6012
rect 22956 5956 23012 6012
rect 23012 5956 23016 6012
rect 22952 5952 23016 5956
rect 23032 6012 23096 6016
rect 23032 5956 23036 6012
rect 23036 5956 23092 6012
rect 23092 5956 23096 6012
rect 23032 5952 23096 5956
rect 23112 6012 23176 6016
rect 23112 5956 23116 6012
rect 23116 5956 23172 6012
rect 23172 5956 23176 6012
rect 23112 5952 23176 5956
rect 23192 6012 23256 6016
rect 23192 5956 23196 6012
rect 23196 5956 23252 6012
rect 23252 5956 23256 6012
rect 23192 5952 23256 5956
rect 20484 5612 20548 5676
rect 7952 5468 8016 5472
rect 7952 5412 7956 5468
rect 7956 5412 8012 5468
rect 8012 5412 8016 5468
rect 7952 5408 8016 5412
rect 8032 5468 8096 5472
rect 8032 5412 8036 5468
rect 8036 5412 8092 5468
rect 8092 5412 8096 5468
rect 8032 5408 8096 5412
rect 8112 5468 8176 5472
rect 8112 5412 8116 5468
rect 8116 5412 8172 5468
rect 8172 5412 8176 5468
rect 8112 5408 8176 5412
rect 8192 5468 8256 5472
rect 8192 5412 8196 5468
rect 8196 5412 8252 5468
rect 8252 5412 8256 5468
rect 8192 5408 8256 5412
rect 17952 5468 18016 5472
rect 17952 5412 17956 5468
rect 17956 5412 18012 5468
rect 18012 5412 18016 5468
rect 17952 5408 18016 5412
rect 18032 5468 18096 5472
rect 18032 5412 18036 5468
rect 18036 5412 18092 5468
rect 18092 5412 18096 5468
rect 18032 5408 18096 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 2952 4924 3016 4928
rect 2952 4868 2956 4924
rect 2956 4868 3012 4924
rect 3012 4868 3016 4924
rect 2952 4864 3016 4868
rect 3032 4924 3096 4928
rect 3032 4868 3036 4924
rect 3036 4868 3092 4924
rect 3092 4868 3096 4924
rect 3032 4864 3096 4868
rect 3112 4924 3176 4928
rect 3112 4868 3116 4924
rect 3116 4868 3172 4924
rect 3172 4868 3176 4924
rect 3112 4864 3176 4868
rect 3192 4924 3256 4928
rect 3192 4868 3196 4924
rect 3196 4868 3252 4924
rect 3252 4868 3256 4924
rect 3192 4864 3256 4868
rect 12952 4924 13016 4928
rect 12952 4868 12956 4924
rect 12956 4868 13012 4924
rect 13012 4868 13016 4924
rect 12952 4864 13016 4868
rect 13032 4924 13096 4928
rect 13032 4868 13036 4924
rect 13036 4868 13092 4924
rect 13092 4868 13096 4924
rect 13032 4864 13096 4868
rect 13112 4924 13176 4928
rect 13112 4868 13116 4924
rect 13116 4868 13172 4924
rect 13172 4868 13176 4924
rect 13112 4864 13176 4868
rect 13192 4924 13256 4928
rect 13192 4868 13196 4924
rect 13196 4868 13252 4924
rect 13252 4868 13256 4924
rect 13192 4864 13256 4868
rect 22952 4924 23016 4928
rect 22952 4868 22956 4924
rect 22956 4868 23012 4924
rect 23012 4868 23016 4924
rect 22952 4864 23016 4868
rect 23032 4924 23096 4928
rect 23032 4868 23036 4924
rect 23036 4868 23092 4924
rect 23092 4868 23096 4924
rect 23032 4864 23096 4868
rect 23112 4924 23176 4928
rect 23112 4868 23116 4924
rect 23116 4868 23172 4924
rect 23172 4868 23176 4924
rect 23112 4864 23176 4868
rect 23192 4924 23256 4928
rect 23192 4868 23196 4924
rect 23196 4868 23252 4924
rect 23252 4868 23256 4924
rect 23192 4864 23256 4868
rect 7952 4380 8016 4384
rect 7952 4324 7956 4380
rect 7956 4324 8012 4380
rect 8012 4324 8016 4380
rect 7952 4320 8016 4324
rect 8032 4380 8096 4384
rect 8032 4324 8036 4380
rect 8036 4324 8092 4380
rect 8092 4324 8096 4380
rect 8032 4320 8096 4324
rect 8112 4380 8176 4384
rect 8112 4324 8116 4380
rect 8116 4324 8172 4380
rect 8172 4324 8176 4380
rect 8112 4320 8176 4324
rect 8192 4380 8256 4384
rect 8192 4324 8196 4380
rect 8196 4324 8252 4380
rect 8252 4324 8256 4380
rect 8192 4320 8256 4324
rect 17952 4380 18016 4384
rect 17952 4324 17956 4380
rect 17956 4324 18012 4380
rect 18012 4324 18016 4380
rect 17952 4320 18016 4324
rect 18032 4380 18096 4384
rect 18032 4324 18036 4380
rect 18036 4324 18092 4380
rect 18092 4324 18096 4380
rect 18032 4320 18096 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 2952 3836 3016 3840
rect 2952 3780 2956 3836
rect 2956 3780 3012 3836
rect 3012 3780 3016 3836
rect 2952 3776 3016 3780
rect 3032 3836 3096 3840
rect 3032 3780 3036 3836
rect 3036 3780 3092 3836
rect 3092 3780 3096 3836
rect 3032 3776 3096 3780
rect 3112 3836 3176 3840
rect 3112 3780 3116 3836
rect 3116 3780 3172 3836
rect 3172 3780 3176 3836
rect 3112 3776 3176 3780
rect 3192 3836 3256 3840
rect 3192 3780 3196 3836
rect 3196 3780 3252 3836
rect 3252 3780 3256 3836
rect 3192 3776 3256 3780
rect 12952 3836 13016 3840
rect 12952 3780 12956 3836
rect 12956 3780 13012 3836
rect 13012 3780 13016 3836
rect 12952 3776 13016 3780
rect 13032 3836 13096 3840
rect 13032 3780 13036 3836
rect 13036 3780 13092 3836
rect 13092 3780 13096 3836
rect 13032 3776 13096 3780
rect 13112 3836 13176 3840
rect 13112 3780 13116 3836
rect 13116 3780 13172 3836
rect 13172 3780 13176 3836
rect 13112 3776 13176 3780
rect 13192 3836 13256 3840
rect 13192 3780 13196 3836
rect 13196 3780 13252 3836
rect 13252 3780 13256 3836
rect 13192 3776 13256 3780
rect 22952 3836 23016 3840
rect 22952 3780 22956 3836
rect 22956 3780 23012 3836
rect 23012 3780 23016 3836
rect 22952 3776 23016 3780
rect 23032 3836 23096 3840
rect 23032 3780 23036 3836
rect 23036 3780 23092 3836
rect 23092 3780 23096 3836
rect 23032 3776 23096 3780
rect 23112 3836 23176 3840
rect 23112 3780 23116 3836
rect 23116 3780 23172 3836
rect 23172 3780 23176 3836
rect 23112 3776 23176 3780
rect 23192 3836 23256 3840
rect 23192 3780 23196 3836
rect 23196 3780 23252 3836
rect 23252 3780 23256 3836
rect 23192 3776 23256 3780
rect 7952 3292 8016 3296
rect 7952 3236 7956 3292
rect 7956 3236 8012 3292
rect 8012 3236 8016 3292
rect 7952 3232 8016 3236
rect 8032 3292 8096 3296
rect 8032 3236 8036 3292
rect 8036 3236 8092 3292
rect 8092 3236 8096 3292
rect 8032 3232 8096 3236
rect 8112 3292 8176 3296
rect 8112 3236 8116 3292
rect 8116 3236 8172 3292
rect 8172 3236 8176 3292
rect 8112 3232 8176 3236
rect 8192 3292 8256 3296
rect 8192 3236 8196 3292
rect 8196 3236 8252 3292
rect 8252 3236 8256 3292
rect 8192 3232 8256 3236
rect 17952 3292 18016 3296
rect 17952 3236 17956 3292
rect 17956 3236 18012 3292
rect 18012 3236 18016 3292
rect 17952 3232 18016 3236
rect 18032 3292 18096 3296
rect 18032 3236 18036 3292
rect 18036 3236 18092 3292
rect 18092 3236 18096 3292
rect 18032 3232 18096 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 2952 2748 3016 2752
rect 2952 2692 2956 2748
rect 2956 2692 3012 2748
rect 3012 2692 3016 2748
rect 2952 2688 3016 2692
rect 3032 2748 3096 2752
rect 3032 2692 3036 2748
rect 3036 2692 3092 2748
rect 3092 2692 3096 2748
rect 3032 2688 3096 2692
rect 3112 2748 3176 2752
rect 3112 2692 3116 2748
rect 3116 2692 3172 2748
rect 3172 2692 3176 2748
rect 3112 2688 3176 2692
rect 3192 2748 3256 2752
rect 3192 2692 3196 2748
rect 3196 2692 3252 2748
rect 3252 2692 3256 2748
rect 3192 2688 3256 2692
rect 12952 2748 13016 2752
rect 12952 2692 12956 2748
rect 12956 2692 13012 2748
rect 13012 2692 13016 2748
rect 12952 2688 13016 2692
rect 13032 2748 13096 2752
rect 13032 2692 13036 2748
rect 13036 2692 13092 2748
rect 13092 2692 13096 2748
rect 13032 2688 13096 2692
rect 13112 2748 13176 2752
rect 13112 2692 13116 2748
rect 13116 2692 13172 2748
rect 13172 2692 13176 2748
rect 13112 2688 13176 2692
rect 13192 2748 13256 2752
rect 13192 2692 13196 2748
rect 13196 2692 13252 2748
rect 13252 2692 13256 2748
rect 13192 2688 13256 2692
rect 22952 2748 23016 2752
rect 22952 2692 22956 2748
rect 22956 2692 23012 2748
rect 23012 2692 23016 2748
rect 22952 2688 23016 2692
rect 23032 2748 23096 2752
rect 23032 2692 23036 2748
rect 23036 2692 23092 2748
rect 23092 2692 23096 2748
rect 23032 2688 23096 2692
rect 23112 2748 23176 2752
rect 23112 2692 23116 2748
rect 23116 2692 23172 2748
rect 23172 2692 23176 2748
rect 23112 2688 23176 2692
rect 23192 2748 23256 2752
rect 23192 2692 23196 2748
rect 23196 2692 23252 2748
rect 23252 2692 23256 2748
rect 23192 2688 23256 2692
rect 7952 2204 8016 2208
rect 7952 2148 7956 2204
rect 7956 2148 8012 2204
rect 8012 2148 8016 2204
rect 7952 2144 8016 2148
rect 8032 2204 8096 2208
rect 8032 2148 8036 2204
rect 8036 2148 8092 2204
rect 8092 2148 8096 2204
rect 8032 2144 8096 2148
rect 8112 2204 8176 2208
rect 8112 2148 8116 2204
rect 8116 2148 8172 2204
rect 8172 2148 8176 2204
rect 8112 2144 8176 2148
rect 8192 2204 8256 2208
rect 8192 2148 8196 2204
rect 8196 2148 8252 2204
rect 8252 2148 8256 2204
rect 8192 2144 8256 2148
rect 17952 2204 18016 2208
rect 17952 2148 17956 2204
rect 17956 2148 18012 2204
rect 18012 2148 18016 2204
rect 17952 2144 18016 2148
rect 18032 2204 18096 2208
rect 18032 2148 18036 2204
rect 18036 2148 18092 2204
rect 18092 2148 18096 2204
rect 18032 2144 18096 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
<< metal4 >>
rect 6499 26076 6565 26077
rect 6499 26012 6500 26076
rect 6564 26012 6565 26076
rect 6499 26011 6565 26012
rect 2944 24512 3264 24528
rect 2944 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3264 24512
rect 2944 23424 3264 24448
rect 2944 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3264 23424
rect 2944 22336 3264 23360
rect 2944 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3264 22336
rect 2944 21248 3264 22272
rect 2944 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3264 21248
rect 2944 20160 3264 21184
rect 2944 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3264 20160
rect 2944 19072 3264 20096
rect 6502 19277 6562 26011
rect 9627 24852 9693 24853
rect 9627 24788 9628 24852
rect 9692 24788 9693 24852
rect 9627 24787 9693 24788
rect 8891 24716 8957 24717
rect 8891 24652 8892 24716
rect 8956 24652 8957 24716
rect 8891 24651 8957 24652
rect 7944 23968 8264 24528
rect 7944 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8264 23968
rect 7944 22880 8264 23904
rect 7944 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8264 22880
rect 7944 21792 8264 22816
rect 7944 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8264 21792
rect 7944 20704 8264 21728
rect 7944 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8264 20704
rect 7944 19616 8264 20640
rect 7944 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8264 19616
rect 6499 19276 6565 19277
rect 6499 19212 6500 19276
rect 6564 19212 6565 19276
rect 6499 19211 6565 19212
rect 2944 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3264 19072
rect 2944 17984 3264 19008
rect 2944 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3264 17984
rect 2944 16896 3264 17920
rect 2944 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3264 16896
rect 2944 15808 3264 16832
rect 2944 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3264 15808
rect 2944 14720 3264 15744
rect 2944 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3264 14720
rect 2944 13632 3264 14656
rect 2944 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3264 13632
rect 2944 12544 3264 13568
rect 2944 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3264 12544
rect 2944 11456 3264 12480
rect 2944 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3264 11456
rect 2944 10368 3264 11392
rect 2944 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3264 10368
rect 2944 9280 3264 10304
rect 2944 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3264 9280
rect 2944 8192 3264 9216
rect 2944 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3264 8192
rect 2944 7104 3264 8128
rect 2944 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3264 7104
rect 2944 6016 3264 7040
rect 2944 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3264 6016
rect 2944 4928 3264 5952
rect 2944 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3264 4928
rect 2944 3840 3264 4864
rect 2944 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3264 3840
rect 2944 2752 3264 3776
rect 2944 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3264 2752
rect 2944 2128 3264 2688
rect 7944 18528 8264 19552
rect 7944 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8264 18528
rect 7944 17440 8264 18464
rect 7944 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8264 17440
rect 7944 16352 8264 17376
rect 8894 16557 8954 24651
rect 9443 23356 9509 23357
rect 9443 23292 9444 23356
rect 9508 23292 9509 23356
rect 9443 23291 9509 23292
rect 8891 16556 8957 16557
rect 8891 16492 8892 16556
rect 8956 16492 8957 16556
rect 8891 16491 8957 16492
rect 7944 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8264 16352
rect 7944 15264 8264 16288
rect 9446 15605 9506 23291
rect 9630 18053 9690 24787
rect 12944 24512 13264 24528
rect 12944 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13264 24512
rect 12019 24308 12085 24309
rect 12019 24244 12020 24308
rect 12084 24244 12085 24308
rect 12019 24243 12085 24244
rect 10363 24036 10429 24037
rect 10363 23972 10364 24036
rect 10428 23972 10429 24036
rect 10363 23971 10429 23972
rect 9627 18052 9693 18053
rect 9627 17988 9628 18052
rect 9692 17988 9693 18052
rect 9627 17987 9693 17988
rect 9443 15604 9509 15605
rect 9443 15540 9444 15604
rect 9508 15540 9509 15604
rect 9443 15539 9509 15540
rect 7944 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8264 15264
rect 7944 14176 8264 15200
rect 10366 15061 10426 23971
rect 11099 22676 11165 22677
rect 11099 22612 11100 22676
rect 11164 22612 11165 22676
rect 11099 22611 11165 22612
rect 11102 17781 11162 22611
rect 11099 17780 11165 17781
rect 11099 17716 11100 17780
rect 11164 17716 11165 17780
rect 11099 17715 11165 17716
rect 10363 15060 10429 15061
rect 10363 14996 10364 15060
rect 10428 14996 10429 15060
rect 10363 14995 10429 14996
rect 7944 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8264 14176
rect 7944 13088 8264 14112
rect 12022 13973 12082 24243
rect 12944 23424 13264 24448
rect 14963 24172 15029 24173
rect 14963 24108 14964 24172
rect 15028 24108 15029 24172
rect 14963 24107 15029 24108
rect 12944 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13264 23424
rect 12387 22812 12453 22813
rect 12387 22748 12388 22812
rect 12452 22810 12453 22812
rect 12571 22812 12637 22813
rect 12571 22810 12572 22812
rect 12452 22750 12572 22810
rect 12452 22748 12453 22750
rect 12387 22747 12453 22748
rect 12571 22748 12572 22750
rect 12636 22748 12637 22812
rect 12571 22747 12637 22748
rect 12944 22336 13264 23360
rect 12944 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13264 22336
rect 12571 21724 12637 21725
rect 12571 21660 12572 21724
rect 12636 21660 12637 21724
rect 12571 21659 12637 21660
rect 12574 21450 12634 21659
rect 12390 21390 12634 21450
rect 12390 21317 12450 21390
rect 12387 21316 12453 21317
rect 12387 21252 12388 21316
rect 12452 21252 12453 21316
rect 12387 21251 12453 21252
rect 12944 21248 13264 22272
rect 13491 21860 13557 21861
rect 13491 21796 13492 21860
rect 13556 21796 13557 21860
rect 13491 21795 13557 21796
rect 12944 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13264 21248
rect 12944 20160 13264 21184
rect 12944 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13264 20160
rect 12944 19072 13264 20096
rect 12944 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13264 19072
rect 12944 17984 13264 19008
rect 12944 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13264 17984
rect 12944 16896 13264 17920
rect 12944 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13264 16896
rect 12944 15808 13264 16832
rect 12944 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13264 15808
rect 12944 14720 13264 15744
rect 12944 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13264 14720
rect 12019 13972 12085 13973
rect 12019 13908 12020 13972
rect 12084 13908 12085 13972
rect 12019 13907 12085 13908
rect 7944 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8264 13088
rect 7944 12000 8264 13024
rect 7944 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8264 12000
rect 7944 10912 8264 11936
rect 7944 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8264 10912
rect 7944 9824 8264 10848
rect 7944 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8264 9824
rect 7944 8736 8264 9760
rect 7944 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8264 8736
rect 7944 7648 8264 8672
rect 7944 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8264 7648
rect 7944 6560 8264 7584
rect 7944 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8264 6560
rect 7944 5472 8264 6496
rect 7944 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8264 5472
rect 7944 4384 8264 5408
rect 7944 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8264 4384
rect 7944 3296 8264 4320
rect 7944 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8264 3296
rect 7944 2208 8264 3232
rect 7944 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8264 2208
rect 7944 2128 8264 2144
rect 12944 13632 13264 14656
rect 12944 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13264 13632
rect 12944 12544 13264 13568
rect 12944 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13264 12544
rect 12944 11456 13264 12480
rect 12944 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13264 11456
rect 12944 10368 13264 11392
rect 12944 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13264 10368
rect 12944 9280 13264 10304
rect 12944 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13264 9280
rect 12944 8192 13264 9216
rect 12944 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13264 8192
rect 12944 7104 13264 8128
rect 13494 7853 13554 21795
rect 13675 20228 13741 20229
rect 13675 20164 13676 20228
rect 13740 20164 13741 20228
rect 13675 20163 13741 20164
rect 13678 13565 13738 20163
rect 14966 15197 15026 24107
rect 17944 23968 18264 24528
rect 17944 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18264 23968
rect 16251 23900 16317 23901
rect 16251 23836 16252 23900
rect 16316 23836 16317 23900
rect 16251 23835 16317 23836
rect 15147 23628 15213 23629
rect 15147 23564 15148 23628
rect 15212 23564 15213 23628
rect 15147 23563 15213 23564
rect 15150 20909 15210 23563
rect 15147 20908 15213 20909
rect 15147 20844 15148 20908
rect 15212 20844 15213 20908
rect 15147 20843 15213 20844
rect 15883 20772 15949 20773
rect 15883 20708 15884 20772
rect 15948 20708 15949 20772
rect 15883 20707 15949 20708
rect 14963 15196 15029 15197
rect 14963 15132 14964 15196
rect 15028 15132 15029 15196
rect 14963 15131 15029 15132
rect 13675 13564 13741 13565
rect 13675 13500 13676 13564
rect 13740 13500 13741 13564
rect 13675 13499 13741 13500
rect 15886 9485 15946 20707
rect 16067 19412 16133 19413
rect 16067 19348 16068 19412
rect 16132 19348 16133 19412
rect 16067 19347 16133 19348
rect 16070 10301 16130 19347
rect 16254 11389 16314 23835
rect 17355 23220 17421 23221
rect 17355 23156 17356 23220
rect 17420 23156 17421 23220
rect 17355 23155 17421 23156
rect 16435 19412 16501 19413
rect 16435 19348 16436 19412
rect 16500 19348 16501 19412
rect 16435 19347 16501 19348
rect 16251 11388 16317 11389
rect 16251 11324 16252 11388
rect 16316 11324 16317 11388
rect 16251 11323 16317 11324
rect 16067 10300 16133 10301
rect 16067 10236 16068 10300
rect 16132 10236 16133 10300
rect 16067 10235 16133 10236
rect 15883 9484 15949 9485
rect 15883 9420 15884 9484
rect 15948 9420 15949 9484
rect 15883 9419 15949 9420
rect 16438 8397 16498 19347
rect 16619 16828 16685 16829
rect 16619 16764 16620 16828
rect 16684 16764 16685 16828
rect 16619 16763 16685 16764
rect 16622 15061 16682 16763
rect 16619 15060 16685 15061
rect 16619 14996 16620 15060
rect 16684 14996 16685 15060
rect 16619 14995 16685 14996
rect 17358 13701 17418 23155
rect 17723 23084 17789 23085
rect 17723 23020 17724 23084
rect 17788 23020 17789 23084
rect 17723 23019 17789 23020
rect 17539 18052 17605 18053
rect 17539 17988 17540 18052
rect 17604 17988 17605 18052
rect 17539 17987 17605 17988
rect 17542 13973 17602 17987
rect 17726 16421 17786 23019
rect 17944 22880 18264 23904
rect 22944 24512 23264 24528
rect 22944 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23264 24512
rect 20115 23492 20181 23493
rect 20115 23428 20116 23492
rect 20180 23428 20181 23492
rect 20115 23427 20181 23428
rect 17944 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18264 22880
rect 17944 21792 18264 22816
rect 17944 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18264 21792
rect 17944 20704 18264 21728
rect 19563 20772 19629 20773
rect 19563 20708 19564 20772
rect 19628 20708 19629 20772
rect 19563 20707 19629 20708
rect 17944 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18264 20704
rect 17944 19616 18264 20640
rect 18459 19820 18525 19821
rect 18459 19756 18460 19820
rect 18524 19756 18525 19820
rect 18459 19755 18525 19756
rect 17944 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18264 19616
rect 17944 18528 18264 19552
rect 17944 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18264 18528
rect 17944 17440 18264 18464
rect 17944 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18264 17440
rect 17723 16420 17789 16421
rect 17723 16356 17724 16420
rect 17788 16356 17789 16420
rect 17723 16355 17789 16356
rect 17944 16352 18264 17376
rect 17944 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18264 16352
rect 17944 15264 18264 16288
rect 17944 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18264 15264
rect 17944 14176 18264 15200
rect 17944 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18264 14176
rect 17539 13972 17605 13973
rect 17539 13908 17540 13972
rect 17604 13908 17605 13972
rect 17539 13907 17605 13908
rect 17355 13700 17421 13701
rect 17355 13636 17356 13700
rect 17420 13636 17421 13700
rect 17355 13635 17421 13636
rect 17723 13564 17789 13565
rect 17723 13500 17724 13564
rect 17788 13500 17789 13564
rect 17723 13499 17789 13500
rect 17726 11661 17786 13499
rect 17944 13088 18264 14112
rect 17944 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18264 13088
rect 17944 12000 18264 13024
rect 17944 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18264 12000
rect 17723 11660 17789 11661
rect 17723 11596 17724 11660
rect 17788 11596 17789 11660
rect 17723 11595 17789 11596
rect 17944 10912 18264 11936
rect 18462 11117 18522 19755
rect 19379 19412 19445 19413
rect 19379 19348 19380 19412
rect 19444 19348 19445 19412
rect 19379 19347 19445 19348
rect 19195 17372 19261 17373
rect 19195 17308 19196 17372
rect 19260 17308 19261 17372
rect 19195 17307 19261 17308
rect 18459 11116 18525 11117
rect 18459 11052 18460 11116
rect 18524 11052 18525 11116
rect 18459 11051 18525 11052
rect 17944 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18264 10912
rect 17944 9824 18264 10848
rect 17944 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18264 9824
rect 17944 8736 18264 9760
rect 17944 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18264 8736
rect 16435 8396 16501 8397
rect 16435 8332 16436 8396
rect 16500 8332 16501 8396
rect 16435 8331 16501 8332
rect 13491 7852 13557 7853
rect 13491 7788 13492 7852
rect 13556 7788 13557 7852
rect 13491 7787 13557 7788
rect 12944 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13264 7104
rect 12944 6016 13264 7040
rect 12944 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13264 6016
rect 12944 4928 13264 5952
rect 12944 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13264 4928
rect 12944 3840 13264 4864
rect 12944 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13264 3840
rect 12944 2752 13264 3776
rect 12944 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13264 2752
rect 12944 2128 13264 2688
rect 17944 7648 18264 8672
rect 19198 7989 19258 17307
rect 19382 15469 19442 19347
rect 19566 16829 19626 20707
rect 19747 20364 19813 20365
rect 19747 20300 19748 20364
rect 19812 20300 19813 20364
rect 19747 20299 19813 20300
rect 19563 16828 19629 16829
rect 19563 16764 19564 16828
rect 19628 16764 19629 16828
rect 19563 16763 19629 16764
rect 19750 15877 19810 20299
rect 19747 15876 19813 15877
rect 19747 15812 19748 15876
rect 19812 15812 19813 15876
rect 19747 15811 19813 15812
rect 19379 15468 19445 15469
rect 19379 15404 19380 15468
rect 19444 15404 19445 15468
rect 19379 15403 19445 15404
rect 20118 11117 20178 23427
rect 22944 23424 23264 24448
rect 22944 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23264 23424
rect 22944 22336 23264 23360
rect 24531 22540 24597 22541
rect 24531 22476 24532 22540
rect 24596 22476 24597 22540
rect 24531 22475 24597 22476
rect 22944 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23264 22336
rect 21035 22132 21101 22133
rect 21035 22068 21036 22132
rect 21100 22068 21101 22132
rect 21035 22067 21101 22068
rect 20851 20772 20917 20773
rect 20851 20708 20852 20772
rect 20916 20708 20917 20772
rect 20851 20707 20917 20708
rect 20667 18596 20733 18597
rect 20667 18532 20668 18596
rect 20732 18532 20733 18596
rect 20667 18531 20733 18532
rect 20670 15741 20730 18531
rect 20667 15740 20733 15741
rect 20667 15676 20668 15740
rect 20732 15676 20733 15740
rect 20667 15675 20733 15676
rect 20483 13836 20549 13837
rect 20483 13772 20484 13836
rect 20548 13772 20549 13836
rect 20483 13771 20549 13772
rect 20115 11116 20181 11117
rect 20115 11052 20116 11116
rect 20180 11052 20181 11116
rect 20115 11051 20181 11052
rect 19195 7988 19261 7989
rect 19195 7924 19196 7988
rect 19260 7924 19261 7988
rect 19195 7923 19261 7924
rect 17944 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18264 7648
rect 17944 6560 18264 7584
rect 17944 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18264 6560
rect 17944 5472 18264 6496
rect 20486 5677 20546 13771
rect 20854 12477 20914 20707
rect 21038 20229 21098 22067
rect 21403 21588 21469 21589
rect 21403 21524 21404 21588
rect 21468 21524 21469 21588
rect 21403 21523 21469 21524
rect 21219 20772 21285 20773
rect 21219 20708 21220 20772
rect 21284 20708 21285 20772
rect 21219 20707 21285 20708
rect 21035 20228 21101 20229
rect 21035 20164 21036 20228
rect 21100 20164 21101 20228
rect 21035 20163 21101 20164
rect 21035 20092 21101 20093
rect 21035 20028 21036 20092
rect 21100 20028 21101 20092
rect 21035 20027 21101 20028
rect 21038 13293 21098 20027
rect 21035 13292 21101 13293
rect 21035 13228 21036 13292
rect 21100 13228 21101 13292
rect 21035 13227 21101 13228
rect 20851 12476 20917 12477
rect 20851 12412 20852 12476
rect 20916 12412 20917 12476
rect 20851 12411 20917 12412
rect 21222 9757 21282 20707
rect 21406 13973 21466 21523
rect 22944 21248 23264 22272
rect 22944 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23264 21248
rect 22691 21044 22757 21045
rect 22691 20980 22692 21044
rect 22756 20980 22757 21044
rect 22691 20979 22757 20980
rect 22694 15333 22754 20979
rect 22944 20160 23264 21184
rect 22944 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23264 20160
rect 22944 19072 23264 20096
rect 22944 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23264 19072
rect 22944 17984 23264 19008
rect 23427 18052 23493 18053
rect 23427 17988 23428 18052
rect 23492 17988 23493 18052
rect 23427 17987 23493 17988
rect 22944 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23264 17984
rect 22944 16896 23264 17920
rect 22944 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23264 16896
rect 22944 15808 23264 16832
rect 22944 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23264 15808
rect 22691 15332 22757 15333
rect 22691 15268 22692 15332
rect 22756 15268 22757 15332
rect 22691 15267 22757 15268
rect 22323 14924 22389 14925
rect 22323 14860 22324 14924
rect 22388 14860 22389 14924
rect 22323 14859 22389 14860
rect 21955 14516 22021 14517
rect 21955 14452 21956 14516
rect 22020 14452 22021 14516
rect 21955 14451 22021 14452
rect 21403 13972 21469 13973
rect 21403 13908 21404 13972
rect 21468 13908 21469 13972
rect 21403 13907 21469 13908
rect 21219 9756 21285 9757
rect 21219 9692 21220 9756
rect 21284 9692 21285 9756
rect 21219 9691 21285 9692
rect 21958 8397 22018 14451
rect 21955 8396 22021 8397
rect 21955 8332 21956 8396
rect 22020 8332 22021 8396
rect 21955 8331 22021 8332
rect 22326 6901 22386 14859
rect 22944 14720 23264 15744
rect 22944 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23264 14720
rect 22944 13632 23264 14656
rect 22944 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23264 13632
rect 22944 12544 23264 13568
rect 22944 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23264 12544
rect 22944 11456 23264 12480
rect 22944 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23264 11456
rect 22944 10368 23264 11392
rect 23430 10709 23490 17987
rect 24534 15605 24594 22475
rect 24531 15604 24597 15605
rect 24531 15540 24532 15604
rect 24596 15540 24597 15604
rect 24531 15539 24597 15540
rect 23427 10708 23493 10709
rect 23427 10644 23428 10708
rect 23492 10644 23493 10708
rect 23427 10643 23493 10644
rect 22944 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23264 10368
rect 22944 9280 23264 10304
rect 22944 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23264 9280
rect 22944 8192 23264 9216
rect 22944 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23264 8192
rect 22944 7104 23264 8128
rect 22944 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23264 7104
rect 22323 6900 22389 6901
rect 22323 6836 22324 6900
rect 22388 6836 22389 6900
rect 22323 6835 22389 6836
rect 22944 6016 23264 7040
rect 22944 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23264 6016
rect 20483 5676 20549 5677
rect 20483 5612 20484 5676
rect 20548 5612 20549 5676
rect 20483 5611 20549 5612
rect 17944 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18264 5472
rect 17944 4384 18264 5408
rect 17944 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18264 4384
rect 17944 3296 18264 4320
rect 17944 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18264 3296
rect 17944 2208 18264 3232
rect 17944 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18264 2208
rect 17944 2128 18264 2144
rect 22944 4928 23264 5952
rect 22944 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23264 4928
rect 22944 3840 23264 4864
rect 22944 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23264 3840
rect 22944 2752 23264 3776
rect 22944 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23264 2752
rect 22944 2128 23264 2688
use sky130_fd_sc_hd__clkbuf_2  _072_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18584 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _073_
timestamp 1676037725
transform 1 0 19872 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _074_
timestamp 1676037725
transform 1 0 21988 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _075_
timestamp 1676037725
transform 1 0 25024 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _076_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24564 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _077_
timestamp 1676037725
transform 1 0 24656 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _078_
timestamp 1676037725
transform 1 0 24656 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _079_
timestamp 1676037725
transform 1 0 24564 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _080_
timestamp 1676037725
transform 1 0 24564 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _081_
timestamp 1676037725
transform 1 0 22632 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _082_
timestamp 1676037725
transform 1 0 21988 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _083_
timestamp 1676037725
transform 1 0 21896 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _084_
timestamp 1676037725
transform 1 0 24656 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _085_
timestamp 1676037725
transform 1 0 24564 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _086_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19412 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _087_
timestamp 1676037725
transform 1 0 20608 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _088_
timestamp 1676037725
transform 1 0 24748 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _089_
timestamp 1676037725
transform 1 0 24748 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _090_
timestamp 1676037725
transform 1 0 23736 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _091_
timestamp 1676037725
transform 1 0 24564 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _092_
timestamp 1676037725
transform 1 0 20700 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _093_
timestamp 1676037725
transform 1 0 21252 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _094_
timestamp 1676037725
transform 1 0 18032 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _095_
timestamp 1676037725
transform 1 0 19964 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _096_
timestamp 1676037725
transform 1 0 15180 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _097_
timestamp 1676037725
transform 1 0 19964 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _098_
timestamp 1676037725
transform 1 0 18032 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _099_
timestamp 1676037725
transform 1 0 19412 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _100_
timestamp 1676037725
transform 1 0 14260 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _101_
timestamp 1676037725
transform 1 0 21344 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _102_
timestamp 1676037725
transform 1 0 14260 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _103_
timestamp 1676037725
transform 1 0 16100 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _104_
timestamp 1676037725
transform 1 0 14260 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _105_
timestamp 1676037725
transform 1 0 15732 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _106_
timestamp 1676037725
transform 1 0 5152 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _107_
timestamp 1676037725
transform 1 0 6532 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _108_
timestamp 1676037725
transform 1 0 5796 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _109_
timestamp 1676037725
transform 1 0 4508 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _110_
timestamp 1676037725
transform 1 0 13432 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _111_
timestamp 1676037725
transform 1 0 15824 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _112_
timestamp 1676037725
transform 1 0 19044 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _113_
timestamp 1676037725
transform 1 0 13432 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _114_
timestamp 1676037725
transform 1 0 6440 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _115_
timestamp 1676037725
transform 1 0 3864 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _116_
timestamp 1676037725
transform 1 0 7728 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _117_
timestamp 1676037725
transform 1 0 7820 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _118_
timestamp 1676037725
transform 1 0 12880 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _119_
timestamp 1676037725
transform 1 0 16928 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _120_
timestamp 1676037725
transform 1 0 19412 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _121_
timestamp 1676037725
transform 1 0 18400 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _122_
timestamp 1676037725
transform 1 0 3220 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _123_
timestamp 1676037725
transform 1 0 5796 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _124_
timestamp 1676037725
transform 1 0 2208 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _125_
timestamp 1676037725
transform 1 0 4508 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _126_
timestamp 1676037725
transform 1 0 7084 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _127_
timestamp 1676037725
transform 1 0 5152 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _128_
timestamp 1676037725
transform 1 0 7084 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _129_
timestamp 1676037725
transform 1 0 9200 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _130_
timestamp 1676037725
transform 1 0 5152 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _131_
timestamp 1676037725
transform 1 0 4508 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17204 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1676037725
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1676037725
transform 1 0 13340 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1676037725
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1676037725
transform 1 0 15272 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1676037725
transform 1 0 17940 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1676037725
transform 1 0 19872 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1676037725
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1676037725
transform 1 0 24840 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1676037725
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1676037725
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__072__A
timestamp 1676037725
transform 1 0 20424 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__073__A
timestamp 1676037725
transform 1 0 21436 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__A
timestamp 1676037725
transform 1 0 23920 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__A
timestamp 1676037725
transform 1 0 25116 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__081__A
timestamp 1676037725
transform 1 0 24012 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__088__A
timestamp 1676037725
transform 1 0 25300 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__A
timestamp 1676037725
transform 1 0 25300 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__A
timestamp 1676037725
transform 1 0 25300 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__A
timestamp 1676037725
transform 1 0 25116 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__100__A
timestamp 1676037725
transform 1 0 13432 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__110__A
timestamp 1676037725
transform 1 0 13248 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__A
timestamp 1676037725
transform 1 0 12788 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__121__A
timestamp 1676037725
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1676037725
transform 1 0 18952 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0__f_prog_clk_A
timestamp 1676037725
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1__f_prog_clk_A
timestamp 1676037725
transform 1 0 15364 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2__f_prog_clk_A
timestamp 1676037725
transform 1 0 11684 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3__f_prog_clk_A
timestamp 1676037725
transform 1 0 16192 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4__f_prog_clk_A
timestamp 1676037725
transform 1 0 21252 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5__f_prog_clk_A
timestamp 1676037725
transform 1 0 21344 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6__f_prog_clk_A
timestamp 1676037725
transform 1 0 21436 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7__f_prog_clk_A
timestamp 1676037725
transform 1 0 24012 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold1_A
timestamp 1676037725
transform 1 0 15180 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold3_A
timestamp 1676037725
transform 1 0 25300 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold4_A
timestamp 1676037725
transform 1 0 6440 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1676037725
transform 1 0 21160 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1676037725
transform 1 0 21528 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1676037725
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1676037725
transform 1 0 13708 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1676037725
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1676037725
transform 1 0 7912 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1676037725
transform 1 0 3772 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1676037725
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1676037725
transform 1 0 9752 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1676037725
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1676037725
transform 1 0 7176 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1676037725
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1676037725
transform 1 0 20884 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1676037725
transform 1 0 21620 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1676037725
transform 1 0 16836 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1676037725
transform 1 0 20792 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1676037725
transform 1 0 15548 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1676037725
transform 1 0 15732 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1676037725
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1676037725
transform 1 0 11040 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1676037725
transform 1 0 10304 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1676037725
transform 1 0 9384 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1676037725
transform 1 0 21344 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1676037725
transform 1 0 22264 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1676037725
transform 1 0 19412 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1676037725
transform 1 0 17020 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1676037725
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1676037725
transform 1 0 25208 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1676037725
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1676037725
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1676037725
transform 1 0 2668 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1676037725
transform 1 0 6256 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1676037725
transform 1 0 16652 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1676037725
transform 1 0 18860 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1676037725
transform 1 0 4232 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1676037725
transform 1 0 16560 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1676037725
transform 1 0 14444 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1676037725
transform 1 0 6532 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1676037725
transform 1 0 6348 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1676037725
transform 1 0 6624 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1676037725
transform 1 0 6716 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1676037725
transform 1 0 2852 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1676037725
transform 1 0 3956 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1676037725
transform 1 0 3956 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1676037725
transform 1 0 6440 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1676037725
transform 1 0 9108 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1676037725
transform 1 0 4784 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1676037725
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1676037725
transform 1 0 1564 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1676037725
transform 1 0 9568 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1676037725
transform 1 0 21160 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1676037725
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1676037725
transform 1 0 8924 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1676037725
transform 1 0 6808 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1676037725
transform 1 0 7176 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1676037725
transform 1 0 11500 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1676037725
transform 1 0 1656 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1676037725
transform 1 0 21252 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1676037725
transform 1 0 7360 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1676037725
transform 1 0 11684 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 1676037725
transform 1 0 6532 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 1676037725
transform 1 0 6532 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 1676037725
transform 1 0 25392 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 1676037725
transform 1 0 25300 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 1676037725
transform 1 0 1656 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input68_A
timestamp 1676037725
transform 1 0 1472 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 1676037725
transform 1 0 2208 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input70_A
timestamp 1676037725
transform 1 0 2116 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output95_A
timestamp 1676037725
transform 1 0 19688 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output103_A
timestamp 1676037725
transform 1 0 2392 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 17480 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21436 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 23828 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 13708 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 11500 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 2392 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 2208 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 6716 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 8924 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 11500 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 24288 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 22908 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 23092 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 25300 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 24196 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 22724 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 22816 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 24196 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 24564 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 25024 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 24012 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 22172 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 21988 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21804 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 20424 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 20240 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21436 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 15732 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 20608 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 21344 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 12052 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1676037725
transform 1 0 14352 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 18860 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 19596 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 24012 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 11684 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 24656 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 20240 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 20056 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 18676 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 16284 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 13432 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 12972 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 11868 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 11040 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 11040 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 11500 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 11040 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 11040 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 12604 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 14904 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 9936 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 12512 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 13616 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 14628 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 16284 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 15732 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 16284 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_0.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 19964 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_2.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 1656 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_2.mux_l2_in_0__A0
timestamp 1676037725
transform 1 0 25208 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_2.sky130_fd_sc_hd__buf_4_0__A
timestamp 1676037725
transform 1 0 4140 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_4.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 21252 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_4.mux_l2_in_0__A0
timestamp 1676037725
transform 1 0 25300 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_6.sky130_fd_sc_hd__buf_4_0__A
timestamp 1676037725
transform 1 0 8096 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_8.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_10.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 25392 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_12.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 21436 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_12.mux_l2_in_0__A0
timestamp 1676037725
transform 1 0 23828 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_14.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 25392 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_16.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 24472 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_18.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 23000 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_34.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 20424 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_48.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 21436 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_50.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 23000 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_0.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 13156 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_0.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 13616 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_0.mux_l1_in_0__S
timestamp 1676037725
transform 1 0 12420 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_0.mux_l1_in_1__S
timestamp 1676037725
transform 1 0 21436 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_2.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 25024 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_2.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_4.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 11684 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_4.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 21896 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_6.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 14996 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_6.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 16192 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_6.sky130_fd_sc_hd__buf_4_0__A
timestamp 1676037725
transform 1 0 4140 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_8.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 21068 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_10.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_12.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_14.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 18860 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_16.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 16008 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_18.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 14812 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_28.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_30.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 20608 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_32.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 19872 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_34.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 17848 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_44.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 15088 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_46.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 18124 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_48.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_50.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 18676 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_50.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 17664 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17112 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_prog_clk
timestamp 1676037725
transform 1 0 9568 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_prog_clk
timestamp 1676037725
transform 1 0 12972 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_prog_clk
timestamp 1676037725
transform 1 0 10396 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_prog_clk
timestamp 1676037725
transform 1 0 12972 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_prog_clk
timestamp 1676037725
transform 1 0 18216 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_prog_clk
timestamp 1676037725
transform 1 0 20792 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_prog_clk
timestamp 1676037725
transform 1 0 18216 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_prog_clk
timestamp 1676037725
transform 1 0 21988 0 -1 18496
box -38 -48 1878 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1676037725
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1676037725
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57
timestamp 1676037725
transform 1 0 6348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6624 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70
timestamp 1676037725
transform 1 0 7544 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1676037725
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1676037725
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1676037725
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1676037725
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1676037725
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1676037725
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1676037725
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1676037725
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1676037725
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1676037725
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1676037725
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1676037725
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1676037725
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_197 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19228 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_201
timestamp 1676037725
transform 1 0 19596 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_204
timestamp 1676037725
transform 1 0 19872 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1676037725
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_225 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21804 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_233
timestamp 1676037725
transform 1 0 22540 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_250
timestamp 1676037725
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1676037725
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_265
timestamp 1676037725
transform 1 0 25484 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1676037725
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1676037725
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1676037725
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1676037725
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1676037725
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_57
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_61
timestamp 1676037725
transform 1 0 6716 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_65
timestamp 1676037725
transform 1 0 7084 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_77
timestamp 1676037725
transform 1 0 8188 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_89
timestamp 1676037725
transform 1 0 9292 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_101
timestamp 1676037725
transform 1 0 10396 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_109
timestamp 1676037725
transform 1 0 11132 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1676037725
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1676037725
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1676037725
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1676037725
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1676037725
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1676037725
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_181
timestamp 1676037725
transform 1 0 17756 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_185
timestamp 1676037725
transform 1 0 18124 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_202
timestamp 1676037725
transform 1 0 19688 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp 1676037725
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_225
timestamp 1676037725
transform 1 0 21804 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_244
timestamp 1676037725
transform 1 0 23552 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_264
timestamp 1676037725
transform 1 0 25392 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1676037725
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1676037725
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1676037725
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1676037725
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1676037725
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1676037725
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1676037725
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1676037725
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1676037725
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1676037725
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1676037725
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1676037725
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1676037725
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1676037725
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1676037725
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1676037725
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1676037725
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1676037725
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1676037725
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1676037725
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_209
timestamp 1676037725
transform 1 0 20332 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_213
timestamp 1676037725
transform 1 0 20700 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_230
timestamp 1676037725
transform 1 0 22264 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_250
timestamp 1676037725
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_253
timestamp 1676037725
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_258
timestamp 1676037725
transform 1 0 24840 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1676037725
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1676037725
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1676037725
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1676037725
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1676037725
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1676037725
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1676037725
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1676037725
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1676037725
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1676037725
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1676037725
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1676037725
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1676037725
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1676037725
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1676037725
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1676037725
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1676037725
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1676037725
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1676037725
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_205
timestamp 1676037725
transform 1 0 19964 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_222
timestamp 1676037725
transform 1 0 21528 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_225
timestamp 1676037725
transform 1 0 21804 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_244
timestamp 1676037725
transform 1 0 23552 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_264
timestamp 1676037725
transform 1 0 25392 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1676037725
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1676037725
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1676037725
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1676037725
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1676037725
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1676037725
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1676037725
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1676037725
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1676037725
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1676037725
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1676037725
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1676037725
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1676037725
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1676037725
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1676037725
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1676037725
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1676037725
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1676037725
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1676037725
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1676037725
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_221
timestamp 1676037725
transform 1 0 21436 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_229
timestamp 1676037725
transform 1 0 22172 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_232
timestamp 1676037725
transform 1 0 22448 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_250
timestamp 1676037725
transform 1 0 24104 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_253
timestamp 1676037725
transform 1 0 24380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_259
timestamp 1676037725
transform 1 0 24932 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_265
timestamp 1676037725
transform 1 0 25484 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1676037725
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1676037725
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1676037725
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1676037725
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1676037725
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1676037725
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1676037725
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1676037725
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1676037725
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1676037725
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1676037725
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1676037725
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1676037725
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1676037725
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1676037725
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1676037725
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1676037725
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1676037725
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1676037725
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1676037725
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1676037725
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1676037725
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_225
timestamp 1676037725
transform 1 0 21804 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_244
timestamp 1676037725
transform 1 0 23552 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_264
timestamp 1676037725
transform 1 0 25392 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1676037725
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1676037725
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1676037725
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1676037725
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1676037725
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1676037725
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1676037725
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1676037725
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1676037725
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1676037725
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1676037725
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1676037725
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1676037725
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1676037725
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1676037725
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1676037725
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1676037725
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1676037725
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1676037725
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_209
timestamp 1676037725
transform 1 0 20332 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_217
timestamp 1676037725
transform 1 0 21068 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_223
timestamp 1676037725
transform 1 0 21620 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_230
timestamp 1676037725
transform 1 0 22264 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_250
timestamp 1676037725
transform 1 0 24104 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_253
timestamp 1676037725
transform 1 0 24380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_6_259
timestamp 1676037725
transform 1 0 24932 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_265
timestamp 1676037725
transform 1 0 25484 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1676037725
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1676037725
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1676037725
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1676037725
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1676037725
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1676037725
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_81
timestamp 1676037725
transform 1 0 8556 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_90
timestamp 1676037725
transform 1 0 9384 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_102
timestamp 1676037725
transform 1 0 10488 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_110
timestamp 1676037725
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1676037725
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1676037725
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1676037725
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1676037725
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1676037725
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1676037725
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1676037725
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1676037725
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1676037725
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1676037725
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_217
timestamp 1676037725
transform 1 0 21068 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_221
timestamp 1676037725
transform 1 0 21436 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_225
timestamp 1676037725
transform 1 0 21804 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_244
timestamp 1676037725
transform 1 0 23552 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_264
timestamp 1676037725
transform 1 0 25392 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1676037725
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1676037725
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1676037725
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1676037725
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1676037725
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1676037725
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1676037725
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1676037725
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1676037725
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1676037725
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1676037725
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1676037725
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1676037725
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1676037725
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1676037725
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1676037725
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1676037725
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1676037725
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1676037725
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_209
timestamp 1676037725
transform 1 0 20332 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_215
timestamp 1676037725
transform 1 0 20884 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_222
timestamp 1676037725
transform 1 0 21528 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_226
timestamp 1676037725
transform 1 0 21896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_230
timestamp 1676037725
transform 1 0 22264 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp 1676037725
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_253
timestamp 1676037725
transform 1 0 24380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_259
timestamp 1676037725
transform 1 0 24932 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_265
timestamp 1676037725
transform 1 0 25484 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1676037725
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1676037725
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1676037725
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1676037725
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1676037725
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1676037725
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1676037725
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1676037725
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1676037725
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1676037725
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1676037725
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1676037725
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1676037725
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1676037725
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1676037725
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1676037725
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1676037725
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1676037725
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1676037725
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_205
timestamp 1676037725
transform 1 0 19964 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_211
timestamp 1676037725
transform 1 0 20516 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_215
timestamp 1676037725
transform 1 0 20884 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_222
timestamp 1676037725
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_225
timestamp 1676037725
transform 1 0 21804 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_244
timestamp 1676037725
transform 1 0 23552 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_264
timestamp 1676037725
transform 1 0 25392 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1676037725
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1676037725
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1676037725
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1676037725
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1676037725
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1676037725
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1676037725
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1676037725
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1676037725
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1676037725
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1676037725
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1676037725
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1676037725
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1676037725
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1676037725
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1676037725
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1676037725
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1676037725
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1676037725
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_197
timestamp 1676037725
transform 1 0 19228 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_203
timestamp 1676037725
transform 1 0 19780 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_209
timestamp 1676037725
transform 1 0 20332 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_216
timestamp 1676037725
transform 1 0 20976 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_223
timestamp 1676037725
transform 1 0 21620 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_230
timestamp 1676037725
transform 1 0 22264 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_250
timestamp 1676037725
transform 1 0 24104 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_253
timestamp 1676037725
transform 1 0 24380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_259
timestamp 1676037725
transform 1 0 24932 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_265
timestamp 1676037725
transform 1 0 25484 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1676037725
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1676037725
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1676037725
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1676037725
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1676037725
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1676037725
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1676037725
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1676037725
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1676037725
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1676037725
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1676037725
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1676037725
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1676037725
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1676037725
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1676037725
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1676037725
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1676037725
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1676037725
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1676037725
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1676037725
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_193
timestamp 1676037725
transform 1 0 18860 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_202
timestamp 1676037725
transform 1 0 19688 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_209
timestamp 1676037725
transform 1 0 20332 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_216
timestamp 1676037725
transform 1 0 20976 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_222
timestamp 1676037725
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_225
timestamp 1676037725
transform 1 0 21804 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_244
timestamp 1676037725
transform 1 0 23552 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_264
timestamp 1676037725
transform 1 0 25392 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1676037725
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1676037725
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1676037725
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1676037725
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1676037725
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1676037725
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1676037725
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1676037725
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1676037725
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1676037725
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_117
timestamp 1676037725
transform 1 0 11868 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1676037725
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1676037725
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1676037725
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1676037725
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1676037725
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1676037725
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1676037725
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_189
timestamp 1676037725
transform 1 0 18492 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_193
timestamp 1676037725
transform 1 0 18860 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_197
timestamp 1676037725
transform 1 0 19228 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_209
timestamp 1676037725
transform 1 0 20332 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_217
timestamp 1676037725
transform 1 0 21068 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_222
timestamp 1676037725
transform 1 0 21528 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_226
timestamp 1676037725
transform 1 0 21896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_230
timestamp 1676037725
transform 1 0 22264 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_250
timestamp 1676037725
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_253
timestamp 1676037725
transform 1 0 24380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_259
timestamp 1676037725
transform 1 0 24932 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_265
timestamp 1676037725
transform 1 0 25484 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1676037725
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1676037725
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1676037725
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1676037725
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1676037725
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1676037725
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1676037725
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1676037725
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1676037725
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1676037725
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1676037725
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1676037725
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1676037725
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1676037725
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1676037725
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1676037725
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1676037725
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1676037725
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1676037725
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_181
timestamp 1676037725
transform 1 0 17756 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_187
timestamp 1676037725
transform 1 0 18308 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_194
timestamp 1676037725
transform 1 0 18952 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_201
timestamp 1676037725
transform 1 0 19596 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_208
timestamp 1676037725
transform 1 0 20240 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_212
timestamp 1676037725
transform 1 0 20608 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_216
timestamp 1676037725
transform 1 0 20976 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_225
timestamp 1676037725
transform 1 0 21804 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_244
timestamp 1676037725
transform 1 0 23552 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_264
timestamp 1676037725
transform 1 0 25392 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1676037725
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1676037725
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1676037725
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1676037725
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1676037725
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1676037725
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1676037725
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1676037725
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1676037725
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1676037725
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1676037725
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1676037725
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1676037725
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1676037725
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1676037725
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1676037725
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1676037725
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1676037725
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_180
timestamp 1676037725
transform 1 0 17664 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1676037725
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_197
timestamp 1676037725
transform 1 0 19228 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_202
timestamp 1676037725
transform 1 0 19688 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_209
timestamp 1676037725
transform 1 0 20332 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_216
timestamp 1676037725
transform 1 0 20976 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_241
timestamp 1676037725
transform 1 0 23276 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_250
timestamp 1676037725
transform 1 0 24104 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1676037725
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_264
timestamp 1676037725
transform 1 0 25392 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1676037725
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1676037725
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1676037725
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1676037725
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1676037725
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1676037725
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1676037725
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1676037725
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1676037725
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1676037725
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1676037725
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1676037725
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1676037725
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1676037725
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1676037725
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_149
timestamp 1676037725
transform 1 0 14812 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_157
timestamp 1676037725
transform 1 0 15548 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_161
timestamp 1676037725
transform 1 0 15916 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_165
timestamp 1676037725
transform 1 0 16284 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1676037725
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_180
timestamp 1676037725
transform 1 0 17664 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_187
timestamp 1676037725
transform 1 0 18308 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_194
timestamp 1676037725
transform 1 0 18952 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_201
timestamp 1676037725
transform 1 0 19596 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_208
timestamp 1676037725
transform 1 0 20240 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_215
timestamp 1676037725
transform 1 0 20884 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 1676037725
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_225
timestamp 1676037725
transform 1 0 21804 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_244
timestamp 1676037725
transform 1 0 23552 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_264
timestamp 1676037725
transform 1 0 25392 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1676037725
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1676037725
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1676037725
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1676037725
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1676037725
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1676037725
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1676037725
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1676037725
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1676037725
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1676037725
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1676037725
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1676037725
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1676037725
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1676037725
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1676037725
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_141
timestamp 1676037725
transform 1 0 14076 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_16_149
timestamp 1676037725
transform 1 0 14812 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_155
timestamp 1676037725
transform 1 0 15364 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_159
timestamp 1676037725
transform 1 0 15732 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_166
timestamp 1676037725
transform 1 0 16376 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_173
timestamp 1676037725
transform 1 0 17020 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_180
timestamp 1676037725
transform 1 0 17664 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_187
timestamp 1676037725
transform 1 0 18308 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1676037725
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_201
timestamp 1676037725
transform 1 0 19596 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_208
timestamp 1676037725
transform 1 0 20240 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_216
timestamp 1676037725
transform 1 0 20976 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_221
timestamp 1676037725
transform 1 0 21436 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_225
timestamp 1676037725
transform 1 0 21804 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_230
timestamp 1676037725
transform 1 0 22264 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_250
timestamp 1676037725
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_253
timestamp 1676037725
transform 1 0 24380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_258
timestamp 1676037725
transform 1 0 24840 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1676037725
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1676037725
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1676037725
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1676037725
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1676037725
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1676037725
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1676037725
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1676037725
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1676037725
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1676037725
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1676037725
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1676037725
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1676037725
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_125
timestamp 1676037725
transform 1 0 12604 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_147
timestamp 1676037725
transform 1 0 14628 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_151
timestamp 1676037725
transform 1 0 14996 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_155
timestamp 1676037725
transform 1 0 15364 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_161
timestamp 1676037725
transform 1 0 15916 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1676037725
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_171
timestamp 1676037725
transform 1 0 16836 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_194
timestamp 1676037725
transform 1 0 18952 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_198
timestamp 1676037725
transform 1 0 19320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_219
timestamp 1676037725
transform 1 0 21252 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1676037725
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_225
timestamp 1676037725
transform 1 0 21804 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_244
timestamp 1676037725
transform 1 0 23552 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_264
timestamp 1676037725
transform 1 0 25392 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1676037725
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1676037725
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1676037725
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1676037725
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1676037725
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1676037725
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1676037725
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1676037725
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1676037725
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1676037725
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1676037725
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1676037725
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1676037725
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_133
timestamp 1676037725
transform 1 0 13340 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1676037725
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_153
timestamp 1676037725
transform 1 0 15180 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_157
timestamp 1676037725
transform 1 0 15548 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_179
timestamp 1676037725
transform 1 0 17572 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_186
timestamp 1676037725
transform 1 0 18216 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1676037725
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_197
timestamp 1676037725
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_219
timestamp 1676037725
transform 1 0 21252 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_226
timestamp 1676037725
transform 1 0 21896 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_250
timestamp 1676037725
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_257
timestamp 1676037725
transform 1 0 24748 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_263
timestamp 1676037725
transform 1 0 25300 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1676037725
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1676037725
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1676037725
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1676037725
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1676037725
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1676037725
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1676037725
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1676037725
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1676037725
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1676037725
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1676037725
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1676037725
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_115
timestamp 1676037725
transform 1 0 11684 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_123
timestamp 1676037725
transform 1 0 12420 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_126
timestamp 1676037725
transform 1 0 12696 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_149
timestamp 1676037725
transform 1 0 14812 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_163
timestamp 1676037725
transform 1 0 16100 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1676037725
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1676037725
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_191
timestamp 1676037725
transform 1 0 18676 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_204
timestamp 1676037725
transform 1 0 19872 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_217
timestamp 1676037725
transform 1 0 21068 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1676037725
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1676037725
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_247
timestamp 1676037725
transform 1 0 23828 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_253
timestamp 1676037725
transform 1 0 24380 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_258
timestamp 1676037725
transform 1 0 24840 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1676037725
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1676037725
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1676037725
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1676037725
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1676037725
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1676037725
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1676037725
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1676037725
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1676037725
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_85
timestamp 1676037725
transform 1 0 8924 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_91
timestamp 1676037725
transform 1 0 9476 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_112
timestamp 1676037725
transform 1 0 11408 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_136
timestamp 1676037725
transform 1 0 13616 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1676037725
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_163
timestamp 1676037725
transform 1 0 16100 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_187
timestamp 1676037725
transform 1 0 18308 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1676037725
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_199
timestamp 1676037725
transform 1 0 19412 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_222
timestamp 1676037725
transform 1 0 21528 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_246
timestamp 1676037725
transform 1 0 23736 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_264
timestamp 1676037725
transform 1 0 25392 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1676037725
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1676037725
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1676037725
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1676037725
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1676037725
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1676037725
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1676037725
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1676037725
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1676037725
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1676037725
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_105
timestamp 1676037725
transform 1 0 10764 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_113
timestamp 1676037725
transform 1 0 11500 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_119
timestamp 1676037725
transform 1 0 12052 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_126
timestamp 1676037725
transform 1 0 12696 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_133
timestamp 1676037725
transform 1 0 13340 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_157
timestamp 1676037725
transform 1 0 15548 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_161
timestamp 1676037725
transform 1 0 15916 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1676037725
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_171
timestamp 1676037725
transform 1 0 16836 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_182
timestamp 1676037725
transform 1 0 17848 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_206
timestamp 1676037725
transform 1 0 20056 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_210
timestamp 1676037725
transform 1 0 20424 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1676037725
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_225
timestamp 1676037725
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_231
timestamp 1676037725
transform 1 0 22356 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_235
timestamp 1676037725
transform 1 0 22724 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_256
timestamp 1676037725
transform 1 0 24656 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_264
timestamp 1676037725
transform 1 0 25392 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1676037725
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1676037725
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1676037725
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1676037725
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1676037725
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1676037725
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1676037725
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1676037725
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1676037725
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1676037725
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_97
timestamp 1676037725
transform 1 0 10028 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_102
timestamp 1676037725
transform 1 0 10488 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_124
timestamp 1676037725
transform 1 0 12512 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_131
timestamp 1676037725
transform 1 0 13156 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1676037725
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1676037725
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_163
timestamp 1676037725
transform 1 0 16100 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_187
timestamp 1676037725
transform 1 0 18308 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1676037725
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1676037725
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_208
timestamp 1676037725
transform 1 0 20240 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_212
timestamp 1676037725
transform 1 0 20608 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_234
timestamp 1676037725
transform 1 0 22632 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_238
timestamp 1676037725
transform 1 0 23000 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_250
timestamp 1676037725
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_253
timestamp 1676037725
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_259
timestamp 1676037725
transform 1 0 24932 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_265
timestamp 1676037725
transform 1 0 25484 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1676037725
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1676037725
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1676037725
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1676037725
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1676037725
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1676037725
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1676037725
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1676037725
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_81
timestamp 1676037725
transform 1 0 8556 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_89
timestamp 1676037725
transform 1 0 9292 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_98
timestamp 1676037725
transform 1 0 10120 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_103
timestamp 1676037725
transform 1 0 10580 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1676037725
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_113
timestamp 1676037725
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_135
timestamp 1676037725
transform 1 0 13524 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_142
timestamp 1676037725
transform 1 0 14168 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_147
timestamp 1676037725
transform 1 0 14628 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_152
timestamp 1676037725
transform 1 0 15088 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_159
timestamp 1676037725
transform 1 0 15732 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1676037725
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_169
timestamp 1676037725
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_191
timestamp 1676037725
transform 1 0 18676 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_196
timestamp 1676037725
transform 1 0 19136 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_218
timestamp 1676037725
transform 1 0 21160 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_225
timestamp 1676037725
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_231
timestamp 1676037725
transform 1 0 22356 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_235
timestamp 1676037725
transform 1 0 22724 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_256
timestamp 1676037725
transform 1 0 24656 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_263
timestamp 1676037725
transform 1 0 25300 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1676037725
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1676037725
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1676037725
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1676037725
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1676037725
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1676037725
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1676037725
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_77
timestamp 1676037725
transform 1 0 8188 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_81
timestamp 1676037725
transform 1 0 8556 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_85
timestamp 1676037725
transform 1 0 8924 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_91
timestamp 1676037725
transform 1 0 9476 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_98
timestamp 1676037725
transform 1 0 10120 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_122
timestamp 1676037725
transform 1 0 12328 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_135
timestamp 1676037725
transform 1 0 13524 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1676037725
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1676037725
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_163
timestamp 1676037725
transform 1 0 16100 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_167
timestamp 1676037725
transform 1 0 16468 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_170
timestamp 1676037725
transform 1 0 16744 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_192
timestamp 1676037725
transform 1 0 18768 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_197
timestamp 1676037725
transform 1 0 19228 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_209
timestamp 1676037725
transform 1 0 20332 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_222
timestamp 1676037725
transform 1 0 21528 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_230
timestamp 1676037725
transform 1 0 22264 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_238
timestamp 1676037725
transform 1 0 23000 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_245
timestamp 1676037725
transform 1 0 23644 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1676037725
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_255
timestamp 1676037725
transform 1 0 24564 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_261
timestamp 1676037725
transform 1 0 25116 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_265
timestamp 1676037725
transform 1 0 25484 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1676037725
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1676037725
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_27
timestamp 1676037725
transform 1 0 3588 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_33
timestamp 1676037725
transform 1 0 4140 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_36
timestamp 1676037725
transform 1 0 4416 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_48
timestamp 1676037725
transform 1 0 5520 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1676037725
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_69
timestamp 1676037725
transform 1 0 7452 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_73
timestamp 1676037725
transform 1 0 7820 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_78
timestamp 1676037725
transform 1 0 8280 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_83
timestamp 1676037725
transform 1 0 8740 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_90
timestamp 1676037725
transform 1 0 9384 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_97
timestamp 1676037725
transform 1 0 10028 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1676037725
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_113
timestamp 1676037725
transform 1 0 11500 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_135
timestamp 1676037725
transform 1 0 13524 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_148
timestamp 1676037725
transform 1 0 14720 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_154
timestamp 1676037725
transform 1 0 15272 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_165
timestamp 1676037725
transform 1 0 16284 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_171
timestamp 1676037725
transform 1 0 16836 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_194
timestamp 1676037725
transform 1 0 18952 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_207
timestamp 1676037725
transform 1 0 20148 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_220
timestamp 1676037725
transform 1 0 21344 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_225
timestamp 1676037725
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_236
timestamp 1676037725
transform 1 0 22816 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_240
timestamp 1676037725
transform 1 0 23184 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_251
timestamp 1676037725
transform 1 0 24196 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_259
timestamp 1676037725
transform 1 0 24932 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_265
timestamp 1676037725
transform 1 0 25484 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1676037725
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1676037725
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1676037725
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp 1676037725
transform 1 0 3772 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_34
timestamp 1676037725
transform 1 0 4232 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_38
timestamp 1676037725
transform 1 0 4600 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_42
timestamp 1676037725
transform 1 0 4968 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_54
timestamp 1676037725
transform 1 0 6072 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_64
timestamp 1676037725
transform 1 0 6992 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_70
timestamp 1676037725
transform 1 0 7544 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_75
timestamp 1676037725
transform 1 0 8004 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 1676037725
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_89
timestamp 1676037725
transform 1 0 9292 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_94
timestamp 1676037725
transform 1 0 9752 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_101
timestamp 1676037725
transform 1 0 10396 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_114
timestamp 1676037725
transform 1 0 11592 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1676037725
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_141
timestamp 1676037725
transform 1 0 14076 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_163
timestamp 1676037725
transform 1 0 16100 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_170
timestamp 1676037725
transform 1 0 16744 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1676037725
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1676037725
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_219
timestamp 1676037725
transform 1 0 21252 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_226
timestamp 1676037725
transform 1 0 21896 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_250
timestamp 1676037725
transform 1 0 24104 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_253
timestamp 1676037725
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_263
timestamp 1676037725
transform 1 0 25300 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1676037725
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1676037725
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_27
timestamp 1676037725
transform 1 0 3588 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_33
timestamp 1676037725
transform 1 0 4140 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_47
timestamp 1676037725
transform 1 0 5428 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1676037725
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_57
timestamp 1676037725
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_62
timestamp 1676037725
transform 1 0 6808 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_69
timestamp 1676037725
transform 1 0 7452 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_76
timestamp 1676037725
transform 1 0 8096 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_80
timestamp 1676037725
transform 1 0 8464 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_84
timestamp 1676037725
transform 1 0 8832 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_108
timestamp 1676037725
transform 1 0 11040 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 1676037725
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_135
timestamp 1676037725
transform 1 0 13524 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_142
timestamp 1676037725
transform 1 0 14168 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_146
timestamp 1676037725
transform 1 0 14536 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_152
timestamp 1676037725
transform 1 0 15088 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_165
timestamp 1676037725
transform 1 0 16284 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1676037725
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_180
timestamp 1676037725
transform 1 0 17664 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_184
timestamp 1676037725
transform 1 0 18032 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_207
timestamp 1676037725
transform 1 0 20148 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_214
timestamp 1676037725
transform 1 0 20792 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_221
timestamp 1676037725
transform 1 0 21436 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_231
timestamp 1676037725
transform 1 0 22356 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_253
timestamp 1676037725
transform 1 0 24380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_261
timestamp 1676037725
transform 1 0 25116 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_265
timestamp 1676037725
transform 1 0 25484 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1676037725
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_15
timestamp 1676037725
transform 1 0 2484 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_26
timestamp 1676037725
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_29
timestamp 1676037725
transform 1 0 3772 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_35
timestamp 1676037725
transform 1 0 4324 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_40
timestamp 1676037725
transform 1 0 4784 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_54
timestamp 1676037725
transform 1 0 6072 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_61
timestamp 1676037725
transform 1 0 6716 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_68
timestamp 1676037725
transform 1 0 7360 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_75
timestamp 1676037725
transform 1 0 8004 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1676037725
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_85
timestamp 1676037725
transform 1 0 8924 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_90
timestamp 1676037725
transform 1 0 9384 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_114
timestamp 1676037725
transform 1 0 11592 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1676037725
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_141
timestamp 1676037725
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_146
timestamp 1676037725
transform 1 0 14536 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_170
timestamp 1676037725
transform 1 0 16744 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_183
timestamp 1676037725
transform 1 0 17940 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_187
timestamp 1676037725
transform 1 0 18308 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_193
timestamp 1676037725
transform 1 0 18860 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1676037725
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_208
timestamp 1676037725
transform 1 0 20240 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_212
timestamp 1676037725
transform 1 0 20608 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_233
timestamp 1676037725
transform 1 0 22540 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_239
timestamp 1676037725
transform 1 0 23092 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_250
timestamp 1676037725
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_264
timestamp 1676037725
transform 1 0 25392 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1676037725
transform 1 0 1380 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_8
timestamp 1676037725
transform 1 0 1840 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_15
timestamp 1676037725
transform 1 0 2484 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_21
timestamp 1676037725
transform 1 0 3036 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_26
timestamp 1676037725
transform 1 0 3496 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_33
timestamp 1676037725
transform 1 0 4140 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_40
timestamp 1676037725
transform 1 0 4784 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_47
timestamp 1676037725
transform 1 0 5428 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_54
timestamp 1676037725
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_57
timestamp 1676037725
transform 1 0 6348 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_62
timestamp 1676037725
transform 1 0 6808 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_67
timestamp 1676037725
transform 1 0 7268 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_74
timestamp 1676037725
transform 1 0 7912 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_81
timestamp 1676037725
transform 1 0 8556 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_105
timestamp 1676037725
transform 1 0 10764 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_113
timestamp 1676037725
transform 1 0 11500 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_125
timestamp 1676037725
transform 1 0 12604 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_149
timestamp 1676037725
transform 1 0 14812 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_162
timestamp 1676037725
transform 1 0 16008 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1676037725
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_180
timestamp 1676037725
transform 1 0 17664 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_193
timestamp 1676037725
transform 1 0 18860 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_206
timestamp 1676037725
transform 1 0 20056 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_219
timestamp 1676037725
transform 1 0 21252 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1676037725
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_225
timestamp 1676037725
transform 1 0 21804 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_247
timestamp 1676037725
transform 1 0 23828 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_253
timestamp 1676037725
transform 1 0 24380 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_264
timestamp 1676037725
transform 1 0 25392 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1676037725
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_7
timestamp 1676037725
transform 1 0 1748 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_12
timestamp 1676037725
transform 1 0 2208 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_19
timestamp 1676037725
transform 1 0 2852 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_26
timestamp 1676037725
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_35
timestamp 1676037725
transform 1 0 4324 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_40
timestamp 1676037725
transform 1 0 4784 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_47
timestamp 1676037725
transform 1 0 5428 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_54
timestamp 1676037725
transform 1 0 6072 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_61
timestamp 1676037725
transform 1 0 6716 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_75
timestamp 1676037725
transform 1 0 8004 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_82
timestamp 1676037725
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_85
timestamp 1676037725
transform 1 0 8924 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_97
timestamp 1676037725
transform 1 0 10028 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_121
timestamp 1676037725
transform 1 0 12236 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_127
timestamp 1676037725
transform 1 0 12788 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1676037725
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_141
timestamp 1676037725
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_152
timestamp 1676037725
transform 1 0 15088 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_176
timestamp 1676037725
transform 1 0 17296 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_182
timestamp 1676037725
transform 1 0 17848 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_193
timestamp 1676037725
transform 1 0 18860 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_197
timestamp 1676037725
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_202
timestamp 1676037725
transform 1 0 19688 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_206
timestamp 1676037725
transform 1 0 20056 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_229
timestamp 1676037725
transform 1 0 22172 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_242
timestamp 1676037725
transform 1 0 23368 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_264
timestamp 1676037725
transform 1 0 25392 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 1676037725
transform 1 0 1380 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_23
timestamp 1676037725
transform 1 0 3220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_29
timestamp 1676037725
transform 1 0 3772 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_33
timestamp 1676037725
transform 1 0 4140 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_47
timestamp 1676037725
transform 1 0 5428 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_54
timestamp 1676037725
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_63
timestamp 1676037725
transform 1 0 6900 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_68
timestamp 1676037725
transform 1 0 7360 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_75
timestamp 1676037725
transform 1 0 8004 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_82
timestamp 1676037725
transform 1 0 8648 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_106
timestamp 1676037725
transform 1 0 10856 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_117
timestamp 1676037725
transform 1 0 11868 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_122
timestamp 1676037725
transform 1 0 12328 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_146
timestamp 1676037725
transform 1 0 14536 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_159
timestamp 1676037725
transform 1 0 15732 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_166
timestamp 1676037725
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_171
timestamp 1676037725
transform 1 0 16836 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_193
timestamp 1676037725
transform 1 0 18860 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_206
timestamp 1676037725
transform 1 0 20056 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_219
timestamp 1676037725
transform 1 0 21252 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1676037725
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_236
timestamp 1676037725
transform 1 0 22816 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_240
timestamp 1676037725
transform 1 0 23184 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_261
timestamp 1676037725
transform 1 0 25116 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_265
timestamp 1676037725
transform 1 0 25484 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_3
timestamp 1676037725
transform 1 0 1380 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_9
timestamp 1676037725
transform 1 0 1932 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_26
timestamp 1676037725
transform 1 0 3496 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_29
timestamp 1676037725
transform 1 0 3772 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_40
timestamp 1676037725
transform 1 0 4784 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_54
timestamp 1676037725
transform 1 0 6072 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_61
timestamp 1676037725
transform 1 0 6716 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_75
timestamp 1676037725
transform 1 0 8004 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_82
timestamp 1676037725
transform 1 0 8648 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_85
timestamp 1676037725
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_90
timestamp 1676037725
transform 1 0 9384 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_97
timestamp 1676037725
transform 1 0 10028 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_110
timestamp 1676037725
transform 1 0 11224 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_134
timestamp 1676037725
transform 1 0 13432 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_141
timestamp 1676037725
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_146
timestamp 1676037725
transform 1 0 14536 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_159
timestamp 1676037725
transform 1 0 15732 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_167
timestamp 1676037725
transform 1 0 16468 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_171
timestamp 1676037725
transform 1 0 16836 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_176
timestamp 1676037725
transform 1 0 17296 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_189
timestamp 1676037725
transform 1 0 18492 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1676037725
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_197
timestamp 1676037725
transform 1 0 19228 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_208
timestamp 1676037725
transform 1 0 20240 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_214
timestamp 1676037725
transform 1 0 20792 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_237
timestamp 1676037725
transform 1 0 22908 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_250
timestamp 1676037725
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_253
timestamp 1676037725
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_264
timestamp 1676037725
transform 1 0 25392 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1676037725
transform 1 0 1380 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_8
timestamp 1676037725
transform 1 0 1840 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_15
timestamp 1676037725
transform 1 0 2484 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_35
timestamp 1676037725
transform 1 0 4324 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_39
timestamp 1676037725
transform 1 0 4692 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_42
timestamp 1676037725
transform 1 0 4968 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_47
timestamp 1676037725
transform 1 0 5428 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 1676037725
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_57
timestamp 1676037725
transform 1 0 6348 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_63
timestamp 1676037725
transform 1 0 6900 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_68
timestamp 1676037725
transform 1 0 7360 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_75
timestamp 1676037725
transform 1 0 8004 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_82
timestamp 1676037725
transform 1 0 8648 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_106
timestamp 1676037725
transform 1 0 10856 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_117
timestamp 1676037725
transform 1 0 11868 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_128
timestamp 1676037725
transform 1 0 12880 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_133
timestamp 1676037725
transform 1 0 13340 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_155
timestamp 1676037725
transform 1 0 15364 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_163
timestamp 1676037725
transform 1 0 16100 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1676037725
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_169
timestamp 1676037725
transform 1 0 16652 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_192
timestamp 1676037725
transform 1 0 18768 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_196
timestamp 1676037725
transform 1 0 19136 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_217
timestamp 1676037725
transform 1 0 21068 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1676037725
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_225
timestamp 1676037725
transform 1 0 21804 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_237
timestamp 1676037725
transform 1 0 22908 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_241
timestamp 1676037725
transform 1 0 23276 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_263
timestamp 1676037725
transform 1 0 25300 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_34_3
timestamp 1676037725
transform 1 0 1380 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_9
timestamp 1676037725
transform 1 0 1932 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_26
timestamp 1676037725
transform 1 0 3496 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_29
timestamp 1676037725
transform 1 0 3772 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_47
timestamp 1676037725
transform 1 0 5428 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_54
timestamp 1676037725
transform 1 0 6072 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_58
timestamp 1676037725
transform 1 0 6440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_61
timestamp 1676037725
transform 1 0 6716 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_79
timestamp 1676037725
transform 1 0 8372 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_87
timestamp 1676037725
transform 1 0 9108 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_92
timestamp 1676037725
transform 1 0 9568 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_105
timestamp 1676037725
transform 1 0 10764 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_129
timestamp 1676037725
transform 1 0 12972 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_133
timestamp 1676037725
transform 1 0 13340 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_138
timestamp 1676037725
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_141
timestamp 1676037725
transform 1 0 14076 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_147
timestamp 1676037725
transform 1 0 14628 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_153
timestamp 1676037725
transform 1 0 15180 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_165
timestamp 1676037725
transform 1 0 16284 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_178
timestamp 1676037725
transform 1 0 17480 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_191
timestamp 1676037725
transform 1 0 18676 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1676037725
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_197
timestamp 1676037725
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_219
timestamp 1676037725
transform 1 0 21252 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_232
timestamp 1676037725
transform 1 0 22448 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_245
timestamp 1676037725
transform 1 0 23644 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1676037725
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_253
timestamp 1676037725
transform 1 0 24380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_264
timestamp 1676037725
transform 1 0 25392 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1676037725
transform 1 0 1380 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_9
timestamp 1676037725
transform 1 0 1932 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_13
timestamp 1676037725
transform 1 0 2300 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_17
timestamp 1676037725
transform 1 0 2668 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_34
timestamp 1676037725
transform 1 0 4232 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_54
timestamp 1676037725
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_57
timestamp 1676037725
transform 1 0 6348 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_62
timestamp 1676037725
transform 1 0 6808 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_82
timestamp 1676037725
transform 1 0 8648 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_106
timestamp 1676037725
transform 1 0 10856 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_119
timestamp 1676037725
transform 1 0 12052 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_130
timestamp 1676037725
transform 1 0 13064 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_136
timestamp 1676037725
transform 1 0 13616 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_147
timestamp 1676037725
transform 1 0 14628 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_160
timestamp 1676037725
transform 1 0 15824 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_171
timestamp 1676037725
transform 1 0 16836 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_182
timestamp 1676037725
transform 1 0 17848 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_206
timestamp 1676037725
transform 1 0 20056 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_219
timestamp 1676037725
transform 1 0 21252 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1676037725
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1676037725
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_236
timestamp 1676037725
transform 1 0 22816 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_240
timestamp 1676037725
transform 1 0 23184 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_262
timestamp 1676037725
transform 1 0 25208 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_3
timestamp 1676037725
transform 1 0 1380 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_8
timestamp 1676037725
transform 1 0 1840 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_26
timestamp 1676037725
transform 1 0 3496 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_29
timestamp 1676037725
transform 1 0 3772 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_41
timestamp 1676037725
transform 1 0 4876 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_45
timestamp 1676037725
transform 1 0 5244 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_62
timestamp 1676037725
transform 1 0 6808 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_82
timestamp 1676037725
transform 1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_87
timestamp 1676037725
transform 1 0 9108 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_92
timestamp 1676037725
transform 1 0 9568 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_96
timestamp 1676037725
transform 1 0 9936 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_100
timestamp 1676037725
transform 1 0 10304 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_124
timestamp 1676037725
transform 1 0 12512 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_36_131
timestamp 1676037725
transform 1 0 13156 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_138
timestamp 1676037725
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_141
timestamp 1676037725
transform 1 0 14076 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_163
timestamp 1676037725
transform 1 0 16100 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_176
timestamp 1676037725
transform 1 0 17296 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_189
timestamp 1676037725
transform 1 0 18492 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1676037725
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_197
timestamp 1676037725
transform 1 0 19228 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_203
timestamp 1676037725
transform 1 0 19780 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_207
timestamp 1676037725
transform 1 0 20148 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_229
timestamp 1676037725
transform 1 0 22172 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_236
timestamp 1676037725
transform 1 0 22816 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_250
timestamp 1676037725
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_253
timestamp 1676037725
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_264
timestamp 1676037725
transform 1 0 25392 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1676037725
transform 1 0 1380 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_9
timestamp 1676037725
transform 1 0 1932 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_16
timestamp 1676037725
transform 1 0 2576 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_34
timestamp 1676037725
transform 1 0 4232 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_54
timestamp 1676037725
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_57
timestamp 1676037725
transform 1 0 6348 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_63
timestamp 1676037725
transform 1 0 6900 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_68
timestamp 1676037725
transform 1 0 7360 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_86
timestamp 1676037725
transform 1 0 9016 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_110
timestamp 1676037725
transform 1 0 11224 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_113
timestamp 1676037725
transform 1 0 11500 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_124
timestamp 1676037725
transform 1 0 12512 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_132
timestamp 1676037725
transform 1 0 13248 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_156
timestamp 1676037725
transform 1 0 15456 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_164
timestamp 1676037725
transform 1 0 16192 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_169
timestamp 1676037725
transform 1 0 16652 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_191
timestamp 1676037725
transform 1 0 18676 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_199
timestamp 1676037725
transform 1 0 19412 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_203
timestamp 1676037725
transform 1 0 19780 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_222
timestamp 1676037725
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_225
timestamp 1676037725
transform 1 0 21804 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_237
timestamp 1676037725
transform 1 0 22908 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_261
timestamp 1676037725
transform 1 0 25116 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_265
timestamp 1676037725
transform 1 0 25484 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_3
timestamp 1676037725
transform 1 0 1380 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_8
timestamp 1676037725
transform 1 0 1840 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_26
timestamp 1676037725
transform 1 0 3496 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_29
timestamp 1676037725
transform 1 0 3772 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_35
timestamp 1676037725
transform 1 0 4324 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_42
timestamp 1676037725
transform 1 0 4968 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_62
timestamp 1676037725
transform 1 0 6808 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_82
timestamp 1676037725
transform 1 0 8648 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_85
timestamp 1676037725
transform 1 0 8924 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_91
timestamp 1676037725
transform 1 0 9476 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_111
timestamp 1676037725
transform 1 0 11316 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_131
timestamp 1676037725
transform 1 0 13156 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_138
timestamp 1676037725
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_141
timestamp 1676037725
transform 1 0 14076 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_147
timestamp 1676037725
transform 1 0 14628 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_171
timestamp 1676037725
transform 1 0 16836 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_184
timestamp 1676037725
transform 1 0 18032 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_192
timestamp 1676037725
transform 1 0 18768 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_197
timestamp 1676037725
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_219
timestamp 1676037725
transform 1 0 21252 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_243
timestamp 1676037725
transform 1 0 23460 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_250
timestamp 1676037725
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_253
timestamp 1676037725
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_264
timestamp 1676037725
transform 1 0 25392 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_3
timestamp 1676037725
transform 1 0 1380 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_9
timestamp 1676037725
transform 1 0 1932 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_16
timestamp 1676037725
transform 1 0 2576 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_34
timestamp 1676037725
transform 1 0 4232 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_54
timestamp 1676037725
transform 1 0 6072 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_57
timestamp 1676037725
transform 1 0 6348 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_69
timestamp 1676037725
transform 1 0 7452 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_73
timestamp 1676037725
transform 1 0 7820 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_90
timestamp 1676037725
transform 1 0 9384 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_110
timestamp 1676037725
transform 1 0 11224 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_117
timestamp 1676037725
transform 1 0 11868 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_135
timestamp 1676037725
transform 1 0 13524 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_139
timestamp 1676037725
transform 1 0 13892 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_150
timestamp 1676037725
transform 1 0 14904 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_155
timestamp 1676037725
transform 1 0 15364 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_166
timestamp 1676037725
transform 1 0 16376 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_169
timestamp 1676037725
transform 1 0 16652 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_180
timestamp 1676037725
transform 1 0 17664 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_204
timestamp 1676037725
transform 1 0 19872 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_210
timestamp 1676037725
transform 1 0 20424 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_222
timestamp 1676037725
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_227
timestamp 1676037725
transform 1 0 21988 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_250
timestamp 1676037725
transform 1 0 24104 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_264
timestamp 1676037725
transform 1 0 25392 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_3
timestamp 1676037725
transform 1 0 1380 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_8
timestamp 1676037725
transform 1 0 1840 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_26
timestamp 1676037725
transform 1 0 3496 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_29
timestamp 1676037725
transform 1 0 3772 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_34
timestamp 1676037725
transform 1 0 4232 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_54
timestamp 1676037725
transform 1 0 6072 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_57
timestamp 1676037725
transform 1 0 6348 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_62
timestamp 1676037725
transform 1 0 6808 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_82
timestamp 1676037725
transform 1 0 8648 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_85
timestamp 1676037725
transform 1 0 8924 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_90
timestamp 1676037725
transform 1 0 9384 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_110
timestamp 1676037725
transform 1 0 11224 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_113
timestamp 1676037725
transform 1 0 11500 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_118
timestamp 1676037725
transform 1 0 11960 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_138
timestamp 1676037725
transform 1 0 13800 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_143
timestamp 1676037725
transform 1 0 14260 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_153
timestamp 1676037725
transform 1 0 15180 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_166
timestamp 1676037725
transform 1 0 16376 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_169
timestamp 1676037725
transform 1 0 16652 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_181
timestamp 1676037725
transform 1 0 17756 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_194
timestamp 1676037725
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_197
timestamp 1676037725
transform 1 0 19228 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_202
timestamp 1676037725
transform 1 0 19688 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_215
timestamp 1676037725
transform 1 0 20884 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_223
timestamp 1676037725
transform 1 0 21620 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_225
timestamp 1676037725
transform 1 0 21804 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_228
timestamp 1676037725
transform 1 0 22080 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_250
timestamp 1676037725
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_253
timestamp 1676037725
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_264
timestamp 1676037725
transform 1 0 25392 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14444 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold2 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20056 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold3
timestamp 1676037725
transform 1 0 24564 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold4 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6808 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold5
timestamp 1676037725
transform 1 0 8648 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1676037725
transform 1 0 6808 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1676037725
transform 1 0 20056 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1676037725
transform 1 0 21252 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1676037725
transform 1 0 8372 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1676037725
transform 1 0 12880 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1676037725
transform 1 0 9476 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1676037725
transform 1 0 8556 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1676037725
transform 1 0 2576 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1676037725
transform 1 0 13064 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1676037725
transform 1 0 10948 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1676037725
transform 1 0 8372 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1676037725
transform 1 0 7176 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1676037725
transform 1 0 16100 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1676037725
transform 1 0 19320 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1676037725
transform 1 0 18676 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1676037725
transform 1 0 18032 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1676037725
transform 1 0 17388 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1676037725
transform 1 0 15088 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1676037725
transform 1 0 15456 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1676037725
transform 1 0 12420 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1676037725
transform 1 0 11776 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1676037725
transform 1 0 10304 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1676037725
transform 1 0 9200 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1676037725
transform 1 0 20700 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1676037725
transform 1 0 21988 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1676037725
transform 1 0 18676 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1676037725
transform 1 0 16744 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1676037725
transform 1 0 18676 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1676037725
transform 1 0 24564 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1676037725
transform 1 0 23368 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1676037725
transform 1 0 16100 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1676037725
transform 1 0 1564 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input33
timestamp 1676037725
transform 1 0 3956 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1676037725
transform 1 0 16100 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1676037725
transform 1 0 18584 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1676037725
transform 1 0 3956 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1676037725
transform 1 0 16468 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1676037725
transform 1 0 14812 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1676037725
transform 1 0 7084 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1676037725
transform 1 0 6440 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1676037725
transform 1 0 7636 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1676037725
transform 1 0 6992 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1676037725
transform 1 0 3220 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1676037725
transform 1 0 4508 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1676037725
transform 1 0 5152 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1676037725
transform 1 0 7084 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1676037725
transform 1 0 9752 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1676037725
transform 1 0 4508 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1676037725
transform 1 0 9108 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1676037725
transform 1 0 1932 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1676037725
transform 1 0 9844 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1676037725
transform 1 0 19412 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1676037725
transform 1 0 16100 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1676037725
transform 1 0 9292 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1676037725
transform 1 0 6532 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input56
timestamp 1676037725
transform 1 0 6532 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1676037725
transform 1 0 9108 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1676037725
transform 1 0 6532 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1676037725
transform 1 0 19412 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1676037725
transform 1 0 7728 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1676037725
transform 1 0 22540 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  input62 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20056 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  input63
timestamp 1676037725
transform 1 0 25024 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input64
timestamp 1676037725
transform 1 0 20608 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input65
timestamp 1676037725
transform 1 0 23184 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input66
timestamp 1676037725
transform 1 0 21988 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input67
timestamp 1676037725
transform 1 0 1564 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input68
timestamp 1676037725
transform 1 0 1564 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input69
timestamp 1676037725
transform 1 0 3956 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input70
timestamp 1676037725
transform 1 0 1564 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_12  output71
timestamp 1676037725
transform 1 0 20056 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output72
timestamp 1676037725
transform 1 0 20056 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output73
timestamp 1676037725
transform 1 0 22080 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output74
timestamp 1676037725
transform 1 0 23920 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output75
timestamp 1676037725
transform 1 0 22632 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output76
timestamp 1676037725
transform 1 0 22080 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output77
timestamp 1676037725
transform 1 0 23920 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output78
timestamp 1676037725
transform 1 0 22632 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output79
timestamp 1676037725
transform 1 0 22080 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output80
timestamp 1676037725
transform 1 0 23920 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output81
timestamp 1676037725
transform 1 0 22632 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output82
timestamp 1676037725
transform 1 0 22080 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output83
timestamp 1676037725
transform 1 0 20792 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output84
timestamp 1676037725
transform 1 0 23920 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output85
timestamp 1676037725
transform 1 0 22632 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output86
timestamp 1676037725
transform 1 0 22080 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output87
timestamp 1676037725
transform 1 0 23920 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output88
timestamp 1676037725
transform 1 0 22080 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output89
timestamp 1676037725
transform 1 0 23920 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output90
timestamp 1676037725
transform 1 0 22632 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output91
timestamp 1676037725
transform 1 0 22080 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output92
timestamp 1676037725
transform 1 0 23920 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output93
timestamp 1676037725
transform 1 0 23920 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output94
timestamp 1676037725
transform 1 0 20056 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output95
timestamp 1676037725
transform 1 0 18216 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output96
timestamp 1676037725
transform 1 0 22632 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output97
timestamp 1676037725
transform 1 0 22080 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output98
timestamp 1676037725
transform 1 0 22632 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output99
timestamp 1676037725
transform 1 0 22080 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output100
timestamp 1676037725
transform 1 0 23920 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output101
timestamp 1676037725
transform 1 0 22632 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output102
timestamp 1676037725
transform 1 0 1748 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output103
timestamp 1676037725
transform 1 0 2760 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output104
timestamp 1676037725
transform 1 0 4600 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output105
timestamp 1676037725
transform 1 0 5336 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output106
timestamp 1676037725
transform 1 0 2024 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output107
timestamp 1676037725
transform 1 0 6900 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output108
timestamp 1676037725
transform 1 0 7176 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output109
timestamp 1676037725
transform 1 0 4600 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output110
timestamp 1676037725
transform 1 0 5336 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output111
timestamp 1676037725
transform 1 0 7176 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output112
timestamp 1676037725
transform 1 0 4600 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output113
timestamp 1676037725
transform 1 0 2024 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output114
timestamp 1676037725
transform 1 0 7544 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output115
timestamp 1676037725
transform 1 0 7176 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output116
timestamp 1676037725
transform 1 0 7176 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output117
timestamp 1676037725
transform 1 0 7912 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output118
timestamp 1676037725
transform 1 0 9844 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output119
timestamp 1676037725
transform 1 0 9752 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output120
timestamp 1676037725
transform 1 0 9752 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output121
timestamp 1676037725
transform 1 0 11684 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output122
timestamp 1676037725
transform 1 0 12052 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output123
timestamp 1676037725
transform 1 0 12328 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output124
timestamp 1676037725
transform 1 0 2024 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output125
timestamp 1676037725
transform 1 0 2852 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output126
timestamp 1676037725
transform 1 0 2024 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output127
timestamp 1676037725
transform 1 0 2760 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output128
timestamp 1676037725
transform 1 0 3956 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output129
timestamp 1676037725
transform 1 0 2760 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output130
timestamp 1676037725
transform 1 0 2024 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output131
timestamp 1676037725
transform 1 0 4600 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 25852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 25852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 25852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 25852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 25852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 25852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 25852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 25852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 25852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 25852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 25852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1676037725
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1676037725
transform -1 0 25852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1676037725
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1676037725
transform -1 0 25852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1676037725
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1676037725
transform -1 0 25852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1676037725
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1676037725
transform -1 0 25852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1676037725
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1676037725
transform -1 0 25852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1676037725
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1676037725
transform -1 0 25852 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1676037725
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1676037725
transform -1 0 25852 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1676037725
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1676037725
transform -1 0 25852 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1676037725
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1676037725
transform -1 0 25852 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1676037725
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1676037725
transform -1 0 25852 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1676037725
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1676037725
transform -1 0 25852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1676037725
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1676037725
transform -1 0 25852 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1676037725
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1676037725
transform -1 0 25852 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1676037725
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1676037725
transform -1 0 25852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1676037725
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1676037725
transform -1 0 25852 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1676037725
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1676037725
transform -1 0 25852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1676037725
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1676037725
transform -1 0 25852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1676037725
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1676037725
transform -1 0 25852 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1676037725
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1676037725
transform -1 0 25852 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1676037725
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1676037725
transform -1 0 25852 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1676037725
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1676037725
transform -1 0 25852 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1676037725
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1676037725
transform -1 0 25852 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1676037725
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1676037725
transform -1 0 25852 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1676037725
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1676037725
transform -1 0 25852 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1676037725
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1676037725
transform -1 0 25852 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1676037725
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1676037725
transform -1 0 25852 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1676037725
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1676037725
transform -1 0 25852 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1676037725
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1676037725
transform -1 0 25852 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1676037725
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1676037725
transform -1 0 25852 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1676037725
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1676037725
transform -1 0 25852 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14904 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 17020 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19228 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 20332 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21620 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22264 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22264 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 23276 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 23368 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 23460 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 23276 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22540 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21068 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 20332 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 20700 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22264 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22816 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22816 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22264 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 21988 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21896 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19688 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19320 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19412 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 18308 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 17112 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 16928 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 16836 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 16468 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 16468 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 15732 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 16836 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 17112 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19412 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19412 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__0_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_1_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21344 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 10028 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 14260 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 15456 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 16928 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19412 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19412 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 18032 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 16836 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 14996 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 13616 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 14260 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 13524 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 12696 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 11592 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11132 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 10672 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 9384 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 9016 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 9016 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 9016 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 8924 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 9200 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 9752 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 11684 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11960 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 11960 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11684 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 10488 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 10672 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 11684 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11776 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 12788 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 14260 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 13708 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 14260 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 14260 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_0.mux_l1_in_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17020 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_0.mux_l1_in_1__159 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23828 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_0.mux_l1_in_1_
timestamp 1676037725
transform 1 0 20424 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_0.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19228 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 24564 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_2.mux_l1_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_2.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_2.mux_l2_in_0__165
timestamp 1676037725
transform 1 0 2208 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 4508 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_4.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16928 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_4.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24564 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_4.mux_l2_in_0__134
timestamp 1676037725
transform 1 0 3864 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 14812 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_6.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_6.mux_l1_in_1_
timestamp 1676037725
transform 1 0 24564 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_6.mux_l1_in_1__139
timestamp 1676037725
transform 1 0 17388 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_6.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 8464 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_8.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15548 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_8.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_8.mux_l2_in_0__140
timestamp 1676037725
transform 1 0 13524 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 17388 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_10.mux_l1_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_10.mux_l2_in_0_
timestamp 1676037725
transform 1 0 23276 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_10.mux_l2_in_0__160
timestamp 1676037725
transform 1 0 16100 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 21988 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_12.mux_l1_in_0_
timestamp 1676037725
transform 1 0 21620 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_12.mux_l2_in_0__161
timestamp 1676037725
transform 1 0 4692 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_12.mux_l2_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 21988 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_14.mux_l1_in_0_
timestamp 1676037725
transform 1 0 22080 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_14.mux_l2_in_0_
timestamp 1676037725
transform 1 0 23368 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_14.mux_l2_in_0__162
timestamp 1676037725
transform 1 0 21988 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 21252 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_16.mux_l1_in_0_
timestamp 1676037725
transform 1 0 23276 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_16.mux_l2_in_0_
timestamp 1676037725
transform 1 0 23276 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_16.mux_l2_in_0__163
timestamp 1676037725
transform 1 0 23828 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19320 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_18.mux_l1_in_0_
timestamp 1676037725
transform 1 0 22540 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_18.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_18.mux_l2_in_0__164
timestamp 1676037725
transform 1 0 20056 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18676 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_28.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20424 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_28.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20700 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_28.mux_l2_in_0__166
timestamp 1676037725
transform 1 0 25024 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 20608 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_30.mux_l1_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_30.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20700 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_30.mux_l2_in_0__167
timestamp 1676037725
transform 1 0 25024 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 21252 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_32.mux_l1_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_32.mux_l2_in_0__132
timestamp 1676037725
transform 1 0 21620 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_32.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19504 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 21988 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_34.mux_l1_in_0_
timestamp 1676037725
transform 1 0 19228 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_34.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19412 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_34.mux_l2_in_0__133
timestamp 1676037725
transform 1 0 18676 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 21160 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_44.mux_l1_in_0_
timestamp 1676037725
transform 1 0 18032 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_44.mux_l2_in_0_
timestamp 1676037725
transform 1 0 17020 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_44.mux_l2_in_0__135
timestamp 1676037725
transform 1 0 17940 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_44.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 20700 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_46.mux_l1_in_0_
timestamp 1676037725
transform 1 0 18032 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_46.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19044 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_46.mux_l2_in_0__136
timestamp 1676037725
transform 1 0 18032 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_46.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 20700 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_48.mux_l1_in_0_
timestamp 1676037725
transform 1 0 19412 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_48.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20240 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_48.mux_l2_in_0__137
timestamp 1676037725
transform 1 0 21620 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_48.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 20608 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_50.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20516 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_50.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_50.mux_l2_in_0__138
timestamp 1676037725
transform 1 0 20056 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_50.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 21344 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_0.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14260 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_0.mux_l1_in_1_
timestamp 1676037725
transform 1 0 19412 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_0.mux_l1_in_1__141
timestamp 1676037725
transform 1 0 20516 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_0.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14904 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 11684 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_2.mux_l1_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_2.mux_l2_in_0_
timestamp 1676037725
transform 1 0 17848 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_2.mux_l2_in_0__147
timestamp 1676037725
transform 1 0 21160 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 13524 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_4.mux_l1_in_0_
timestamp 1676037725
transform 1 0 22816 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_4.mux_l2_in_0_
timestamp 1676037725
transform 1 0 18124 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_4.mux_l2_in_0__152
timestamp 1676037725
transform 1 0 15456 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 3956 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_6.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14996 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_6.mux_l1_in_1_
timestamp 1676037725
transform 1 0 15548 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_6.mux_l1_in_1__157
timestamp 1676037725
transform 1 0 5152 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_6.mux_l2_in_0_
timestamp 1676037725
transform 1 0 17204 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 3864 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_8.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20424 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_8.mux_l2_in_0__158
timestamp 1676037725
transform 1 0 19412 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_8.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14076 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 5796 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_10.mux_l1_in_0_
timestamp 1676037725
transform 1 0 17664 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_10.mux_l2_in_0_
timestamp 1676037725
transform 1 0 13800 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_10.mux_l2_in_0__142
timestamp 1676037725
transform 1 0 14260 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 8372 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_12.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16652 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_12.mux_l2_in_0__143
timestamp 1676037725
transform 1 0 10028 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_12.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12236 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 3220 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_14.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16468 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_14.mux_l2_in_0__144
timestamp 1676037725
transform 1 0 4692 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_14.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11684 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 9108 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_16.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15456 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_16.mux_l2_in_0_
timestamp 1676037725
transform 1 0 9936 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_16.mux_l2_in_0__145
timestamp 1676037725
transform 1 0 7728 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 8280 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_18.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14904 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_18.mux_l2_in_0_
timestamp 1676037725
transform 1 0 10396 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_18.mux_l2_in_0__146
timestamp 1676037725
transform 1 0 8372 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 5796 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_28.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15180 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_28.mux_l2_in_0__148
timestamp 1676037725
transform 1 0 9108 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_28.mux_l2_in_0_
timestamp 1676037725
transform 1 0 9200 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 1564 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_30.mux_l1_in_0_
timestamp 1676037725
transform 1 0 17664 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_30.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12052 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_30.mux_l2_in_0__149
timestamp 1676037725
transform 1 0 9292 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 6532 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_32.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_32.mux_l2_in_0__150
timestamp 1676037725
transform 1 0 12052 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_32.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11776 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 8372 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_34.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15456 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_34.mux_l2_in_0__151
timestamp 1676037725
transform 1 0 9752 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_34.mux_l2_in_0_
timestamp 1676037725
transform 1 0 10764 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 5796 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_44.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15456 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_44.mux_l2_in_0__153
timestamp 1676037725
transform 1 0 10120 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_44.mux_l2_in_0_
timestamp 1676037725
transform 1 0 10396 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_44.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 7084 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_46.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_46.mux_l2_in_0__154
timestamp 1676037725
transform 1 0 13892 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_46.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12696 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_46.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 7728 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_48.mux_l1_in_0_
timestamp 1676037725
transform 1 0 19320 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_48.mux_l2_in_0_
timestamp 1676037725
transform 1 0 13892 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_48.mux_l2_in_0__155
timestamp 1676037725
transform 1 0 13892 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_48.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 8372 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_50.mux_l1_in_0_
timestamp 1676037725
transform 1 0 17112 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_50.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12972 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_50.mux_l2_in_0__156
timestamp 1676037725
transform 1 0 14260 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_50.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 6440 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1676037725
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1676037725
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1676037725
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1676037725
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1676037725
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1676037725
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1676037725
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1676037725
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1676037725
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1676037725
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1676037725
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1676037725
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1676037725
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1676037725
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1676037725
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1676037725
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1676037725
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1676037725
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1676037725
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1676037725
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1676037725
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1676037725
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1676037725
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1676037725
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1676037725
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1676037725
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1676037725
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1676037725
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1676037725
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1676037725
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1676037725
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1676037725
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1676037725
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1676037725
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1676037725
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1676037725
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1676037725
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1676037725
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1676037725
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1676037725
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1676037725
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1676037725
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1676037725
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1676037725
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1676037725
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1676037725
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1676037725
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1676037725
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1676037725
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1676037725
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1676037725
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1676037725
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1676037725
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1676037725
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1676037725
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1676037725
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1676037725
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1676037725
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1676037725
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1676037725
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1676037725
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1676037725
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1676037725
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1676037725
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1676037725
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1676037725
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1676037725
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1676037725
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1676037725
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1676037725
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1676037725
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1676037725
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1676037725
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1676037725
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1676037725
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1676037725
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1676037725
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1676037725
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1676037725
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1676037725
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1676037725
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1676037725
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1676037725
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1676037725
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1676037725
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1676037725
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1676037725
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1676037725
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1676037725
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1676037725
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1676037725
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1676037725
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1676037725
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1676037725
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1676037725
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1676037725
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1676037725
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1676037725
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1676037725
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1676037725
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1676037725
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1676037725
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1676037725
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1676037725
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1676037725
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1676037725
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1676037725
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1676037725
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1676037725
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1676037725
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1676037725
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1676037725
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1676037725
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1676037725
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1676037725
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1676037725
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1676037725
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1676037725
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1676037725
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1676037725
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1676037725
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1676037725
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1676037725
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1676037725
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1676037725
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1676037725
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1676037725
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1676037725
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1676037725
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1676037725
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1676037725
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1676037725
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1676037725
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1676037725
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1676037725
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1676037725
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1676037725
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1676037725
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1676037725
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1676037725
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1676037725
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1676037725
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1676037725
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1676037725
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1676037725
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1676037725
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1676037725
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1676037725
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1676037725
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1676037725
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1676037725
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1676037725
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1676037725
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1676037725
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1676037725
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1676037725
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1676037725
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1676037725
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1676037725
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1676037725
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1676037725
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1676037725
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1676037725
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1676037725
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1676037725
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1676037725
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1676037725
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1676037725
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1676037725
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1676037725
transform 1 0 6256 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1676037725
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1676037725
transform 1 0 11408 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1676037725
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1676037725
transform 1 0 16560 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1676037725
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1676037725
transform 1 0 21712 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1676037725
transform 1 0 24288 0 1 23936
box -38 -48 130 592
<< labels >>
flabel metal4 s 7944 2128 8264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 17944 2128 18264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2944 2128 3264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 12944 2128 13264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 22944 2128 23264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 6734 0 6790 800 0 FreeSans 224 90 0 0 ccff_head
port 2 nsew signal input
flabel metal3 s 26200 280 27000 400 0 FreeSans 480 0 0 0 ccff_tail
port 3 nsew signal tristate
flabel metal3 s 26200 12928 27000 13048 0 FreeSans 480 0 0 0 chanx_right_in[0]
port 4 nsew signal input
flabel metal3 s 26200 17008 27000 17128 0 FreeSans 480 0 0 0 chanx_right_in[10]
port 5 nsew signal input
flabel metal3 s 26200 17416 27000 17536 0 FreeSans 480 0 0 0 chanx_right_in[11]
port 6 nsew signal input
flabel metal3 s 26200 17824 27000 17944 0 FreeSans 480 0 0 0 chanx_right_in[12]
port 7 nsew signal input
flabel metal3 s 26200 18232 27000 18352 0 FreeSans 480 0 0 0 chanx_right_in[13]
port 8 nsew signal input
flabel metal3 s 26200 18640 27000 18760 0 FreeSans 480 0 0 0 chanx_right_in[14]
port 9 nsew signal input
flabel metal3 s 26200 19048 27000 19168 0 FreeSans 480 0 0 0 chanx_right_in[15]
port 10 nsew signal input
flabel metal3 s 26200 19456 27000 19576 0 FreeSans 480 0 0 0 chanx_right_in[16]
port 11 nsew signal input
flabel metal3 s 26200 19864 27000 19984 0 FreeSans 480 0 0 0 chanx_right_in[17]
port 12 nsew signal input
flabel metal3 s 26200 20272 27000 20392 0 FreeSans 480 0 0 0 chanx_right_in[18]
port 13 nsew signal input
flabel metal3 s 26200 20680 27000 20800 0 FreeSans 480 0 0 0 chanx_right_in[19]
port 14 nsew signal input
flabel metal3 s 26200 13336 27000 13456 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 15 nsew signal input
flabel metal3 s 26200 21088 27000 21208 0 FreeSans 480 0 0 0 chanx_right_in[20]
port 16 nsew signal input
flabel metal3 s 26200 21496 27000 21616 0 FreeSans 480 0 0 0 chanx_right_in[21]
port 17 nsew signal input
flabel metal3 s 26200 21904 27000 22024 0 FreeSans 480 0 0 0 chanx_right_in[22]
port 18 nsew signal input
flabel metal3 s 26200 22312 27000 22432 0 FreeSans 480 0 0 0 chanx_right_in[23]
port 19 nsew signal input
flabel metal3 s 26200 22720 27000 22840 0 FreeSans 480 0 0 0 chanx_right_in[24]
port 20 nsew signal input
flabel metal3 s 26200 23128 27000 23248 0 FreeSans 480 0 0 0 chanx_right_in[25]
port 21 nsew signal input
flabel metal3 s 26200 23536 27000 23656 0 FreeSans 480 0 0 0 chanx_right_in[26]
port 22 nsew signal input
flabel metal3 s 26200 23944 27000 24064 0 FreeSans 480 0 0 0 chanx_right_in[27]
port 23 nsew signal input
flabel metal3 s 26200 24352 27000 24472 0 FreeSans 480 0 0 0 chanx_right_in[28]
port 24 nsew signal input
flabel metal3 s 26200 24760 27000 24880 0 FreeSans 480 0 0 0 chanx_right_in[29]
port 25 nsew signal input
flabel metal3 s 26200 13744 27000 13864 0 FreeSans 480 0 0 0 chanx_right_in[2]
port 26 nsew signal input
flabel metal3 s 26200 14152 27000 14272 0 FreeSans 480 0 0 0 chanx_right_in[3]
port 27 nsew signal input
flabel metal3 s 26200 14560 27000 14680 0 FreeSans 480 0 0 0 chanx_right_in[4]
port 28 nsew signal input
flabel metal3 s 26200 14968 27000 15088 0 FreeSans 480 0 0 0 chanx_right_in[5]
port 29 nsew signal input
flabel metal3 s 26200 15376 27000 15496 0 FreeSans 480 0 0 0 chanx_right_in[6]
port 30 nsew signal input
flabel metal3 s 26200 15784 27000 15904 0 FreeSans 480 0 0 0 chanx_right_in[7]
port 31 nsew signal input
flabel metal3 s 26200 16192 27000 16312 0 FreeSans 480 0 0 0 chanx_right_in[8]
port 32 nsew signal input
flabel metal3 s 26200 16600 27000 16720 0 FreeSans 480 0 0 0 chanx_right_in[9]
port 33 nsew signal input
flabel metal3 s 26200 688 27000 808 0 FreeSans 480 0 0 0 chanx_right_out[0]
port 34 nsew signal tristate
flabel metal3 s 26200 4768 27000 4888 0 FreeSans 480 0 0 0 chanx_right_out[10]
port 35 nsew signal tristate
flabel metal3 s 26200 5176 27000 5296 0 FreeSans 480 0 0 0 chanx_right_out[11]
port 36 nsew signal tristate
flabel metal3 s 26200 5584 27000 5704 0 FreeSans 480 0 0 0 chanx_right_out[12]
port 37 nsew signal tristate
flabel metal3 s 26200 5992 27000 6112 0 FreeSans 480 0 0 0 chanx_right_out[13]
port 38 nsew signal tristate
flabel metal3 s 26200 6400 27000 6520 0 FreeSans 480 0 0 0 chanx_right_out[14]
port 39 nsew signal tristate
flabel metal3 s 26200 6808 27000 6928 0 FreeSans 480 0 0 0 chanx_right_out[15]
port 40 nsew signal tristate
flabel metal3 s 26200 7216 27000 7336 0 FreeSans 480 0 0 0 chanx_right_out[16]
port 41 nsew signal tristate
flabel metal3 s 26200 7624 27000 7744 0 FreeSans 480 0 0 0 chanx_right_out[17]
port 42 nsew signal tristate
flabel metal3 s 26200 8032 27000 8152 0 FreeSans 480 0 0 0 chanx_right_out[18]
port 43 nsew signal tristate
flabel metal3 s 26200 8440 27000 8560 0 FreeSans 480 0 0 0 chanx_right_out[19]
port 44 nsew signal tristate
flabel metal3 s 26200 1096 27000 1216 0 FreeSans 480 0 0 0 chanx_right_out[1]
port 45 nsew signal tristate
flabel metal3 s 26200 8848 27000 8968 0 FreeSans 480 0 0 0 chanx_right_out[20]
port 46 nsew signal tristate
flabel metal3 s 26200 9256 27000 9376 0 FreeSans 480 0 0 0 chanx_right_out[21]
port 47 nsew signal tristate
flabel metal3 s 26200 9664 27000 9784 0 FreeSans 480 0 0 0 chanx_right_out[22]
port 48 nsew signal tristate
flabel metal3 s 26200 10072 27000 10192 0 FreeSans 480 0 0 0 chanx_right_out[23]
port 49 nsew signal tristate
flabel metal3 s 26200 10480 27000 10600 0 FreeSans 480 0 0 0 chanx_right_out[24]
port 50 nsew signal tristate
flabel metal3 s 26200 10888 27000 11008 0 FreeSans 480 0 0 0 chanx_right_out[25]
port 51 nsew signal tristate
flabel metal3 s 26200 11296 27000 11416 0 FreeSans 480 0 0 0 chanx_right_out[26]
port 52 nsew signal tristate
flabel metal3 s 26200 11704 27000 11824 0 FreeSans 480 0 0 0 chanx_right_out[27]
port 53 nsew signal tristate
flabel metal3 s 26200 12112 27000 12232 0 FreeSans 480 0 0 0 chanx_right_out[28]
port 54 nsew signal tristate
flabel metal3 s 26200 12520 27000 12640 0 FreeSans 480 0 0 0 chanx_right_out[29]
port 55 nsew signal tristate
flabel metal3 s 26200 1504 27000 1624 0 FreeSans 480 0 0 0 chanx_right_out[2]
port 56 nsew signal tristate
flabel metal3 s 26200 1912 27000 2032 0 FreeSans 480 0 0 0 chanx_right_out[3]
port 57 nsew signal tristate
flabel metal3 s 26200 2320 27000 2440 0 FreeSans 480 0 0 0 chanx_right_out[4]
port 58 nsew signal tristate
flabel metal3 s 26200 2728 27000 2848 0 FreeSans 480 0 0 0 chanx_right_out[5]
port 59 nsew signal tristate
flabel metal3 s 26200 3136 27000 3256 0 FreeSans 480 0 0 0 chanx_right_out[6]
port 60 nsew signal tristate
flabel metal3 s 26200 3544 27000 3664 0 FreeSans 480 0 0 0 chanx_right_out[7]
port 61 nsew signal tristate
flabel metal3 s 26200 3952 27000 4072 0 FreeSans 480 0 0 0 chanx_right_out[8]
port 62 nsew signal tristate
flabel metal3 s 26200 4360 27000 4480 0 FreeSans 480 0 0 0 chanx_right_out[9]
port 63 nsew signal tristate
flabel metal2 s 12714 26200 12770 27000 0 FreeSans 224 90 0 0 chany_top_in[0]
port 64 nsew signal input
flabel metal2 s 16394 26200 16450 27000 0 FreeSans 224 90 0 0 chany_top_in[10]
port 65 nsew signal input
flabel metal2 s 16762 26200 16818 27000 0 FreeSans 224 90 0 0 chany_top_in[11]
port 66 nsew signal input
flabel metal2 s 17130 26200 17186 27000 0 FreeSans 224 90 0 0 chany_top_in[12]
port 67 nsew signal input
flabel metal2 s 17498 26200 17554 27000 0 FreeSans 224 90 0 0 chany_top_in[13]
port 68 nsew signal input
flabel metal2 s 17866 26200 17922 27000 0 FreeSans 224 90 0 0 chany_top_in[14]
port 69 nsew signal input
flabel metal2 s 18234 26200 18290 27000 0 FreeSans 224 90 0 0 chany_top_in[15]
port 70 nsew signal input
flabel metal2 s 18602 26200 18658 27000 0 FreeSans 224 90 0 0 chany_top_in[16]
port 71 nsew signal input
flabel metal2 s 18970 26200 19026 27000 0 FreeSans 224 90 0 0 chany_top_in[17]
port 72 nsew signal input
flabel metal2 s 19338 26200 19394 27000 0 FreeSans 224 90 0 0 chany_top_in[18]
port 73 nsew signal input
flabel metal2 s 19706 26200 19762 27000 0 FreeSans 224 90 0 0 chany_top_in[19]
port 74 nsew signal input
flabel metal2 s 13082 26200 13138 27000 0 FreeSans 224 90 0 0 chany_top_in[1]
port 75 nsew signal input
flabel metal2 s 20074 26200 20130 27000 0 FreeSans 224 90 0 0 chany_top_in[20]
port 76 nsew signal input
flabel metal2 s 20442 26200 20498 27000 0 FreeSans 224 90 0 0 chany_top_in[21]
port 77 nsew signal input
flabel metal2 s 20810 26200 20866 27000 0 FreeSans 224 90 0 0 chany_top_in[22]
port 78 nsew signal input
flabel metal2 s 21178 26200 21234 27000 0 FreeSans 224 90 0 0 chany_top_in[23]
port 79 nsew signal input
flabel metal2 s 21546 26200 21602 27000 0 FreeSans 224 90 0 0 chany_top_in[24]
port 80 nsew signal input
flabel metal2 s 21914 26200 21970 27000 0 FreeSans 224 90 0 0 chany_top_in[25]
port 81 nsew signal input
flabel metal2 s 22282 26200 22338 27000 0 FreeSans 224 90 0 0 chany_top_in[26]
port 82 nsew signal input
flabel metal2 s 22650 26200 22706 27000 0 FreeSans 224 90 0 0 chany_top_in[27]
port 83 nsew signal input
flabel metal2 s 23018 26200 23074 27000 0 FreeSans 224 90 0 0 chany_top_in[28]
port 84 nsew signal input
flabel metal2 s 23386 26200 23442 27000 0 FreeSans 224 90 0 0 chany_top_in[29]
port 85 nsew signal input
flabel metal2 s 13450 26200 13506 27000 0 FreeSans 224 90 0 0 chany_top_in[2]
port 86 nsew signal input
flabel metal2 s 13818 26200 13874 27000 0 FreeSans 224 90 0 0 chany_top_in[3]
port 87 nsew signal input
flabel metal2 s 14186 26200 14242 27000 0 FreeSans 224 90 0 0 chany_top_in[4]
port 88 nsew signal input
flabel metal2 s 14554 26200 14610 27000 0 FreeSans 224 90 0 0 chany_top_in[5]
port 89 nsew signal input
flabel metal2 s 14922 26200 14978 27000 0 FreeSans 224 90 0 0 chany_top_in[6]
port 90 nsew signal input
flabel metal2 s 15290 26200 15346 27000 0 FreeSans 224 90 0 0 chany_top_in[7]
port 91 nsew signal input
flabel metal2 s 15658 26200 15714 27000 0 FreeSans 224 90 0 0 chany_top_in[8]
port 92 nsew signal input
flabel metal2 s 16026 26200 16082 27000 0 FreeSans 224 90 0 0 chany_top_in[9]
port 93 nsew signal input
flabel metal2 s 1674 26200 1730 27000 0 FreeSans 224 90 0 0 chany_top_out[0]
port 94 nsew signal tristate
flabel metal2 s 5354 26200 5410 27000 0 FreeSans 224 90 0 0 chany_top_out[10]
port 95 nsew signal tristate
flabel metal2 s 5722 26200 5778 27000 0 FreeSans 224 90 0 0 chany_top_out[11]
port 96 nsew signal tristate
flabel metal2 s 6090 26200 6146 27000 0 FreeSans 224 90 0 0 chany_top_out[12]
port 97 nsew signal tristate
flabel metal2 s 6458 26200 6514 27000 0 FreeSans 224 90 0 0 chany_top_out[13]
port 98 nsew signal tristate
flabel metal2 s 6826 26200 6882 27000 0 FreeSans 224 90 0 0 chany_top_out[14]
port 99 nsew signal tristate
flabel metal2 s 7194 26200 7250 27000 0 FreeSans 224 90 0 0 chany_top_out[15]
port 100 nsew signal tristate
flabel metal2 s 7562 26200 7618 27000 0 FreeSans 224 90 0 0 chany_top_out[16]
port 101 nsew signal tristate
flabel metal2 s 7930 26200 7986 27000 0 FreeSans 224 90 0 0 chany_top_out[17]
port 102 nsew signal tristate
flabel metal2 s 8298 26200 8354 27000 0 FreeSans 224 90 0 0 chany_top_out[18]
port 103 nsew signal tristate
flabel metal2 s 8666 26200 8722 27000 0 FreeSans 224 90 0 0 chany_top_out[19]
port 104 nsew signal tristate
flabel metal2 s 2042 26200 2098 27000 0 FreeSans 224 90 0 0 chany_top_out[1]
port 105 nsew signal tristate
flabel metal2 s 9034 26200 9090 27000 0 FreeSans 224 90 0 0 chany_top_out[20]
port 106 nsew signal tristate
flabel metal2 s 9402 26200 9458 27000 0 FreeSans 224 90 0 0 chany_top_out[21]
port 107 nsew signal tristate
flabel metal2 s 9770 26200 9826 27000 0 FreeSans 224 90 0 0 chany_top_out[22]
port 108 nsew signal tristate
flabel metal2 s 10138 26200 10194 27000 0 FreeSans 224 90 0 0 chany_top_out[23]
port 109 nsew signal tristate
flabel metal2 s 10506 26200 10562 27000 0 FreeSans 224 90 0 0 chany_top_out[24]
port 110 nsew signal tristate
flabel metal2 s 10874 26200 10930 27000 0 FreeSans 224 90 0 0 chany_top_out[25]
port 111 nsew signal tristate
flabel metal2 s 11242 26200 11298 27000 0 FreeSans 224 90 0 0 chany_top_out[26]
port 112 nsew signal tristate
flabel metal2 s 11610 26200 11666 27000 0 FreeSans 224 90 0 0 chany_top_out[27]
port 113 nsew signal tristate
flabel metal2 s 11978 26200 12034 27000 0 FreeSans 224 90 0 0 chany_top_out[28]
port 114 nsew signal tristate
flabel metal2 s 12346 26200 12402 27000 0 FreeSans 224 90 0 0 chany_top_out[29]
port 115 nsew signal tristate
flabel metal2 s 2410 26200 2466 27000 0 FreeSans 224 90 0 0 chany_top_out[2]
port 116 nsew signal tristate
flabel metal2 s 2778 26200 2834 27000 0 FreeSans 224 90 0 0 chany_top_out[3]
port 117 nsew signal tristate
flabel metal2 s 3146 26200 3202 27000 0 FreeSans 224 90 0 0 chany_top_out[4]
port 118 nsew signal tristate
flabel metal2 s 3514 26200 3570 27000 0 FreeSans 224 90 0 0 chany_top_out[5]
port 119 nsew signal tristate
flabel metal2 s 3882 26200 3938 27000 0 FreeSans 224 90 0 0 chany_top_out[6]
port 120 nsew signal tristate
flabel metal2 s 4250 26200 4306 27000 0 FreeSans 224 90 0 0 chany_top_out[7]
port 121 nsew signal tristate
flabel metal2 s 4618 26200 4674 27000 0 FreeSans 224 90 0 0 chany_top_out[8]
port 122 nsew signal tristate
flabel metal2 s 4986 26200 5042 27000 0 FreeSans 224 90 0 0 chany_top_out[9]
port 123 nsew signal tristate
flabel metal2 s 20166 0 20222 800 0 FreeSans 224 90 0 0 prog_clk
port 124 nsew signal input
flabel metal2 s 24490 26200 24546 27000 0 FreeSans 224 90 0 0 prog_reset
port 125 nsew signal input
flabel metal2 s 24858 26200 24914 27000 0 FreeSans 224 90 0 0 reset
port 126 nsew signal input
flabel metal3 s 26200 25168 27000 25288 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
port 127 nsew signal input
flabel metal3 s 26200 25576 27000 25696 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
port 128 nsew signal input
flabel metal3 s 26200 25984 27000 26104 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
port 129 nsew signal input
flabel metal3 s 26200 26392 27000 26512 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
port 130 nsew signal input
flabel metal2 s 25226 26200 25282 27000 0 FreeSans 224 90 0 0 test_enable
port 131 nsew signal input
flabel metal3 s 0 22584 800 22704 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
port 132 nsew signal input
flabel metal3 s 0 23672 800 23792 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
port 133 nsew signal input
flabel metal3 s 0 24760 800 24880 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
port 134 nsew signal input
flabel metal3 s 0 25848 800 25968 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
port 135 nsew signal input
rlabel metal1 13478 23936 13478 23936 0 VGND
rlabel metal1 13478 24480 13478 24480 0 VPWR
rlabel metal1 6670 2278 6670 2278 0 ccff_head
rlabel metal3 24894 340 24894 340 0 ccff_tail
rlabel metal2 22126 8789 22126 8789 0 chanx_right_in[0]
rlabel metal1 21666 7378 21666 7378 0 chanx_right_in[10]
rlabel metal2 21114 17612 21114 17612 0 chanx_right_in[11]
rlabel metal1 13938 15674 13938 15674 0 chanx_right_in[12]
rlabel metal1 15594 18904 15594 18904 0 chanx_right_in[13]
rlabel metal2 17158 17833 17158 17833 0 chanx_right_in[14]
rlabel via2 3910 18683 3910 18683 0 chanx_right_in[15]
rlabel metal1 13294 13872 13294 13872 0 chanx_right_in[16]
rlabel metal2 14122 14586 14122 14586 0 chanx_right_in[17]
rlabel metal2 15870 15640 15870 15640 0 chanx_right_in[18]
rlabel metal2 15134 19669 15134 19669 0 chanx_right_in[19]
rlabel metal1 17802 11526 17802 11526 0 chanx_right_in[1]
rlabel metal1 21298 12750 21298 12750 0 chanx_right_in[20]
rlabel metal2 21666 13860 21666 13860 0 chanx_right_in[21]
rlabel metal2 18676 12852 18676 12852 0 chanx_right_in[22]
rlabel metal2 21436 12852 21436 12852 0 chanx_right_in[23]
rlabel metal3 18423 13260 18423 13260 0 chanx_right_in[24]
rlabel metal3 16537 13668 16537 13668 0 chanx_right_in[25]
rlabel metal2 13570 14161 13570 14161 0 chanx_right_in[26]
rlabel via2 12006 13923 12006 13923 0 chanx_right_in[27]
rlabel metal2 17710 24344 17710 24344 0 chanx_right_in[28]
rlabel metal2 18446 23698 18446 23698 0 chanx_right_in[29]
rlabel metal2 22034 13175 22034 13175 0 chanx_right_in[2]
rlabel metal1 22310 5678 22310 5678 0 chanx_right_in[3]
rlabel metal1 19136 13294 19136 13294 0 chanx_right_in[4]
rlabel metal2 17204 13668 17204 13668 0 chanx_right_in[5]
rlabel metal3 19734 13396 19734 13396 0 chanx_right_in[6]
rlabel metal1 25024 11322 25024 11322 0 chanx_right_in[7]
rlabel metal1 24702 15674 24702 15674 0 chanx_right_in[8]
rlabel metal1 19642 13226 19642 13226 0 chanx_right_in[9]
rlabel metal2 25070 1853 25070 1853 0 chanx_right_out[0]
rlabel metal1 24104 5270 24104 5270 0 chanx_right_out[10]
rlabel metal2 24794 4641 24794 4641 0 chanx_right_out[11]
rlabel metal3 25676 5644 25676 5644 0 chanx_right_out[12]
rlabel metal1 24104 6358 24104 6358 0 chanx_right_out[13]
rlabel metal2 24702 5797 24702 5797 0 chanx_right_out[14]
rlabel metal1 24380 6834 24380 6834 0 chanx_right_out[15]
rlabel metal1 24104 7446 24104 7446 0 chanx_right_out[16]
rlabel metal3 25584 7684 25584 7684 0 chanx_right_out[17]
rlabel metal1 24426 7922 24426 7922 0 chanx_right_out[18]
rlabel metal1 24104 8534 24104 8534 0 chanx_right_out[19]
rlabel metal3 24250 1156 24250 1156 0 chanx_right_out[1]
rlabel metal2 24702 8109 24702 8109 0 chanx_right_out[20]
rlabel metal1 24380 9010 24380 9010 0 chanx_right_out[21]
rlabel metal2 23322 9673 23322 9673 0 chanx_right_out[22]
rlabel metal2 24610 9265 24610 9265 0 chanx_right_out[23]
rlabel metal1 24104 10710 24104 10710 0 chanx_right_out[24]
rlabel metal2 24794 10217 24794 10217 0 chanx_right_out[25]
rlabel metal1 24380 11186 24380 11186 0 chanx_right_out[26]
rlabel metal1 24104 11798 24104 11798 0 chanx_right_out[27]
rlabel metal2 24702 11373 24702 11373 0 chanx_right_out[28]
rlabel metal3 25768 12580 25768 12580 0 chanx_right_out[29]
rlabel metal2 22126 2805 22126 2805 0 chanx_right_out[2]
rlabel metal1 20792 2618 20792 2618 0 chanx_right_out[3]
rlabel metal3 25676 2380 25676 2380 0 chanx_right_out[4]
rlabel metal1 24104 3094 24104 3094 0 chanx_right_out[5]
rlabel metal3 25676 3196 25676 3196 0 chanx_right_out[6]
rlabel metal1 23322 4012 23322 4012 0 chanx_right_out[7]
rlabel metal2 25162 3553 25162 3553 0 chanx_right_out[8]
rlabel metal3 25676 4420 25676 4420 0 chanx_right_out[9]
rlabel metal3 12604 22304 12604 22304 0 chany_top_in[0]
rlabel metal2 12466 23375 12466 23375 0 chany_top_in[10]
rlabel metal2 16698 20366 16698 20366 0 chany_top_in[11]
rlabel metal1 18860 17646 18860 17646 0 chany_top_in[12]
rlabel metal2 17526 25493 17526 25493 0 chany_top_in[13]
rlabel metal1 16698 16490 16698 16490 0 chany_top_in[14]
rlabel metal1 15502 14994 15502 14994 0 chany_top_in[15]
rlabel metal3 15548 23256 15548 23256 0 chany_top_in[16]
rlabel metal2 18998 26173 18998 26173 0 chany_top_in[17]
rlabel metal3 17388 22848 17388 22848 0 chany_top_in[18]
rlabel metal2 19734 25442 19734 25442 0 chany_top_in[19]
rlabel metal3 12995 22780 12995 22780 0 chany_top_in[1]
rlabel metal2 19826 25024 19826 25024 0 chany_top_in[20]
rlabel metal2 13386 19312 13386 19312 0 chany_top_in[21]
rlabel metal2 20838 25561 20838 25561 0 chany_top_in[22]
rlabel metal3 13892 16796 13892 16796 0 chany_top_in[23]
rlabel metal2 21429 26316 21429 26316 0 chany_top_in[24]
rlabel via1 9338 16762 9338 16762 0 chany_top_in[25]
rlabel metal1 1932 18734 1932 18734 0 chany_top_in[26]
rlabel metal1 10166 15470 10166 15470 0 chany_top_in[27]
rlabel metal3 21459 20740 21459 20740 0 chany_top_in[28]
rlabel metal3 16905 14076 16905 14076 0 chany_top_in[29]
rlabel metal2 13478 24218 13478 24218 0 chany_top_in[2]
rlabel metal1 12742 22406 12742 22406 0 chany_top_in[3]
rlabel metal1 12650 23086 12650 23086 0 chany_top_in[4]
rlabel metal2 14582 24932 14582 24932 0 chany_top_in[5]
rlabel metal2 6762 23732 6762 23732 0 chany_top_in[6]
rlabel metal1 20470 20230 20470 20230 0 chany_top_in[7]
rlabel metal2 14214 18496 14214 18496 0 chany_top_in[8]
rlabel metal2 20194 21862 20194 21862 0 chany_top_in[9]
rlabel metal1 2070 19278 2070 19278 0 chany_top_out[0]
rlabel metal1 4692 23766 4692 23766 0 chany_top_out[10]
rlabel metal2 5750 24490 5750 24490 0 chany_top_out[11]
rlabel metal2 6118 24184 6118 24184 0 chany_top_out[12]
rlabel metal1 4876 24242 4876 24242 0 chany_top_out[13]
rlabel metal1 7176 20978 7176 20978 0 chany_top_out[14]
rlabel metal1 7498 21454 7498 21454 0 chany_top_out[15]
rlabel metal1 6624 23766 6624 23766 0 chany_top_out[16]
rlabel metal1 7130 23154 7130 23154 0 chany_top_out[17]
rlabel metal2 8326 24184 8326 24184 0 chany_top_out[18]
rlabel metal2 5842 24446 5842 24446 0 chany_top_out[19]
rlabel metal1 2300 19890 2300 19890 0 chany_top_out[1]
rlabel metal2 8786 24497 8786 24497 0 chany_top_out[20]
rlabel metal1 8326 23188 8326 23188 0 chany_top_out[21]
rlabel metal1 8970 24242 8970 24242 0 chany_top_out[22]
rlabel metal1 9660 23766 9660 23766 0 chany_top_out[23]
rlabel metal2 10534 24728 10534 24728 0 chany_top_out[24]
rlabel metal2 10902 25034 10902 25034 0 chany_top_out[25]
rlabel metal2 10994 24531 10994 24531 0 chany_top_out[26]
rlabel metal1 11914 23154 11914 23154 0 chany_top_out[27]
rlabel metal2 12006 24966 12006 24966 0 chany_top_out[28]
rlabel metal1 12834 24276 12834 24276 0 chany_top_out[29]
rlabel metal2 2714 24888 2714 24888 0 chany_top_out[2]
rlabel metal1 3220 26418 3220 26418 0 chany_top_out[3]
rlabel metal2 3029 26316 3029 26316 0 chany_top_out[4]
rlabel metal2 3542 23878 3542 23878 0 chany_top_out[5]
rlabel metal1 4324 20978 4324 20978 0 chany_top_out[6]
rlabel metal1 4140 22678 4140 22678 0 chany_top_out[7]
rlabel metal1 3956 23154 3956 23154 0 chany_top_out[8]
rlabel metal2 5067 26316 5067 26316 0 chany_top_out[9]
rlabel metal1 21758 18326 21758 18326 0 clknet_0_prog_clk
rlabel metal1 10488 13158 10488 13158 0 clknet_3_0__leaf_prog_clk
rlabel metal1 15042 15538 15042 15538 0 clknet_3_1__leaf_prog_clk
rlabel metal2 9062 20978 9062 20978 0 clknet_3_2__leaf_prog_clk
rlabel metal1 14076 22066 14076 22066 0 clknet_3_3__leaf_prog_clk
rlabel metal1 19458 14042 19458 14042 0 clknet_3_4__leaf_prog_clk
rlabel metal1 19596 13294 19596 13294 0 clknet_3_5__leaf_prog_clk
rlabel metal1 20378 18700 20378 18700 0 clknet_3_6__leaf_prog_clk
rlabel metal1 21413 17714 21413 17714 0 clknet_3_7__leaf_prog_clk
rlabel metal2 6854 4726 6854 4726 0 net1
rlabel metal4 16652 15912 16652 15912 0 net10
rlabel metal1 24196 3026 24196 3026 0 net100
rlabel metal2 22678 5745 22678 5745 0 net101
rlabel metal2 3818 20451 3818 20451 0 net102
rlabel via2 19458 22491 19458 22491 0 net103
rlabel metal3 12834 21284 12834 21284 0 net104
rlabel metal1 5980 17850 5980 17850 0 net105
rlabel metal1 3082 24174 3082 24174 0 net106
rlabel metal1 7452 17850 7452 17850 0 net107
rlabel metal1 7636 17306 7636 17306 0 net108
rlabel metal1 12765 22746 12765 22746 0 net109
rlabel metal2 20470 23273 20470 23273 0 net11
rlabel via3 15203 20876 15203 20876 0 net110
rlabel metal3 12604 21488 12604 21488 0 net111
rlabel metal2 19090 24055 19090 24055 0 net112
rlabel metal1 2254 19788 2254 19788 0 net113
rlabel metal1 3266 18836 3266 18836 0 net114
rlabel metal1 5888 18938 5888 18938 0 net115
rlabel metal1 3128 20570 3128 20570 0 net116
rlabel metal1 4876 19346 4876 19346 0 net117
rlabel metal1 7498 18802 7498 18802 0 net118
rlabel metal1 5382 19890 5382 19890 0 net119
rlabel metal1 13386 17816 13386 17816 0 net12
rlabel metal1 7452 19890 7452 19890 0 net120
rlabel metal1 11730 23018 11730 23018 0 net121
rlabel metal2 9476 19924 9476 19924 0 net122
rlabel metal1 11684 19686 11684 19686 0 net123
rlabel metal1 2254 20842 2254 20842 0 net124
rlabel metal2 15962 20281 15962 20281 0 net125
rlabel metal1 2254 21930 2254 21930 0 net126
rlabel metal1 2990 21556 2990 21556 0 net127
rlabel metal1 5796 18394 5796 18394 0 net128
rlabel metal1 4094 18122 4094 18122 0 net129
rlabel metal1 14444 20910 14444 20910 0 net13
rlabel metal2 2254 22916 2254 22916 0 net130
rlabel metal2 16054 22253 16054 22253 0 net131
rlabel metal1 20792 15402 20792 15402 0 net132
rlabel metal1 19274 14314 19274 14314 0 net133
rlabel metal1 3818 18394 3818 18394 0 net134
rlabel metal1 17710 12274 17710 12274 0 net135
rlabel metal1 18998 12818 18998 12818 0 net136
rlabel metal1 21390 12138 21390 12138 0 net137
rlabel metal1 23966 9962 23966 9962 0 net138
rlabel metal1 18538 16422 18538 16422 0 net139
rlabel via3 15893 20740 15893 20740 0 net14
rlabel metal1 14720 14586 14720 14586 0 net140
rlabel metal2 20562 18530 20562 18530 0 net141
rlabel metal1 14260 19822 14260 19822 0 net142
rlabel metal2 10074 21760 10074 21760 0 net143
rlabel metal1 8418 22746 8418 22746 0 net144
rlabel metal2 7774 20740 7774 20740 0 net145
rlabel metal1 9614 19754 9614 19754 0 net146
rlabel metal1 20562 17238 20562 17238 0 net147
rlabel metal1 9384 18734 9384 18734 0 net148
rlabel metal2 12466 20672 12466 20672 0 net149
rlabel metal1 17112 21930 17112 21930 0 net15
rlabel metal1 12144 18394 12144 18394 0 net150
rlabel metal1 11040 16558 11040 16558 0 net151
rlabel via2 15318 15147 15318 15147 0 net152
rlabel metal1 10488 16218 10488 16218 0 net153
rlabel metal1 13478 15470 13478 15470 0 net154
rlabel metal2 13938 15606 13938 15606 0 net155
rlabel metal1 14030 17714 14030 17714 0 net156
rlabel metal2 5198 22848 5198 22848 0 net157
rlabel metal2 19366 23936 19366 23936 0 net158
rlabel metal2 20838 19924 20838 19924 0 net159
rlabel metal3 17779 19788 17779 19788 0 net16
rlabel metal1 20562 14280 20562 14280 0 net160
rlabel metal2 18906 13940 18906 13940 0 net161
rlabel metal2 22034 8976 22034 8976 0 net162
rlabel metal1 23782 10098 23782 10098 0 net163
rlabel metal1 20102 7956 20102 7956 0 net164
rlabel via2 2254 18309 2254 18309 0 net165
rlabel metal1 25070 12342 25070 12342 0 net166
rlabel metal1 24012 14926 24012 14926 0 net167
rlabel metal1 20194 24140 20194 24140 0 net168
rlabel metal1 11829 8874 11829 8874 0 net169
rlabel via3 17549 13940 17549 13940 0 net17
rlabel metal1 16008 17714 16008 17714 0 net170
rlabel metal1 7268 2618 7268 2618 0 net171
rlabel metal1 9844 8874 9844 8874 0 net172
rlabel metal3 18883 12444 18883 12444 0 net18
rlabel metal1 15640 23630 15640 23630 0 net19
rlabel metal3 16353 19380 16353 19380 0 net2
rlabel metal1 12512 14042 12512 14042 0 net20
rlabel metal1 25576 11254 25576 11254 0 net21
rlabel metal1 16422 14824 16422 14824 0 net22
rlabel metal1 12834 22474 12834 22474 0 net23
rlabel metal3 15985 19380 15985 19380 0 net24
rlabel metal1 18078 17646 18078 17646 0 net25
rlabel metal1 18906 13498 18906 13498 0 net26
rlabel metal1 17112 17170 17112 17170 0 net27
rlabel metal1 18262 9350 18262 9350 0 net28
rlabel metal2 24610 11475 24610 11475 0 net29
rlabel metal2 13570 21879 13570 21879 0 net3
rlabel metal2 16008 20434 16008 20434 0 net30
rlabel metal1 16284 14042 16284 14042 0 net31
rlabel metal2 17526 20961 17526 20961 0 net32
rlabel metal3 17020 14484 17020 14484 0 net33
rlabel metal1 20654 14824 20654 14824 0 net34
rlabel metal1 18630 17544 18630 17544 0 net35
rlabel metal2 19734 17731 19734 17731 0 net36
rlabel metal2 16514 16150 16514 16150 0 net37
rlabel metal2 21942 18853 21942 18853 0 net38
rlabel metal1 21022 18326 21022 18326 0 net39
rlabel metal2 8418 17408 8418 17408 0 net4
rlabel metal2 6762 15895 6762 15895 0 net40
rlabel metal2 7682 17629 7682 17629 0 net41
rlabel via2 7038 18139 7038 18139 0 net42
rlabel metal1 5497 12410 5497 12410 0 net43
rlabel metal2 6854 16813 6854 16813 0 net44
rlabel metal2 8142 18785 8142 18785 0 net45
rlabel metal2 21942 17901 21942 17901 0 net46
rlabel metal1 22908 20434 22908 20434 0 net47
rlabel metal3 18860 21148 18860 21148 0 net48
rlabel metal1 25622 11322 25622 11322 0 net49
rlabel metal1 13156 14586 13156 14586 0 net5
rlabel metal2 1978 21998 1978 21998 0 net50
rlabel metal2 17342 24276 17342 24276 0 net51
rlabel metal2 19458 10625 19458 10625 0 net52
rlabel via2 1794 24157 1794 24157 0 net53
rlabel metal1 19596 11118 19596 11118 0 net54
rlabel metal2 19458 14399 19458 14399 0 net55
rlabel metal1 25714 14586 25714 14586 0 net56
rlabel metal1 20654 16014 20654 16014 0 net57
rlabel metal1 20010 17646 20010 17646 0 net58
rlabel metal1 18998 18598 18998 18598 0 net59
rlabel metal2 14674 18088 14674 18088 0 net6
rlabel metal1 18400 18190 18400 18190 0 net60
rlabel metal1 23092 21862 23092 21862 0 net61
rlabel metal2 20286 23358 20286 23358 0 net62
rlabel metal1 17664 21522 17664 21522 0 net63
rlabel metal2 18446 18972 18446 18972 0 net64
rlabel metal3 20700 21488 20700 21488 0 net65
rlabel metal2 20930 17782 20930 17782 0 net66
rlabel metal1 13708 19754 13708 19754 0 net67
rlabel metal1 8464 20978 8464 20978 0 net68
rlabel metal1 15916 20978 15916 20978 0 net69
rlabel metal1 9062 16966 9062 16966 0 net7
rlabel metal2 1794 21216 1794 21216 0 net70
rlabel metal1 20470 2414 20470 2414 0 net71
rlabel metal1 20056 3026 20056 3026 0 net72
rlabel metal1 22402 5202 22402 5202 0 net73
rlabel metal1 24656 4114 24656 4114 0 net74
rlabel metal1 23184 5678 23184 5678 0 net75
rlabel metal1 23552 8806 23552 8806 0 net76
rlabel metal1 23368 5202 23368 5202 0 net77
rlabel metal1 22678 6800 22678 6800 0 net78
rlabel metal1 22310 7344 22310 7344 0 net79
rlabel via2 2622 18853 2622 18853 0 net8
rlabel metal1 23828 6290 23828 6290 0 net80
rlabel metal1 22862 7820 22862 7820 0 net81
rlabel metal1 22126 8432 22126 8432 0 net82
rlabel metal1 20470 3502 20470 3502 0 net83
rlabel metal1 23184 7378 23184 7378 0 net84
rlabel metal1 21436 6630 21436 6630 0 net85
rlabel metal1 22126 9588 22126 9588 0 net86
rlabel metal1 23092 8466 23092 8466 0 net87
rlabel metal1 22126 10676 22126 10676 0 net88
rlabel metal2 23966 10030 23966 10030 0 net89
rlabel metal1 13386 14042 13386 14042 0 net9
rlabel metal1 18078 9452 18078 9452 0 net90
rlabel metal2 22218 10166 22218 10166 0 net91
rlabel metal2 23966 10846 23966 10846 0 net92
rlabel metal1 23966 11696 23966 11696 0 net93
rlabel metal2 20286 4879 20286 4879 0 net94
rlabel metal1 19136 3026 19136 3026 0 net95
rlabel metal1 23736 2414 23736 2414 0 net96
rlabel metal1 22954 3026 22954 3026 0 net97
rlabel metal1 23184 3502 23184 3502 0 net98
rlabel metal1 22770 4114 22770 4114 0 net99
rlabel metal2 18998 15606 18998 15606 0 prog_clk
rlabel metal1 24518 16558 24518 16558 0 prog_reset
rlabel metal2 6578 21325 6578 21325 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal2 20654 24140 20654 24140 0 right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal2 23230 21726 23230 21726 0 right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal1 25622 9146 25622 9146 0 right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal2 15226 16626 15226 16626 0 sb_0__0_.mem_right_track_0.ccff_head
rlabel metal2 19918 19822 19918 19822 0 sb_0__0_.mem_right_track_0.ccff_tail
rlabel metal1 17204 19278 17204 19278 0 sb_0__0_.mem_right_track_0.mem_out\[0\]
rlabel metal2 25254 19516 25254 19516 0 sb_0__0_.mem_right_track_10.ccff_head
rlabel metal2 21390 19550 21390 19550 0 sb_0__0_.mem_right_track_10.ccff_tail
rlabel metal2 25070 18224 25070 18224 0 sb_0__0_.mem_right_track_10.mem_out\[0\]
rlabel metal2 22218 17170 22218 17170 0 sb_0__0_.mem_right_track_12.ccff_tail
rlabel via1 20746 19669 20746 19669 0 sb_0__0_.mem_right_track_12.mem_out\[0\]
rlabel metal2 23966 15572 23966 15572 0 sb_0__0_.mem_right_track_14.ccff_tail
rlabel metal1 22586 17850 22586 17850 0 sb_0__0_.mem_right_track_14.mem_out\[0\]
rlabel metal1 23598 12274 23598 12274 0 sb_0__0_.mem_right_track_16.ccff_tail
rlabel metal1 24564 15130 24564 15130 0 sb_0__0_.mem_right_track_16.mem_out\[0\]
rlabel metal1 23506 12954 23506 12954 0 sb_0__0_.mem_right_track_18.ccff_tail
rlabel metal1 23230 12070 23230 12070 0 sb_0__0_.mem_right_track_18.mem_out\[0\]
rlabel metal1 22908 22066 22908 22066 0 sb_0__0_.mem_right_track_2.ccff_tail
rlabel metal1 20792 21930 20792 21930 0 sb_0__0_.mem_right_track_2.mem_out\[0\]
rlabel metal2 21298 14382 21298 14382 0 sb_0__0_.mem_right_track_28.ccff_tail
rlabel metal1 20010 13192 20010 13192 0 sb_0__0_.mem_right_track_28.mem_out\[0\]
rlabel metal1 21160 16762 21160 16762 0 sb_0__0_.mem_right_track_30.ccff_tail
rlabel metal1 20325 16762 20325 16762 0 sb_0__0_.mem_right_track_30.mem_out\[0\]
rlabel metal2 18906 15980 18906 15980 0 sb_0__0_.mem_right_track_32.ccff_tail
rlabel metal1 20148 17306 20148 17306 0 sb_0__0_.mem_right_track_32.mem_out\[0\]
rlabel metal2 18630 14620 18630 14620 0 sb_0__0_.mem_right_track_34.ccff_tail
rlabel metal1 17158 15096 17158 15096 0 sb_0__0_.mem_right_track_34.mem_out\[0\]
rlabel metal1 25346 18190 25346 18190 0 sb_0__0_.mem_right_track_4.ccff_tail
rlabel metal2 22586 23460 22586 23460 0 sb_0__0_.mem_right_track_4.mem_out\[0\]
rlabel metal1 17296 13158 17296 13158 0 sb_0__0_.mem_right_track_44.ccff_tail
rlabel metal1 18492 14518 18492 14518 0 sb_0__0_.mem_right_track_44.mem_out\[0\]
rlabel metal1 19136 12682 19136 12682 0 sb_0__0_.mem_right_track_46.ccff_tail
rlabel metal1 17158 12920 17158 12920 0 sb_0__0_.mem_right_track_46.mem_out\[0\]
rlabel metal1 20654 12682 20654 12682 0 sb_0__0_.mem_right_track_48.ccff_tail
rlabel metal2 19780 14212 19780 14212 0 sb_0__0_.mem_right_track_48.mem_out\[0\]
rlabel metal1 21436 11594 21436 11594 0 sb_0__0_.mem_right_track_50.mem_out\[0\]
rlabel metal1 24380 22406 24380 22406 0 sb_0__0_.mem_right_track_6.ccff_tail
rlabel metal1 17526 23562 17526 23562 0 sb_0__0_.mem_right_track_6.mem_out\[0\]
rlabel metal1 16422 21454 16422 21454 0 sb_0__0_.mem_right_track_8.mem_out\[0\]
rlabel metal1 15916 18666 15916 18666 0 sb_0__0_.mem_top_track_0.ccff_tail
rlabel metal1 20516 19890 20516 19890 0 sb_0__0_.mem_top_track_0.mem_out\[0\]
rlabel metal1 15088 22746 15088 22746 0 sb_0__0_.mem_top_track_10.ccff_head
rlabel metal1 14490 20230 14490 20230 0 sb_0__0_.mem_top_track_10.ccff_tail
rlabel metal1 15686 21862 15686 21862 0 sb_0__0_.mem_top_track_10.mem_out\[0\]
rlabel metal1 11960 20978 11960 20978 0 sb_0__0_.mem_top_track_12.ccff_tail
rlabel metal1 14536 19482 14536 19482 0 sb_0__0_.mem_top_track_12.mem_out\[0\]
rlabel metal2 12466 22270 12466 22270 0 sb_0__0_.mem_top_track_14.ccff_tail
rlabel metal1 12880 21114 12880 21114 0 sb_0__0_.mem_top_track_14.mem_out\[0\]
rlabel metal2 10534 20672 10534 20672 0 sb_0__0_.mem_top_track_16.ccff_tail
rlabel metal2 11178 21964 11178 21964 0 sb_0__0_.mem_top_track_16.mem_out\[0\]
rlabel metal2 10810 18768 10810 18768 0 sb_0__0_.mem_top_track_18.ccff_tail
rlabel metal2 10810 19754 10810 19754 0 sb_0__0_.mem_top_track_18.mem_out\[0\]
rlabel metal1 19136 20978 19136 20978 0 sb_0__0_.mem_top_track_2.ccff_tail
rlabel metal1 18032 20366 18032 20366 0 sb_0__0_.mem_top_track_2.mem_out\[0\]
rlabel metal2 10074 17340 10074 17340 0 sb_0__0_.mem_top_track_28.ccff_tail
rlabel metal1 15778 18122 15778 18122 0 sb_0__0_.mem_top_track_28.mem_out\[0\]
rlabel metal2 12834 19040 12834 19040 0 sb_0__0_.mem_top_track_30.ccff_tail
rlabel metal2 17940 19482 17940 19482 0 sb_0__0_.mem_top_track_30.mem_out\[0\]
rlabel metal2 12374 17306 12374 17306 0 sb_0__0_.mem_top_track_32.ccff_tail
rlabel metal1 15134 17510 15134 17510 0 sb_0__0_.mem_top_track_32.mem_out\[0\]
rlabel metal2 12282 15028 12282 15028 0 sb_0__0_.mem_top_track_34.ccff_tail
rlabel metal1 13800 16014 13800 16014 0 sb_0__0_.mem_top_track_34.mem_out\[0\]
rlabel metal1 18262 23630 18262 23630 0 sb_0__0_.mem_top_track_4.ccff_tail
rlabel metal1 20976 21046 20976 21046 0 sb_0__0_.mem_top_track_4.mem_out\[0\]
rlabel metal2 11086 15572 11086 15572 0 sb_0__0_.mem_top_track_44.ccff_tail
rlabel metal2 15410 15402 15410 15402 0 sb_0__0_.mem_top_track_44.mem_out\[0\]
rlabel metal1 14398 13226 14398 13226 0 sb_0__0_.mem_top_track_46.ccff_tail
rlabel metal1 13984 13430 13984 13430 0 sb_0__0_.mem_top_track_46.mem_out\[0\]
rlabel metal2 14582 15232 14582 15232 0 sb_0__0_.mem_top_track_48.ccff_tail
rlabel metal1 16192 13498 16192 13498 0 sb_0__0_.mem_top_track_48.mem_out\[0\]
rlabel metal1 16146 14518 16146 14518 0 sb_0__0_.mem_top_track_50.mem_out\[0\]
rlabel metal1 16560 23154 16560 23154 0 sb_0__0_.mem_top_track_6.ccff_tail
rlabel metal1 17894 22542 17894 22542 0 sb_0__0_.mem_top_track_6.mem_out\[0\]
rlabel metal1 17250 23290 17250 23290 0 sb_0__0_.mem_top_track_8.mem_out\[0\]
rlabel metal1 21574 7888 21574 7888 0 sb_0__0_.mux_right_track_0.out
rlabel metal1 19412 19346 19412 19346 0 sb_0__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20056 19482 20056 19482 0 sb_0__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19320 19482 19320 19482 0 sb_0__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 22034 6664 22034 6664 0 sb_0__0_.mux_right_track_10.out
rlabel metal1 24196 21862 24196 21862 0 sb_0__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal3 22287 6868 22287 6868 0 sb_0__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20240 9554 20240 9554 0 sb_0__0_.mux_right_track_12.out
rlabel metal1 22402 16218 22402 16218 0 sb_0__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22264 11118 22264 11118 0 sb_0__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19688 10098 19688 10098 0 sb_0__0_.mux_right_track_14.out
rlabel metal1 23368 16014 23368 16014 0 sb_0__0_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21482 10608 21482 10608 0 sb_0__0_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21252 6766 21252 6766 0 sb_0__0_.mux_right_track_16.out
rlabel metal1 23690 14450 23690 14450 0 sb_0__0_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 20608 13362 20608 13362 0 sb_0__0_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20378 7854 20378 7854 0 sb_0__0_.mux_right_track_18.out
rlabel metal1 25208 13294 25208 13294 0 sb_0__0_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 21574 11356 21574 11356 0 sb_0__0_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 13892 12274 13892 12274 0 sb_0__0_.mux_right_track_2.out
rlabel metal1 24840 24106 24840 24106 0 sb_0__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal3 18492 19448 18492 19448 0 sb_0__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 20838 8602 20838 8602 0 sb_0__0_.mux_right_track_28.out
rlabel metal1 20838 14042 20838 14042 0 sb_0__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20792 10642 20792 10642 0 sb_0__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19458 9044 19458 9044 0 sb_0__0_.mux_right_track_30.out
rlabel metal1 21252 15334 21252 15334 0 sb_0__0_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20976 15606 20976 15606 0 sb_0__0_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21988 8058 21988 8058 0 sb_0__0_.mux_right_track_32.out
rlabel metal2 20010 18428 20010 18428 0 sb_0__0_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal3 20861 14484 20861 14484 0 sb_0__0_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24150 7854 24150 7854 0 sb_0__0_.mux_right_track_34.out
rlabel metal2 19918 16218 19918 16218 0 sb_0__0_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19734 14586 19734 14586 0 sb_0__0_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 17250 8466 17250 8466 0 sb_0__0_.mux_right_track_4.out
rlabel metal2 17112 20876 17112 20876 0 sb_0__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 21206 18071 21206 18071 0 sb_0__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 23414 6698 23414 6698 0 sb_0__0_.mux_right_track_44.out
rlabel metal2 17526 16048 17526 16048 0 sb_0__0_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18216 9622 18216 9622 0 sb_0__0_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24656 5678 24656 5678 0 sb_0__0_.mux_right_track_46.out
rlabel metal1 18998 12750 18998 12750 0 sb_0__0_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19458 12614 19458 12614 0 sb_0__0_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24150 4590 24150 4590 0 sb_0__0_.mux_right_track_48.out
rlabel metal1 20148 12954 20148 12954 0 sb_0__0_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 20286 12517 20286 12517 0 sb_0__0_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24702 3502 24702 3502 0 sb_0__0_.mux_right_track_50.out
rlabel metal1 25162 9962 25162 9962 0 sb_0__0_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 21758 7956 21758 7956 0 sb_0__0_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 13386 9554 13386 9554 0 sb_0__0_.mux_right_track_6.out
rlabel metal1 19458 22984 19458 22984 0 sb_0__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 24794 17850 24794 17850 0 sb_0__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 8694 16048 8694 16048 0 sb_0__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 18814 10234 18814 10234 0 sb_0__0_.mux_right_track_8.out
rlabel metal3 17089 20604 17089 20604 0 sb_0__0_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 17618 10353 17618 10353 0 sb_0__0_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 4554 17068 4554 17068 0 sb_0__0_.mux_top_track_0.out
rlabel metal2 14306 19176 14306 19176 0 sb_0__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17020 19482 17020 19482 0 sb_0__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14904 19482 14904 19482 0 sb_0__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 7774 18734 7774 18734 0 sb_0__0_.mux_top_track_10.out
rlabel metal2 17710 21726 17710 21726 0 sb_0__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 8602 20502 8602 20502 0 sb_0__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 3312 17850 3312 17850 0 sb_0__0_.mux_top_track_12.out
rlabel metal1 16652 21114 16652 21114 0 sb_0__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 3450 17170 3450 17170 0 sb_0__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 2438 20366 2438 20366 0 sb_0__0_.mux_top_track_14.out
rlabel metal1 16192 22134 16192 22134 0 sb_0__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 11178 19652 11178 19652 0 sb_0__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 7176 18394 7176 18394 0 sb_0__0_.mux_top_track_16.out
rlabel metal1 10442 21046 10442 21046 0 sb_0__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 8510 19652 8510 19652 0 sb_0__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 3818 18734 3818 18734 0 sb_0__0_.mux_top_track_18.out
rlabel metal1 10902 19958 10902 19958 0 sb_0__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 8832 20026 8832 20026 0 sb_0__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 5198 17748 5198 17748 0 sb_0__0_.mux_top_track_2.out
rlabel metal1 18354 21046 18354 21046 0 sb_0__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17894 20808 17894 20808 0 sb_0__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 4094 20264 4094 20264 0 sb_0__0_.mux_top_track_28.out
rlabel metal1 14904 18394 14904 18394 0 sb_0__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 1794 20468 1794 20468 0 sb_0__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 7222 21318 7222 21318 0 sb_0__0_.mux_top_track_30.out
rlabel metal1 15594 19958 15594 19958 0 sb_0__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 11868 20230 11868 20230 0 sb_0__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 8372 18938 8372 18938 0 sb_0__0_.mux_top_track_32.out
rlabel metal1 15686 18190 15686 18190 0 sb_0__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 11822 18156 11822 18156 0 sb_0__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 6440 17646 6440 17646 0 sb_0__0_.mux_top_track_34.out
rlabel metal2 15042 16864 15042 16864 0 sb_0__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 10810 16218 10810 16218 0 sb_0__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 8372 23086 8372 23086 0 sb_0__0_.mux_top_track_4.out
rlabel metal1 18952 24038 18952 24038 0 sb_0__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 18170 24616 18170 24616 0 sb_0__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 4738 18292 4738 18292 0 sb_0__0_.mux_top_track_44.out
rlabel metal1 13202 16218 13202 16218 0 sb_0__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 9660 15878 9660 15878 0 sb_0__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 6486 18258 6486 18258 0 sb_0__0_.mux_top_track_46.out
rlabel metal1 13202 15572 13202 15572 0 sb_0__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 11178 15504 11178 15504 0 sb_0__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 7590 19482 7590 19482 0 sb_0__0_.mux_top_track_48.out
rlabel metal1 17894 15946 17894 15946 0 sb_0__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13110 15368 13110 15368 0 sb_0__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 5474 18258 5474 18258 0 sb_0__0_.mux_top_track_50.out
rlabel metal1 15318 17850 15318 17850 0 sb_0__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 9706 19159 9706 19159 0 sb_0__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 3956 17306 3956 17306 0 sb_0__0_.mux_top_track_6.out
rlabel metal2 15042 22134 15042 22134 0 sb_0__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17204 23086 17204 23086 0 sb_0__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 4094 17238 4094 17238 0 sb_0__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 5842 19652 5842 19652 0 sb_0__0_.mux_top_track_8.out
rlabel metal2 20470 21607 20470 21607 0 sb_0__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 14122 24276 14122 24276 0 sb_0__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 1472 22610 1472 22610 0 top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal1 1426 23698 1426 23698 0 top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal2 3450 23749 3450 23749 0 top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal1 1932 21590 1932 21590 0 top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
<< properties >>
string FIXED_BBOX 0 0 27000 27000
<< end >>
