magic
tech sky130A
magscale 1 2
timestamp 1656242501
<< viali >>
rect 5549 20553 5583 20587
rect 5917 20553 5951 20587
rect 6561 20553 6595 20587
rect 9321 20553 9355 20587
rect 11253 20553 11287 20587
rect 15945 20553 15979 20587
rect 16865 20553 16899 20587
rect 17601 20553 17635 20587
rect 18613 20553 18647 20587
rect 19441 20553 19475 20587
rect 20821 20553 20855 20587
rect 4813 20485 4847 20519
rect 1685 20417 1719 20451
rect 2697 20417 2731 20451
rect 3801 20417 3835 20451
rect 5181 20417 5215 20451
rect 5733 20417 5767 20451
rect 6101 20417 6135 20451
rect 6377 20417 6411 20451
rect 6929 20417 6963 20451
rect 7205 20417 7239 20451
rect 7481 20417 7515 20451
rect 7941 20417 7975 20451
rect 8033 20417 8067 20451
rect 8493 20417 8527 20451
rect 8585 20417 8619 20451
rect 9045 20417 9079 20451
rect 9505 20417 9539 20451
rect 9781 20417 9815 20451
rect 9873 20417 9907 20451
rect 10517 20417 10551 20451
rect 11069 20417 11103 20451
rect 11713 20417 11747 20451
rect 12725 20417 12759 20451
rect 12817 20417 12851 20451
rect 13737 20417 13771 20451
rect 15025 20417 15059 20451
rect 15393 20417 15427 20451
rect 15761 20417 15795 20451
rect 16129 20417 16163 20451
rect 16681 20417 16715 20451
rect 17049 20417 17083 20451
rect 17417 20417 17451 20451
rect 17785 20417 17819 20451
rect 18153 20417 18187 20451
rect 18797 20417 18831 20451
rect 19257 20417 19291 20451
rect 19625 20417 19659 20451
rect 19993 20417 20027 20451
rect 20361 20417 20395 20451
rect 21005 20417 21039 20451
rect 21097 20417 21131 20451
rect 21465 20417 21499 20451
rect 2421 20349 2455 20383
rect 3341 20349 3375 20383
rect 3617 20349 3651 20383
rect 4077 20349 4111 20383
rect 10241 20349 10275 20383
rect 10425 20349 10459 20383
rect 12449 20349 12483 20383
rect 13093 20349 13127 20383
rect 14657 20349 14691 20383
rect 14933 20349 14967 20383
rect 7757 20281 7791 20315
rect 10885 20281 10919 20315
rect 15209 20281 15243 20315
rect 16313 20281 16347 20315
rect 17233 20281 17267 20315
rect 18337 20281 18371 20315
rect 19809 20281 19843 20315
rect 20545 20281 20579 20315
rect 1501 20213 1535 20247
rect 4905 20213 4939 20247
rect 5365 20213 5399 20247
rect 6837 20213 6871 20247
rect 7113 20213 7147 20247
rect 7389 20213 7423 20247
rect 7665 20213 7699 20247
rect 8217 20213 8251 20247
rect 8309 20213 8343 20247
rect 8769 20213 8803 20247
rect 9229 20213 9263 20247
rect 9597 20213 9631 20247
rect 10057 20213 10091 20247
rect 11529 20213 11563 20247
rect 13921 20213 13955 20247
rect 15577 20213 15611 20247
rect 17969 20213 18003 20247
rect 18981 20213 19015 20247
rect 20177 20213 20211 20247
rect 21281 20213 21315 20247
rect 1869 20009 1903 20043
rect 2237 20009 2271 20043
rect 3065 20009 3099 20043
rect 3617 20009 3651 20043
rect 8401 20009 8435 20043
rect 9689 20009 9723 20043
rect 10609 20009 10643 20043
rect 13645 20009 13679 20043
rect 15117 20009 15151 20043
rect 15853 20009 15887 20043
rect 16865 20009 16899 20043
rect 17417 20009 17451 20043
rect 17785 20009 17819 20043
rect 18429 20009 18463 20043
rect 18889 20009 18923 20043
rect 19901 20009 19935 20043
rect 20269 20009 20303 20043
rect 21005 20009 21039 20043
rect 3433 19941 3467 19975
rect 4169 19941 4203 19975
rect 4813 19941 4847 19975
rect 7389 19941 7423 19975
rect 10517 19941 10551 19975
rect 13921 19941 13955 19975
rect 16589 19941 16623 19975
rect 19441 19941 19475 19975
rect 20729 19941 20763 19975
rect 2789 19873 2823 19907
rect 7481 19873 7515 19907
rect 7849 19873 7883 19907
rect 9045 19873 9079 19907
rect 9965 19873 9999 19907
rect 14657 19873 14691 19907
rect 1685 19805 1719 19839
rect 2053 19805 2087 19839
rect 2421 19805 2455 19839
rect 2605 19805 2639 19839
rect 2881 19805 2915 19839
rect 3249 19805 3283 19839
rect 3985 19805 4019 19839
rect 4261 19805 4295 19839
rect 4629 19805 4663 19839
rect 4997 19805 5031 19839
rect 5733 19805 5767 19839
rect 6009 19805 6043 19839
rect 11989 19805 12023 19839
rect 12449 19805 12483 19839
rect 12725 19805 12759 19839
rect 13461 19805 13495 19839
rect 13737 19805 13771 19839
rect 14933 19805 14967 19839
rect 15485 19805 15519 19839
rect 16037 19805 16071 19839
rect 16313 19805 16347 19839
rect 16405 19805 16439 19839
rect 16681 19805 16715 19839
rect 17141 19805 17175 19839
rect 17233 19805 17267 19839
rect 17509 19805 17543 19839
rect 17969 19805 18003 19839
rect 18061 19805 18095 19839
rect 18613 19805 18647 19839
rect 18705 19805 18739 19839
rect 19257 19805 19291 19839
rect 19533 19805 19567 19839
rect 20085 19805 20119 19839
rect 20453 19805 20487 19839
rect 20545 19805 20579 19839
rect 21189 19805 21223 19839
rect 21281 19805 21315 19839
rect 3801 19737 3835 19771
rect 6254 19737 6288 19771
rect 8033 19737 8067 19771
rect 8493 19737 8527 19771
rect 9321 19737 9355 19771
rect 10149 19737 10183 19771
rect 11744 19737 11778 19771
rect 14473 19737 14507 19771
rect 15577 19737 15611 19771
rect 19073 19737 19107 19771
rect 1501 19669 1535 19703
rect 4445 19669 4479 19703
rect 7941 19669 7975 19703
rect 9229 19669 9263 19703
rect 10057 19669 10091 19703
rect 12081 19669 12115 19703
rect 14105 19669 14139 19703
rect 14565 19669 14599 19703
rect 15301 19669 15335 19703
rect 16129 19669 16163 19703
rect 16957 19669 16991 19703
rect 17693 19669 17727 19703
rect 18245 19669 18279 19703
rect 19717 19669 19751 19703
rect 21465 19669 21499 19703
rect 2145 19465 2179 19499
rect 2421 19465 2455 19499
rect 2881 19465 2915 19499
rect 2973 19465 3007 19499
rect 3249 19465 3283 19499
rect 3709 19465 3743 19499
rect 3985 19465 4019 19499
rect 4353 19465 4387 19499
rect 12633 19465 12667 19499
rect 12817 19465 12851 19499
rect 13369 19465 13403 19499
rect 15025 19465 15059 19499
rect 15393 19465 15427 19499
rect 15669 19465 15703 19499
rect 15945 19465 15979 19499
rect 16497 19465 16531 19499
rect 17509 19465 17543 19499
rect 18153 19465 18187 19499
rect 18613 19465 18647 19499
rect 18889 19465 18923 19499
rect 19349 19465 19383 19499
rect 20269 19465 20303 19499
rect 20729 19465 20763 19499
rect 21097 19465 21131 19499
rect 5825 19397 5859 19431
rect 8309 19397 8343 19431
rect 17785 19397 17819 19431
rect 1685 19329 1719 19363
rect 2053 19329 2087 19363
rect 2329 19329 2363 19363
rect 2605 19329 2639 19363
rect 2697 19329 2731 19363
rect 3157 19329 3191 19363
rect 3433 19329 3467 19363
rect 3525 19329 3559 19363
rect 3801 19329 3835 19363
rect 4997 19329 5031 19363
rect 5733 19329 5767 19363
rect 7582 19329 7616 19363
rect 7849 19329 7883 19363
rect 7941 19333 7975 19367
rect 8401 19329 8435 19363
rect 8668 19329 8702 19363
rect 9965 19329 9999 19363
rect 10232 19329 10266 19363
rect 11989 19329 12023 19363
rect 14482 19329 14516 19363
rect 14841 19329 14875 19363
rect 15209 19329 15243 19363
rect 15485 19329 15519 19363
rect 15761 19329 15795 19363
rect 16313 19329 16347 19363
rect 17141 19329 17175 19363
rect 17877 19329 17911 19363
rect 18337 19329 18371 19363
rect 18429 19329 18463 19363
rect 18705 19329 18739 19363
rect 18981 19329 19015 19363
rect 19717 19329 19751 19363
rect 19993 19329 20027 19363
rect 20453 19329 20487 19363
rect 20545 19329 20579 19363
rect 20913 19329 20947 19363
rect 21281 19329 21315 19363
rect 4721 19261 4755 19295
rect 4905 19261 4939 19295
rect 5641 19261 5675 19295
rect 11621 19261 11655 19295
rect 11713 19261 11747 19295
rect 13001 19261 13035 19295
rect 14749 19261 14783 19295
rect 16865 19261 16899 19295
rect 17049 19261 17083 19295
rect 19165 19261 19199 19295
rect 1869 19193 1903 19227
rect 4537 19193 4571 19227
rect 6469 19193 6503 19227
rect 9781 19193 9815 19227
rect 16037 19193 16071 19227
rect 18061 19193 18095 19227
rect 19533 19193 19567 19227
rect 19901 19193 19935 19227
rect 1501 19125 1535 19159
rect 4169 19125 4203 19159
rect 5365 19125 5399 19159
rect 6193 19125 6227 19159
rect 8125 19125 8159 19159
rect 11345 19125 11379 19159
rect 13277 19125 13311 19159
rect 20177 19125 20211 19159
rect 21465 19125 21499 19159
rect 1961 18921 1995 18955
rect 2973 18921 3007 18955
rect 4905 18921 4939 18955
rect 7205 18921 7239 18955
rect 11529 18921 11563 18955
rect 13553 18921 13587 18955
rect 13645 18921 13679 18955
rect 13921 18921 13955 18955
rect 15485 18921 15519 18955
rect 17509 18921 17543 18955
rect 20545 18921 20579 18955
rect 21097 18921 21131 18955
rect 4077 18853 4111 18887
rect 6377 18853 6411 18887
rect 7389 18853 7423 18887
rect 9781 18853 9815 18887
rect 11253 18853 11287 18887
rect 13277 18853 13311 18887
rect 16589 18853 16623 18887
rect 17601 18853 17635 18887
rect 18521 18853 18555 18887
rect 20821 18853 20855 18887
rect 2421 18785 2455 18819
rect 2513 18785 2547 18819
rect 4353 18785 4387 18819
rect 5825 18785 5859 18819
rect 6653 18785 6687 18819
rect 9229 18785 9263 18819
rect 16957 18785 16991 18819
rect 18153 18785 18187 18819
rect 20085 18785 20119 18819
rect 1685 18717 1719 18751
rect 2145 18717 2179 18751
rect 3341 18717 3375 18751
rect 3801 18717 3835 18751
rect 6745 18717 6779 18751
rect 8769 18717 8803 18751
rect 9873 18717 9907 18751
rect 11805 18717 11839 18751
rect 11897 18717 11931 18751
rect 13369 18717 13403 18751
rect 14105 18717 14139 18751
rect 14372 18717 14406 18751
rect 17969 18717 18003 18751
rect 20361 18717 20395 18751
rect 20637 18717 20671 18751
rect 20913 18717 20947 18751
rect 21281 18717 21315 18751
rect 1777 18649 1811 18683
rect 2605 18649 2639 18683
rect 3065 18649 3099 18683
rect 4445 18649 4479 18683
rect 5549 18649 5583 18683
rect 6009 18649 6043 18683
rect 6837 18649 6871 18683
rect 8524 18649 8558 18683
rect 10129 18649 10163 18683
rect 12142 18649 12176 18683
rect 17049 18649 17083 18683
rect 17141 18649 17175 18683
rect 1501 18581 1535 18615
rect 3525 18581 3559 18615
rect 4537 18581 4571 18615
rect 4997 18581 5031 18615
rect 5181 18581 5215 18615
rect 5917 18581 5951 18615
rect 9321 18581 9355 18615
rect 9413 18581 9447 18615
rect 11437 18581 11471 18615
rect 18061 18581 18095 18615
rect 20269 18581 20303 18615
rect 21465 18581 21499 18615
rect 1961 18377 1995 18411
rect 2421 18377 2455 18411
rect 3433 18377 3467 18411
rect 3893 18377 3927 18411
rect 4077 18377 4111 18411
rect 4537 18377 4571 18411
rect 4905 18377 4939 18411
rect 5549 18377 5583 18411
rect 6101 18377 6135 18411
rect 6561 18377 6595 18411
rect 8033 18377 8067 18411
rect 11161 18377 11195 18411
rect 11989 18377 12023 18411
rect 12449 18377 12483 18411
rect 16129 18377 16163 18411
rect 17601 18377 17635 18411
rect 20729 18377 20763 18411
rect 3065 18309 3099 18343
rect 5733 18309 5767 18343
rect 7674 18309 7708 18343
rect 8585 18309 8619 18343
rect 9496 18309 9530 18343
rect 11069 18309 11103 18343
rect 13461 18309 13495 18343
rect 1685 18241 1719 18275
rect 2145 18241 2179 18275
rect 2237 18241 2271 18275
rect 2513 18241 2547 18275
rect 3617 18241 3651 18275
rect 7941 18241 7975 18275
rect 8309 18241 8343 18275
rect 8953 18241 8987 18275
rect 9137 18241 9171 18275
rect 9229 18241 9263 18275
rect 12081 18241 12115 18275
rect 14677 18241 14711 18275
rect 14933 18241 14967 18275
rect 15761 18241 15795 18275
rect 17417 18241 17451 18275
rect 20545 18241 20579 18275
rect 21005 18241 21039 18275
rect 21281 18241 21315 18275
rect 10701 18173 10735 18207
rect 11805 18173 11839 18207
rect 15485 18173 15519 18207
rect 15669 18173 15703 18207
rect 18429 18173 18463 18207
rect 1777 18105 1811 18139
rect 2881 18105 2915 18139
rect 5917 18105 5951 18139
rect 6469 18105 6503 18139
rect 8677 18105 8711 18139
rect 17785 18105 17819 18139
rect 20821 18105 20855 18139
rect 1501 18037 1535 18071
rect 2697 18037 2731 18071
rect 3341 18037 3375 18071
rect 10609 18037 10643 18071
rect 13553 18037 13587 18071
rect 18061 18037 18095 18071
rect 21465 18037 21499 18071
rect 2145 17833 2179 17867
rect 2421 17833 2455 17867
rect 2605 17833 2639 17867
rect 5641 17833 5675 17867
rect 7481 17833 7515 17867
rect 7757 17833 7791 17867
rect 7941 17833 7975 17867
rect 8769 17833 8803 17867
rect 9045 17833 9079 17867
rect 9413 17833 9447 17867
rect 10425 17833 10459 17867
rect 13645 17833 13679 17867
rect 16589 17833 16623 17867
rect 19993 17833 20027 17867
rect 9229 17765 9263 17799
rect 16497 17765 16531 17799
rect 8217 17697 8251 17731
rect 9689 17697 9723 17731
rect 9873 17697 9907 17731
rect 11345 17697 11379 17731
rect 12173 17697 12207 17731
rect 13093 17697 13127 17731
rect 17141 17697 17175 17731
rect 17969 17697 18003 17731
rect 18797 17697 18831 17731
rect 1685 17629 1719 17663
rect 2053 17629 2087 17663
rect 2329 17629 2363 17663
rect 7113 17629 7147 17663
rect 8309 17629 8343 17663
rect 13829 17629 13863 17663
rect 14289 17629 14323 17663
rect 15761 17629 15795 17663
rect 16313 17629 16347 17663
rect 18613 17629 18647 17663
rect 19809 17629 19843 17663
rect 20913 17629 20947 17663
rect 21281 17629 21315 17663
rect 2789 17561 2823 17595
rect 6846 17561 6880 17595
rect 7297 17561 7331 17595
rect 8401 17561 8435 17595
rect 12449 17561 12483 17595
rect 13277 17561 13311 17595
rect 15494 17561 15528 17595
rect 17785 17561 17819 17595
rect 18705 17561 18739 17595
rect 1501 17493 1535 17527
rect 1869 17493 1903 17527
rect 5733 17493 5767 17527
rect 9965 17493 9999 17527
rect 10333 17493 10367 17527
rect 11069 17493 11103 17527
rect 11437 17493 11471 17527
rect 11529 17493 11563 17527
rect 11897 17493 11931 17527
rect 12357 17493 12391 17527
rect 12817 17493 12851 17527
rect 13185 17493 13219 17527
rect 14381 17493 14415 17527
rect 16957 17493 16991 17527
rect 17049 17493 17083 17527
rect 17417 17493 17451 17527
rect 17877 17493 17911 17527
rect 18245 17493 18279 17527
rect 21097 17493 21131 17527
rect 21465 17493 21499 17527
rect 9689 17289 9723 17323
rect 10057 17289 10091 17323
rect 11345 17289 11379 17323
rect 16681 17289 16715 17323
rect 17969 17289 18003 17323
rect 19901 17289 19935 17323
rect 6920 17221 6954 17255
rect 8484 17221 8518 17255
rect 12081 17221 12115 17255
rect 16129 17221 16163 17255
rect 18337 17221 18371 17255
rect 1685 17153 1719 17187
rect 4169 17153 4203 17187
rect 4261 17153 4295 17187
rect 4813 17153 4847 17187
rect 5080 17153 5114 17187
rect 6561 17153 6595 17187
rect 6653 17153 6687 17187
rect 11989 17153 12023 17187
rect 12449 17153 12483 17187
rect 12716 17153 12750 17187
rect 15045 17153 15079 17187
rect 15301 17153 15335 17187
rect 17049 17153 17083 17187
rect 17877 17153 17911 17187
rect 19717 17153 19751 17187
rect 21281 17153 21315 17187
rect 4445 17085 4479 17119
rect 8217 17085 8251 17119
rect 10149 17085 10183 17119
rect 10333 17085 10367 17119
rect 10609 17085 10643 17119
rect 12173 17085 12207 17119
rect 15853 17085 15887 17119
rect 16037 17085 16071 17119
rect 17141 17085 17175 17119
rect 17325 17085 17359 17119
rect 18061 17085 18095 17119
rect 13829 17017 13863 17051
rect 17509 17017 17543 17051
rect 1501 16949 1535 16983
rect 3801 16949 3835 16983
rect 6193 16949 6227 16983
rect 8033 16949 8067 16983
rect 9597 16949 9631 16983
rect 11621 16949 11655 16983
rect 13921 16949 13955 16983
rect 16497 16949 16531 16983
rect 21465 16949 21499 16983
rect 2237 16745 2271 16779
rect 4537 16745 4571 16779
rect 6377 16745 6411 16779
rect 6561 16745 6595 16779
rect 8217 16745 8251 16779
rect 9321 16745 9355 16779
rect 11805 16745 11839 16779
rect 13829 16745 13863 16779
rect 17233 16745 17267 16779
rect 18245 16745 18279 16779
rect 20637 16745 20671 16779
rect 13277 16677 13311 16711
rect 13553 16677 13587 16711
rect 16129 16677 16163 16711
rect 17417 16677 17451 16711
rect 2697 16609 2731 16643
rect 2881 16609 2915 16643
rect 3985 16609 4019 16643
rect 6653 16609 6687 16643
rect 10793 16609 10827 16643
rect 11897 16609 11931 16643
rect 14105 16609 14139 16643
rect 16589 16609 16623 16643
rect 17969 16609 18003 16643
rect 18705 16609 18739 16643
rect 18889 16609 18923 16643
rect 20085 16609 20119 16643
rect 1685 16541 1719 16575
rect 2053 16541 2087 16575
rect 4077 16541 4111 16575
rect 6909 16541 6943 16575
rect 10526 16541 10560 16575
rect 10885 16541 10919 16575
rect 12153 16541 12187 16575
rect 13369 16541 13403 16575
rect 17877 16541 17911 16575
rect 20453 16541 20487 16575
rect 20729 16541 20763 16575
rect 21189 16541 21223 16575
rect 21281 16541 21315 16575
rect 2973 16473 3007 16507
rect 3433 16473 3467 16507
rect 14350 16473 14384 16507
rect 1501 16405 1535 16439
rect 2421 16405 2455 16439
rect 3341 16405 3375 16439
rect 4169 16405 4203 16439
rect 8033 16405 8067 16439
rect 9413 16405 9447 16439
rect 11069 16405 11103 16439
rect 15485 16405 15519 16439
rect 16405 16405 16439 16439
rect 16773 16405 16807 16439
rect 16865 16405 16899 16439
rect 17785 16405 17819 16439
rect 18613 16405 18647 16439
rect 20269 16405 20303 16439
rect 20913 16405 20947 16439
rect 21005 16405 21039 16439
rect 21465 16405 21499 16439
rect 2145 16201 2179 16235
rect 2421 16201 2455 16235
rect 3617 16201 3651 16235
rect 4813 16201 4847 16235
rect 6193 16201 6227 16235
rect 9873 16201 9907 16235
rect 10977 16201 11011 16235
rect 11345 16201 11379 16235
rect 13737 16201 13771 16235
rect 17141 16201 17175 16235
rect 17601 16201 17635 16235
rect 20545 16201 20579 16235
rect 20821 16201 20855 16235
rect 3157 16133 3191 16167
rect 3801 16133 3835 16167
rect 18061 16133 18095 16167
rect 18521 16133 18555 16167
rect 1685 16065 1719 16099
rect 2053 16065 2087 16099
rect 2329 16065 2363 16099
rect 2605 16065 2639 16099
rect 2789 16065 2823 16099
rect 3249 16065 3283 16099
rect 5181 16065 5215 16099
rect 6377 16065 6411 16099
rect 6633 16065 6667 16099
rect 9505 16065 9539 16099
rect 12081 16065 12115 16099
rect 13829 16065 13863 16099
rect 14085 16065 14119 16099
rect 17969 16065 18003 16099
rect 20361 16065 20395 16099
rect 20637 16065 20671 16099
rect 20913 16065 20947 16099
rect 21281 16065 21315 16099
rect 2973 15997 3007 16031
rect 5273 15997 5307 16031
rect 5365 15997 5399 16031
rect 9229 15997 9263 16031
rect 9413 15997 9447 16031
rect 10701 15997 10735 16031
rect 10885 15997 10919 16031
rect 12173 15997 12207 16031
rect 12265 15997 12299 16031
rect 17233 15997 17267 16031
rect 17325 15997 17359 16031
rect 18153 15997 18187 16031
rect 1869 15929 1903 15963
rect 11713 15929 11747 15963
rect 16405 15929 16439 15963
rect 16773 15929 16807 15963
rect 18613 15929 18647 15963
rect 21097 15929 21131 15963
rect 1501 15861 1535 15895
rect 7757 15861 7791 15895
rect 9965 15861 9999 15895
rect 12541 15861 12575 15895
rect 15209 15861 15243 15895
rect 20177 15861 20211 15895
rect 21465 15861 21499 15895
rect 1961 15657 1995 15691
rect 2237 15657 2271 15691
rect 5457 15657 5491 15691
rect 6285 15657 6319 15691
rect 8953 15657 8987 15691
rect 10057 15657 10091 15691
rect 10885 15657 10919 15691
rect 11805 15657 11839 15691
rect 11989 15657 12023 15691
rect 13829 15657 13863 15691
rect 15577 15657 15611 15691
rect 17049 15657 17083 15691
rect 20269 15657 20303 15691
rect 21005 15657 21039 15691
rect 21465 15657 21499 15691
rect 2513 15589 2547 15623
rect 7849 15589 7883 15623
rect 6101 15521 6135 15555
rect 9505 15521 9539 15555
rect 10609 15521 10643 15555
rect 11345 15521 11379 15555
rect 11437 15521 11471 15555
rect 12633 15521 12667 15555
rect 14105 15521 14139 15555
rect 17601 15521 17635 15555
rect 18429 15521 18463 15555
rect 20729 15521 20763 15555
rect 1685 15453 1719 15487
rect 2145 15453 2179 15487
rect 2421 15453 2455 15487
rect 2697 15453 2731 15487
rect 2881 15453 2915 15487
rect 7665 15453 7699 15487
rect 9321 15453 9355 15487
rect 12357 15453 12391 15487
rect 12449 15453 12483 15487
rect 16957 15453 16991 15487
rect 17417 15453 17451 15487
rect 20085 15453 20119 15487
rect 20821 15453 20855 15487
rect 21281 15453 21315 15487
rect 3065 15385 3099 15419
rect 5825 15385 5859 15419
rect 7420 15385 7454 15419
rect 9413 15385 9447 15419
rect 9965 15385 9999 15419
rect 10425 15385 10459 15419
rect 11253 15385 11287 15419
rect 14372 15385 14406 15419
rect 16712 15385 16746 15419
rect 18337 15385 18371 15419
rect 1501 15317 1535 15351
rect 4537 15317 4571 15351
rect 5917 15317 5951 15351
rect 10517 15317 10551 15351
rect 15485 15317 15519 15351
rect 17509 15317 17543 15351
rect 17877 15317 17911 15351
rect 18245 15317 18279 15351
rect 18705 15317 18739 15351
rect 1777 15113 1811 15147
rect 2053 15113 2087 15147
rect 2697 15113 2731 15147
rect 3065 15113 3099 15147
rect 5181 15113 5215 15147
rect 6193 15113 6227 15147
rect 6653 15113 6687 15147
rect 9597 15113 9631 15147
rect 11253 15113 11287 15147
rect 13737 15113 13771 15147
rect 15393 15113 15427 15147
rect 17325 15113 17359 15147
rect 18613 15113 18647 15147
rect 20729 15113 20763 15147
rect 21005 15113 21039 15147
rect 5273 15045 5307 15079
rect 6469 15045 6503 15079
rect 8585 15045 8619 15079
rect 17877 15045 17911 15079
rect 1685 14977 1719 15011
rect 1961 14977 1995 15011
rect 2237 14977 2271 15011
rect 2605 14977 2639 15011
rect 2881 14977 2915 15011
rect 4353 14977 4387 15011
rect 7869 14977 7903 15011
rect 8125 14977 8159 15011
rect 8493 14977 8527 15011
rect 9781 14977 9815 15011
rect 10048 14977 10082 15011
rect 12653 14977 12687 15011
rect 12909 14977 12943 15011
rect 14953 14977 14987 15011
rect 15209 14977 15243 15011
rect 18981 14977 19015 15011
rect 20545 14977 20579 15011
rect 20821 14977 20855 15011
rect 21281 14977 21315 15011
rect 4445 14909 4479 14943
rect 4629 14909 4663 14943
rect 5365 14909 5399 14943
rect 8309 14909 8343 14943
rect 17049 14909 17083 14943
rect 17233 14909 17267 14943
rect 19073 14909 19107 14943
rect 19165 14909 19199 14943
rect 2421 14841 2455 14875
rect 3985 14841 4019 14875
rect 11161 14841 11195 14875
rect 17693 14841 17727 14875
rect 1501 14773 1535 14807
rect 4813 14773 4847 14807
rect 6745 14773 6779 14807
rect 8953 14773 8987 14807
rect 11529 14773 11563 14807
rect 13829 14773 13863 14807
rect 21189 14773 21223 14807
rect 21465 14773 21499 14807
rect 2881 14569 2915 14603
rect 4537 14569 4571 14603
rect 9137 14569 9171 14603
rect 10701 14569 10735 14603
rect 11345 14569 11379 14603
rect 13829 14569 13863 14603
rect 14105 14569 14139 14603
rect 16865 14569 16899 14603
rect 19257 14569 19291 14603
rect 12909 14501 12943 14535
rect 20821 14501 20855 14535
rect 3985 14433 4019 14467
rect 5825 14433 5859 14467
rect 7849 14433 7883 14467
rect 9321 14433 9355 14467
rect 11529 14433 11563 14467
rect 15485 14433 15519 14467
rect 16221 14433 16255 14467
rect 19809 14433 19843 14467
rect 1685 14365 1719 14399
rect 2053 14365 2087 14399
rect 3065 14365 3099 14399
rect 4169 14365 4203 14399
rect 5549 14365 5583 14399
rect 7389 14365 7423 14399
rect 7941 14365 7975 14399
rect 8033 14365 8067 14399
rect 15218 14365 15252 14399
rect 16497 14365 16531 14399
rect 18889 14365 18923 14399
rect 19625 14365 19659 14399
rect 20637 14365 20671 14399
rect 20913 14365 20947 14399
rect 21281 14365 21315 14399
rect 5641 14297 5675 14331
rect 7122 14297 7156 14331
rect 9588 14297 9622 14331
rect 11774 14297 11808 14331
rect 19717 14297 19751 14331
rect 1501 14229 1535 14263
rect 1869 14229 1903 14263
rect 4077 14229 4111 14263
rect 5181 14229 5215 14263
rect 6009 14229 6043 14263
rect 8401 14229 8435 14263
rect 16405 14229 16439 14263
rect 17601 14229 17635 14263
rect 18705 14229 18739 14263
rect 19073 14229 19107 14263
rect 20085 14229 20119 14263
rect 21097 14229 21131 14263
rect 21465 14229 21499 14263
rect 1869 14025 1903 14059
rect 4537 14025 4571 14059
rect 4905 14025 4939 14059
rect 5365 14025 5399 14059
rect 5917 14025 5951 14059
rect 6193 14025 6227 14059
rect 8309 14025 8343 14059
rect 9873 14025 9907 14059
rect 13185 14025 13219 14059
rect 14013 14025 14047 14059
rect 16681 14025 16715 14059
rect 18245 14025 18279 14059
rect 18705 14025 18739 14059
rect 19073 14025 19107 14059
rect 19165 14025 19199 14059
rect 19533 14025 19567 14059
rect 4077 13957 4111 13991
rect 4629 13957 4663 13991
rect 10232 13957 10266 13991
rect 1685 13889 1719 13923
rect 2053 13889 2087 13923
rect 2145 13889 2179 13923
rect 4169 13889 4203 13923
rect 5273 13889 5307 13923
rect 6377 13889 6411 13923
rect 6644 13889 6678 13923
rect 8493 13889 8527 13923
rect 8760 13889 8794 13923
rect 9965 13889 9999 13923
rect 12817 13889 12851 13923
rect 14197 13889 14231 13923
rect 14464 13889 14498 13923
rect 17049 13889 17083 13923
rect 17877 13889 17911 13923
rect 21281 13889 21315 13923
rect 3985 13821 4019 13855
rect 5457 13821 5491 13855
rect 12541 13821 12575 13855
rect 12725 13821 12759 13855
rect 15853 13821 15887 13855
rect 17141 13821 17175 13855
rect 17233 13821 17267 13855
rect 17601 13821 17635 13855
rect 17785 13821 17819 13855
rect 18429 13821 18463 13855
rect 18613 13821 18647 13855
rect 19625 13821 19659 13855
rect 19717 13821 19751 13855
rect 15577 13753 15611 13787
rect 21189 13753 21223 13787
rect 1501 13685 1535 13719
rect 7757 13685 7791 13719
rect 11345 13685 11379 13719
rect 16037 13685 16071 13719
rect 21465 13685 21499 13719
rect 1869 13481 1903 13515
rect 4077 13481 4111 13515
rect 6193 13481 6227 13515
rect 7849 13481 7883 13515
rect 8677 13481 8711 13515
rect 10425 13481 10459 13515
rect 11161 13481 11195 13515
rect 12817 13481 12851 13515
rect 18245 13481 18279 13515
rect 21005 13481 21039 13515
rect 21281 13481 21315 13515
rect 1593 13413 1627 13447
rect 10333 13413 10367 13447
rect 15853 13413 15887 13447
rect 16681 13413 16715 13447
rect 4721 13345 4755 13379
rect 7757 13345 7791 13379
rect 8401 13345 8435 13379
rect 8953 13345 8987 13379
rect 13461 13345 13495 13379
rect 14381 13345 14415 13379
rect 15485 13345 15519 13379
rect 15577 13345 15611 13379
rect 16405 13345 16439 13379
rect 17233 13345 17267 13379
rect 17601 13345 17635 13379
rect 18981 13345 19015 13379
rect 1409 13277 1443 13311
rect 1685 13277 1719 13311
rect 2053 13277 2087 13311
rect 7501 13277 7535 13311
rect 8309 13277 8343 13311
rect 12725 13277 12759 13311
rect 14565 13277 14599 13311
rect 16221 13277 16255 13311
rect 17877 13277 17911 13311
rect 19257 13277 19291 13311
rect 20821 13277 20855 13311
rect 21097 13277 21131 13311
rect 21557 13277 21591 13311
rect 9220 13209 9254 13243
rect 12458 13209 12492 13243
rect 13277 13209 13311 13243
rect 14473 13209 14507 13243
rect 15393 13209 15427 13243
rect 2237 13141 2271 13175
rect 4445 13141 4479 13175
rect 4537 13141 4571 13175
rect 6377 13141 6411 13175
rect 8217 13141 8251 13175
rect 11345 13141 11379 13175
rect 13185 13141 13219 13175
rect 14933 13141 14967 13175
rect 15025 13141 15059 13175
rect 16313 13141 16347 13175
rect 17049 13141 17083 13175
rect 17141 13141 17175 13175
rect 17785 13141 17819 13175
rect 19441 13141 19475 13175
rect 20729 13141 20763 13175
rect 21373 13141 21407 13175
rect 2329 12937 2363 12971
rect 3433 12937 3467 12971
rect 3985 12937 4019 12971
rect 5365 12937 5399 12971
rect 8309 12937 8343 12971
rect 8861 12937 8895 12971
rect 9505 12937 9539 12971
rect 9597 12937 9631 12971
rect 9965 12937 9999 12971
rect 10333 12937 10367 12971
rect 11805 12937 11839 12971
rect 11897 12937 11931 12971
rect 12265 12937 12299 12971
rect 16957 12937 16991 12971
rect 17509 12937 17543 12971
rect 19073 12937 19107 12971
rect 19993 12937 20027 12971
rect 21005 12937 21039 12971
rect 2973 12869 3007 12903
rect 5917 12869 5951 12903
rect 7490 12869 7524 12903
rect 8769 12869 8803 12903
rect 14565 12869 14599 12903
rect 16221 12869 16255 12903
rect 16497 12869 16531 12903
rect 17877 12869 17911 12903
rect 2513 12801 2547 12835
rect 3065 12801 3099 12835
rect 3893 12801 3927 12835
rect 5825 12801 5859 12835
rect 7757 12801 7791 12835
rect 10425 12801 10459 12835
rect 12633 12801 12667 12835
rect 12725 12801 12759 12835
rect 12992 12801 13026 12835
rect 15770 12801 15804 12835
rect 16037 12801 16071 12835
rect 17049 12801 17083 12835
rect 18705 12801 18739 12835
rect 19809 12801 19843 12835
rect 20821 12801 20855 12835
rect 21097 12801 21131 12835
rect 21465 12801 21499 12835
rect 1961 12733 1995 12767
rect 2237 12733 2271 12767
rect 2881 12733 2915 12767
rect 4169 12733 4203 12767
rect 4905 12733 4939 12767
rect 6101 12733 6135 12767
rect 8033 12733 8067 12767
rect 8953 12733 8987 12767
rect 9413 12733 9447 12767
rect 10149 12733 10183 12767
rect 11713 12733 11747 12767
rect 16773 12733 16807 12767
rect 17969 12733 18003 12767
rect 18061 12733 18095 12767
rect 18429 12733 18463 12767
rect 18613 12733 18647 12767
rect 20269 12733 20303 12767
rect 3525 12665 3559 12699
rect 5457 12665 5491 12699
rect 8401 12665 8435 12699
rect 10793 12665 10827 12699
rect 14657 12665 14691 12699
rect 17417 12665 17451 12699
rect 21281 12665 21315 12699
rect 6377 12597 6411 12631
rect 10885 12597 10919 12631
rect 14105 12597 14139 12631
rect 2145 12393 2179 12427
rect 2789 12393 2823 12427
rect 3893 12393 3927 12427
rect 4445 12393 4479 12427
rect 7113 12393 7147 12427
rect 9781 12393 9815 12427
rect 13185 12393 13219 12427
rect 18613 12393 18647 12427
rect 19257 12393 19291 12427
rect 21373 12393 21407 12427
rect 1685 12325 1719 12359
rect 8769 12325 8803 12359
rect 15485 12325 15519 12359
rect 21189 12325 21223 12359
rect 2605 12257 2639 12291
rect 3249 12257 3283 12291
rect 3433 12257 3467 12291
rect 5089 12257 5123 12291
rect 7665 12257 7699 12291
rect 8125 12257 8159 12291
rect 8309 12257 8343 12291
rect 9229 12257 9263 12291
rect 9321 12257 9355 12291
rect 10057 12257 10091 12291
rect 11253 12257 11287 12291
rect 12633 12257 12667 12291
rect 12725 12257 12759 12291
rect 16865 12257 16899 12291
rect 17509 12257 17543 12291
rect 17969 12257 18003 12291
rect 19809 12257 19843 12291
rect 20637 12257 20671 12291
rect 1501 12189 1535 12223
rect 2329 12189 2363 12223
rect 3157 12189 3191 12223
rect 3985 12189 4019 12223
rect 4813 12189 4847 12223
rect 6193 12189 6227 12223
rect 6469 12189 6503 12223
rect 7481 12189 7515 12223
rect 8401 12189 8435 12223
rect 10241 12189 10275 12223
rect 11529 12189 11563 12223
rect 14105 12189 14139 12223
rect 18705 12189 18739 12223
rect 20453 12189 20487 12223
rect 1869 12121 1903 12155
rect 2421 12121 2455 12155
rect 9413 12121 9447 12155
rect 11161 12121 11195 12155
rect 12817 12121 12851 12155
rect 14372 12121 14406 12155
rect 19625 12121 19659 12155
rect 20545 12121 20579 12155
rect 21005 12121 21039 12155
rect 21465 12121 21499 12155
rect 1961 12053 1995 12087
rect 4905 12053 4939 12087
rect 6009 12053 6043 12087
rect 7573 12053 7607 12087
rect 10149 12053 10183 12087
rect 10609 12053 10643 12087
rect 10701 12053 10735 12087
rect 11069 12053 11103 12087
rect 12173 12053 12207 12087
rect 12265 12053 12299 12087
rect 13921 12053 13955 12087
rect 16957 12053 16991 12087
rect 17325 12053 17359 12087
rect 17417 12053 17451 12087
rect 18153 12053 18187 12087
rect 18245 12053 18279 12087
rect 19717 12053 19751 12087
rect 20085 12053 20119 12087
rect 1869 11849 1903 11883
rect 2329 11849 2363 11883
rect 5733 11849 5767 11883
rect 8953 11849 8987 11883
rect 10885 11849 10919 11883
rect 14289 11849 14323 11883
rect 16957 11849 16991 11883
rect 17509 11849 17543 11883
rect 18337 11849 18371 11883
rect 18797 11849 18831 11883
rect 19165 11849 19199 11883
rect 20361 11849 20395 11883
rect 21373 11849 21407 11883
rect 2605 11781 2639 11815
rect 12164 11781 12198 11815
rect 17969 11781 18003 11815
rect 19533 11781 19567 11815
rect 1501 11713 1535 11747
rect 2053 11713 2087 11747
rect 2145 11713 2179 11747
rect 2421 11713 2455 11747
rect 6377 11713 6411 11747
rect 6644 11713 6678 11747
rect 8217 11713 8251 11747
rect 9137 11713 9171 11747
rect 9404 11713 9438 11747
rect 10977 11713 11011 11747
rect 15413 11713 15447 11747
rect 17049 11713 17083 11747
rect 17877 11713 17911 11747
rect 18705 11713 18739 11747
rect 21281 11713 21315 11747
rect 21557 11713 21591 11747
rect 1685 11645 1719 11679
rect 5825 11645 5859 11679
rect 6009 11645 6043 11679
rect 8309 11645 8343 11679
rect 8401 11645 8435 11679
rect 10793 11645 10827 11679
rect 11897 11645 11931 11679
rect 15669 11645 15703 11679
rect 16865 11645 16899 11679
rect 18061 11645 18095 11679
rect 18889 11645 18923 11679
rect 19625 11645 19659 11679
rect 19809 11645 19843 11679
rect 19993 11645 20027 11679
rect 20729 11645 20763 11679
rect 7757 11577 7791 11611
rect 10517 11577 10551 11611
rect 11345 11577 11379 11611
rect 14105 11577 14139 11611
rect 17417 11577 17451 11611
rect 20913 11577 20947 11611
rect 5365 11509 5399 11543
rect 7849 11509 7883 11543
rect 8677 11509 8711 11543
rect 11713 11509 11747 11543
rect 13277 11509 13311 11543
rect 21097 11509 21131 11543
rect 1961 11305 1995 11339
rect 7297 11305 7331 11339
rect 10701 11305 10735 11339
rect 15853 11305 15887 11339
rect 17141 11305 17175 11339
rect 17325 11305 17359 11339
rect 19257 11305 19291 11339
rect 20177 11305 20211 11339
rect 1685 11237 1719 11271
rect 8769 11237 8803 11271
rect 13737 11237 13771 11271
rect 15485 11237 15519 11271
rect 20637 11237 20671 11271
rect 2697 11169 2731 11203
rect 4445 11169 4479 11203
rect 5089 11169 5123 11203
rect 10885 11169 10919 11203
rect 12357 11169 12391 11203
rect 16221 11169 16255 11203
rect 16589 11169 16623 11203
rect 19809 11169 19843 11203
rect 20913 11169 20947 11203
rect 1777 11101 1811 11135
rect 2513 11101 2547 11135
rect 4169 11101 4203 11135
rect 4813 11101 4847 11135
rect 5825 11101 5859 11135
rect 5917 11101 5951 11135
rect 7389 11101 7423 11135
rect 8953 11101 8987 11135
rect 9220 11101 9254 11135
rect 11152 11101 11186 11135
rect 13921 11101 13955 11135
rect 14105 11101 14139 11135
rect 18797 11101 18831 11135
rect 18981 11101 19015 11135
rect 19625 11101 19659 11135
rect 20821 11101 20855 11135
rect 21281 11101 21315 11135
rect 21465 11101 21499 11135
rect 1501 11033 1535 11067
rect 2881 11033 2915 11067
rect 4629 11033 4663 11067
rect 6162 11033 6196 11067
rect 7656 11033 7690 11067
rect 12624 11033 12658 11067
rect 14350 11033 14384 11067
rect 15761 11033 15795 11067
rect 16681 11033 16715 11067
rect 16773 11033 16807 11067
rect 19717 11033 19751 11067
rect 20545 11033 20579 11067
rect 21097 11033 21131 11067
rect 2053 10965 2087 10999
rect 2421 10965 2455 10999
rect 3801 10965 3835 10999
rect 4261 10965 4295 10999
rect 10333 10965 10367 10999
rect 12265 10965 12299 10999
rect 1777 10761 1811 10795
rect 2237 10761 2271 10795
rect 2329 10761 2363 10795
rect 2789 10761 2823 10795
rect 3801 10761 3835 10795
rect 10333 10761 10367 10795
rect 10793 10761 10827 10795
rect 12265 10761 12299 10795
rect 14197 10761 14231 10795
rect 17693 10761 17727 10795
rect 18061 10761 18095 10795
rect 18521 10761 18555 10795
rect 19809 10761 19843 10795
rect 20085 10761 20119 10795
rect 20821 10761 20855 10795
rect 7490 10693 7524 10727
rect 9220 10693 9254 10727
rect 15402 10693 15436 10727
rect 1869 10625 1903 10659
rect 2697 10625 2731 10659
rect 4629 10625 4663 10659
rect 4721 10625 4755 10659
rect 5365 10625 5399 10659
rect 10701 10625 10735 10659
rect 17325 10625 17359 10659
rect 18153 10625 18187 10659
rect 19441 10625 19475 10659
rect 19901 10625 19935 10659
rect 20177 10625 20211 10659
rect 20729 10625 20763 10659
rect 21465 10625 21499 10659
rect 1685 10557 1719 10591
rect 2973 10557 3007 10591
rect 3893 10557 3927 10591
rect 4077 10557 4111 10591
rect 4813 10557 4847 10591
rect 7757 10557 7791 10591
rect 8953 10557 8987 10591
rect 10517 10557 10551 10591
rect 15669 10557 15703 10591
rect 17049 10557 17083 10591
rect 17233 10557 17267 10591
rect 17969 10557 18003 10591
rect 19257 10557 19291 10591
rect 19349 10557 19383 10591
rect 20913 10557 20947 10591
rect 6193 10489 6227 10523
rect 11161 10489 11195 10523
rect 21281 10489 21315 10523
rect 3433 10421 3467 10455
rect 4261 10421 4295 10455
rect 5181 10421 5215 10455
rect 6377 10421 6411 10455
rect 7849 10421 7883 10455
rect 8585 10421 8619 10455
rect 8769 10421 8803 10455
rect 14289 10421 14323 10455
rect 18981 10421 19015 10455
rect 20361 10421 20395 10455
rect 2329 10217 2363 10251
rect 2789 10217 2823 10251
rect 3985 10217 4019 10251
rect 10333 10217 10367 10251
rect 17417 10217 17451 10251
rect 18337 10217 18371 10251
rect 19993 10217 20027 10251
rect 21189 10217 21223 10251
rect 21373 10217 21407 10251
rect 1685 10149 1719 10183
rect 5733 10149 5767 10183
rect 13093 10149 13127 10183
rect 18245 10149 18279 10183
rect 2053 10081 2087 10115
rect 3341 10081 3375 10115
rect 4629 10081 4663 10115
rect 9781 10081 9815 10115
rect 15669 10081 15703 10115
rect 16589 10081 16623 10115
rect 16865 10081 16899 10115
rect 18889 10081 18923 10115
rect 19349 10081 19383 10115
rect 20637 10081 20671 10115
rect 20729 10081 20763 10115
rect 1501 10013 1535 10047
rect 2145 10013 2179 10047
rect 2421 10013 2455 10047
rect 3157 10013 3191 10047
rect 4445 10013 4479 10047
rect 4905 10013 4939 10047
rect 5457 10013 5491 10047
rect 5641 10013 5675 10047
rect 7113 10013 7147 10047
rect 11621 10013 11655 10047
rect 11713 10013 11747 10047
rect 14197 10013 14231 10047
rect 16957 10013 16991 10047
rect 18705 10013 18739 10047
rect 19533 10013 19567 10047
rect 21005 10013 21039 10047
rect 21465 10013 21499 10047
rect 1869 9945 1903 9979
rect 2605 9945 2639 9979
rect 3249 9945 3283 9979
rect 6868 9945 6902 9979
rect 11958 9945 11992 9979
rect 15402 9945 15436 9979
rect 4353 9877 4387 9911
rect 9873 9877 9907 9911
rect 9965 9877 9999 9911
rect 14289 9877 14323 9911
rect 17049 9877 17083 9911
rect 18797 9877 18831 9911
rect 19625 9877 19659 9911
rect 20177 9877 20211 9911
rect 20545 9877 20579 9911
rect 2329 9673 2363 9707
rect 3249 9673 3283 9707
rect 4813 9673 4847 9707
rect 17417 9673 17451 9707
rect 19441 9673 19475 9707
rect 19901 9673 19935 9707
rect 20637 9673 20671 9707
rect 4077 9605 4111 9639
rect 10140 9605 10174 9639
rect 18153 9605 18187 9639
rect 2789 9537 2823 9571
rect 5926 9537 5960 9571
rect 7490 9537 7524 9571
rect 7757 9537 7791 9571
rect 8217 9537 8251 9571
rect 8473 9537 8507 9571
rect 14729 9537 14763 9571
rect 18245 9537 18279 9571
rect 19073 9537 19107 9571
rect 21281 9537 21315 9571
rect 1409 9469 1443 9503
rect 1685 9469 1719 9503
rect 3341 9469 3375 9503
rect 3433 9469 3467 9503
rect 4169 9469 4203 9503
rect 4353 9469 4387 9503
rect 6193 9469 6227 9503
rect 9873 9469 9907 9503
rect 14473 9469 14507 9503
rect 17141 9469 17175 9503
rect 17325 9469 17359 9503
rect 18061 9469 18095 9503
rect 18889 9469 18923 9503
rect 18981 9469 19015 9503
rect 19993 9469 20027 9503
rect 20085 9469 20119 9503
rect 21557 9469 21591 9503
rect 15945 9401 15979 9435
rect 16957 9401 16991 9435
rect 17785 9401 17819 9435
rect 18613 9401 18647 9435
rect 19533 9401 19567 9435
rect 2605 9333 2639 9367
rect 2881 9333 2915 9367
rect 3709 9333 3743 9367
rect 6377 9333 6411 9367
rect 7941 9333 7975 9367
rect 8033 9333 8067 9367
rect 9597 9333 9631 9367
rect 9781 9333 9815 9367
rect 11253 9333 11287 9367
rect 14289 9333 14323 9367
rect 15853 9333 15887 9367
rect 2421 9129 2455 9163
rect 6285 9129 6319 9163
rect 15485 9129 15519 9163
rect 19257 9129 19291 9163
rect 20637 9129 20671 9163
rect 7849 9061 7883 9095
rect 8769 9061 8803 9095
rect 9045 9061 9079 9095
rect 16957 9061 16991 9095
rect 17969 9061 18003 9095
rect 20361 9061 20395 9095
rect 1961 8993 1995 9027
rect 2881 8993 2915 9027
rect 3065 8993 3099 9027
rect 8401 8993 8435 9027
rect 17601 8993 17635 9027
rect 18521 8993 18555 9027
rect 19901 8993 19935 9027
rect 21005 8993 21039 9027
rect 2237 8925 2271 8959
rect 3249 8925 3283 8959
rect 4905 8925 4939 8959
rect 6377 8925 6411 8959
rect 8217 8925 8251 8959
rect 10250 8925 10284 8959
rect 10517 8925 10551 8959
rect 10609 8925 10643 8959
rect 10865 8925 10899 8959
rect 13205 8925 13239 8959
rect 13461 8925 13495 8959
rect 14105 8925 14139 8959
rect 15577 8925 15611 8959
rect 15844 8925 15878 8959
rect 20453 8925 20487 8959
rect 20729 8925 20763 8959
rect 5172 8857 5206 8891
rect 6622 8857 6656 8891
rect 14372 8857 14406 8891
rect 17509 8857 17543 8891
rect 20177 8857 20211 8891
rect 2789 8789 2823 8823
rect 7757 8789 7791 8823
rect 8309 8789 8343 8823
rect 9137 8789 9171 8823
rect 11989 8789 12023 8823
rect 12081 8789 12115 8823
rect 13829 8789 13863 8823
rect 17049 8789 17083 8823
rect 17417 8789 17451 8823
rect 18613 8789 18647 8823
rect 18705 8789 18739 8823
rect 19073 8789 19107 8823
rect 19625 8789 19659 8823
rect 19717 8789 19751 8823
rect 1593 8585 1627 8619
rect 2421 8585 2455 8619
rect 2881 8585 2915 8619
rect 3249 8585 3283 8619
rect 3801 8585 3835 8619
rect 4261 8585 4295 8619
rect 11345 8585 11379 8619
rect 13461 8585 13495 8619
rect 17417 8585 17451 8619
rect 17969 8585 18003 8619
rect 18889 8585 18923 8619
rect 19533 8585 19567 8619
rect 19993 8585 20027 8619
rect 20821 8585 20855 8619
rect 3617 8517 3651 8551
rect 6469 8517 6503 8551
rect 6653 8517 6687 8551
rect 7205 8517 7239 8551
rect 10333 8517 10367 8551
rect 10885 8517 10919 8551
rect 12348 8517 12382 8551
rect 16230 8517 16264 8551
rect 21189 8517 21223 8551
rect 1409 8449 1443 8483
rect 2053 8449 2087 8483
rect 4169 8449 4203 8483
rect 8410 8449 8444 8483
rect 8677 8449 8711 8483
rect 8769 8449 8803 8483
rect 9025 8449 9059 8483
rect 10977 8449 11011 8483
rect 14769 8449 14803 8483
rect 15025 8449 15059 8483
rect 16497 8449 16531 8483
rect 17049 8449 17083 8483
rect 17877 8449 17911 8483
rect 18337 8449 18371 8483
rect 18797 8449 18831 8483
rect 19073 8449 19107 8483
rect 20361 8449 20395 8483
rect 1777 8381 1811 8415
rect 1961 8381 1995 8415
rect 2605 8381 2639 8415
rect 2789 8381 2823 8415
rect 3341 8381 3375 8415
rect 4353 8381 4387 8415
rect 10701 8381 10735 8415
rect 11805 8381 11839 8415
rect 12081 8381 12115 8415
rect 16773 8381 16807 8415
rect 16957 8381 16991 8415
rect 18153 8381 18187 8415
rect 19625 8381 19659 8415
rect 19717 8381 19751 8415
rect 20453 8381 20487 8415
rect 20545 8381 20579 8415
rect 21281 8381 21315 8415
rect 21373 8381 21407 8415
rect 7297 8313 7331 8347
rect 10149 8313 10183 8347
rect 10517 8313 10551 8347
rect 13645 8313 13679 8347
rect 15117 8313 15151 8347
rect 19165 8313 19199 8347
rect 11989 8245 12023 8279
rect 17509 8245 17543 8279
rect 1409 8041 1443 8075
rect 2421 8041 2455 8075
rect 2513 8041 2547 8075
rect 3525 8041 3559 8075
rect 11069 8041 11103 8075
rect 17141 8041 17175 8075
rect 19625 8041 19659 8075
rect 20545 8041 20579 8075
rect 21373 8041 21407 8075
rect 21557 8041 21591 8075
rect 4353 7973 4387 8007
rect 5273 7973 5307 8007
rect 5641 7973 5675 8007
rect 7389 7973 7423 8007
rect 9689 7973 9723 8007
rect 11161 7973 11195 8007
rect 14105 7973 14139 8007
rect 1869 7905 1903 7939
rect 3157 7905 3191 7939
rect 4997 7905 5031 7939
rect 9137 7905 9171 7939
rect 10517 7905 10551 7939
rect 16497 7905 16531 7939
rect 16589 7905 16623 7939
rect 17693 7905 17727 7939
rect 18613 7905 18647 7939
rect 20177 7905 20211 7939
rect 20729 7905 20763 7939
rect 2053 7837 2087 7871
rect 5549 7837 5583 7871
rect 7021 7837 7055 7871
rect 7297 7837 7331 7871
rect 8769 7837 8803 7871
rect 9229 7837 9263 7871
rect 10609 7837 10643 7871
rect 10701 7837 10735 7871
rect 12541 7837 12575 7871
rect 13461 7837 13495 7871
rect 13829 7837 13863 7871
rect 15485 7837 15519 7871
rect 15577 7837 15611 7871
rect 16681 7837 16715 7871
rect 21005 7837 21039 7871
rect 1961 7769 1995 7803
rect 2881 7769 2915 7803
rect 3433 7769 3467 7803
rect 3801 7769 3835 7803
rect 6776 7769 6810 7803
rect 8502 7769 8536 7803
rect 12296 7769 12330 7803
rect 15218 7769 15252 7803
rect 17601 7769 17635 7803
rect 18337 7769 18371 7803
rect 20913 7769 20947 7803
rect 2973 7701 3007 7735
rect 4721 7701 4755 7735
rect 4813 7701 4847 7735
rect 9321 7701 9355 7735
rect 17049 7701 17083 7735
rect 17509 7701 17543 7735
rect 17969 7701 18003 7735
rect 18429 7701 18463 7735
rect 19993 7701 20027 7735
rect 20085 7701 20119 7735
rect 3157 7497 3191 7531
rect 3525 7497 3559 7531
rect 4261 7497 4295 7531
rect 4629 7497 4663 7531
rect 5089 7497 5123 7531
rect 5457 7497 5491 7531
rect 8953 7497 8987 7531
rect 9413 7497 9447 7531
rect 9965 7497 9999 7531
rect 10333 7497 10367 7531
rect 10701 7497 10735 7531
rect 11253 7497 11287 7531
rect 16865 7497 16899 7531
rect 17233 7497 17267 7531
rect 18153 7497 18187 7531
rect 20637 7497 20671 7531
rect 4721 7429 4755 7463
rect 6009 7429 6043 7463
rect 10793 7429 10827 7463
rect 17325 7429 17359 7463
rect 18521 7429 18555 7463
rect 18613 7429 18647 7463
rect 2789 7361 2823 7395
rect 3249 7361 3283 7395
rect 3709 7361 3743 7395
rect 8585 7361 8619 7395
rect 9045 7361 9079 7395
rect 9873 7361 9907 7395
rect 20453 7361 20487 7395
rect 21005 7361 21039 7395
rect 1961 7293 1995 7327
rect 2237 7293 2271 7327
rect 2513 7293 2547 7327
rect 2697 7293 2731 7327
rect 4813 7293 4847 7327
rect 5549 7293 5583 7327
rect 5733 7293 5767 7327
rect 8769 7293 8803 7327
rect 10057 7293 10091 7327
rect 10885 7293 10919 7327
rect 17417 7293 17451 7327
rect 18705 7293 18739 7327
rect 20177 7293 20211 7327
rect 20729 7293 20763 7327
rect 9505 7225 9539 7259
rect 3893 7157 3927 7191
rect 8217 7157 8251 7191
rect 17785 7157 17819 7191
rect 20269 7157 20303 7191
rect 4997 6953 5031 6987
rect 9689 6953 9723 6987
rect 1961 6885 1995 6919
rect 20913 6885 20947 6919
rect 2605 6817 2639 6851
rect 3525 6817 3559 6851
rect 3985 6817 4019 6851
rect 4445 6817 4479 6851
rect 5641 6817 5675 6851
rect 6469 6817 6503 6851
rect 9045 6817 9079 6851
rect 10425 6817 10459 6851
rect 12541 6817 12575 6851
rect 20361 6817 20395 6851
rect 21281 6817 21315 6851
rect 1501 6749 1535 6783
rect 1777 6749 1811 6783
rect 2421 6749 2455 6783
rect 4537 6749 4571 6783
rect 6377 6749 6411 6783
rect 20545 6749 20579 6783
rect 20821 6749 20855 6783
rect 21097 6749 21131 6783
rect 21465 6749 21499 6783
rect 3801 6681 3835 6715
rect 5457 6681 5491 6715
rect 6285 6681 6319 6715
rect 6745 6681 6779 6715
rect 9781 6681 9815 6715
rect 12817 6681 12851 6715
rect 13277 6681 13311 6715
rect 20177 6681 20211 6715
rect 1593 6613 1627 6647
rect 2053 6613 2087 6647
rect 2513 6613 2547 6647
rect 2881 6613 2915 6647
rect 3249 6613 3283 6647
rect 3341 6613 3375 6647
rect 4629 6613 4663 6647
rect 5089 6613 5123 6647
rect 5549 6613 5583 6647
rect 5917 6613 5951 6647
rect 9229 6613 9263 6647
rect 9321 6613 9355 6647
rect 12725 6613 12759 6647
rect 13185 6613 13219 6647
rect 20637 6613 20671 6647
rect 2605 6409 2639 6443
rect 3157 6409 3191 6443
rect 3525 6409 3559 6443
rect 4905 6409 4939 6443
rect 5273 6409 5307 6443
rect 11713 6409 11747 6443
rect 12725 6409 12759 6443
rect 14197 6409 14231 6443
rect 14657 6409 14691 6443
rect 15485 6409 15519 6443
rect 3065 6341 3099 6375
rect 3985 6341 4019 6375
rect 12081 6341 12115 6375
rect 15393 6341 15427 6375
rect 15945 6341 15979 6375
rect 13093 6273 13127 6307
rect 14565 6273 14599 6307
rect 21005 6273 21039 6307
rect 1961 6205 1995 6239
rect 2237 6205 2271 6239
rect 2329 6205 2363 6239
rect 2973 6205 3007 6239
rect 4077 6205 4111 6239
rect 4169 6205 4203 6239
rect 5365 6205 5399 6239
rect 5457 6205 5491 6239
rect 5825 6205 5859 6239
rect 12173 6205 12207 6239
rect 12265 6205 12299 6239
rect 13185 6205 13219 6239
rect 13369 6205 13403 6239
rect 14105 6205 14139 6239
rect 14749 6205 14783 6239
rect 15577 6205 15611 6239
rect 20637 6205 20671 6239
rect 20729 6205 20763 6239
rect 15025 6137 15059 6171
rect 3617 6069 3651 6103
rect 1777 5865 1811 5899
rect 3341 5865 3375 5899
rect 5365 5865 5399 5899
rect 21097 5865 21131 5899
rect 2421 5729 2455 5763
rect 2789 5729 2823 5763
rect 4721 5729 4755 5763
rect 14565 5729 14599 5763
rect 20821 5729 20855 5763
rect 1409 5661 1443 5695
rect 21005 5661 21039 5695
rect 21281 5661 21315 5695
rect 21557 5661 21591 5695
rect 2237 5593 2271 5627
rect 2973 5593 3007 5627
rect 4905 5593 4939 5627
rect 1593 5525 1627 5559
rect 2145 5525 2179 5559
rect 2881 5525 2915 5559
rect 4997 5525 5031 5559
rect 21373 5525 21407 5559
rect 1593 5321 1627 5355
rect 2421 5321 2455 5355
rect 2789 5321 2823 5355
rect 21373 5321 21407 5355
rect 2053 5253 2087 5287
rect 1409 5185 1443 5219
rect 2881 5185 2915 5219
rect 21281 5185 21315 5219
rect 21557 5185 21591 5219
rect 1869 5117 1903 5151
rect 1961 5117 1995 5151
rect 2513 5049 2547 5083
rect 1593 4777 1627 4811
rect 2145 4777 2179 4811
rect 1869 4709 1903 4743
rect 21005 4641 21039 4675
rect 1409 4573 1443 4607
rect 1685 4573 1719 4607
rect 1961 4573 1995 4607
rect 2237 4573 2271 4607
rect 20637 4573 20671 4607
rect 20729 4573 20763 4607
rect 1685 4233 1719 4267
rect 21097 4233 21131 4267
rect 1869 4165 1903 4199
rect 1409 4097 1443 4131
rect 2053 4097 2087 4131
rect 21005 4097 21039 4131
rect 21281 4097 21315 4131
rect 21557 4097 21591 4131
rect 20821 4029 20855 4063
rect 1593 3961 1627 3995
rect 21373 3961 21407 3995
rect 1593 3689 1627 3723
rect 21373 3689 21407 3723
rect 1409 3485 1443 3519
rect 1685 3485 1719 3519
rect 21281 3485 21315 3519
rect 21557 3485 21591 3519
rect 1869 3349 1903 3383
rect 1593 3145 1627 3179
rect 1869 3145 1903 3179
rect 2145 3145 2179 3179
rect 6193 3145 6227 3179
rect 21373 3145 21407 3179
rect 1409 3009 1443 3043
rect 1685 3009 1719 3043
rect 1961 3009 1995 3043
rect 6009 3009 6043 3043
rect 9137 3009 9171 3043
rect 17049 3009 17083 3043
rect 21005 3009 21039 3043
rect 21281 3009 21315 3043
rect 21557 3009 21591 3043
rect 2421 2941 2455 2975
rect 20821 2941 20855 2975
rect 8953 2873 8987 2907
rect 16865 2873 16899 2907
rect 21097 2873 21131 2907
rect 2237 2805 2271 2839
rect 2513 2601 2547 2635
rect 11529 2601 11563 2635
rect 16129 2601 16163 2635
rect 20729 2601 20763 2635
rect 21097 2601 21131 2635
rect 20269 2533 20303 2567
rect 1961 2465 1995 2499
rect 20453 2465 20487 2499
rect 2237 2397 2271 2431
rect 2329 2397 2363 2431
rect 2605 2397 2639 2431
rect 7205 2397 7239 2431
rect 11713 2397 11747 2431
rect 16313 2397 16347 2431
rect 20913 2397 20947 2431
rect 21281 2397 21315 2431
rect 21557 2397 21591 2431
rect 2789 2329 2823 2363
rect 7021 2261 7055 2295
rect 11805 2261 11839 2295
rect 16037 2261 16071 2295
rect 20637 2261 20671 2295
rect 21373 2261 21407 2295
<< metal1 >>
rect 8938 20816 8944 20868
rect 8996 20856 9002 20868
rect 15562 20856 15568 20868
rect 8996 20828 15568 20856
rect 8996 20816 9002 20828
rect 15562 20816 15568 20828
rect 15620 20816 15626 20868
rect 1104 20698 22056 20720
rect 1104 20646 6148 20698
rect 6200 20646 6212 20698
rect 6264 20646 6276 20698
rect 6328 20646 6340 20698
rect 6392 20646 6404 20698
rect 6456 20646 11346 20698
rect 11398 20646 11410 20698
rect 11462 20646 11474 20698
rect 11526 20646 11538 20698
rect 11590 20646 11602 20698
rect 11654 20646 16544 20698
rect 16596 20646 16608 20698
rect 16660 20646 16672 20698
rect 16724 20646 16736 20698
rect 16788 20646 16800 20698
rect 16852 20646 21742 20698
rect 21794 20646 21806 20698
rect 21858 20646 21870 20698
rect 21922 20646 21934 20698
rect 21986 20646 21998 20698
rect 22050 20646 22056 20698
rect 1104 20624 22056 20646
rect 5534 20584 5540 20596
rect 5495 20556 5540 20584
rect 5534 20544 5540 20556
rect 5592 20544 5598 20596
rect 5718 20544 5724 20596
rect 5776 20584 5782 20596
rect 5905 20587 5963 20593
rect 5905 20584 5917 20587
rect 5776 20556 5917 20584
rect 5776 20544 5782 20556
rect 5905 20553 5917 20556
rect 5951 20553 5963 20587
rect 5905 20547 5963 20553
rect 5994 20544 6000 20596
rect 6052 20584 6058 20596
rect 6549 20587 6607 20593
rect 6549 20584 6561 20587
rect 6052 20556 6561 20584
rect 6052 20544 6058 20556
rect 6549 20553 6561 20556
rect 6595 20553 6607 20587
rect 6549 20547 6607 20553
rect 7374 20544 7380 20596
rect 7432 20584 7438 20596
rect 8938 20584 8944 20596
rect 7432 20556 8944 20584
rect 7432 20544 7438 20556
rect 8938 20544 8944 20556
rect 8996 20544 9002 20596
rect 9030 20544 9036 20596
rect 9088 20544 9094 20596
rect 9214 20544 9220 20596
rect 9272 20584 9278 20596
rect 9309 20587 9367 20593
rect 9309 20584 9321 20587
rect 9272 20556 9321 20584
rect 9272 20544 9278 20556
rect 9309 20553 9321 20556
rect 9355 20553 9367 20587
rect 9766 20584 9772 20596
rect 9309 20547 9367 20553
rect 9416 20556 9772 20584
rect 4246 20476 4252 20528
rect 4304 20516 4310 20528
rect 4522 20516 4528 20528
rect 4304 20488 4528 20516
rect 4304 20476 4310 20488
rect 4522 20476 4528 20488
rect 4580 20516 4586 20528
rect 4801 20519 4859 20525
rect 4801 20516 4813 20519
rect 4580 20488 4813 20516
rect 4580 20476 4586 20488
rect 4801 20485 4813 20488
rect 4847 20485 4859 20519
rect 5442 20516 5448 20528
rect 4801 20479 4859 20485
rect 5184 20488 5448 20516
rect 1670 20448 1676 20460
rect 1631 20420 1676 20448
rect 1670 20408 1676 20420
rect 1728 20408 1734 20460
rect 2038 20408 2044 20460
rect 2096 20448 2102 20460
rect 2685 20451 2743 20457
rect 2685 20448 2697 20451
rect 2096 20420 2697 20448
rect 2096 20408 2102 20420
rect 2685 20417 2697 20420
rect 2731 20417 2743 20451
rect 2685 20411 2743 20417
rect 2866 20408 2872 20460
rect 2924 20448 2930 20460
rect 2924 20420 3464 20448
rect 2924 20408 2930 20420
rect 2409 20383 2467 20389
rect 2409 20349 2421 20383
rect 2455 20349 2467 20383
rect 2409 20343 2467 20349
rect 2424 20312 2452 20343
rect 3234 20340 3240 20392
rect 3292 20380 3298 20392
rect 3329 20383 3387 20389
rect 3329 20380 3341 20383
rect 3292 20352 3341 20380
rect 3292 20340 3298 20352
rect 3329 20349 3341 20352
rect 3375 20349 3387 20383
rect 3436 20380 3464 20420
rect 3510 20408 3516 20460
rect 3568 20448 3574 20460
rect 5184 20457 5212 20488
rect 5442 20476 5448 20488
rect 5500 20516 5506 20528
rect 6822 20516 6828 20528
rect 5500 20488 6828 20516
rect 5500 20476 5506 20488
rect 6822 20476 6828 20488
rect 6880 20476 6886 20528
rect 7006 20476 7012 20528
rect 7064 20516 7070 20528
rect 7558 20516 7564 20528
rect 7064 20488 7564 20516
rect 7064 20476 7070 20488
rect 3789 20451 3847 20457
rect 3789 20448 3801 20451
rect 3568 20420 3801 20448
rect 3568 20408 3574 20420
rect 3789 20417 3801 20420
rect 3835 20417 3847 20451
rect 3789 20411 3847 20417
rect 5169 20451 5227 20457
rect 5169 20417 5181 20451
rect 5215 20417 5227 20451
rect 5169 20411 5227 20417
rect 5534 20408 5540 20460
rect 5592 20448 5598 20460
rect 5721 20451 5779 20457
rect 5721 20448 5733 20451
rect 5592 20420 5733 20448
rect 5592 20408 5598 20420
rect 5721 20417 5733 20420
rect 5767 20417 5779 20451
rect 5721 20411 5779 20417
rect 5810 20408 5816 20460
rect 5868 20448 5874 20460
rect 6089 20451 6147 20457
rect 6089 20448 6101 20451
rect 5868 20420 6101 20448
rect 5868 20408 5874 20420
rect 6089 20417 6101 20420
rect 6135 20417 6147 20451
rect 6362 20448 6368 20460
rect 6323 20420 6368 20448
rect 6089 20411 6147 20417
rect 6362 20408 6368 20420
rect 6420 20408 6426 20460
rect 6917 20451 6975 20457
rect 6917 20417 6929 20451
rect 6963 20448 6975 20451
rect 7098 20448 7104 20460
rect 6963 20420 7104 20448
rect 6963 20417 6975 20420
rect 6917 20411 6975 20417
rect 7098 20408 7104 20420
rect 7156 20408 7162 20460
rect 7208 20457 7236 20488
rect 7558 20476 7564 20488
rect 7616 20476 7622 20528
rect 8294 20516 8300 20528
rect 7944 20488 8300 20516
rect 7193 20451 7251 20457
rect 7193 20417 7205 20451
rect 7239 20417 7251 20451
rect 7193 20411 7251 20417
rect 7469 20451 7527 20457
rect 7469 20417 7481 20451
rect 7515 20448 7527 20451
rect 7834 20448 7840 20460
rect 7515 20420 7840 20448
rect 7515 20417 7527 20420
rect 7469 20411 7527 20417
rect 7834 20408 7840 20420
rect 7892 20408 7898 20460
rect 7944 20457 7972 20488
rect 8294 20476 8300 20488
rect 8352 20476 8358 20528
rect 9048 20516 9076 20544
rect 8496 20488 9076 20516
rect 7929 20451 7987 20457
rect 7929 20417 7941 20451
rect 7975 20417 7987 20451
rect 7929 20411 7987 20417
rect 8018 20408 8024 20460
rect 8076 20448 8082 20460
rect 8386 20448 8392 20460
rect 8076 20420 8392 20448
rect 8076 20408 8082 20420
rect 8386 20408 8392 20420
rect 8444 20408 8450 20460
rect 8496 20457 8524 20488
rect 8481 20451 8539 20457
rect 8481 20417 8493 20451
rect 8527 20417 8539 20451
rect 8481 20411 8539 20417
rect 8573 20451 8631 20457
rect 8573 20417 8585 20451
rect 8619 20417 8631 20451
rect 8573 20411 8631 20417
rect 9033 20451 9091 20457
rect 9033 20417 9045 20451
rect 9079 20448 9091 20451
rect 9416 20448 9444 20556
rect 9766 20544 9772 20556
rect 9824 20544 9830 20596
rect 10502 20544 10508 20596
rect 10560 20544 10566 20596
rect 11241 20587 11299 20593
rect 11241 20553 11253 20587
rect 11287 20584 11299 20587
rect 15933 20587 15991 20593
rect 15933 20584 15945 20587
rect 11287 20556 15424 20584
rect 11287 20553 11299 20556
rect 11241 20547 11299 20553
rect 10520 20516 10548 20544
rect 9784 20488 10548 20516
rect 9079 20420 9444 20448
rect 9493 20451 9551 20457
rect 9079 20417 9091 20420
rect 9033 20411 9091 20417
rect 9493 20417 9505 20451
rect 9539 20448 9551 20451
rect 9582 20448 9588 20460
rect 9539 20420 9588 20448
rect 9539 20417 9551 20420
rect 9493 20411 9551 20417
rect 3605 20383 3663 20389
rect 3605 20380 3617 20383
rect 3436 20352 3617 20380
rect 3329 20343 3387 20349
rect 3605 20349 3617 20352
rect 3651 20380 3663 20383
rect 3970 20380 3976 20392
rect 3651 20352 3976 20380
rect 3651 20349 3663 20352
rect 3605 20343 3663 20349
rect 3970 20340 3976 20352
rect 4028 20340 4034 20392
rect 4065 20383 4123 20389
rect 4065 20349 4077 20383
rect 4111 20380 4123 20383
rect 4338 20380 4344 20392
rect 4111 20352 4344 20380
rect 4111 20349 4123 20352
rect 4065 20343 4123 20349
rect 4338 20340 4344 20352
rect 4396 20340 4402 20392
rect 4706 20340 4712 20392
rect 4764 20380 4770 20392
rect 8110 20380 8116 20392
rect 4764 20352 8116 20380
rect 4764 20340 4770 20352
rect 8110 20340 8116 20352
rect 8168 20340 8174 20392
rect 8588 20324 8616 20411
rect 9582 20408 9588 20420
rect 9640 20408 9646 20460
rect 9784 20457 9812 20488
rect 13078 20476 13084 20528
rect 13136 20476 13142 20528
rect 15102 20516 15108 20528
rect 13832 20488 15108 20516
rect 9769 20451 9827 20457
rect 9769 20417 9781 20451
rect 9815 20417 9827 20451
rect 9769 20411 9827 20417
rect 9858 20408 9864 20460
rect 9916 20448 9922 20460
rect 10505 20451 10563 20457
rect 10505 20448 10517 20451
rect 9916 20420 9961 20448
rect 10060 20420 10517 20448
rect 9916 20408 9922 20420
rect 8662 20340 8668 20392
rect 8720 20380 8726 20392
rect 10060 20380 10088 20420
rect 10505 20417 10517 20420
rect 10551 20417 10563 20451
rect 11054 20448 11060 20460
rect 11015 20420 11060 20448
rect 10505 20411 10563 20417
rect 11054 20408 11060 20420
rect 11112 20408 11118 20460
rect 11238 20408 11244 20460
rect 11296 20448 11302 20460
rect 11701 20451 11759 20457
rect 11701 20448 11713 20451
rect 11296 20420 11713 20448
rect 11296 20408 11302 20420
rect 11701 20417 11713 20420
rect 11747 20417 11759 20451
rect 11701 20411 11759 20417
rect 11974 20408 11980 20460
rect 12032 20448 12038 20460
rect 12250 20448 12256 20460
rect 12032 20420 12256 20448
rect 12032 20408 12038 20420
rect 12250 20408 12256 20420
rect 12308 20448 12314 20460
rect 12713 20451 12771 20457
rect 12713 20448 12725 20451
rect 12308 20420 12725 20448
rect 12308 20408 12314 20420
rect 12713 20417 12725 20420
rect 12759 20417 12771 20451
rect 12713 20411 12771 20417
rect 12802 20408 12808 20460
rect 12860 20448 12866 20460
rect 13096 20448 13124 20476
rect 13630 20448 13636 20460
rect 12860 20420 12905 20448
rect 13096 20420 13636 20448
rect 12860 20408 12866 20420
rect 13630 20408 13636 20420
rect 13688 20448 13694 20460
rect 13725 20451 13783 20457
rect 13725 20448 13737 20451
rect 13688 20420 13737 20448
rect 13688 20408 13694 20420
rect 13725 20417 13737 20420
rect 13771 20417 13783 20451
rect 13725 20411 13783 20417
rect 10226 20380 10232 20392
rect 8720 20352 10088 20380
rect 10187 20352 10232 20380
rect 8720 20340 8726 20352
rect 10226 20340 10232 20352
rect 10284 20340 10290 20392
rect 10410 20380 10416 20392
rect 10371 20352 10416 20380
rect 10410 20340 10416 20352
rect 10468 20340 10474 20392
rect 12437 20383 12495 20389
rect 12437 20349 12449 20383
rect 12483 20380 12495 20383
rect 12526 20380 12532 20392
rect 12483 20352 12532 20380
rect 12483 20349 12495 20352
rect 12437 20343 12495 20349
rect 12526 20340 12532 20352
rect 12584 20340 12590 20392
rect 12986 20340 12992 20392
rect 13044 20380 13050 20392
rect 13081 20383 13139 20389
rect 13081 20380 13093 20383
rect 13044 20352 13093 20380
rect 13044 20340 13050 20352
rect 13081 20349 13093 20352
rect 13127 20349 13139 20383
rect 13832 20380 13860 20488
rect 15102 20476 15108 20488
rect 15160 20476 15166 20528
rect 14274 20408 14280 20460
rect 14332 20448 14338 20460
rect 15013 20451 15071 20457
rect 15013 20448 15025 20451
rect 14332 20420 15025 20448
rect 14332 20408 14338 20420
rect 15013 20417 15025 20420
rect 15059 20417 15071 20451
rect 15013 20411 15071 20417
rect 15194 20408 15200 20460
rect 15252 20408 15258 20460
rect 15396 20457 15424 20556
rect 15488 20556 15945 20584
rect 15381 20451 15439 20457
rect 15381 20417 15393 20451
rect 15427 20417 15439 20451
rect 15381 20411 15439 20417
rect 13081 20343 13139 20349
rect 13740 20352 13860 20380
rect 2682 20312 2688 20324
rect 2424 20284 2688 20312
rect 2682 20272 2688 20284
rect 2740 20272 2746 20324
rect 5718 20272 5724 20324
rect 5776 20312 5782 20324
rect 7745 20315 7803 20321
rect 7745 20312 7757 20315
rect 5776 20284 7757 20312
rect 5776 20272 5782 20284
rect 7745 20281 7757 20284
rect 7791 20281 7803 20315
rect 8570 20312 8576 20324
rect 8483 20284 8576 20312
rect 7745 20275 7803 20281
rect 8570 20272 8576 20284
rect 8628 20312 8634 20324
rect 9398 20312 9404 20324
rect 8628 20284 9404 20312
rect 8628 20272 8634 20284
rect 9398 20272 9404 20284
rect 9456 20272 9462 20324
rect 9674 20272 9680 20324
rect 9732 20312 9738 20324
rect 9858 20312 9864 20324
rect 9732 20284 9864 20312
rect 9732 20272 9738 20284
rect 9858 20272 9864 20284
rect 9916 20312 9922 20324
rect 10778 20312 10784 20324
rect 9916 20284 10784 20312
rect 9916 20272 9922 20284
rect 10778 20272 10784 20284
rect 10836 20272 10842 20324
rect 10873 20315 10931 20321
rect 10873 20281 10885 20315
rect 10919 20312 10931 20315
rect 13740 20312 13768 20352
rect 13906 20340 13912 20392
rect 13964 20380 13970 20392
rect 14458 20380 14464 20392
rect 13964 20352 14464 20380
rect 13964 20340 13970 20352
rect 14458 20340 14464 20352
rect 14516 20340 14522 20392
rect 14645 20383 14703 20389
rect 14645 20349 14657 20383
rect 14691 20380 14703 20383
rect 14734 20380 14740 20392
rect 14691 20352 14740 20380
rect 14691 20349 14703 20352
rect 14645 20343 14703 20349
rect 14734 20340 14740 20352
rect 14792 20340 14798 20392
rect 14826 20340 14832 20392
rect 14884 20380 14890 20392
rect 14921 20383 14979 20389
rect 14921 20380 14933 20383
rect 14884 20352 14933 20380
rect 14884 20340 14890 20352
rect 14921 20349 14933 20352
rect 14967 20349 14979 20383
rect 15212 20380 15240 20408
rect 15488 20380 15516 20556
rect 15933 20553 15945 20556
rect 15979 20553 15991 20587
rect 15933 20547 15991 20553
rect 16022 20544 16028 20596
rect 16080 20584 16086 20596
rect 16853 20587 16911 20593
rect 16853 20584 16865 20587
rect 16080 20556 16865 20584
rect 16080 20544 16086 20556
rect 16853 20553 16865 20556
rect 16899 20553 16911 20587
rect 16853 20547 16911 20553
rect 16942 20544 16948 20596
rect 17000 20584 17006 20596
rect 17589 20587 17647 20593
rect 17589 20584 17601 20587
rect 17000 20556 17601 20584
rect 17000 20544 17006 20556
rect 17589 20553 17601 20556
rect 17635 20553 17647 20587
rect 17589 20547 17647 20553
rect 17954 20544 17960 20596
rect 18012 20584 18018 20596
rect 18601 20587 18659 20593
rect 18601 20584 18613 20587
rect 18012 20556 18613 20584
rect 18012 20544 18018 20556
rect 18601 20553 18613 20556
rect 18647 20553 18659 20587
rect 18601 20547 18659 20553
rect 18690 20544 18696 20596
rect 18748 20584 18754 20596
rect 19429 20587 19487 20593
rect 19429 20584 19441 20587
rect 18748 20556 19441 20584
rect 18748 20544 18754 20556
rect 19429 20553 19441 20556
rect 19475 20553 19487 20587
rect 19429 20547 19487 20553
rect 20070 20544 20076 20596
rect 20128 20584 20134 20596
rect 20809 20587 20867 20593
rect 20809 20584 20821 20587
rect 20128 20556 20821 20584
rect 20128 20544 20134 20556
rect 20809 20553 20821 20556
rect 20855 20553 20867 20587
rect 20809 20547 20867 20553
rect 15562 20476 15568 20528
rect 15620 20516 15626 20528
rect 19058 20516 19064 20528
rect 15620 20488 19064 20516
rect 15620 20476 15626 20488
rect 19058 20476 19064 20488
rect 19116 20476 19122 20528
rect 19444 20488 21128 20516
rect 15654 20408 15660 20460
rect 15712 20448 15718 20460
rect 15749 20451 15807 20457
rect 15749 20448 15761 20451
rect 15712 20420 15761 20448
rect 15712 20408 15718 20420
rect 15749 20417 15761 20420
rect 15795 20417 15807 20451
rect 16114 20448 16120 20460
rect 16075 20420 16120 20448
rect 15749 20411 15807 20417
rect 16114 20408 16120 20420
rect 16172 20408 16178 20460
rect 16206 20408 16212 20460
rect 16264 20448 16270 20460
rect 16669 20451 16727 20457
rect 16669 20448 16681 20451
rect 16264 20420 16681 20448
rect 16264 20408 16270 20420
rect 16669 20417 16681 20420
rect 16715 20417 16727 20451
rect 16669 20411 16727 20417
rect 16850 20408 16856 20460
rect 16908 20448 16914 20460
rect 17037 20451 17095 20457
rect 17037 20448 17049 20451
rect 16908 20420 17049 20448
rect 16908 20408 16914 20420
rect 17037 20417 17049 20420
rect 17083 20417 17095 20451
rect 17402 20448 17408 20460
rect 17363 20420 17408 20448
rect 17037 20411 17095 20417
rect 17402 20408 17408 20420
rect 17460 20408 17466 20460
rect 17770 20448 17776 20460
rect 17731 20420 17776 20448
rect 17770 20408 17776 20420
rect 17828 20408 17834 20460
rect 18138 20448 18144 20460
rect 18099 20420 18144 20448
rect 18138 20408 18144 20420
rect 18196 20408 18202 20460
rect 18785 20451 18843 20457
rect 18785 20417 18797 20451
rect 18831 20448 18843 20451
rect 18874 20448 18880 20460
rect 18831 20420 18880 20448
rect 18831 20417 18843 20420
rect 18785 20411 18843 20417
rect 18874 20408 18880 20420
rect 18932 20408 18938 20460
rect 18966 20408 18972 20460
rect 19024 20448 19030 20460
rect 19245 20451 19303 20457
rect 19245 20448 19257 20451
rect 19024 20420 19257 20448
rect 19024 20408 19030 20420
rect 19245 20417 19257 20420
rect 19291 20417 19303 20451
rect 19245 20411 19303 20417
rect 19444 20380 19472 20488
rect 19610 20448 19616 20460
rect 19571 20420 19616 20448
rect 19610 20408 19616 20420
rect 19668 20408 19674 20460
rect 19978 20448 19984 20460
rect 19939 20420 19984 20448
rect 19978 20408 19984 20420
rect 20036 20408 20042 20460
rect 20346 20448 20352 20460
rect 20307 20420 20352 20448
rect 20346 20408 20352 20420
rect 20404 20408 20410 20460
rect 21100 20457 21128 20488
rect 20993 20451 21051 20457
rect 20993 20417 21005 20451
rect 21039 20417 21051 20451
rect 20993 20411 21051 20417
rect 21085 20451 21143 20457
rect 21085 20417 21097 20451
rect 21131 20417 21143 20451
rect 21085 20411 21143 20417
rect 15212 20352 15516 20380
rect 18984 20352 19472 20380
rect 14921 20343 14979 20349
rect 10919 20284 13768 20312
rect 10919 20281 10931 20284
rect 10873 20275 10931 20281
rect 13814 20272 13820 20324
rect 13872 20312 13878 20324
rect 15197 20315 15255 20321
rect 15197 20312 15209 20315
rect 13872 20284 15209 20312
rect 13872 20272 13878 20284
rect 15197 20281 15209 20284
rect 15243 20281 15255 20315
rect 15197 20275 15255 20281
rect 15286 20272 15292 20324
rect 15344 20312 15350 20324
rect 16301 20315 16359 20321
rect 16301 20312 16313 20315
rect 15344 20284 16313 20312
rect 15344 20272 15350 20284
rect 16301 20281 16313 20284
rect 16347 20281 16359 20315
rect 16301 20275 16359 20281
rect 16574 20272 16580 20324
rect 16632 20312 16638 20324
rect 17221 20315 17279 20321
rect 17221 20312 17233 20315
rect 16632 20284 17233 20312
rect 16632 20272 16638 20284
rect 17221 20281 17233 20284
rect 17267 20281 17279 20315
rect 17221 20275 17279 20281
rect 17494 20272 17500 20324
rect 17552 20312 17558 20324
rect 18325 20315 18383 20321
rect 18325 20312 18337 20315
rect 17552 20284 18337 20312
rect 17552 20272 17558 20284
rect 18325 20281 18337 20284
rect 18371 20281 18383 20315
rect 18325 20275 18383 20281
rect 1486 20244 1492 20256
rect 1447 20216 1492 20244
rect 1486 20204 1492 20216
rect 1544 20204 1550 20256
rect 4890 20244 4896 20256
rect 4851 20216 4896 20244
rect 4890 20204 4896 20216
rect 4948 20204 4954 20256
rect 5258 20204 5264 20256
rect 5316 20244 5322 20256
rect 5353 20247 5411 20253
rect 5353 20244 5365 20247
rect 5316 20216 5365 20244
rect 5316 20204 5322 20216
rect 5353 20213 5365 20216
rect 5399 20213 5411 20247
rect 6822 20244 6828 20256
rect 6783 20216 6828 20244
rect 5353 20207 5411 20213
rect 6822 20204 6828 20216
rect 6880 20204 6886 20256
rect 7101 20247 7159 20253
rect 7101 20213 7113 20247
rect 7147 20244 7159 20247
rect 7190 20244 7196 20256
rect 7147 20216 7196 20244
rect 7147 20213 7159 20216
rect 7101 20207 7159 20213
rect 7190 20204 7196 20216
rect 7248 20204 7254 20256
rect 7377 20247 7435 20253
rect 7377 20213 7389 20247
rect 7423 20244 7435 20247
rect 7466 20244 7472 20256
rect 7423 20216 7472 20244
rect 7423 20213 7435 20216
rect 7377 20207 7435 20213
rect 7466 20204 7472 20216
rect 7524 20204 7530 20256
rect 7650 20244 7656 20256
rect 7611 20216 7656 20244
rect 7650 20204 7656 20216
rect 7708 20204 7714 20256
rect 8202 20244 8208 20256
rect 8163 20216 8208 20244
rect 8202 20204 8208 20216
rect 8260 20204 8266 20256
rect 8294 20204 8300 20256
rect 8352 20244 8358 20256
rect 8352 20216 8397 20244
rect 8352 20204 8358 20216
rect 8478 20204 8484 20256
rect 8536 20244 8542 20256
rect 8757 20247 8815 20253
rect 8757 20244 8769 20247
rect 8536 20216 8769 20244
rect 8536 20204 8542 20216
rect 8757 20213 8769 20216
rect 8803 20213 8815 20247
rect 8757 20207 8815 20213
rect 9217 20247 9275 20253
rect 9217 20213 9229 20247
rect 9263 20244 9275 20247
rect 9306 20244 9312 20256
rect 9263 20216 9312 20244
rect 9263 20213 9275 20216
rect 9217 20207 9275 20213
rect 9306 20204 9312 20216
rect 9364 20204 9370 20256
rect 9490 20204 9496 20256
rect 9548 20244 9554 20256
rect 9585 20247 9643 20253
rect 9585 20244 9597 20247
rect 9548 20216 9597 20244
rect 9548 20204 9554 20216
rect 9585 20213 9597 20216
rect 9631 20213 9643 20247
rect 9585 20207 9643 20213
rect 9950 20204 9956 20256
rect 10008 20244 10014 20256
rect 10045 20247 10103 20253
rect 10045 20244 10057 20247
rect 10008 20216 10057 20244
rect 10008 20204 10014 20216
rect 10045 20213 10057 20216
rect 10091 20213 10103 20247
rect 10045 20207 10103 20213
rect 11517 20247 11575 20253
rect 11517 20213 11529 20247
rect 11563 20244 11575 20247
rect 12158 20244 12164 20256
rect 11563 20216 12164 20244
rect 11563 20213 11575 20216
rect 11517 20207 11575 20213
rect 12158 20204 12164 20216
rect 12216 20204 12222 20256
rect 13906 20244 13912 20256
rect 13867 20216 13912 20244
rect 13906 20204 13912 20216
rect 13964 20204 13970 20256
rect 14182 20204 14188 20256
rect 14240 20244 14246 20256
rect 15565 20247 15623 20253
rect 15565 20244 15577 20247
rect 14240 20216 15577 20244
rect 14240 20204 14246 20216
rect 15565 20213 15577 20216
rect 15611 20213 15623 20247
rect 15565 20207 15623 20213
rect 17126 20204 17132 20256
rect 17184 20244 17190 20256
rect 17957 20247 18015 20253
rect 17957 20244 17969 20247
rect 17184 20216 17969 20244
rect 17184 20204 17190 20216
rect 17957 20213 17969 20216
rect 18003 20213 18015 20247
rect 17957 20207 18015 20213
rect 18690 20204 18696 20256
rect 18748 20244 18754 20256
rect 18984 20253 19012 20352
rect 19702 20340 19708 20392
rect 19760 20380 19766 20392
rect 21008 20380 21036 20411
rect 21358 20408 21364 20460
rect 21416 20448 21422 20460
rect 21453 20451 21511 20457
rect 21453 20448 21465 20451
rect 21416 20420 21465 20448
rect 21416 20408 21422 20420
rect 21453 20417 21465 20420
rect 21499 20417 21511 20451
rect 21453 20411 21511 20417
rect 21376 20380 21404 20408
rect 19760 20352 20576 20380
rect 21008 20352 21404 20380
rect 19760 20340 19766 20352
rect 19334 20272 19340 20324
rect 19392 20312 19398 20324
rect 20548 20321 20576 20352
rect 19797 20315 19855 20321
rect 19797 20312 19809 20315
rect 19392 20284 19809 20312
rect 19392 20272 19398 20284
rect 19797 20281 19809 20284
rect 19843 20281 19855 20315
rect 19797 20275 19855 20281
rect 20533 20315 20591 20321
rect 20533 20281 20545 20315
rect 20579 20281 20591 20315
rect 20533 20275 20591 20281
rect 18969 20247 19027 20253
rect 18969 20244 18981 20247
rect 18748 20216 18981 20244
rect 18748 20204 18754 20216
rect 18969 20213 18981 20216
rect 19015 20213 19027 20247
rect 18969 20207 19027 20213
rect 19426 20204 19432 20256
rect 19484 20244 19490 20256
rect 20165 20247 20223 20253
rect 20165 20244 20177 20247
rect 19484 20216 20177 20244
rect 19484 20204 19490 20216
rect 20165 20213 20177 20216
rect 20211 20213 20223 20247
rect 20165 20207 20223 20213
rect 20438 20204 20444 20256
rect 20496 20244 20502 20256
rect 21269 20247 21327 20253
rect 21269 20244 21281 20247
rect 20496 20216 21281 20244
rect 20496 20204 20502 20216
rect 21269 20213 21281 20216
rect 21315 20213 21327 20247
rect 21269 20207 21327 20213
rect 1104 20154 21896 20176
rect 1104 20102 3549 20154
rect 3601 20102 3613 20154
rect 3665 20102 3677 20154
rect 3729 20102 3741 20154
rect 3793 20102 3805 20154
rect 3857 20102 8747 20154
rect 8799 20102 8811 20154
rect 8863 20102 8875 20154
rect 8927 20102 8939 20154
rect 8991 20102 9003 20154
rect 9055 20102 13945 20154
rect 13997 20102 14009 20154
rect 14061 20102 14073 20154
rect 14125 20102 14137 20154
rect 14189 20102 14201 20154
rect 14253 20102 19143 20154
rect 19195 20102 19207 20154
rect 19259 20102 19271 20154
rect 19323 20102 19335 20154
rect 19387 20102 19399 20154
rect 19451 20102 21896 20154
rect 1104 20080 21896 20102
rect 1854 20040 1860 20052
rect 1815 20012 1860 20040
rect 1854 20000 1860 20012
rect 1912 20000 1918 20052
rect 2225 20043 2283 20049
rect 2225 20009 2237 20043
rect 2271 20040 2283 20043
rect 2774 20040 2780 20052
rect 2271 20012 2780 20040
rect 2271 20009 2283 20012
rect 2225 20003 2283 20009
rect 2774 20000 2780 20012
rect 2832 20000 2838 20052
rect 3050 20040 3056 20052
rect 3011 20012 3056 20040
rect 3050 20000 3056 20012
rect 3108 20000 3114 20052
rect 3234 20000 3240 20052
rect 3292 20040 3298 20052
rect 3510 20040 3516 20052
rect 3292 20012 3516 20040
rect 3292 20000 3298 20012
rect 3510 20000 3516 20012
rect 3568 20000 3574 20052
rect 3605 20043 3663 20049
rect 3605 20009 3617 20043
rect 3651 20040 3663 20043
rect 7098 20040 7104 20052
rect 3651 20012 7104 20040
rect 3651 20009 3663 20012
rect 3605 20003 3663 20009
rect 7098 20000 7104 20012
rect 7156 20000 7162 20052
rect 8389 20043 8447 20049
rect 8389 20009 8401 20043
rect 8435 20040 8447 20043
rect 8662 20040 8668 20052
rect 8435 20012 8668 20040
rect 8435 20009 8447 20012
rect 8389 20003 8447 20009
rect 8662 20000 8668 20012
rect 8720 20000 8726 20052
rect 9677 20043 9735 20049
rect 9677 20009 9689 20043
rect 9723 20040 9735 20043
rect 10410 20040 10416 20052
rect 9723 20012 10416 20040
rect 9723 20009 9735 20012
rect 9677 20003 9735 20009
rect 10410 20000 10416 20012
rect 10468 20000 10474 20052
rect 10594 20040 10600 20052
rect 10555 20012 10600 20040
rect 10594 20000 10600 20012
rect 10652 20000 10658 20052
rect 13633 20043 13691 20049
rect 13633 20009 13645 20043
rect 13679 20040 13691 20043
rect 14274 20040 14280 20052
rect 13679 20012 14280 20040
rect 13679 20009 13691 20012
rect 13633 20003 13691 20009
rect 14274 20000 14280 20012
rect 14332 20000 14338 20052
rect 14550 20000 14556 20052
rect 14608 20040 14614 20052
rect 15105 20043 15163 20049
rect 15105 20040 15117 20043
rect 14608 20012 15117 20040
rect 14608 20000 14614 20012
rect 15105 20009 15117 20012
rect 15151 20009 15163 20043
rect 15105 20003 15163 20009
rect 15746 20000 15752 20052
rect 15804 20040 15810 20052
rect 15841 20043 15899 20049
rect 15841 20040 15853 20043
rect 15804 20012 15853 20040
rect 15804 20000 15810 20012
rect 15841 20009 15853 20012
rect 15887 20009 15899 20043
rect 16850 20040 16856 20052
rect 15841 20003 15899 20009
rect 15948 20012 16712 20040
rect 16811 20012 16856 20040
rect 3421 19975 3479 19981
rect 3421 19941 3433 19975
rect 3467 19941 3479 19975
rect 3421 19935 3479 19941
rect 4157 19975 4215 19981
rect 4157 19941 4169 19975
rect 4203 19972 4215 19975
rect 4706 19972 4712 19984
rect 4203 19944 4712 19972
rect 4203 19941 4215 19944
rect 4157 19935 4215 19941
rect 2777 19907 2835 19913
rect 2777 19873 2789 19907
rect 2823 19904 2835 19907
rect 3436 19904 3464 19935
rect 4706 19932 4712 19944
rect 4764 19932 4770 19984
rect 4801 19975 4859 19981
rect 4801 19941 4813 19975
rect 4847 19941 4859 19975
rect 4801 19935 4859 19941
rect 7377 19975 7435 19981
rect 7377 19941 7389 19975
rect 7423 19972 7435 19975
rect 7558 19972 7564 19984
rect 7423 19944 7564 19972
rect 7423 19941 7435 19944
rect 7377 19935 7435 19941
rect 4816 19904 4844 19935
rect 7558 19932 7564 19944
rect 7616 19932 7622 19984
rect 8478 19932 8484 19984
rect 8536 19972 8542 19984
rect 9398 19972 9404 19984
rect 8536 19944 9404 19972
rect 8536 19932 8542 19944
rect 9398 19932 9404 19944
rect 9456 19932 9462 19984
rect 9582 19932 9588 19984
rect 9640 19972 9646 19984
rect 10134 19972 10140 19984
rect 9640 19944 10140 19972
rect 9640 19932 9646 19944
rect 10134 19932 10140 19944
rect 10192 19932 10198 19984
rect 10505 19975 10563 19981
rect 10505 19941 10517 19975
rect 10551 19972 10563 19975
rect 10870 19972 10876 19984
rect 10551 19944 10876 19972
rect 10551 19941 10563 19944
rect 10505 19935 10563 19941
rect 10870 19932 10876 19944
rect 10928 19932 10934 19984
rect 13909 19975 13967 19981
rect 13909 19941 13921 19975
rect 13955 19972 13967 19975
rect 13955 19944 14964 19972
rect 13955 19941 13967 19944
rect 13909 19935 13967 19941
rect 2823 19876 3372 19904
rect 3436 19876 4752 19904
rect 4816 19876 6132 19904
rect 2823 19873 2835 19876
rect 2777 19867 2835 19873
rect 1673 19839 1731 19845
rect 1673 19805 1685 19839
rect 1719 19805 1731 19839
rect 1673 19799 1731 19805
rect 2041 19839 2099 19845
rect 2041 19805 2053 19839
rect 2087 19836 2099 19839
rect 2222 19836 2228 19848
rect 2087 19808 2228 19836
rect 2087 19805 2099 19808
rect 2041 19799 2099 19805
rect 1688 19768 1716 19799
rect 2222 19796 2228 19808
rect 2280 19796 2286 19848
rect 2409 19839 2467 19845
rect 2409 19805 2421 19839
rect 2455 19805 2467 19839
rect 2409 19799 2467 19805
rect 2314 19768 2320 19780
rect 1688 19740 2320 19768
rect 2314 19728 2320 19740
rect 2372 19728 2378 19780
rect 2424 19768 2452 19799
rect 2498 19796 2504 19848
rect 2556 19836 2562 19848
rect 2593 19839 2651 19845
rect 2593 19836 2605 19839
rect 2556 19808 2605 19836
rect 2556 19796 2562 19808
rect 2593 19805 2605 19808
rect 2639 19805 2651 19839
rect 2866 19836 2872 19848
rect 2827 19808 2872 19836
rect 2593 19799 2651 19805
rect 2866 19796 2872 19808
rect 2924 19796 2930 19848
rect 3142 19796 3148 19848
rect 3200 19836 3206 19848
rect 3237 19839 3295 19845
rect 3237 19836 3249 19839
rect 3200 19808 3249 19836
rect 3200 19796 3206 19808
rect 3237 19805 3249 19808
rect 3283 19805 3295 19839
rect 3237 19799 3295 19805
rect 2424 19740 2774 19768
rect 1486 19700 1492 19712
rect 1447 19672 1492 19700
rect 1486 19660 1492 19672
rect 1544 19660 1550 19712
rect 2746 19700 2774 19740
rect 3234 19700 3240 19712
rect 2746 19672 3240 19700
rect 3234 19660 3240 19672
rect 3292 19660 3298 19712
rect 3344 19700 3372 19876
rect 3878 19796 3884 19848
rect 3936 19836 3942 19848
rect 3973 19839 4031 19845
rect 3973 19836 3985 19839
rect 3936 19808 3985 19836
rect 3936 19796 3942 19808
rect 3973 19805 3985 19808
rect 4019 19805 4031 19839
rect 4246 19836 4252 19848
rect 4207 19808 4252 19836
rect 3973 19799 4031 19805
rect 4246 19796 4252 19808
rect 4304 19796 4310 19848
rect 4614 19836 4620 19848
rect 4575 19808 4620 19836
rect 4614 19796 4620 19808
rect 4672 19796 4678 19848
rect 4724 19836 4752 19876
rect 4982 19836 4988 19848
rect 4724 19808 4844 19836
rect 4943 19808 4988 19836
rect 3789 19771 3847 19777
rect 3789 19737 3801 19771
rect 3835 19768 3847 19771
rect 4706 19768 4712 19780
rect 3835 19740 4712 19768
rect 3835 19737 3847 19740
rect 3789 19731 3847 19737
rect 4706 19728 4712 19740
rect 4764 19728 4770 19780
rect 4154 19700 4160 19712
rect 3344 19672 4160 19700
rect 4154 19660 4160 19672
rect 4212 19660 4218 19712
rect 4430 19700 4436 19712
rect 4391 19672 4436 19700
rect 4430 19660 4436 19672
rect 4488 19660 4494 19712
rect 4816 19700 4844 19808
rect 4982 19796 4988 19808
rect 5040 19796 5046 19848
rect 5721 19839 5779 19845
rect 5721 19805 5733 19839
rect 5767 19836 5779 19839
rect 5994 19836 6000 19848
rect 5767 19808 6000 19836
rect 5767 19805 5779 19808
rect 5721 19799 5779 19805
rect 5994 19796 6000 19808
rect 6052 19796 6058 19848
rect 6104 19836 6132 19876
rect 7282 19864 7288 19916
rect 7340 19904 7346 19916
rect 7469 19907 7527 19913
rect 7469 19904 7481 19907
rect 7340 19876 7481 19904
rect 7340 19864 7346 19876
rect 7469 19873 7481 19876
rect 7515 19873 7527 19907
rect 7469 19867 7527 19873
rect 7837 19907 7895 19913
rect 7837 19873 7849 19907
rect 7883 19904 7895 19907
rect 9033 19907 9091 19913
rect 9033 19904 9045 19907
rect 7883 19876 9045 19904
rect 7883 19873 7895 19876
rect 7837 19867 7895 19873
rect 9033 19873 9045 19876
rect 9079 19904 9091 19907
rect 9766 19904 9772 19916
rect 9079 19876 9772 19904
rect 9079 19873 9091 19876
rect 9033 19867 9091 19873
rect 9766 19864 9772 19876
rect 9824 19864 9830 19916
rect 9953 19907 10011 19913
rect 9953 19873 9965 19907
rect 9999 19904 10011 19907
rect 10042 19904 10048 19916
rect 9999 19876 10048 19904
rect 9999 19873 10011 19876
rect 9953 19867 10011 19873
rect 10042 19864 10048 19876
rect 10100 19864 10106 19916
rect 10226 19864 10232 19916
rect 10284 19904 10290 19916
rect 10778 19904 10784 19916
rect 10284 19876 10784 19904
rect 10284 19864 10290 19876
rect 10778 19864 10784 19876
rect 10836 19864 10842 19916
rect 12066 19864 12072 19916
rect 12124 19904 12130 19916
rect 13354 19904 13360 19916
rect 12124 19876 13360 19904
rect 12124 19864 12130 19876
rect 13354 19864 13360 19876
rect 13412 19904 13418 19916
rect 14645 19907 14703 19913
rect 14645 19904 14657 19907
rect 13412 19876 14657 19904
rect 13412 19864 13418 19876
rect 14645 19873 14657 19876
rect 14691 19873 14703 19907
rect 14645 19867 14703 19873
rect 6104 19808 6776 19836
rect 4890 19728 4896 19780
rect 4948 19768 4954 19780
rect 4948 19740 5580 19768
rect 4948 19728 4954 19740
rect 5166 19700 5172 19712
rect 4816 19672 5172 19700
rect 5166 19660 5172 19672
rect 5224 19660 5230 19712
rect 5552 19700 5580 19740
rect 5626 19728 5632 19780
rect 5684 19768 5690 19780
rect 6242 19771 6300 19777
rect 6242 19768 6254 19771
rect 5684 19740 6254 19768
rect 5684 19728 5690 19740
rect 6242 19737 6254 19740
rect 6288 19737 6300 19771
rect 6748 19768 6776 19808
rect 6822 19796 6828 19848
rect 6880 19836 6886 19848
rect 9674 19836 9680 19848
rect 6880 19808 9680 19836
rect 6880 19796 6886 19808
rect 9674 19796 9680 19808
rect 9732 19796 9738 19848
rect 10318 19836 10324 19848
rect 10060 19808 10324 19836
rect 7742 19768 7748 19780
rect 6748 19740 7748 19768
rect 6242 19731 6300 19737
rect 7742 19728 7748 19740
rect 7800 19728 7806 19780
rect 8021 19771 8079 19777
rect 8021 19737 8033 19771
rect 8067 19768 8079 19771
rect 8481 19771 8539 19777
rect 8481 19768 8493 19771
rect 8067 19740 8493 19768
rect 8067 19737 8079 19740
rect 8021 19731 8079 19737
rect 8481 19737 8493 19740
rect 8527 19737 8539 19771
rect 8481 19731 8539 19737
rect 8938 19728 8944 19780
rect 8996 19768 9002 19780
rect 9309 19771 9367 19777
rect 9309 19768 9321 19771
rect 8996 19740 9321 19768
rect 8996 19728 9002 19740
rect 9309 19737 9321 19740
rect 9355 19737 9367 19771
rect 9309 19731 9367 19737
rect 9398 19728 9404 19780
rect 9456 19768 9462 19780
rect 10060 19768 10088 19808
rect 10318 19796 10324 19808
rect 10376 19796 10382 19848
rect 11882 19796 11888 19848
rect 11940 19836 11946 19848
rect 11977 19839 12035 19845
rect 11977 19836 11989 19839
rect 11940 19808 11989 19836
rect 11940 19796 11946 19808
rect 11977 19805 11989 19808
rect 12023 19805 12035 19839
rect 11977 19799 12035 19805
rect 12434 19796 12440 19848
rect 12492 19836 12498 19848
rect 12618 19836 12624 19848
rect 12492 19808 12624 19836
rect 12492 19796 12498 19808
rect 12618 19796 12624 19808
rect 12676 19796 12682 19848
rect 12710 19796 12716 19848
rect 12768 19836 12774 19848
rect 13446 19836 13452 19848
rect 12768 19808 12813 19836
rect 13407 19808 13452 19836
rect 12768 19796 12774 19808
rect 13446 19796 13452 19808
rect 13504 19796 13510 19848
rect 13538 19796 13544 19848
rect 13596 19836 13602 19848
rect 13725 19839 13783 19845
rect 13725 19836 13737 19839
rect 13596 19808 13737 19836
rect 13596 19796 13602 19808
rect 13725 19805 13737 19808
rect 13771 19805 13783 19839
rect 13725 19799 13783 19805
rect 13814 19796 13820 19848
rect 13872 19836 13878 19848
rect 14826 19836 14832 19848
rect 13872 19808 14832 19836
rect 13872 19796 13878 19808
rect 14826 19796 14832 19808
rect 14884 19796 14890 19848
rect 14936 19845 14964 19944
rect 15194 19932 15200 19984
rect 15252 19972 15258 19984
rect 15948 19972 15976 20012
rect 15252 19944 15976 19972
rect 16577 19975 16635 19981
rect 15252 19932 15258 19944
rect 16577 19941 16589 19975
rect 16623 19941 16635 19975
rect 16684 19972 16712 20012
rect 16850 20000 16856 20012
rect 16908 20000 16914 20052
rect 17402 20040 17408 20052
rect 17363 20012 17408 20040
rect 17402 20000 17408 20012
rect 17460 20000 17466 20052
rect 17770 20040 17776 20052
rect 17731 20012 17776 20040
rect 17770 20000 17776 20012
rect 17828 20000 17834 20052
rect 18230 20000 18236 20052
rect 18288 20040 18294 20052
rect 18417 20043 18475 20049
rect 18417 20040 18429 20043
rect 18288 20012 18429 20040
rect 18288 20000 18294 20012
rect 18417 20009 18429 20012
rect 18463 20009 18475 20043
rect 18874 20040 18880 20052
rect 18835 20012 18880 20040
rect 18417 20003 18475 20009
rect 18874 20000 18880 20012
rect 18932 20000 18938 20052
rect 19886 20040 19892 20052
rect 19847 20012 19892 20040
rect 19886 20000 19892 20012
rect 19944 20000 19950 20052
rect 20254 20040 20260 20052
rect 20215 20012 20260 20040
rect 20254 20000 20260 20012
rect 20312 20000 20318 20052
rect 20806 20000 20812 20052
rect 20864 20040 20870 20052
rect 20993 20043 21051 20049
rect 20993 20040 21005 20043
rect 20864 20012 21005 20040
rect 20864 20000 20870 20012
rect 20993 20009 21005 20012
rect 21039 20009 21051 20043
rect 20993 20003 21051 20009
rect 19429 19975 19487 19981
rect 16684 19944 17540 19972
rect 16577 19935 16635 19941
rect 15010 19864 15016 19916
rect 15068 19904 15074 19916
rect 16114 19904 16120 19916
rect 15068 19876 16120 19904
rect 15068 19864 15074 19876
rect 16114 19864 16120 19876
rect 16172 19864 16178 19916
rect 14921 19839 14979 19845
rect 14921 19805 14933 19839
rect 14967 19805 14979 19839
rect 14921 19799 14979 19805
rect 15286 19796 15292 19848
rect 15344 19836 15350 19848
rect 15473 19839 15531 19845
rect 15473 19836 15485 19839
rect 15344 19808 15485 19836
rect 15344 19796 15350 19808
rect 15473 19805 15485 19808
rect 15519 19805 15531 19839
rect 15473 19799 15531 19805
rect 16025 19839 16083 19845
rect 16025 19805 16037 19839
rect 16071 19805 16083 19839
rect 16298 19836 16304 19848
rect 16259 19808 16304 19836
rect 16025 19799 16083 19805
rect 11790 19777 11796 19780
rect 9456 19740 10088 19768
rect 10137 19771 10195 19777
rect 9456 19728 9462 19740
rect 10137 19737 10149 19771
rect 10183 19768 10195 19771
rect 11732 19771 11796 19777
rect 10183 19740 10732 19768
rect 10183 19737 10195 19740
rect 10137 19731 10195 19737
rect 7006 19700 7012 19712
rect 5552 19672 7012 19700
rect 7006 19660 7012 19672
rect 7064 19660 7070 19712
rect 7374 19660 7380 19712
rect 7432 19700 7438 19712
rect 7929 19703 7987 19709
rect 7929 19700 7941 19703
rect 7432 19672 7941 19700
rect 7432 19660 7438 19672
rect 7929 19669 7941 19672
rect 7975 19669 7987 19703
rect 7929 19663 7987 19669
rect 8110 19660 8116 19712
rect 8168 19700 8174 19712
rect 9030 19700 9036 19712
rect 8168 19672 9036 19700
rect 8168 19660 8174 19672
rect 9030 19660 9036 19672
rect 9088 19700 9094 19712
rect 9217 19703 9275 19709
rect 9217 19700 9229 19703
rect 9088 19672 9229 19700
rect 9088 19660 9094 19672
rect 9217 19669 9229 19672
rect 9263 19669 9275 19703
rect 9217 19663 9275 19669
rect 9674 19660 9680 19712
rect 9732 19700 9738 19712
rect 10045 19703 10103 19709
rect 10045 19700 10057 19703
rect 9732 19672 10057 19700
rect 9732 19660 9738 19672
rect 10045 19669 10057 19672
rect 10091 19669 10103 19703
rect 10704 19700 10732 19740
rect 11732 19737 11744 19771
rect 11778 19737 11796 19771
rect 11732 19731 11796 19737
rect 11790 19728 11796 19731
rect 11848 19728 11854 19780
rect 12342 19728 12348 19780
rect 12400 19768 12406 19780
rect 14461 19771 14519 19777
rect 14461 19768 14473 19771
rect 12400 19740 14473 19768
rect 12400 19728 12406 19740
rect 14461 19737 14473 19740
rect 14507 19768 14519 19771
rect 14844 19768 14872 19796
rect 15565 19771 15623 19777
rect 15565 19768 15577 19771
rect 14507 19740 14780 19768
rect 14844 19740 15577 19768
rect 14507 19737 14519 19740
rect 14461 19731 14519 19737
rect 12069 19703 12127 19709
rect 12069 19700 12081 19703
rect 10704 19672 12081 19700
rect 10045 19663 10103 19669
rect 12069 19669 12081 19672
rect 12115 19669 12127 19703
rect 12069 19663 12127 19669
rect 13170 19660 13176 19712
rect 13228 19700 13234 19712
rect 14093 19703 14151 19709
rect 14093 19700 14105 19703
rect 13228 19672 14105 19700
rect 13228 19660 13234 19672
rect 14093 19669 14105 19672
rect 14139 19669 14151 19703
rect 14093 19663 14151 19669
rect 14550 19660 14556 19712
rect 14608 19700 14614 19712
rect 14752 19700 14780 19740
rect 15565 19737 15577 19740
rect 15611 19737 15623 19771
rect 16040 19768 16068 19799
rect 16298 19796 16304 19808
rect 16356 19796 16362 19848
rect 16390 19796 16396 19848
rect 16448 19836 16454 19848
rect 16592 19836 16620 19935
rect 16669 19839 16727 19845
rect 16669 19836 16681 19839
rect 16448 19808 16493 19836
rect 16592 19808 16681 19836
rect 16448 19796 16454 19808
rect 16669 19805 16681 19808
rect 16715 19805 16727 19839
rect 16669 19799 16727 19805
rect 16942 19796 16948 19848
rect 17000 19836 17006 19848
rect 17129 19839 17187 19845
rect 17129 19836 17141 19839
rect 17000 19808 17141 19836
rect 17000 19796 17006 19808
rect 17129 19805 17141 19808
rect 17175 19805 17187 19839
rect 17129 19799 17187 19805
rect 17218 19796 17224 19848
rect 17276 19836 17282 19848
rect 17512 19845 17540 19944
rect 19429 19941 19441 19975
rect 19475 19941 19487 19975
rect 19429 19935 19487 19941
rect 20717 19975 20775 19981
rect 20717 19941 20729 19975
rect 20763 19972 20775 19975
rect 21174 19972 21180 19984
rect 20763 19944 21180 19972
rect 20763 19941 20775 19944
rect 20717 19935 20775 19941
rect 19444 19904 19472 19935
rect 21174 19932 21180 19944
rect 21232 19932 21238 19984
rect 19444 19876 20576 19904
rect 17497 19839 17555 19845
rect 17276 19808 17321 19836
rect 17276 19796 17282 19808
rect 17497 19805 17509 19839
rect 17543 19805 17555 19839
rect 17957 19839 18015 19845
rect 17957 19836 17969 19839
rect 17497 19799 17555 19805
rect 17696 19808 17969 19836
rect 16040 19740 16988 19768
rect 15565 19731 15623 19737
rect 14826 19700 14832 19712
rect 14608 19672 14653 19700
rect 14752 19672 14832 19700
rect 14608 19660 14614 19672
rect 14826 19660 14832 19672
rect 14884 19660 14890 19712
rect 14918 19660 14924 19712
rect 14976 19700 14982 19712
rect 15289 19703 15347 19709
rect 15289 19700 15301 19703
rect 14976 19672 15301 19700
rect 14976 19660 14982 19672
rect 15289 19669 15301 19672
rect 15335 19669 15347 19703
rect 15289 19663 15347 19669
rect 15746 19660 15752 19712
rect 15804 19700 15810 19712
rect 16960 19709 16988 19740
rect 17696 19709 17724 19808
rect 17957 19805 17969 19808
rect 18003 19805 18015 19839
rect 17957 19799 18015 19805
rect 18046 19796 18052 19848
rect 18104 19836 18110 19848
rect 18598 19836 18604 19848
rect 18104 19808 18149 19836
rect 18559 19808 18604 19836
rect 18104 19796 18110 19808
rect 18598 19796 18604 19808
rect 18656 19796 18662 19848
rect 18693 19839 18751 19845
rect 18693 19805 18705 19839
rect 18739 19805 18751 19839
rect 18693 19799 18751 19805
rect 18708 19768 18736 19799
rect 18782 19796 18788 19848
rect 18840 19836 18846 19848
rect 19245 19839 19303 19845
rect 19245 19836 19257 19839
rect 18840 19808 19257 19836
rect 18840 19796 18846 19808
rect 19245 19805 19257 19808
rect 19291 19805 19303 19839
rect 19245 19799 19303 19805
rect 19521 19839 19579 19845
rect 19521 19805 19533 19839
rect 19567 19836 19579 19839
rect 19702 19836 19708 19848
rect 19567 19808 19708 19836
rect 19567 19805 19579 19808
rect 19521 19799 19579 19805
rect 18248 19740 18736 19768
rect 19061 19771 19119 19777
rect 18248 19709 18276 19740
rect 19061 19737 19073 19771
rect 19107 19768 19119 19771
rect 19536 19768 19564 19799
rect 19702 19796 19708 19808
rect 19760 19796 19766 19848
rect 20073 19839 20131 19845
rect 20073 19805 20085 19839
rect 20119 19836 20131 19839
rect 20254 19836 20260 19848
rect 20119 19808 20260 19836
rect 20119 19805 20131 19808
rect 20073 19799 20131 19805
rect 20254 19796 20260 19808
rect 20312 19796 20318 19848
rect 20548 19845 20576 19876
rect 20441 19839 20499 19845
rect 20441 19805 20453 19839
rect 20487 19805 20499 19839
rect 20441 19799 20499 19805
rect 20533 19839 20591 19845
rect 20533 19805 20545 19839
rect 20579 19805 20591 19839
rect 20533 19799 20591 19805
rect 19107 19740 19564 19768
rect 20456 19768 20484 19799
rect 20990 19796 20996 19848
rect 21048 19836 21054 19848
rect 21177 19839 21235 19845
rect 21177 19836 21189 19839
rect 21048 19808 21189 19836
rect 21048 19796 21054 19808
rect 21177 19805 21189 19808
rect 21223 19805 21235 19839
rect 21177 19799 21235 19805
rect 21269 19839 21327 19845
rect 21269 19805 21281 19839
rect 21315 19805 21327 19839
rect 21269 19799 21327 19805
rect 20714 19768 20720 19780
rect 20456 19740 20720 19768
rect 19107 19737 19119 19740
rect 19061 19731 19119 19737
rect 20714 19728 20720 19740
rect 20772 19728 20778 19780
rect 16117 19703 16175 19709
rect 16117 19700 16129 19703
rect 15804 19672 16129 19700
rect 15804 19660 15810 19672
rect 16117 19669 16129 19672
rect 16163 19669 16175 19703
rect 16117 19663 16175 19669
rect 16945 19703 17003 19709
rect 16945 19669 16957 19703
rect 16991 19669 17003 19703
rect 16945 19663 17003 19669
rect 17681 19703 17739 19709
rect 17681 19669 17693 19703
rect 17727 19669 17739 19703
rect 17681 19663 17739 19669
rect 18233 19703 18291 19709
rect 18233 19669 18245 19703
rect 18279 19669 18291 19703
rect 18233 19663 18291 19669
rect 19705 19703 19763 19709
rect 19705 19669 19717 19703
rect 19751 19700 19763 19703
rect 19794 19700 19800 19712
rect 19751 19672 19800 19700
rect 19751 19669 19763 19672
rect 19705 19663 19763 19669
rect 19794 19660 19800 19672
rect 19852 19660 19858 19712
rect 20162 19660 20168 19712
rect 20220 19700 20226 19712
rect 21284 19700 21312 19799
rect 21450 19700 21456 19712
rect 20220 19672 21312 19700
rect 21411 19672 21456 19700
rect 20220 19660 20226 19672
rect 21450 19660 21456 19672
rect 21508 19660 21514 19712
rect 1104 19610 22056 19632
rect 1104 19558 6148 19610
rect 6200 19558 6212 19610
rect 6264 19558 6276 19610
rect 6328 19558 6340 19610
rect 6392 19558 6404 19610
rect 6456 19558 11346 19610
rect 11398 19558 11410 19610
rect 11462 19558 11474 19610
rect 11526 19558 11538 19610
rect 11590 19558 11602 19610
rect 11654 19558 16544 19610
rect 16596 19558 16608 19610
rect 16660 19558 16672 19610
rect 16724 19558 16736 19610
rect 16788 19558 16800 19610
rect 16852 19558 21742 19610
rect 21794 19558 21806 19610
rect 21858 19558 21870 19610
rect 21922 19558 21934 19610
rect 21986 19558 21998 19610
rect 22050 19558 22056 19610
rect 1104 19536 22056 19558
rect 2133 19499 2191 19505
rect 2133 19465 2145 19499
rect 2179 19465 2191 19499
rect 2133 19459 2191 19465
rect 2148 19428 2176 19459
rect 2314 19456 2320 19508
rect 2372 19496 2378 19508
rect 2409 19499 2467 19505
rect 2409 19496 2421 19499
rect 2372 19468 2421 19496
rect 2372 19456 2378 19468
rect 2409 19465 2421 19468
rect 2455 19465 2467 19499
rect 2866 19496 2872 19508
rect 2827 19468 2872 19496
rect 2409 19459 2467 19465
rect 2866 19456 2872 19468
rect 2924 19456 2930 19508
rect 2961 19499 3019 19505
rect 2961 19465 2973 19499
rect 3007 19465 3019 19499
rect 3234 19496 3240 19508
rect 3195 19468 3240 19496
rect 2961 19459 3019 19465
rect 1688 19400 2176 19428
rect 1688 19369 1716 19400
rect 2222 19388 2228 19440
rect 2280 19428 2286 19440
rect 2976 19428 3004 19459
rect 3234 19456 3240 19468
rect 3292 19456 3298 19508
rect 3326 19456 3332 19508
rect 3384 19496 3390 19508
rect 3697 19499 3755 19505
rect 3697 19496 3709 19499
rect 3384 19468 3709 19496
rect 3384 19456 3390 19468
rect 3697 19465 3709 19468
rect 3743 19465 3755 19499
rect 3970 19496 3976 19508
rect 3931 19468 3976 19496
rect 3697 19459 3755 19465
rect 3970 19456 3976 19468
rect 4028 19456 4034 19508
rect 4341 19499 4399 19505
rect 4341 19465 4353 19499
rect 4387 19496 4399 19499
rect 4982 19496 4988 19508
rect 4387 19468 4988 19496
rect 4387 19465 4399 19468
rect 4341 19459 4399 19465
rect 4982 19456 4988 19468
rect 5040 19456 5046 19508
rect 5074 19456 5080 19508
rect 5132 19496 5138 19508
rect 7926 19496 7932 19508
rect 5132 19468 7932 19496
rect 5132 19456 5138 19468
rect 7926 19456 7932 19468
rect 7984 19456 7990 19508
rect 8478 19456 8484 19508
rect 8536 19496 8542 19508
rect 9214 19496 9220 19508
rect 8536 19468 9220 19496
rect 8536 19456 8542 19468
rect 9214 19456 9220 19468
rect 9272 19456 9278 19508
rect 9674 19456 9680 19508
rect 9732 19496 9738 19508
rect 12342 19496 12348 19508
rect 9732 19468 12348 19496
rect 9732 19456 9738 19468
rect 12342 19456 12348 19468
rect 12400 19456 12406 19508
rect 12618 19496 12624 19508
rect 12579 19468 12624 19496
rect 12618 19456 12624 19468
rect 12676 19456 12682 19508
rect 12802 19496 12808 19508
rect 12763 19468 12808 19496
rect 12802 19456 12808 19468
rect 12860 19456 12866 19508
rect 13354 19496 13360 19508
rect 13315 19468 13360 19496
rect 13354 19456 13360 19468
rect 13412 19456 13418 19508
rect 15010 19496 15016 19508
rect 14971 19468 15016 19496
rect 15010 19456 15016 19468
rect 15068 19456 15074 19508
rect 15381 19499 15439 19505
rect 15381 19465 15393 19499
rect 15427 19465 15439 19499
rect 15654 19496 15660 19508
rect 15615 19468 15660 19496
rect 15381 19459 15439 19465
rect 2280 19400 3004 19428
rect 2280 19388 2286 19400
rect 3050 19388 3056 19440
rect 3108 19428 3114 19440
rect 5813 19431 5871 19437
rect 5813 19428 5825 19431
rect 3108 19400 3556 19428
rect 3108 19388 3114 19400
rect 1673 19363 1731 19369
rect 1673 19329 1685 19363
rect 1719 19329 1731 19363
rect 2038 19360 2044 19372
rect 1999 19332 2044 19360
rect 1673 19323 1731 19329
rect 2038 19320 2044 19332
rect 2096 19320 2102 19372
rect 2314 19360 2320 19372
rect 2227 19332 2320 19360
rect 2314 19320 2320 19332
rect 2372 19360 2378 19372
rect 2593 19363 2651 19369
rect 2372 19332 2544 19360
rect 2372 19320 2378 19332
rect 1854 19224 1860 19236
rect 1815 19196 1860 19224
rect 1854 19184 1860 19196
rect 1912 19184 1918 19236
rect 1486 19156 1492 19168
rect 1447 19128 1492 19156
rect 1486 19116 1492 19128
rect 1544 19116 1550 19168
rect 2516 19156 2544 19332
rect 2593 19329 2605 19363
rect 2639 19329 2651 19363
rect 2593 19323 2651 19329
rect 2685 19363 2743 19369
rect 2685 19329 2697 19363
rect 2731 19360 2743 19363
rect 2958 19360 2964 19372
rect 2731 19332 2964 19360
rect 2731 19329 2743 19332
rect 2685 19323 2743 19329
rect 2608 19292 2636 19323
rect 2958 19320 2964 19332
rect 3016 19320 3022 19372
rect 3145 19363 3203 19369
rect 3145 19329 3157 19363
rect 3191 19360 3203 19363
rect 3234 19360 3240 19372
rect 3191 19332 3240 19360
rect 3191 19329 3203 19332
rect 3145 19323 3203 19329
rect 3234 19320 3240 19332
rect 3292 19320 3298 19372
rect 3326 19320 3332 19372
rect 3384 19360 3390 19372
rect 3528 19369 3556 19400
rect 3620 19400 5825 19428
rect 3421 19363 3479 19369
rect 3421 19360 3433 19363
rect 3384 19332 3433 19360
rect 3384 19320 3390 19332
rect 3421 19329 3433 19332
rect 3467 19329 3479 19363
rect 3421 19323 3479 19329
rect 3513 19363 3571 19369
rect 3513 19329 3525 19363
rect 3559 19329 3571 19363
rect 3513 19323 3571 19329
rect 2866 19292 2872 19304
rect 2608 19264 2872 19292
rect 2866 19252 2872 19264
rect 2924 19252 2930 19304
rect 3620 19292 3648 19400
rect 5813 19397 5825 19400
rect 5859 19428 5871 19431
rect 5902 19428 5908 19440
rect 5859 19400 5908 19428
rect 5859 19397 5871 19400
rect 5813 19391 5871 19397
rect 5902 19388 5908 19400
rect 5960 19388 5966 19440
rect 7098 19388 7104 19440
rect 7156 19428 7162 19440
rect 7156 19400 7788 19428
rect 7156 19388 7162 19400
rect 3786 19360 3792 19372
rect 3747 19332 3792 19360
rect 3786 19320 3792 19332
rect 3844 19320 3850 19372
rect 3970 19320 3976 19372
rect 4028 19360 4034 19372
rect 4985 19363 5043 19369
rect 4985 19360 4997 19363
rect 4028 19332 4997 19360
rect 4028 19320 4034 19332
rect 4985 19329 4997 19332
rect 5031 19329 5043 19363
rect 4985 19323 5043 19329
rect 5166 19320 5172 19372
rect 5224 19360 5230 19372
rect 5721 19363 5779 19369
rect 5721 19360 5733 19363
rect 5224 19332 5733 19360
rect 5224 19320 5230 19332
rect 5721 19329 5733 19332
rect 5767 19360 5779 19363
rect 6730 19360 6736 19372
rect 5767 19332 6736 19360
rect 5767 19329 5779 19332
rect 5721 19323 5779 19329
rect 6730 19320 6736 19332
rect 6788 19320 6794 19372
rect 7558 19320 7564 19372
rect 7616 19369 7622 19372
rect 7616 19360 7628 19369
rect 7760 19364 7788 19400
rect 8294 19388 8300 19440
rect 8352 19428 8358 19440
rect 11882 19428 11888 19440
rect 8352 19400 11888 19428
rect 8352 19388 8358 19400
rect 7837 19364 7895 19369
rect 7760 19363 7895 19364
rect 7616 19332 7661 19360
rect 7760 19336 7849 19363
rect 7616 19323 7628 19332
rect 7837 19329 7849 19336
rect 7883 19329 7895 19363
rect 7837 19323 7895 19329
rect 7929 19367 7987 19373
rect 7929 19333 7941 19367
rect 7975 19333 7987 19367
rect 7929 19327 7987 19333
rect 7616 19320 7622 19323
rect 3528 19264 3648 19292
rect 3528 19224 3556 19264
rect 4154 19252 4160 19304
rect 4212 19292 4218 19304
rect 4338 19292 4344 19304
rect 4212 19264 4344 19292
rect 4212 19252 4218 19264
rect 4338 19252 4344 19264
rect 4396 19252 4402 19304
rect 4706 19292 4712 19304
rect 4667 19264 4712 19292
rect 4706 19252 4712 19264
rect 4764 19252 4770 19304
rect 4890 19292 4896 19304
rect 4851 19264 4896 19292
rect 4890 19252 4896 19264
rect 4948 19252 4954 19304
rect 5626 19292 5632 19304
rect 5587 19264 5632 19292
rect 5626 19252 5632 19264
rect 5684 19252 5690 19304
rect 7944 19292 7972 19327
rect 8110 19320 8116 19372
rect 8168 19344 8174 19372
rect 8404 19369 8432 19400
rect 8662 19369 8668 19372
rect 8389 19363 8447 19369
rect 8168 19320 8294 19344
rect 8389 19329 8401 19363
rect 8435 19360 8447 19363
rect 8435 19332 8469 19360
rect 8435 19329 8447 19332
rect 8389 19323 8447 19329
rect 8656 19323 8668 19369
rect 8720 19360 8726 19372
rect 8720 19332 8756 19360
rect 8662 19320 8668 19323
rect 8720 19320 8726 19332
rect 9030 19320 9036 19372
rect 9088 19360 9094 19372
rect 9968 19369 9996 19400
rect 11882 19388 11888 19400
rect 11940 19388 11946 19440
rect 15396 19428 15424 19459
rect 15654 19456 15660 19468
rect 15712 19456 15718 19508
rect 15933 19499 15991 19505
rect 15933 19465 15945 19499
rect 15979 19496 15991 19499
rect 16206 19496 16212 19508
rect 15979 19468 16212 19496
rect 15979 19465 15991 19468
rect 15933 19459 15991 19465
rect 16206 19456 16212 19468
rect 16264 19456 16270 19508
rect 16485 19499 16543 19505
rect 16485 19465 16497 19499
rect 16531 19496 16543 19499
rect 17218 19496 17224 19508
rect 16531 19468 17224 19496
rect 16531 19465 16543 19468
rect 16485 19459 16543 19465
rect 17218 19456 17224 19468
rect 17276 19456 17282 19508
rect 17497 19499 17555 19505
rect 17497 19465 17509 19499
rect 17543 19465 17555 19499
rect 18138 19496 18144 19508
rect 18099 19468 18144 19496
rect 17497 19459 17555 19465
rect 13740 19400 15056 19428
rect 15396 19400 15792 19428
rect 9953 19363 10011 19369
rect 9088 19344 9444 19360
rect 9499 19344 9619 19360
rect 9088 19332 9619 19344
rect 9088 19320 9094 19332
rect 8128 19316 8294 19320
rect 9416 19316 9527 19332
rect 7852 19264 7972 19292
rect 2746 19196 3556 19224
rect 2746 19156 2774 19196
rect 3602 19184 3608 19236
rect 3660 19224 3666 19236
rect 4525 19227 4583 19233
rect 3660 19196 4476 19224
rect 3660 19184 3666 19196
rect 4154 19156 4160 19168
rect 2516 19128 2774 19156
rect 4115 19128 4160 19156
rect 4154 19116 4160 19128
rect 4212 19116 4218 19168
rect 4448 19156 4476 19196
rect 4525 19193 4537 19227
rect 4571 19224 4583 19227
rect 5994 19224 6000 19236
rect 4571 19196 6000 19224
rect 4571 19193 4583 19196
rect 4525 19187 4583 19193
rect 5994 19184 6000 19196
rect 6052 19184 6058 19236
rect 6457 19227 6515 19233
rect 6457 19193 6469 19227
rect 6503 19224 6515 19227
rect 6638 19224 6644 19236
rect 6503 19196 6644 19224
rect 6503 19193 6515 19196
rect 6457 19187 6515 19193
rect 6638 19184 6644 19196
rect 6696 19184 6702 19236
rect 4798 19156 4804 19168
rect 4448 19128 4804 19156
rect 4798 19116 4804 19128
rect 4856 19116 4862 19168
rect 5350 19156 5356 19168
rect 5311 19128 5356 19156
rect 5350 19116 5356 19128
rect 5408 19116 5414 19168
rect 6178 19156 6184 19168
rect 6139 19128 6184 19156
rect 6178 19116 6184 19128
rect 6236 19116 6242 19168
rect 6546 19116 6552 19168
rect 6604 19156 6610 19168
rect 7852 19156 7880 19264
rect 7926 19156 7932 19168
rect 6604 19128 7932 19156
rect 6604 19116 6610 19128
rect 7926 19116 7932 19128
rect 7984 19116 7990 19168
rect 8110 19156 8116 19168
rect 8071 19128 8116 19156
rect 8110 19116 8116 19128
rect 8168 19116 8174 19168
rect 8266 19156 8294 19316
rect 9591 19292 9619 19332
rect 9953 19329 9965 19363
rect 9999 19329 10011 19363
rect 9953 19323 10011 19329
rect 10042 19320 10048 19372
rect 10100 19360 10106 19372
rect 10220 19363 10278 19369
rect 10220 19360 10232 19363
rect 10100 19332 10232 19360
rect 10100 19320 10106 19332
rect 10220 19329 10232 19332
rect 10266 19360 10278 19363
rect 11974 19360 11980 19372
rect 10266 19332 11836 19360
rect 11935 19332 11980 19360
rect 10266 19329 10278 19332
rect 10220 19323 10278 19329
rect 11609 19295 11667 19301
rect 9591 19264 9996 19292
rect 9766 19184 9772 19236
rect 9824 19224 9830 19236
rect 9824 19196 9869 19224
rect 9824 19184 9830 19196
rect 9674 19156 9680 19168
rect 8266 19128 9680 19156
rect 9674 19116 9680 19128
rect 9732 19116 9738 19168
rect 9968 19156 9996 19264
rect 11609 19261 11621 19295
rect 11655 19292 11667 19295
rect 11698 19292 11704 19304
rect 11655 19264 11704 19292
rect 11655 19261 11667 19264
rect 11609 19255 11667 19261
rect 11698 19252 11704 19264
rect 11756 19252 11762 19304
rect 11808 19292 11836 19332
rect 11974 19320 11980 19332
rect 12032 19320 12038 19372
rect 12066 19320 12072 19372
rect 12124 19360 12130 19372
rect 12124 19332 12204 19360
rect 12124 19320 12130 19332
rect 12176 19292 12204 19332
rect 11808 19264 12204 19292
rect 12250 19252 12256 19304
rect 12308 19292 12314 19304
rect 12989 19295 13047 19301
rect 12989 19292 13001 19295
rect 12308 19264 13001 19292
rect 12308 19252 12314 19264
rect 12989 19261 13001 19264
rect 13035 19261 13047 19295
rect 12989 19255 13047 19261
rect 10962 19184 10968 19236
rect 11020 19224 11026 19236
rect 13740 19224 13768 19400
rect 14458 19320 14464 19372
rect 14516 19369 14522 19372
rect 14516 19360 14528 19369
rect 14829 19364 14887 19369
rect 14918 19364 14924 19372
rect 14829 19363 14924 19364
rect 14516 19332 14561 19360
rect 14516 19323 14528 19332
rect 14829 19329 14841 19363
rect 14875 19336 14924 19363
rect 14875 19329 14887 19336
rect 14829 19323 14887 19329
rect 14516 19320 14522 19323
rect 14918 19320 14924 19336
rect 14976 19320 14982 19372
rect 14737 19295 14795 19301
rect 14737 19261 14749 19295
rect 14783 19261 14795 19295
rect 15028 19292 15056 19400
rect 15194 19360 15200 19372
rect 15155 19332 15200 19360
rect 15194 19320 15200 19332
rect 15252 19320 15258 19372
rect 15473 19363 15531 19369
rect 15473 19329 15485 19363
rect 15519 19360 15531 19363
rect 15654 19360 15660 19372
rect 15519 19332 15660 19360
rect 15519 19329 15531 19332
rect 15473 19323 15531 19329
rect 15654 19320 15660 19332
rect 15712 19320 15718 19372
rect 15764 19369 15792 19400
rect 15749 19363 15807 19369
rect 15749 19329 15761 19363
rect 15795 19329 15807 19363
rect 15749 19323 15807 19329
rect 15838 19320 15844 19372
rect 15896 19360 15902 19372
rect 16301 19363 16359 19369
rect 16301 19360 16313 19363
rect 15896 19332 16313 19360
rect 15896 19320 15902 19332
rect 16301 19329 16313 19332
rect 16347 19329 16359 19363
rect 17126 19360 17132 19372
rect 17087 19332 17132 19360
rect 16301 19323 16359 19329
rect 17126 19320 17132 19332
rect 17184 19320 17190 19372
rect 17512 19360 17540 19459
rect 18138 19456 18144 19468
rect 18196 19456 18202 19508
rect 18598 19496 18604 19508
rect 18559 19468 18604 19496
rect 18598 19456 18604 19468
rect 18656 19456 18662 19508
rect 18877 19499 18935 19505
rect 18877 19465 18889 19499
rect 18923 19496 18935 19499
rect 18966 19496 18972 19508
rect 18923 19468 18972 19496
rect 18923 19465 18935 19468
rect 18877 19459 18935 19465
rect 18966 19456 18972 19468
rect 19024 19456 19030 19508
rect 19058 19456 19064 19508
rect 19116 19496 19122 19508
rect 19337 19499 19395 19505
rect 19337 19496 19349 19499
rect 19116 19468 19349 19496
rect 19116 19456 19122 19468
rect 19337 19465 19349 19468
rect 19383 19496 19395 19499
rect 19978 19496 19984 19508
rect 19383 19468 19984 19496
rect 19383 19465 19395 19468
rect 19337 19459 19395 19465
rect 19978 19456 19984 19468
rect 20036 19456 20042 19508
rect 20254 19496 20260 19508
rect 20215 19468 20260 19496
rect 20254 19456 20260 19468
rect 20312 19456 20318 19508
rect 20717 19499 20775 19505
rect 20717 19465 20729 19499
rect 20763 19496 20775 19499
rect 20898 19496 20904 19508
rect 20763 19468 20904 19496
rect 20763 19465 20775 19468
rect 20717 19459 20775 19465
rect 20898 19456 20904 19468
rect 20956 19456 20962 19508
rect 21082 19496 21088 19508
rect 21043 19468 21088 19496
rect 21082 19456 21088 19468
rect 21140 19456 21146 19508
rect 17773 19431 17831 19437
rect 17773 19397 17785 19431
rect 17819 19428 17831 19431
rect 17954 19428 17960 19440
rect 17819 19400 17960 19428
rect 17819 19397 17831 19400
rect 17773 19391 17831 19397
rect 17954 19388 17960 19400
rect 18012 19388 18018 19440
rect 19794 19388 19800 19440
rect 19852 19428 19858 19440
rect 19852 19400 20576 19428
rect 19852 19388 19858 19400
rect 17865 19363 17923 19369
rect 17865 19360 17877 19363
rect 17512 19332 17877 19360
rect 17865 19329 17877 19332
rect 17911 19329 17923 19363
rect 18325 19363 18383 19369
rect 18325 19360 18337 19363
rect 17865 19323 17923 19329
rect 18064 19332 18337 19360
rect 16390 19292 16396 19304
rect 15028 19264 16396 19292
rect 14737 19255 14795 19261
rect 11020 19196 13768 19224
rect 11020 19184 11026 19196
rect 11146 19156 11152 19168
rect 9968 19128 11152 19156
rect 11146 19116 11152 19128
rect 11204 19116 11210 19168
rect 11333 19159 11391 19165
rect 11333 19125 11345 19159
rect 11379 19156 11391 19159
rect 11790 19156 11796 19168
rect 11379 19128 11796 19156
rect 11379 19125 11391 19128
rect 11333 19119 11391 19125
rect 11790 19116 11796 19128
rect 11848 19116 11854 19168
rect 13265 19159 13323 19165
rect 13265 19125 13277 19159
rect 13311 19156 13323 19159
rect 14366 19156 14372 19168
rect 13311 19128 14372 19156
rect 13311 19125 13323 19128
rect 13265 19119 13323 19125
rect 14366 19116 14372 19128
rect 14424 19156 14430 19168
rect 14752 19156 14780 19255
rect 16390 19252 16396 19264
rect 16448 19252 16454 19304
rect 16850 19292 16856 19304
rect 16811 19264 16856 19292
rect 16850 19252 16856 19264
rect 16908 19252 16914 19304
rect 17034 19292 17040 19304
rect 16995 19264 17040 19292
rect 17034 19252 17040 19264
rect 17092 19252 17098 19304
rect 14826 19184 14832 19236
rect 14884 19224 14890 19236
rect 16022 19224 16028 19236
rect 14884 19196 16028 19224
rect 14884 19184 14890 19196
rect 16022 19184 16028 19196
rect 16080 19184 16086 19236
rect 18064 19233 18092 19332
rect 18325 19329 18337 19332
rect 18371 19329 18383 19363
rect 18325 19323 18383 19329
rect 18414 19320 18420 19372
rect 18472 19360 18478 19372
rect 18693 19363 18751 19369
rect 18472 19332 18517 19360
rect 18472 19320 18478 19332
rect 18693 19329 18705 19363
rect 18739 19360 18751 19363
rect 18874 19360 18880 19372
rect 18739 19332 18880 19360
rect 18739 19329 18751 19332
rect 18693 19323 18751 19329
rect 18874 19320 18880 19332
rect 18932 19360 18938 19372
rect 18969 19363 19027 19369
rect 18969 19360 18981 19363
rect 18932 19332 18981 19360
rect 18932 19320 18938 19332
rect 18969 19329 18981 19332
rect 19015 19329 19027 19363
rect 18969 19323 19027 19329
rect 19518 19320 19524 19372
rect 19576 19360 19582 19372
rect 19705 19363 19763 19369
rect 19705 19360 19717 19363
rect 19576 19332 19717 19360
rect 19576 19320 19582 19332
rect 19705 19329 19717 19332
rect 19751 19329 19763 19363
rect 19978 19360 19984 19372
rect 19939 19332 19984 19360
rect 19705 19323 19763 19329
rect 19978 19320 19984 19332
rect 20036 19320 20042 19372
rect 20548 19369 20576 19400
rect 20441 19363 20499 19369
rect 20441 19329 20453 19363
rect 20487 19329 20499 19363
rect 20441 19323 20499 19329
rect 20533 19363 20591 19369
rect 20533 19329 20545 19363
rect 20579 19329 20591 19363
rect 20898 19360 20904 19372
rect 20859 19332 20904 19360
rect 20533 19323 20591 19329
rect 18230 19252 18236 19304
rect 18288 19292 18294 19304
rect 19153 19295 19211 19301
rect 19153 19292 19165 19295
rect 18288 19264 19165 19292
rect 18288 19252 18294 19264
rect 19153 19261 19165 19264
rect 19199 19292 19211 19295
rect 20456 19292 20484 19323
rect 20898 19320 20904 19332
rect 20956 19320 20962 19372
rect 21266 19360 21272 19372
rect 21227 19332 21272 19360
rect 21266 19320 21272 19332
rect 21324 19320 21330 19372
rect 19199 19264 20484 19292
rect 19199 19261 19211 19264
rect 19153 19255 19211 19261
rect 18049 19227 18107 19233
rect 18049 19193 18061 19227
rect 18095 19193 18107 19227
rect 18049 19187 18107 19193
rect 18138 19184 18144 19236
rect 18196 19224 18202 19236
rect 19518 19224 19524 19236
rect 18196 19196 19524 19224
rect 18196 19184 18202 19196
rect 19518 19184 19524 19196
rect 19576 19184 19582 19236
rect 19889 19227 19947 19233
rect 19889 19193 19901 19227
rect 19935 19224 19947 19227
rect 20806 19224 20812 19236
rect 19935 19196 20812 19224
rect 19935 19193 19947 19196
rect 19889 19187 19947 19193
rect 20806 19184 20812 19196
rect 20864 19184 20870 19236
rect 20162 19156 20168 19168
rect 14424 19128 14780 19156
rect 20123 19128 20168 19156
rect 14424 19116 14430 19128
rect 20162 19116 20168 19128
rect 20220 19116 20226 19168
rect 21450 19156 21456 19168
rect 21411 19128 21456 19156
rect 21450 19116 21456 19128
rect 21508 19116 21514 19168
rect 1104 19066 21896 19088
rect 1104 19014 3549 19066
rect 3601 19014 3613 19066
rect 3665 19014 3677 19066
rect 3729 19014 3741 19066
rect 3793 19014 3805 19066
rect 3857 19014 8747 19066
rect 8799 19014 8811 19066
rect 8863 19014 8875 19066
rect 8927 19014 8939 19066
rect 8991 19014 9003 19066
rect 9055 19014 13945 19066
rect 13997 19014 14009 19066
rect 14061 19014 14073 19066
rect 14125 19014 14137 19066
rect 14189 19014 14201 19066
rect 14253 19014 19143 19066
rect 19195 19014 19207 19066
rect 19259 19014 19271 19066
rect 19323 19014 19335 19066
rect 19387 19014 19399 19066
rect 19451 19014 21896 19066
rect 1104 18992 21896 19014
rect 1949 18955 2007 18961
rect 1949 18921 1961 18955
rect 1995 18952 2007 18955
rect 2038 18952 2044 18964
rect 1995 18924 2044 18952
rect 1995 18921 2007 18924
rect 1949 18915 2007 18921
rect 2038 18912 2044 18924
rect 2096 18912 2102 18964
rect 2406 18912 2412 18964
rect 2464 18952 2470 18964
rect 2961 18955 3019 18961
rect 2464 18924 2636 18952
rect 2464 18912 2470 18924
rect 1854 18844 1860 18896
rect 1912 18884 1918 18896
rect 1912 18856 2544 18884
rect 1912 18844 1918 18856
rect 1762 18776 1768 18828
rect 1820 18816 1826 18828
rect 2406 18816 2412 18828
rect 1820 18788 2268 18816
rect 2367 18788 2412 18816
rect 1820 18776 1826 18788
rect 1673 18751 1731 18757
rect 1673 18717 1685 18751
rect 1719 18748 1731 18751
rect 2038 18748 2044 18760
rect 1719 18720 2044 18748
rect 1719 18717 1731 18720
rect 1673 18711 1731 18717
rect 2038 18708 2044 18720
rect 2096 18708 2102 18760
rect 2133 18751 2191 18757
rect 2133 18717 2145 18751
rect 2179 18717 2191 18751
rect 2240 18748 2268 18788
rect 2406 18776 2412 18788
rect 2464 18776 2470 18828
rect 2516 18825 2544 18856
rect 2501 18819 2559 18825
rect 2501 18785 2513 18819
rect 2547 18785 2559 18819
rect 2608 18816 2636 18924
rect 2961 18921 2973 18955
rect 3007 18952 3019 18955
rect 3970 18952 3976 18964
rect 3007 18924 3976 18952
rect 3007 18921 3019 18924
rect 2961 18915 3019 18921
rect 3970 18912 3976 18924
rect 4028 18912 4034 18964
rect 4890 18952 4896 18964
rect 4851 18924 4896 18952
rect 4890 18912 4896 18924
rect 4948 18912 4954 18964
rect 6638 18952 6644 18964
rect 5184 18924 6644 18952
rect 2682 18844 2688 18896
rect 2740 18884 2746 18896
rect 3234 18884 3240 18896
rect 2740 18856 3240 18884
rect 2740 18844 2746 18856
rect 3234 18844 3240 18856
rect 3292 18844 3298 18896
rect 3326 18844 3332 18896
rect 3384 18884 3390 18896
rect 4065 18887 4123 18893
rect 4065 18884 4077 18887
rect 3384 18856 4077 18884
rect 3384 18844 3390 18856
rect 4065 18853 4077 18856
rect 4111 18884 4123 18887
rect 4982 18884 4988 18896
rect 4111 18856 4988 18884
rect 4111 18853 4123 18856
rect 4065 18847 4123 18853
rect 4982 18844 4988 18856
rect 5040 18844 5046 18896
rect 4341 18819 4399 18825
rect 4341 18816 4353 18819
rect 2608 18788 4353 18816
rect 2501 18779 2559 18785
rect 4341 18785 4353 18788
rect 4387 18816 4399 18819
rect 5184 18816 5212 18924
rect 6638 18912 6644 18924
rect 6696 18912 6702 18964
rect 7193 18955 7251 18961
rect 7193 18921 7205 18955
rect 7239 18952 7251 18955
rect 10962 18952 10968 18964
rect 7239 18924 10968 18952
rect 7239 18921 7251 18924
rect 7193 18915 7251 18921
rect 10962 18912 10968 18924
rect 11020 18912 11026 18964
rect 11422 18912 11428 18964
rect 11480 18952 11486 18964
rect 11517 18955 11575 18961
rect 11517 18952 11529 18955
rect 11480 18924 11529 18952
rect 11480 18912 11486 18924
rect 11517 18921 11529 18924
rect 11563 18921 11575 18955
rect 11517 18915 11575 18921
rect 13446 18912 13452 18964
rect 13504 18952 13510 18964
rect 13541 18955 13599 18961
rect 13541 18952 13553 18955
rect 13504 18924 13553 18952
rect 13504 18912 13510 18924
rect 13541 18921 13553 18924
rect 13587 18921 13599 18955
rect 13541 18915 13599 18921
rect 13630 18912 13636 18964
rect 13688 18952 13694 18964
rect 13909 18955 13967 18961
rect 13688 18924 13733 18952
rect 13688 18912 13694 18924
rect 13909 18921 13921 18955
rect 13955 18952 13967 18955
rect 14090 18952 14096 18964
rect 13955 18924 14096 18952
rect 13955 18921 13967 18924
rect 13909 18915 13967 18921
rect 14090 18912 14096 18924
rect 14148 18952 14154 18964
rect 14366 18952 14372 18964
rect 14148 18924 14372 18952
rect 14148 18912 14154 18924
rect 14366 18912 14372 18924
rect 14424 18912 14430 18964
rect 14458 18912 14464 18964
rect 14516 18952 14522 18964
rect 15473 18955 15531 18961
rect 15473 18952 15485 18955
rect 14516 18924 15485 18952
rect 14516 18912 14522 18924
rect 15473 18921 15485 18924
rect 15519 18952 15531 18955
rect 16850 18952 16856 18964
rect 15519 18924 16856 18952
rect 15519 18921 15531 18924
rect 15473 18915 15531 18921
rect 16850 18912 16856 18924
rect 16908 18912 16914 18964
rect 17034 18912 17040 18964
rect 17092 18952 17098 18964
rect 17497 18955 17555 18961
rect 17497 18952 17509 18955
rect 17092 18924 17509 18952
rect 17092 18912 17098 18924
rect 17497 18921 17509 18924
rect 17543 18921 17555 18955
rect 17497 18915 17555 18921
rect 20533 18955 20591 18961
rect 20533 18921 20545 18955
rect 20579 18952 20591 18955
rect 20898 18952 20904 18964
rect 20579 18924 20904 18952
rect 20579 18921 20591 18924
rect 20533 18915 20591 18921
rect 20898 18912 20904 18924
rect 20956 18912 20962 18964
rect 21085 18955 21143 18961
rect 21085 18921 21097 18955
rect 21131 18952 21143 18955
rect 21542 18952 21548 18964
rect 21131 18924 21548 18952
rect 21131 18921 21143 18924
rect 21085 18915 21143 18921
rect 21542 18912 21548 18924
rect 21600 18912 21606 18964
rect 5626 18844 5632 18896
rect 5684 18884 5690 18896
rect 6270 18884 6276 18896
rect 5684 18856 6276 18884
rect 5684 18844 5690 18856
rect 5828 18825 5856 18856
rect 6270 18844 6276 18856
rect 6328 18844 6334 18896
rect 6365 18887 6423 18893
rect 6365 18853 6377 18887
rect 6411 18853 6423 18887
rect 6365 18847 6423 18853
rect 4387 18788 5212 18816
rect 5813 18819 5871 18825
rect 4387 18785 4399 18788
rect 4341 18779 4399 18785
rect 5813 18785 5825 18819
rect 5859 18785 5871 18819
rect 6380 18816 6408 18847
rect 6454 18844 6460 18896
rect 6512 18884 6518 18896
rect 7377 18887 7435 18893
rect 7377 18884 7389 18887
rect 6512 18856 7389 18884
rect 6512 18844 6518 18856
rect 7377 18853 7389 18856
rect 7423 18853 7435 18887
rect 7377 18847 7435 18853
rect 8763 18856 9619 18884
rect 6546 18816 6552 18828
rect 6380 18788 6552 18816
rect 5813 18779 5871 18785
rect 6546 18776 6552 18788
rect 6604 18776 6610 18828
rect 6641 18819 6699 18825
rect 6641 18785 6653 18819
rect 6687 18816 6699 18819
rect 7558 18816 7564 18828
rect 6687 18788 7564 18816
rect 6687 18785 6699 18788
rect 6641 18779 6699 18785
rect 7558 18776 7564 18788
rect 7616 18776 7622 18828
rect 8763 18816 8791 18856
rect 8671 18788 8791 18816
rect 9217 18819 9275 18825
rect 3329 18751 3387 18757
rect 3329 18748 3341 18751
rect 2240 18720 3341 18748
rect 2133 18711 2191 18717
rect 3329 18717 3341 18720
rect 3375 18748 3387 18751
rect 3789 18751 3847 18757
rect 3789 18748 3801 18751
rect 3375 18720 3801 18748
rect 3375 18717 3387 18720
rect 3329 18711 3387 18717
rect 3789 18717 3801 18720
rect 3835 18717 3847 18751
rect 3789 18711 3847 18717
rect 1765 18683 1823 18689
rect 1765 18649 1777 18683
rect 1811 18680 1823 18683
rect 2148 18680 2176 18711
rect 3970 18708 3976 18760
rect 4028 18748 4034 18760
rect 4028 18720 6132 18748
rect 4028 18708 4034 18720
rect 2593 18683 2651 18689
rect 1811 18652 2544 18680
rect 1811 18649 1823 18652
rect 1765 18643 1823 18649
rect 1486 18612 1492 18624
rect 1447 18584 1492 18612
rect 1486 18572 1492 18584
rect 1544 18572 1550 18624
rect 2516 18612 2544 18652
rect 2593 18649 2605 18683
rect 2639 18680 2651 18683
rect 3053 18683 3111 18689
rect 3053 18680 3065 18683
rect 2639 18652 3065 18680
rect 2639 18649 2651 18652
rect 2593 18643 2651 18649
rect 3053 18649 3065 18652
rect 3099 18649 3111 18683
rect 4430 18680 4436 18692
rect 3053 18643 3111 18649
rect 3160 18652 3740 18680
rect 4391 18652 4436 18680
rect 3160 18612 3188 18652
rect 3510 18612 3516 18624
rect 2516 18584 3188 18612
rect 3471 18584 3516 18612
rect 3510 18572 3516 18584
rect 3568 18572 3574 18624
rect 3712 18612 3740 18652
rect 4430 18640 4436 18652
rect 4488 18640 4494 18692
rect 5537 18683 5595 18689
rect 5537 18649 5549 18683
rect 5583 18680 5595 18683
rect 5997 18683 6055 18689
rect 5997 18680 6009 18683
rect 5583 18652 6009 18680
rect 5583 18649 5595 18652
rect 5537 18643 5595 18649
rect 5997 18649 6009 18652
rect 6043 18649 6055 18683
rect 6104 18680 6132 18720
rect 6178 18708 6184 18760
rect 6236 18748 6242 18760
rect 6733 18751 6791 18757
rect 6733 18748 6745 18751
rect 6236 18720 6745 18748
rect 6236 18708 6242 18720
rect 6733 18717 6745 18720
rect 6779 18717 6791 18751
rect 8671 18748 8699 18788
rect 9217 18785 9229 18819
rect 9263 18785 9275 18819
rect 9217 18779 9275 18785
rect 6733 18711 6791 18717
rect 6912 18720 8699 18748
rect 6104 18652 6500 18680
rect 5997 18643 6055 18649
rect 4525 18615 4583 18621
rect 4525 18612 4537 18615
rect 3712 18584 4537 18612
rect 4525 18581 4537 18584
rect 4571 18612 4583 18615
rect 4798 18612 4804 18624
rect 4571 18584 4804 18612
rect 4571 18581 4583 18584
rect 4525 18575 4583 18581
rect 4798 18572 4804 18584
rect 4856 18612 4862 18624
rect 4985 18615 5043 18621
rect 4985 18612 4997 18615
rect 4856 18584 4997 18612
rect 4856 18572 4862 18584
rect 4985 18581 4997 18584
rect 5031 18581 5043 18615
rect 5166 18612 5172 18624
rect 5127 18584 5172 18612
rect 4985 18575 5043 18581
rect 5166 18572 5172 18584
rect 5224 18612 5230 18624
rect 5905 18615 5963 18621
rect 5905 18612 5917 18615
rect 5224 18584 5917 18612
rect 5224 18572 5230 18584
rect 5905 18581 5917 18584
rect 5951 18581 5963 18615
rect 6472 18612 6500 18652
rect 6546 18640 6552 18692
rect 6604 18680 6610 18692
rect 6825 18683 6883 18689
rect 6825 18680 6837 18683
rect 6604 18652 6837 18680
rect 6604 18640 6610 18652
rect 6825 18649 6837 18652
rect 6871 18649 6883 18683
rect 6825 18643 6883 18649
rect 6912 18612 6940 18720
rect 8754 18708 8760 18760
rect 8812 18748 8818 18760
rect 9232 18748 9260 18779
rect 9490 18748 9496 18760
rect 8812 18720 8857 18748
rect 9232 18720 9496 18748
rect 8812 18708 8818 18720
rect 9490 18708 9496 18720
rect 9548 18708 9554 18760
rect 8512 18683 8570 18689
rect 8512 18649 8524 18683
rect 8558 18680 8570 18683
rect 9214 18680 9220 18692
rect 8558 18652 9220 18680
rect 8558 18649 8570 18652
rect 8512 18643 8570 18649
rect 9214 18640 9220 18652
rect 9272 18640 9278 18692
rect 6472 18584 6940 18612
rect 5905 18575 5963 18581
rect 9030 18572 9036 18624
rect 9088 18612 9094 18624
rect 9309 18615 9367 18621
rect 9309 18612 9321 18615
rect 9088 18584 9321 18612
rect 9088 18572 9094 18584
rect 9309 18581 9321 18584
rect 9355 18581 9367 18615
rect 9309 18575 9367 18581
rect 9401 18615 9459 18621
rect 9401 18581 9413 18615
rect 9447 18612 9459 18615
rect 9591 18612 9619 18856
rect 9674 18844 9680 18896
rect 9732 18884 9738 18896
rect 9769 18887 9827 18893
rect 9769 18884 9781 18887
rect 9732 18856 9781 18884
rect 9732 18844 9738 18856
rect 9769 18853 9781 18856
rect 9815 18853 9827 18887
rect 9769 18847 9827 18853
rect 11241 18887 11299 18893
rect 11241 18853 11253 18887
rect 11287 18884 11299 18887
rect 11330 18884 11336 18896
rect 11287 18856 11336 18884
rect 11287 18853 11299 18856
rect 11241 18847 11299 18853
rect 11330 18844 11336 18856
rect 11388 18844 11394 18896
rect 13265 18887 13323 18893
rect 13265 18853 13277 18887
rect 13311 18853 13323 18887
rect 16574 18884 16580 18896
rect 16535 18856 16580 18884
rect 13265 18847 13323 18853
rect 13280 18816 13308 18847
rect 16574 18844 16580 18856
rect 16632 18844 16638 18896
rect 17126 18844 17132 18896
rect 17184 18884 17190 18896
rect 17589 18887 17647 18893
rect 17589 18884 17601 18887
rect 17184 18856 17601 18884
rect 17184 18844 17190 18856
rect 17589 18853 17601 18856
rect 17635 18853 17647 18887
rect 17589 18847 17647 18853
rect 18509 18887 18567 18893
rect 18509 18853 18521 18887
rect 18555 18884 18567 18887
rect 20809 18887 20867 18893
rect 18555 18856 20760 18884
rect 18555 18853 18567 18856
rect 18509 18847 18567 18853
rect 16945 18819 17003 18825
rect 13280 18788 14228 18816
rect 9861 18751 9919 18757
rect 9861 18717 9873 18751
rect 9907 18748 9919 18751
rect 11793 18751 11851 18757
rect 11793 18748 11805 18751
rect 9907 18720 11805 18748
rect 9907 18717 9919 18720
rect 9861 18711 9919 18717
rect 11793 18717 11805 18720
rect 11839 18748 11851 18751
rect 11882 18748 11888 18760
rect 11839 18720 11888 18748
rect 11839 18717 11851 18720
rect 11793 18711 11851 18717
rect 11882 18708 11888 18720
rect 11940 18748 11946 18760
rect 12434 18748 12440 18760
rect 11940 18720 12440 18748
rect 11940 18708 11946 18720
rect 12434 18708 12440 18720
rect 12492 18708 12498 18760
rect 13262 18708 13268 18760
rect 13320 18748 13326 18760
rect 13357 18751 13415 18757
rect 13357 18748 13369 18751
rect 13320 18720 13369 18748
rect 13320 18708 13326 18720
rect 13357 18717 13369 18720
rect 13403 18717 13415 18751
rect 14090 18748 14096 18760
rect 14051 18720 14096 18748
rect 13357 18711 13415 18717
rect 14090 18708 14096 18720
rect 14148 18708 14154 18760
rect 14200 18748 14228 18788
rect 16945 18785 16957 18819
rect 16991 18816 17003 18819
rect 18141 18819 18199 18825
rect 18141 18816 18153 18819
rect 16991 18788 18153 18816
rect 16991 18785 17003 18788
rect 16945 18779 17003 18785
rect 18141 18785 18153 18788
rect 18187 18785 18199 18819
rect 18141 18779 18199 18785
rect 14360 18751 14418 18757
rect 14360 18748 14372 18751
rect 14200 18720 14372 18748
rect 14360 18717 14372 18720
rect 14406 18748 14418 18751
rect 16960 18748 16988 18779
rect 17954 18748 17960 18760
rect 14406 18720 16988 18748
rect 17915 18720 17960 18748
rect 14406 18717 14418 18720
rect 14360 18711 14418 18717
rect 17954 18708 17960 18720
rect 18012 18708 18018 18760
rect 9766 18640 9772 18692
rect 9824 18680 9830 18692
rect 10117 18683 10175 18689
rect 10117 18680 10129 18683
rect 9824 18652 10129 18680
rect 9824 18640 9830 18652
rect 10117 18649 10129 18652
rect 10163 18649 10175 18683
rect 10117 18643 10175 18649
rect 10704 18652 11284 18680
rect 10704 18612 10732 18652
rect 9447 18584 10732 18612
rect 11256 18612 11284 18652
rect 11330 18640 11336 18692
rect 11388 18680 11394 18692
rect 12130 18683 12188 18689
rect 12130 18680 12142 18683
rect 11388 18652 12142 18680
rect 11388 18640 11394 18652
rect 12130 18649 12142 18652
rect 12176 18649 12188 18683
rect 12130 18643 12188 18649
rect 16574 18640 16580 18692
rect 16632 18680 16638 18692
rect 17037 18683 17095 18689
rect 17037 18680 17049 18683
rect 16632 18652 17049 18680
rect 16632 18640 16638 18652
rect 17037 18649 17049 18652
rect 17083 18649 17095 18683
rect 17037 18643 17095 18649
rect 17129 18683 17187 18689
rect 17129 18649 17141 18683
rect 17175 18680 17187 18683
rect 17218 18680 17224 18692
rect 17175 18652 17224 18680
rect 17175 18649 17187 18652
rect 17129 18643 17187 18649
rect 17218 18640 17224 18652
rect 17276 18680 17282 18692
rect 18524 18680 18552 18847
rect 20073 18819 20131 18825
rect 20073 18785 20085 18819
rect 20119 18816 20131 18819
rect 20732 18816 20760 18856
rect 20809 18853 20821 18887
rect 20855 18884 20867 18887
rect 21266 18884 21272 18896
rect 20855 18856 21272 18884
rect 20855 18853 20867 18856
rect 20809 18847 20867 18853
rect 21266 18844 21272 18856
rect 21324 18844 21330 18896
rect 22278 18816 22284 18828
rect 20119 18788 20668 18816
rect 20732 18788 22284 18816
rect 20119 18785 20131 18788
rect 20073 18779 20131 18785
rect 20640 18760 20668 18788
rect 22278 18776 22284 18788
rect 22336 18776 22342 18828
rect 20349 18751 20407 18757
rect 20349 18717 20361 18751
rect 20395 18717 20407 18751
rect 20622 18748 20628 18760
rect 20583 18720 20628 18748
rect 20349 18711 20407 18717
rect 17276 18652 18552 18680
rect 17276 18640 17282 18652
rect 20364 18624 20392 18711
rect 20622 18708 20628 18720
rect 20680 18708 20686 18760
rect 20806 18708 20812 18760
rect 20864 18748 20870 18760
rect 20901 18751 20959 18757
rect 20901 18748 20913 18751
rect 20864 18720 20913 18748
rect 20864 18708 20870 18720
rect 20901 18717 20913 18720
rect 20947 18717 20959 18751
rect 21266 18748 21272 18760
rect 21227 18720 21272 18748
rect 20901 18711 20959 18717
rect 21266 18708 21272 18720
rect 21324 18708 21330 18760
rect 11425 18615 11483 18621
rect 11425 18612 11437 18615
rect 11256 18584 11437 18612
rect 9447 18581 9459 18584
rect 9401 18575 9459 18581
rect 11425 18581 11437 18584
rect 11471 18612 11483 18615
rect 13446 18612 13452 18624
rect 11471 18584 13452 18612
rect 11471 18581 11483 18584
rect 11425 18575 11483 18581
rect 13446 18572 13452 18584
rect 13504 18572 13510 18624
rect 18049 18615 18107 18621
rect 18049 18581 18061 18615
rect 18095 18612 18107 18615
rect 18322 18612 18328 18624
rect 18095 18584 18328 18612
rect 18095 18581 18107 18584
rect 18049 18575 18107 18581
rect 18322 18572 18328 18584
rect 18380 18572 18386 18624
rect 20257 18615 20315 18621
rect 20257 18581 20269 18615
rect 20303 18612 20315 18615
rect 20346 18612 20352 18624
rect 20303 18584 20352 18612
rect 20303 18581 20315 18584
rect 20257 18575 20315 18581
rect 20346 18572 20352 18584
rect 20404 18572 20410 18624
rect 21450 18612 21456 18624
rect 21411 18584 21456 18612
rect 21450 18572 21456 18584
rect 21508 18572 21514 18624
rect 1104 18522 22056 18544
rect 1104 18470 6148 18522
rect 6200 18470 6212 18522
rect 6264 18470 6276 18522
rect 6328 18470 6340 18522
rect 6392 18470 6404 18522
rect 6456 18470 11346 18522
rect 11398 18470 11410 18522
rect 11462 18470 11474 18522
rect 11526 18470 11538 18522
rect 11590 18470 11602 18522
rect 11654 18470 16544 18522
rect 16596 18470 16608 18522
rect 16660 18470 16672 18522
rect 16724 18470 16736 18522
rect 16788 18470 16800 18522
rect 16852 18470 21742 18522
rect 21794 18470 21806 18522
rect 21858 18470 21870 18522
rect 21922 18470 21934 18522
rect 21986 18470 21998 18522
rect 22050 18470 22056 18522
rect 1104 18448 22056 18470
rect 1670 18368 1676 18420
rect 1728 18408 1734 18420
rect 1949 18411 2007 18417
rect 1949 18408 1961 18411
rect 1728 18380 1961 18408
rect 1728 18368 1734 18380
rect 1949 18377 1961 18380
rect 1995 18377 2007 18411
rect 1949 18371 2007 18377
rect 2409 18411 2467 18417
rect 2409 18377 2421 18411
rect 2455 18408 2467 18411
rect 2682 18408 2688 18420
rect 2455 18380 2688 18408
rect 2455 18377 2467 18380
rect 2409 18371 2467 18377
rect 2682 18368 2688 18380
rect 2740 18368 2746 18420
rect 3142 18368 3148 18420
rect 3200 18408 3206 18420
rect 3421 18411 3479 18417
rect 3421 18408 3433 18411
rect 3200 18380 3433 18408
rect 3200 18368 3206 18380
rect 3421 18377 3433 18380
rect 3467 18377 3479 18411
rect 3878 18408 3884 18420
rect 3839 18380 3884 18408
rect 3421 18371 3479 18377
rect 3878 18368 3884 18380
rect 3936 18368 3942 18420
rect 4062 18408 4068 18420
rect 4023 18380 4068 18408
rect 4062 18368 4068 18380
rect 4120 18368 4126 18420
rect 4522 18408 4528 18420
rect 4483 18380 4528 18408
rect 4522 18368 4528 18380
rect 4580 18368 4586 18420
rect 4614 18368 4620 18420
rect 4672 18408 4678 18420
rect 4893 18411 4951 18417
rect 4893 18408 4905 18411
rect 4672 18380 4905 18408
rect 4672 18368 4678 18380
rect 4893 18377 4905 18380
rect 4939 18377 4951 18411
rect 4893 18371 4951 18377
rect 5442 18368 5448 18420
rect 5500 18408 5506 18420
rect 5537 18411 5595 18417
rect 5537 18408 5549 18411
rect 5500 18380 5549 18408
rect 5500 18368 5506 18380
rect 5537 18377 5549 18380
rect 5583 18377 5595 18411
rect 5537 18371 5595 18377
rect 5902 18368 5908 18420
rect 5960 18408 5966 18420
rect 6089 18411 6147 18417
rect 6089 18408 6101 18411
rect 5960 18380 6101 18408
rect 5960 18368 5966 18380
rect 6089 18377 6101 18380
rect 6135 18377 6147 18411
rect 6089 18371 6147 18377
rect 6549 18411 6607 18417
rect 6549 18377 6561 18411
rect 6595 18408 6607 18411
rect 6595 18380 7788 18408
rect 6595 18377 6607 18380
rect 6549 18371 6607 18377
rect 1394 18300 1400 18352
rect 1452 18340 1458 18352
rect 1452 18312 2268 18340
rect 1452 18300 1458 18312
rect 1673 18275 1731 18281
rect 1673 18241 1685 18275
rect 1719 18272 1731 18275
rect 1946 18272 1952 18284
rect 1719 18244 1952 18272
rect 1719 18241 1731 18244
rect 1673 18235 1731 18241
rect 1946 18232 1952 18244
rect 2004 18232 2010 18284
rect 2240 18281 2268 18312
rect 2958 18300 2964 18352
rect 3016 18340 3022 18352
rect 3053 18343 3111 18349
rect 3053 18340 3065 18343
rect 3016 18312 3065 18340
rect 3016 18300 3022 18312
rect 3053 18309 3065 18312
rect 3099 18340 3111 18343
rect 3970 18340 3976 18352
rect 3099 18312 3976 18340
rect 3099 18309 3111 18312
rect 3053 18303 3111 18309
rect 3970 18300 3976 18312
rect 4028 18300 4034 18352
rect 5721 18343 5779 18349
rect 5721 18309 5733 18343
rect 5767 18340 5779 18343
rect 5810 18340 5816 18352
rect 5767 18312 5816 18340
rect 5767 18309 5779 18312
rect 5721 18303 5779 18309
rect 5810 18300 5816 18312
rect 5868 18300 5874 18352
rect 2133 18275 2191 18281
rect 2133 18241 2145 18275
rect 2179 18241 2191 18275
rect 2133 18235 2191 18241
rect 2225 18275 2283 18281
rect 2225 18241 2237 18275
rect 2271 18241 2283 18275
rect 2225 18235 2283 18241
rect 1302 18096 1308 18148
rect 1360 18136 1366 18148
rect 1765 18139 1823 18145
rect 1765 18136 1777 18139
rect 1360 18108 1777 18136
rect 1360 18096 1366 18108
rect 1765 18105 1777 18108
rect 1811 18136 1823 18139
rect 1854 18136 1860 18148
rect 1811 18108 1860 18136
rect 1811 18105 1823 18108
rect 1765 18099 1823 18105
rect 1854 18096 1860 18108
rect 1912 18096 1918 18148
rect 2148 18136 2176 18235
rect 2406 18232 2412 18284
rect 2464 18272 2470 18284
rect 2501 18275 2559 18281
rect 2501 18272 2513 18275
rect 2464 18244 2513 18272
rect 2464 18232 2470 18244
rect 2501 18241 2513 18244
rect 2547 18241 2559 18275
rect 2501 18235 2559 18241
rect 3418 18232 3424 18284
rect 3476 18272 3482 18284
rect 3605 18275 3663 18281
rect 3605 18272 3617 18275
rect 3476 18244 3617 18272
rect 3476 18232 3482 18244
rect 3605 18241 3617 18244
rect 3651 18241 3663 18275
rect 3605 18235 3663 18241
rect 4706 18164 4712 18216
rect 4764 18204 4770 18216
rect 6564 18204 6592 18371
rect 6638 18300 6644 18352
rect 6696 18340 6702 18352
rect 7662 18343 7720 18349
rect 7662 18340 7674 18343
rect 6696 18312 7674 18340
rect 6696 18300 6702 18312
rect 7662 18309 7674 18312
rect 7708 18309 7720 18343
rect 7760 18340 7788 18380
rect 7926 18368 7932 18420
rect 7984 18408 7990 18420
rect 8021 18411 8079 18417
rect 8021 18408 8033 18411
rect 7984 18380 8033 18408
rect 7984 18368 7990 18380
rect 8021 18377 8033 18380
rect 8067 18377 8079 18411
rect 8662 18408 8668 18420
rect 8021 18371 8079 18377
rect 8128 18380 8668 18408
rect 8128 18340 8156 18380
rect 8662 18368 8668 18380
rect 8720 18368 8726 18420
rect 9582 18368 9588 18420
rect 9640 18408 9646 18420
rect 11149 18411 11207 18417
rect 11149 18408 11161 18411
rect 9640 18380 11161 18408
rect 9640 18368 9646 18380
rect 11149 18377 11161 18380
rect 11195 18377 11207 18411
rect 11149 18371 11207 18377
rect 11977 18411 12035 18417
rect 11977 18377 11989 18411
rect 12023 18408 12035 18411
rect 12437 18411 12495 18417
rect 12023 18380 12296 18408
rect 12023 18377 12035 18380
rect 11977 18371 12035 18377
rect 8570 18340 8576 18352
rect 7760 18312 8156 18340
rect 8531 18312 8576 18340
rect 7662 18303 7720 18309
rect 8570 18300 8576 18312
rect 8628 18300 8634 18352
rect 9490 18349 9496 18352
rect 9484 18340 9496 18349
rect 9403 18312 9496 18340
rect 9484 18303 9496 18312
rect 9548 18340 9554 18352
rect 10226 18340 10232 18352
rect 9548 18312 10232 18340
rect 9490 18300 9496 18303
rect 9548 18300 9554 18312
rect 10226 18300 10232 18312
rect 10284 18340 10290 18352
rect 10594 18340 10600 18352
rect 10284 18312 10600 18340
rect 10284 18300 10290 18312
rect 10594 18300 10600 18312
rect 10652 18300 10658 18352
rect 11057 18343 11115 18349
rect 11057 18340 11069 18343
rect 10796 18312 11069 18340
rect 7929 18275 7987 18281
rect 7929 18241 7941 18275
rect 7975 18272 7987 18275
rect 8297 18275 8355 18281
rect 8297 18272 8309 18275
rect 7975 18244 8309 18272
rect 7975 18241 7987 18244
rect 7929 18235 7987 18241
rect 8297 18241 8309 18244
rect 8343 18272 8355 18275
rect 8754 18272 8760 18284
rect 8343 18244 8760 18272
rect 8343 18241 8355 18244
rect 8297 18235 8355 18241
rect 8754 18232 8760 18244
rect 8812 18272 8818 18284
rect 8941 18275 8999 18281
rect 8941 18272 8953 18275
rect 8812 18244 8953 18272
rect 8812 18232 8818 18244
rect 8941 18241 8953 18244
rect 8987 18272 8999 18275
rect 9125 18275 9183 18281
rect 9125 18272 9137 18275
rect 8987 18244 9137 18272
rect 8987 18241 8999 18244
rect 8941 18235 8999 18241
rect 9125 18241 9137 18244
rect 9171 18272 9183 18275
rect 9217 18275 9275 18281
rect 9217 18272 9229 18275
rect 9171 18244 9229 18272
rect 9171 18241 9183 18244
rect 9125 18235 9183 18241
rect 9217 18241 9229 18244
rect 9263 18272 9275 18275
rect 10796 18272 10824 18312
rect 11057 18309 11069 18312
rect 11103 18340 11115 18343
rect 11882 18340 11888 18352
rect 11103 18312 11888 18340
rect 11103 18309 11115 18312
rect 11057 18303 11115 18309
rect 11882 18300 11888 18312
rect 11940 18300 11946 18352
rect 9263 18244 10824 18272
rect 9263 18241 9275 18244
rect 9217 18235 9275 18241
rect 10870 18232 10876 18284
rect 10928 18272 10934 18284
rect 12069 18275 12127 18281
rect 12069 18272 12081 18275
rect 10928 18244 12081 18272
rect 10928 18232 10934 18244
rect 12069 18241 12081 18244
rect 12115 18241 12127 18275
rect 12268 18272 12296 18380
rect 12437 18377 12449 18411
rect 12483 18408 12495 18411
rect 16117 18411 16175 18417
rect 12483 18380 15240 18408
rect 12483 18377 12495 18380
rect 12437 18371 12495 18377
rect 13449 18343 13507 18349
rect 13449 18309 13461 18343
rect 13495 18340 13507 18343
rect 14366 18340 14372 18352
rect 13495 18312 14372 18340
rect 13495 18309 13507 18312
rect 13449 18303 13507 18309
rect 13170 18272 13176 18284
rect 12268 18244 13176 18272
rect 12069 18235 12127 18241
rect 13170 18232 13176 18244
rect 13228 18232 13234 18284
rect 10686 18204 10692 18216
rect 4764 18176 6592 18204
rect 10647 18176 10692 18204
rect 4764 18164 4770 18176
rect 10686 18164 10692 18176
rect 10744 18164 10750 18216
rect 11790 18204 11796 18216
rect 11751 18176 11796 18204
rect 11790 18164 11796 18176
rect 11848 18164 11854 18216
rect 12434 18164 12440 18216
rect 12492 18204 12498 18216
rect 13464 18204 13492 18303
rect 14366 18300 14372 18312
rect 14424 18340 14430 18352
rect 15212 18340 15240 18380
rect 16117 18377 16129 18411
rect 16163 18408 16175 18411
rect 16298 18408 16304 18420
rect 16163 18380 16304 18408
rect 16163 18377 16175 18380
rect 16117 18371 16175 18377
rect 16298 18368 16304 18380
rect 16356 18368 16362 18420
rect 17589 18411 17647 18417
rect 17589 18377 17601 18411
rect 17635 18408 17647 18411
rect 18414 18408 18420 18420
rect 17635 18380 18420 18408
rect 17635 18377 17647 18380
rect 17589 18371 17647 18377
rect 18414 18368 18420 18380
rect 18472 18368 18478 18420
rect 20717 18411 20775 18417
rect 20717 18377 20729 18411
rect 20763 18408 20775 18411
rect 21266 18408 21272 18420
rect 20763 18380 21272 18408
rect 20763 18377 20775 18380
rect 20717 18371 20775 18377
rect 21266 18368 21272 18380
rect 21324 18368 21330 18420
rect 18046 18340 18052 18352
rect 14424 18312 14964 18340
rect 15212 18312 18052 18340
rect 14424 18300 14430 18312
rect 14665 18275 14723 18281
rect 14665 18241 14677 18275
rect 14711 18272 14723 18275
rect 14826 18272 14832 18284
rect 14711 18244 14832 18272
rect 14711 18241 14723 18244
rect 14665 18235 14723 18241
rect 14826 18232 14832 18244
rect 14884 18232 14890 18284
rect 14936 18281 14964 18312
rect 18046 18300 18052 18312
rect 18104 18300 18110 18352
rect 14921 18275 14979 18281
rect 14921 18241 14933 18275
rect 14967 18241 14979 18275
rect 15746 18272 15752 18284
rect 15707 18244 15752 18272
rect 14921 18235 14979 18241
rect 15746 18232 15752 18244
rect 15804 18232 15810 18284
rect 17402 18272 17408 18284
rect 17363 18244 17408 18272
rect 17402 18232 17408 18244
rect 17460 18232 17466 18284
rect 20530 18272 20536 18284
rect 20491 18244 20536 18272
rect 20530 18232 20536 18244
rect 20588 18232 20594 18284
rect 20993 18275 21051 18281
rect 20993 18241 21005 18275
rect 21039 18241 21051 18275
rect 20993 18235 21051 18241
rect 15473 18207 15531 18213
rect 15473 18204 15485 18207
rect 12492 18176 13492 18204
rect 14936 18176 15485 18204
rect 12492 18164 12498 18176
rect 2498 18136 2504 18148
rect 2148 18108 2504 18136
rect 2498 18096 2504 18108
rect 2556 18096 2562 18148
rect 2866 18136 2872 18148
rect 2779 18108 2872 18136
rect 2866 18096 2872 18108
rect 2924 18136 2930 18148
rect 3142 18136 3148 18148
rect 2924 18108 3148 18136
rect 2924 18096 2930 18108
rect 3142 18096 3148 18108
rect 3200 18096 3206 18148
rect 3234 18096 3240 18148
rect 3292 18136 3298 18148
rect 5905 18139 5963 18145
rect 3292 18108 5856 18136
rect 3292 18096 3298 18108
rect 1486 18068 1492 18080
rect 1447 18040 1492 18068
rect 1486 18028 1492 18040
rect 1544 18028 1550 18080
rect 2682 18068 2688 18080
rect 2643 18040 2688 18068
rect 2682 18028 2688 18040
rect 2740 18028 2746 18080
rect 3326 18068 3332 18080
rect 3239 18040 3332 18068
rect 3326 18028 3332 18040
rect 3384 18068 3390 18080
rect 4062 18068 4068 18080
rect 3384 18040 4068 18068
rect 3384 18028 3390 18040
rect 4062 18028 4068 18040
rect 4120 18028 4126 18080
rect 5828 18068 5856 18108
rect 5905 18105 5917 18139
rect 5951 18136 5963 18139
rect 5994 18136 6000 18148
rect 5951 18108 6000 18136
rect 5951 18105 5963 18108
rect 5905 18099 5963 18105
rect 5994 18096 6000 18108
rect 6052 18136 6058 18148
rect 6457 18139 6515 18145
rect 6457 18136 6469 18139
rect 6052 18108 6469 18136
rect 6052 18096 6058 18108
rect 6457 18105 6469 18108
rect 6503 18136 6515 18139
rect 6638 18136 6644 18148
rect 6503 18108 6644 18136
rect 6503 18105 6515 18108
rect 6457 18099 6515 18105
rect 6638 18096 6644 18108
rect 6696 18096 6702 18148
rect 8294 18096 8300 18148
rect 8352 18136 8358 18148
rect 8665 18139 8723 18145
rect 8665 18136 8677 18139
rect 8352 18108 8677 18136
rect 8352 18096 8358 18108
rect 8665 18105 8677 18108
rect 8711 18105 8723 18139
rect 8665 18099 8723 18105
rect 9030 18068 9036 18080
rect 5828 18040 9036 18068
rect 9030 18028 9036 18040
rect 9088 18068 9094 18080
rect 9490 18068 9496 18080
rect 9088 18040 9496 18068
rect 9088 18028 9094 18040
rect 9490 18028 9496 18040
rect 9548 18028 9554 18080
rect 10502 18028 10508 18080
rect 10560 18068 10566 18080
rect 10597 18071 10655 18077
rect 10597 18068 10609 18071
rect 10560 18040 10609 18068
rect 10560 18028 10566 18040
rect 10597 18037 10609 18040
rect 10643 18037 10655 18071
rect 10597 18031 10655 18037
rect 12802 18028 12808 18080
rect 12860 18068 12866 18080
rect 13541 18071 13599 18077
rect 13541 18068 13553 18071
rect 12860 18040 13553 18068
rect 12860 18028 12866 18040
rect 13541 18037 13553 18040
rect 13587 18068 13599 18071
rect 14936 18068 14964 18176
rect 15473 18173 15485 18176
rect 15519 18173 15531 18207
rect 15473 18167 15531 18173
rect 15562 18164 15568 18216
rect 15620 18204 15626 18216
rect 15657 18207 15715 18213
rect 15657 18204 15669 18207
rect 15620 18176 15669 18204
rect 15620 18164 15626 18176
rect 15657 18173 15669 18176
rect 15703 18173 15715 18207
rect 18414 18204 18420 18216
rect 18375 18176 18420 18204
rect 15657 18167 15715 18173
rect 18414 18164 18420 18176
rect 18472 18164 18478 18216
rect 19886 18164 19892 18216
rect 19944 18204 19950 18216
rect 21008 18204 21036 18235
rect 21174 18232 21180 18284
rect 21232 18272 21238 18284
rect 21269 18275 21327 18281
rect 21269 18272 21281 18275
rect 21232 18244 21281 18272
rect 21232 18232 21238 18244
rect 21269 18241 21281 18244
rect 21315 18241 21327 18275
rect 21269 18235 21327 18241
rect 19944 18176 21036 18204
rect 19944 18164 19950 18176
rect 17773 18139 17831 18145
rect 17773 18105 17785 18139
rect 17819 18136 17831 18139
rect 18322 18136 18328 18148
rect 17819 18108 18328 18136
rect 17819 18105 17831 18108
rect 17773 18099 17831 18105
rect 18322 18096 18328 18108
rect 18380 18096 18386 18148
rect 20714 18096 20720 18148
rect 20772 18136 20778 18148
rect 20809 18139 20867 18145
rect 20809 18136 20821 18139
rect 20772 18108 20821 18136
rect 20772 18096 20778 18108
rect 20809 18105 20821 18108
rect 20855 18105 20867 18139
rect 20809 18099 20867 18105
rect 18046 18068 18052 18080
rect 13587 18040 14964 18068
rect 18007 18040 18052 18068
rect 13587 18037 13599 18040
rect 13541 18031 13599 18037
rect 18046 18028 18052 18040
rect 18104 18028 18110 18080
rect 21450 18068 21456 18080
rect 21411 18040 21456 18068
rect 21450 18028 21456 18040
rect 21508 18028 21514 18080
rect 1104 17978 21896 18000
rect 1104 17926 3549 17978
rect 3601 17926 3613 17978
rect 3665 17926 3677 17978
rect 3729 17926 3741 17978
rect 3793 17926 3805 17978
rect 3857 17926 8747 17978
rect 8799 17926 8811 17978
rect 8863 17926 8875 17978
rect 8927 17926 8939 17978
rect 8991 17926 9003 17978
rect 9055 17926 13945 17978
rect 13997 17926 14009 17978
rect 14061 17926 14073 17978
rect 14125 17926 14137 17978
rect 14189 17926 14201 17978
rect 14253 17926 19143 17978
rect 19195 17926 19207 17978
rect 19259 17926 19271 17978
rect 19323 17926 19335 17978
rect 19387 17926 19399 17978
rect 19451 17926 21896 17978
rect 1104 17904 21896 17926
rect 2038 17824 2044 17876
rect 2096 17864 2102 17876
rect 2133 17867 2191 17873
rect 2133 17864 2145 17867
rect 2096 17836 2145 17864
rect 2096 17824 2102 17836
rect 2133 17833 2145 17836
rect 2179 17833 2191 17867
rect 2133 17827 2191 17833
rect 2314 17824 2320 17876
rect 2372 17864 2378 17876
rect 2409 17867 2467 17873
rect 2409 17864 2421 17867
rect 2372 17836 2421 17864
rect 2372 17824 2378 17836
rect 2409 17833 2421 17836
rect 2455 17833 2467 17867
rect 2590 17864 2596 17876
rect 2551 17836 2596 17864
rect 2409 17827 2467 17833
rect 2424 17728 2452 17827
rect 2590 17824 2596 17836
rect 2648 17824 2654 17876
rect 5629 17867 5687 17873
rect 5629 17833 5641 17867
rect 5675 17864 5687 17867
rect 5994 17864 6000 17876
rect 5675 17836 6000 17864
rect 5675 17833 5687 17836
rect 5629 17827 5687 17833
rect 5994 17824 6000 17836
rect 6052 17824 6058 17876
rect 6914 17824 6920 17876
rect 6972 17864 6978 17876
rect 7374 17864 7380 17876
rect 6972 17836 7380 17864
rect 6972 17824 6978 17836
rect 7374 17824 7380 17836
rect 7432 17864 7438 17876
rect 7469 17867 7527 17873
rect 7469 17864 7481 17867
rect 7432 17836 7481 17864
rect 7432 17824 7438 17836
rect 7469 17833 7481 17836
rect 7515 17833 7527 17867
rect 7469 17827 7527 17833
rect 7745 17867 7803 17873
rect 7745 17833 7757 17867
rect 7791 17864 7803 17867
rect 7834 17864 7840 17876
rect 7791 17836 7840 17864
rect 7791 17833 7803 17836
rect 7745 17827 7803 17833
rect 7834 17824 7840 17836
rect 7892 17824 7898 17876
rect 7929 17867 7987 17873
rect 7929 17833 7941 17867
rect 7975 17864 7987 17867
rect 8386 17864 8392 17876
rect 7975 17836 8392 17864
rect 7975 17833 7987 17836
rect 7929 17827 7987 17833
rect 8386 17824 8392 17836
rect 8444 17824 8450 17876
rect 8754 17864 8760 17876
rect 8715 17836 8760 17864
rect 8754 17824 8760 17836
rect 8812 17824 8818 17876
rect 9033 17867 9091 17873
rect 9033 17833 9045 17867
rect 9079 17864 9091 17867
rect 9122 17864 9128 17876
rect 9079 17836 9128 17864
rect 9079 17833 9091 17836
rect 9033 17827 9091 17833
rect 9122 17824 9128 17836
rect 9180 17824 9186 17876
rect 9401 17867 9459 17873
rect 9401 17833 9413 17867
rect 9447 17864 9459 17867
rect 9858 17864 9864 17876
rect 9447 17836 9864 17864
rect 9447 17833 9459 17836
rect 9401 17827 9459 17833
rect 9858 17824 9864 17836
rect 9916 17824 9922 17876
rect 10410 17864 10416 17876
rect 10371 17836 10416 17864
rect 10410 17824 10416 17836
rect 10468 17824 10474 17876
rect 11146 17824 11152 17876
rect 11204 17864 11210 17876
rect 12066 17864 12072 17876
rect 11204 17836 12072 17864
rect 11204 17824 11210 17836
rect 12066 17824 12072 17836
rect 12124 17824 12130 17876
rect 12618 17824 12624 17876
rect 12676 17864 12682 17876
rect 13633 17867 13691 17873
rect 12676 17836 13308 17864
rect 12676 17824 12682 17836
rect 8018 17756 8024 17808
rect 8076 17796 8082 17808
rect 9217 17799 9275 17805
rect 9217 17796 9229 17799
rect 8076 17768 9229 17796
rect 8076 17756 8082 17768
rect 9217 17765 9229 17768
rect 9263 17765 9275 17799
rect 10502 17796 10508 17808
rect 9217 17759 9275 17765
rect 9692 17768 10508 17796
rect 2590 17728 2596 17740
rect 2424 17700 2596 17728
rect 2590 17688 2596 17700
rect 2648 17688 2654 17740
rect 8202 17728 8208 17740
rect 8163 17700 8208 17728
rect 8202 17688 8208 17700
rect 8260 17688 8266 17740
rect 9692 17737 9720 17768
rect 10502 17756 10508 17768
rect 10560 17756 10566 17808
rect 11514 17796 11520 17808
rect 11256 17768 11520 17796
rect 11256 17740 11284 17768
rect 11514 17756 11520 17768
rect 11572 17756 11578 17808
rect 13280 17796 13308 17836
rect 13633 17833 13645 17867
rect 13679 17864 13691 17867
rect 15562 17864 15568 17876
rect 13679 17836 15568 17864
rect 13679 17833 13691 17836
rect 13633 17827 13691 17833
rect 15562 17824 15568 17836
rect 15620 17824 15626 17876
rect 15746 17824 15752 17876
rect 15804 17864 15810 17876
rect 16577 17867 16635 17873
rect 16577 17864 16589 17867
rect 15804 17836 16589 17864
rect 15804 17824 15810 17836
rect 16577 17833 16589 17836
rect 16623 17833 16635 17867
rect 16577 17827 16635 17833
rect 19981 17867 20039 17873
rect 19981 17833 19993 17867
rect 20027 17864 20039 17867
rect 20530 17864 20536 17876
rect 20027 17836 20536 17864
rect 20027 17833 20039 17836
rect 19981 17827 20039 17833
rect 20530 17824 20536 17836
rect 20588 17824 20594 17876
rect 14550 17796 14556 17808
rect 13280 17768 14556 17796
rect 14550 17756 14556 17768
rect 14608 17756 14614 17808
rect 16485 17799 16543 17805
rect 16485 17765 16497 17799
rect 16531 17796 16543 17799
rect 16942 17796 16948 17808
rect 16531 17768 16948 17796
rect 16531 17765 16543 17768
rect 16485 17759 16543 17765
rect 16942 17756 16948 17768
rect 17000 17756 17006 17808
rect 17494 17756 17500 17808
rect 17552 17796 17558 17808
rect 17552 17768 18828 17796
rect 17552 17756 17558 17768
rect 18800 17740 18828 17768
rect 9677 17731 9735 17737
rect 9677 17697 9689 17731
rect 9723 17697 9735 17731
rect 9677 17691 9735 17697
rect 9766 17688 9772 17740
rect 9824 17728 9830 17740
rect 9861 17731 9919 17737
rect 9861 17728 9873 17731
rect 9824 17700 9873 17728
rect 9824 17688 9830 17700
rect 9861 17697 9873 17700
rect 9907 17697 9919 17731
rect 9861 17691 9919 17697
rect 10042 17688 10048 17740
rect 10100 17728 10106 17740
rect 11238 17728 11244 17740
rect 10100 17700 11244 17728
rect 10100 17688 10106 17700
rect 11238 17688 11244 17700
rect 11296 17688 11302 17740
rect 11333 17731 11391 17737
rect 11333 17697 11345 17731
rect 11379 17728 11391 17731
rect 11698 17728 11704 17740
rect 11379 17700 11704 17728
rect 11379 17697 11391 17700
rect 11333 17691 11391 17697
rect 11698 17688 11704 17700
rect 11756 17728 11762 17740
rect 12158 17728 12164 17740
rect 11756 17700 12164 17728
rect 11756 17688 11762 17700
rect 12158 17688 12164 17700
rect 12216 17688 12222 17740
rect 13081 17731 13139 17737
rect 13081 17697 13093 17731
rect 13127 17728 13139 17731
rect 13998 17728 14004 17740
rect 13127 17700 14004 17728
rect 13127 17697 13139 17700
rect 13081 17691 13139 17697
rect 13998 17688 14004 17700
rect 14056 17688 14062 17740
rect 15838 17688 15844 17740
rect 15896 17728 15902 17740
rect 17129 17731 17187 17737
rect 17129 17728 17141 17731
rect 15896 17700 17141 17728
rect 15896 17688 15902 17700
rect 17129 17697 17141 17700
rect 17175 17697 17187 17731
rect 17129 17691 17187 17697
rect 17586 17688 17592 17740
rect 17644 17728 17650 17740
rect 17957 17731 18015 17737
rect 17957 17728 17969 17731
rect 17644 17700 17969 17728
rect 17644 17688 17650 17700
rect 17957 17697 17969 17700
rect 18003 17697 18015 17731
rect 18782 17728 18788 17740
rect 18695 17700 18788 17728
rect 17957 17691 18015 17697
rect 18782 17688 18788 17700
rect 18840 17688 18846 17740
rect 1578 17620 1584 17672
rect 1636 17660 1642 17672
rect 1673 17663 1731 17669
rect 1673 17660 1685 17663
rect 1636 17632 1685 17660
rect 1636 17620 1642 17632
rect 1673 17629 1685 17632
rect 1719 17629 1731 17663
rect 2038 17660 2044 17672
rect 1999 17632 2044 17660
rect 1673 17623 1731 17629
rect 2038 17620 2044 17632
rect 2096 17620 2102 17672
rect 2314 17660 2320 17672
rect 2275 17632 2320 17660
rect 2314 17620 2320 17632
rect 2372 17620 2378 17672
rect 7101 17663 7159 17669
rect 7101 17629 7113 17663
rect 7147 17629 7159 17663
rect 7101 17623 7159 17629
rect 2222 17552 2228 17604
rect 2280 17592 2286 17604
rect 2777 17595 2835 17601
rect 2777 17592 2789 17595
rect 2280 17564 2789 17592
rect 2280 17552 2286 17564
rect 2777 17561 2789 17564
rect 2823 17561 2835 17595
rect 2777 17555 2835 17561
rect 6822 17552 6828 17604
rect 6880 17601 6886 17604
rect 6880 17592 6892 17601
rect 7116 17592 7144 17623
rect 7650 17620 7656 17672
rect 7708 17660 7714 17672
rect 8018 17660 8024 17672
rect 7708 17632 8024 17660
rect 7708 17620 7714 17632
rect 8018 17620 8024 17632
rect 8076 17660 8082 17672
rect 8297 17663 8355 17669
rect 8297 17660 8309 17663
rect 8076 17632 8309 17660
rect 8076 17620 8082 17632
rect 8297 17629 8309 17632
rect 8343 17629 8355 17663
rect 8297 17623 8355 17629
rect 8754 17620 8760 17672
rect 8812 17660 8818 17672
rect 8812 17632 13676 17660
rect 8812 17620 8818 17632
rect 7285 17595 7343 17601
rect 7285 17592 7297 17595
rect 6880 17564 6925 17592
rect 7116 17564 7297 17592
rect 6880 17555 6892 17564
rect 6880 17552 6886 17555
rect 1486 17524 1492 17536
rect 1447 17496 1492 17524
rect 1486 17484 1492 17496
rect 1544 17484 1550 17536
rect 1854 17524 1860 17536
rect 1815 17496 1860 17524
rect 1854 17484 1860 17496
rect 1912 17484 1918 17536
rect 5074 17484 5080 17536
rect 5132 17524 5138 17536
rect 5721 17527 5779 17533
rect 5721 17524 5733 17527
rect 5132 17496 5733 17524
rect 5132 17484 5138 17496
rect 5721 17493 5733 17496
rect 5767 17493 5779 17527
rect 5721 17487 5779 17493
rect 6638 17484 6644 17536
rect 6696 17524 6702 17536
rect 7116 17524 7144 17564
rect 7285 17561 7297 17564
rect 7331 17592 7343 17595
rect 8202 17592 8208 17604
rect 7331 17564 8208 17592
rect 7331 17561 7343 17564
rect 7285 17555 7343 17561
rect 8202 17552 8208 17564
rect 8260 17552 8266 17604
rect 8389 17595 8447 17601
rect 8389 17561 8401 17595
rect 8435 17592 8447 17595
rect 8570 17592 8576 17604
rect 8435 17564 8576 17592
rect 8435 17561 8447 17564
rect 8389 17555 8447 17561
rect 8570 17552 8576 17564
rect 8628 17592 8634 17604
rect 9398 17592 9404 17604
rect 8628 17564 9404 17592
rect 8628 17552 8634 17564
rect 9398 17552 9404 17564
rect 9456 17552 9462 17604
rect 11974 17592 11980 17604
rect 9600 17564 11980 17592
rect 6696 17496 7144 17524
rect 6696 17484 6702 17496
rect 7742 17484 7748 17536
rect 7800 17524 7806 17536
rect 9600 17524 9628 17564
rect 11974 17552 11980 17564
rect 12032 17592 12038 17604
rect 12437 17595 12495 17601
rect 12437 17592 12449 17595
rect 12032 17564 12449 17592
rect 12032 17552 12038 17564
rect 12437 17561 12449 17564
rect 12483 17592 12495 17595
rect 12618 17592 12624 17604
rect 12483 17564 12624 17592
rect 12483 17561 12495 17564
rect 12437 17555 12495 17561
rect 12618 17552 12624 17564
rect 12676 17552 12682 17604
rect 13265 17595 13323 17601
rect 13265 17592 13277 17595
rect 12820 17564 13277 17592
rect 7800 17496 9628 17524
rect 7800 17484 7806 17496
rect 9674 17484 9680 17536
rect 9732 17524 9738 17536
rect 9953 17527 10011 17533
rect 9953 17524 9965 17527
rect 9732 17496 9965 17524
rect 9732 17484 9738 17496
rect 9953 17493 9965 17496
rect 9999 17493 10011 17527
rect 9953 17487 10011 17493
rect 10134 17484 10140 17536
rect 10192 17524 10198 17536
rect 10321 17527 10379 17533
rect 10321 17524 10333 17527
rect 10192 17496 10333 17524
rect 10192 17484 10198 17496
rect 10321 17493 10333 17496
rect 10367 17493 10379 17527
rect 10321 17487 10379 17493
rect 10594 17484 10600 17536
rect 10652 17524 10658 17536
rect 10962 17524 10968 17536
rect 10652 17496 10968 17524
rect 10652 17484 10658 17496
rect 10962 17484 10968 17496
rect 11020 17524 11026 17536
rect 11057 17527 11115 17533
rect 11057 17524 11069 17527
rect 11020 17496 11069 17524
rect 11020 17484 11026 17496
rect 11057 17493 11069 17496
rect 11103 17524 11115 17527
rect 11425 17527 11483 17533
rect 11425 17524 11437 17527
rect 11103 17496 11437 17524
rect 11103 17493 11115 17496
rect 11057 17487 11115 17493
rect 11425 17493 11437 17496
rect 11471 17493 11483 17527
rect 11425 17487 11483 17493
rect 11514 17484 11520 17536
rect 11572 17524 11578 17536
rect 11572 17496 11617 17524
rect 11572 17484 11578 17496
rect 11790 17484 11796 17536
rect 11848 17524 11854 17536
rect 11885 17527 11943 17533
rect 11885 17524 11897 17527
rect 11848 17496 11897 17524
rect 11848 17484 11854 17496
rect 11885 17493 11897 17496
rect 11931 17493 11943 17527
rect 11885 17487 11943 17493
rect 12066 17484 12072 17536
rect 12124 17524 12130 17536
rect 12820 17533 12848 17564
rect 13265 17561 13277 17564
rect 13311 17561 13323 17595
rect 13648 17592 13676 17632
rect 13722 17620 13728 17672
rect 13780 17660 13786 17672
rect 13817 17663 13875 17669
rect 13817 17660 13829 17663
rect 13780 17632 13829 17660
rect 13780 17620 13786 17632
rect 13817 17629 13829 17632
rect 13863 17660 13875 17663
rect 14277 17663 14335 17669
rect 14277 17660 14289 17663
rect 13863 17632 14289 17660
rect 13863 17629 13875 17632
rect 13817 17623 13875 17629
rect 14277 17629 14289 17632
rect 14323 17660 14335 17663
rect 15746 17660 15752 17672
rect 14323 17632 15752 17660
rect 14323 17629 14335 17632
rect 14277 17623 14335 17629
rect 15746 17620 15752 17632
rect 15804 17620 15810 17672
rect 16298 17660 16304 17672
rect 16259 17632 16304 17660
rect 16298 17620 16304 17632
rect 16356 17620 16362 17672
rect 18046 17620 18052 17672
rect 18104 17660 18110 17672
rect 18104 17632 18368 17660
rect 18104 17620 18110 17632
rect 13648 17564 15424 17592
rect 13265 17555 13323 17561
rect 12345 17527 12403 17533
rect 12345 17524 12357 17527
rect 12124 17496 12357 17524
rect 12124 17484 12130 17496
rect 12345 17493 12357 17496
rect 12391 17493 12403 17527
rect 12345 17487 12403 17493
rect 12805 17527 12863 17533
rect 12805 17493 12817 17527
rect 12851 17493 12863 17527
rect 13170 17524 13176 17536
rect 13131 17496 13176 17524
rect 12805 17487 12863 17493
rect 13170 17484 13176 17496
rect 13228 17484 13234 17536
rect 14366 17524 14372 17536
rect 14327 17496 14372 17524
rect 14366 17484 14372 17496
rect 14424 17484 14430 17536
rect 15396 17524 15424 17564
rect 15470 17552 15476 17604
rect 15528 17601 15534 17604
rect 15528 17592 15540 17601
rect 17678 17592 17684 17604
rect 15528 17564 15573 17592
rect 16776 17564 17684 17592
rect 15528 17555 15540 17564
rect 15528 17552 15534 17555
rect 16776 17524 16804 17564
rect 17678 17552 17684 17564
rect 17736 17552 17742 17604
rect 17773 17595 17831 17601
rect 17773 17561 17785 17595
rect 17819 17592 17831 17595
rect 18340 17592 18368 17632
rect 18414 17620 18420 17672
rect 18472 17660 18478 17672
rect 18601 17663 18659 17669
rect 18601 17660 18613 17663
rect 18472 17632 18613 17660
rect 18472 17620 18478 17632
rect 18601 17629 18613 17632
rect 18647 17629 18659 17663
rect 19794 17660 19800 17672
rect 19755 17632 19800 17660
rect 18601 17623 18659 17629
rect 19794 17620 19800 17632
rect 19852 17620 19858 17672
rect 20622 17620 20628 17672
rect 20680 17660 20686 17672
rect 20901 17663 20959 17669
rect 20901 17660 20913 17663
rect 20680 17632 20913 17660
rect 20680 17620 20686 17632
rect 20901 17629 20913 17632
rect 20947 17629 20959 17663
rect 21266 17660 21272 17672
rect 21227 17632 21272 17660
rect 20901 17623 20959 17629
rect 21266 17620 21272 17632
rect 21324 17620 21330 17672
rect 18693 17595 18751 17601
rect 18693 17592 18705 17595
rect 17819 17564 18276 17592
rect 18340 17564 18705 17592
rect 17819 17561 17831 17564
rect 17773 17555 17831 17561
rect 16942 17524 16948 17536
rect 15396 17496 16804 17524
rect 16903 17496 16948 17524
rect 16942 17484 16948 17496
rect 17000 17484 17006 17536
rect 17037 17527 17095 17533
rect 17037 17493 17049 17527
rect 17083 17524 17095 17527
rect 17218 17524 17224 17536
rect 17083 17496 17224 17524
rect 17083 17493 17095 17496
rect 17037 17487 17095 17493
rect 17218 17484 17224 17496
rect 17276 17484 17282 17536
rect 17402 17524 17408 17536
rect 17363 17496 17408 17524
rect 17402 17484 17408 17496
rect 17460 17484 17466 17536
rect 17865 17527 17923 17533
rect 17865 17493 17877 17527
rect 17911 17524 17923 17527
rect 18138 17524 18144 17536
rect 17911 17496 18144 17524
rect 17911 17493 17923 17496
rect 17865 17487 17923 17493
rect 18138 17484 18144 17496
rect 18196 17484 18202 17536
rect 18248 17533 18276 17564
rect 18693 17561 18705 17564
rect 18739 17561 18751 17595
rect 18693 17555 18751 17561
rect 18233 17527 18291 17533
rect 18233 17493 18245 17527
rect 18279 17493 18291 17527
rect 21082 17524 21088 17536
rect 21043 17496 21088 17524
rect 18233 17487 18291 17493
rect 21082 17484 21088 17496
rect 21140 17484 21146 17536
rect 21450 17524 21456 17536
rect 21411 17496 21456 17524
rect 21450 17484 21456 17496
rect 21508 17484 21514 17536
rect 1104 17434 22056 17456
rect 1104 17382 6148 17434
rect 6200 17382 6212 17434
rect 6264 17382 6276 17434
rect 6328 17382 6340 17434
rect 6392 17382 6404 17434
rect 6456 17382 11346 17434
rect 11398 17382 11410 17434
rect 11462 17382 11474 17434
rect 11526 17382 11538 17434
rect 11590 17382 11602 17434
rect 11654 17382 16544 17434
rect 16596 17382 16608 17434
rect 16660 17382 16672 17434
rect 16724 17382 16736 17434
rect 16788 17382 16800 17434
rect 16852 17382 21742 17434
rect 21794 17382 21806 17434
rect 21858 17382 21870 17434
rect 21922 17382 21934 17434
rect 21986 17382 21998 17434
rect 22050 17382 22056 17434
rect 1104 17360 22056 17382
rect 4338 17280 4344 17332
rect 4396 17320 4402 17332
rect 9398 17320 9404 17332
rect 4396 17292 9404 17320
rect 4396 17280 4402 17292
rect 9398 17280 9404 17292
rect 9456 17280 9462 17332
rect 9674 17320 9680 17332
rect 9635 17292 9680 17320
rect 9674 17280 9680 17292
rect 9732 17280 9738 17332
rect 10045 17323 10103 17329
rect 10045 17289 10057 17323
rect 10091 17320 10103 17323
rect 10686 17320 10692 17332
rect 10091 17292 10692 17320
rect 10091 17289 10103 17292
rect 10045 17283 10103 17289
rect 10686 17280 10692 17292
rect 10744 17280 10750 17332
rect 11333 17323 11391 17329
rect 11333 17289 11345 17323
rect 11379 17320 11391 17323
rect 11882 17320 11888 17332
rect 11379 17292 11888 17320
rect 11379 17289 11391 17292
rect 11333 17283 11391 17289
rect 11882 17280 11888 17292
rect 11940 17280 11946 17332
rect 14550 17280 14556 17332
rect 14608 17320 14614 17332
rect 14826 17320 14832 17332
rect 14608 17292 14832 17320
rect 14608 17280 14614 17292
rect 14826 17280 14832 17292
rect 14884 17320 14890 17332
rect 15838 17320 15844 17332
rect 14884 17292 15844 17320
rect 14884 17280 14890 17292
rect 15838 17280 15844 17292
rect 15896 17280 15902 17332
rect 16298 17280 16304 17332
rect 16356 17320 16362 17332
rect 16669 17323 16727 17329
rect 16669 17320 16681 17323
rect 16356 17292 16681 17320
rect 16356 17280 16362 17292
rect 16669 17289 16681 17292
rect 16715 17289 16727 17323
rect 16669 17283 16727 17289
rect 17678 17280 17684 17332
rect 17736 17320 17742 17332
rect 17957 17323 18015 17329
rect 17957 17320 17969 17323
rect 17736 17292 17969 17320
rect 17736 17280 17742 17292
rect 17957 17289 17969 17292
rect 18003 17289 18015 17323
rect 19886 17320 19892 17332
rect 19847 17292 19892 17320
rect 17957 17283 18015 17289
rect 19886 17280 19892 17292
rect 19944 17280 19950 17332
rect 6908 17255 6966 17261
rect 4816 17224 6592 17252
rect 1673 17187 1731 17193
rect 1673 17153 1685 17187
rect 1719 17184 1731 17187
rect 2222 17184 2228 17196
rect 1719 17156 2228 17184
rect 1719 17153 1731 17156
rect 1673 17147 1731 17153
rect 2222 17144 2228 17156
rect 2280 17144 2286 17196
rect 4154 17184 4160 17196
rect 4115 17156 4160 17184
rect 4154 17144 4160 17156
rect 4212 17144 4218 17196
rect 4249 17187 4307 17193
rect 4249 17153 4261 17187
rect 4295 17184 4307 17187
rect 4706 17184 4712 17196
rect 4295 17156 4712 17184
rect 4295 17153 4307 17156
rect 4249 17147 4307 17153
rect 4706 17144 4712 17156
rect 4764 17144 4770 17196
rect 4816 17193 4844 17224
rect 5074 17193 5080 17196
rect 4801 17187 4859 17193
rect 4801 17153 4813 17187
rect 4847 17153 4859 17187
rect 5068 17184 5080 17193
rect 5035 17156 5080 17184
rect 4801 17147 4859 17153
rect 5068 17147 5080 17156
rect 5132 17184 5138 17196
rect 5350 17184 5356 17196
rect 5132 17156 5356 17184
rect 5074 17144 5080 17147
rect 5132 17144 5138 17156
rect 5350 17144 5356 17156
rect 5408 17144 5414 17196
rect 6564 17193 6592 17224
rect 6908 17221 6920 17255
rect 6954 17252 6966 17255
rect 7558 17252 7564 17264
rect 6954 17224 7564 17252
rect 6954 17221 6966 17224
rect 6908 17215 6966 17221
rect 7558 17212 7564 17224
rect 7616 17212 7622 17264
rect 8472 17255 8530 17261
rect 8472 17221 8484 17255
rect 8518 17252 8530 17255
rect 11606 17252 11612 17264
rect 8518 17224 11612 17252
rect 8518 17221 8530 17224
rect 8472 17215 8530 17221
rect 11606 17212 11612 17224
rect 11664 17212 11670 17264
rect 12066 17252 12072 17264
rect 12027 17224 12072 17252
rect 12066 17212 12072 17224
rect 12124 17212 12130 17264
rect 16117 17255 16175 17261
rect 16117 17221 16129 17255
rect 16163 17252 16175 17255
rect 17402 17252 17408 17264
rect 16163 17224 17408 17252
rect 16163 17221 16175 17224
rect 16117 17215 16175 17221
rect 17402 17212 17408 17224
rect 17460 17212 17466 17264
rect 17770 17212 17776 17264
rect 17828 17252 17834 17264
rect 18325 17255 18383 17261
rect 18325 17252 18337 17255
rect 17828 17224 18337 17252
rect 17828 17212 17834 17224
rect 18325 17221 18337 17224
rect 18371 17221 18383 17255
rect 18325 17215 18383 17221
rect 6549 17187 6607 17193
rect 6549 17153 6561 17187
rect 6595 17184 6607 17187
rect 6638 17184 6644 17196
rect 6595 17156 6644 17184
rect 6595 17153 6607 17156
rect 6549 17147 6607 17153
rect 6638 17144 6644 17156
rect 6696 17144 6702 17196
rect 6730 17144 6736 17196
rect 6788 17184 6794 17196
rect 6788 17156 8064 17184
rect 6788 17144 6794 17156
rect 4433 17119 4491 17125
rect 4433 17085 4445 17119
rect 4479 17085 4491 17119
rect 4433 17079 4491 17085
rect 1486 16980 1492 16992
rect 1447 16952 1492 16980
rect 1486 16940 1492 16952
rect 1544 16940 1550 16992
rect 3234 16940 3240 16992
rect 3292 16980 3298 16992
rect 3789 16983 3847 16989
rect 3789 16980 3801 16983
rect 3292 16952 3801 16980
rect 3292 16940 3298 16952
rect 3789 16949 3801 16952
rect 3835 16949 3847 16983
rect 4448 16980 4476 17079
rect 8036 17048 8064 17156
rect 8294 17144 8300 17196
rect 8352 17184 8358 17196
rect 11790 17184 11796 17196
rect 8352 17156 11796 17184
rect 8352 17144 8358 17156
rect 11790 17144 11796 17156
rect 11848 17144 11854 17196
rect 11974 17184 11980 17196
rect 11935 17156 11980 17184
rect 11974 17144 11980 17156
rect 12032 17144 12038 17196
rect 12434 17144 12440 17196
rect 12492 17184 12498 17196
rect 12704 17187 12762 17193
rect 12492 17156 12537 17184
rect 12492 17144 12498 17156
rect 12704 17153 12716 17187
rect 12750 17184 12762 17187
rect 13078 17184 13084 17196
rect 12750 17156 13084 17184
rect 12750 17153 12762 17156
rect 12704 17147 12762 17153
rect 13078 17144 13084 17156
rect 13136 17144 13142 17196
rect 15033 17187 15091 17193
rect 15033 17153 15045 17187
rect 15079 17184 15091 17187
rect 15194 17184 15200 17196
rect 15079 17156 15200 17184
rect 15079 17153 15091 17156
rect 15033 17147 15091 17153
rect 15194 17144 15200 17156
rect 15252 17144 15258 17196
rect 15289 17187 15347 17193
rect 15289 17153 15301 17187
rect 15335 17184 15347 17187
rect 15746 17184 15752 17196
rect 15335 17156 15752 17184
rect 15335 17153 15347 17156
rect 15289 17147 15347 17153
rect 15746 17144 15752 17156
rect 15804 17144 15810 17196
rect 17034 17184 17040 17196
rect 16995 17156 17040 17184
rect 17034 17144 17040 17156
rect 17092 17144 17098 17196
rect 17862 17184 17868 17196
rect 17823 17156 17868 17184
rect 17862 17144 17868 17156
rect 17920 17144 17926 17196
rect 18230 17144 18236 17196
rect 18288 17184 18294 17196
rect 19705 17187 19763 17193
rect 19705 17184 19717 17187
rect 18288 17156 19717 17184
rect 18288 17144 18294 17156
rect 19705 17153 19717 17156
rect 19751 17153 19763 17187
rect 19705 17147 19763 17153
rect 20530 17144 20536 17196
rect 20588 17184 20594 17196
rect 21269 17187 21327 17193
rect 21269 17184 21281 17187
rect 20588 17156 21281 17184
rect 20588 17144 20594 17156
rect 21269 17153 21281 17156
rect 21315 17153 21327 17187
rect 21269 17147 21327 17153
rect 8202 17116 8208 17128
rect 8163 17088 8208 17116
rect 8202 17076 8208 17088
rect 8260 17076 8266 17128
rect 9766 17076 9772 17128
rect 9824 17116 9830 17128
rect 10137 17119 10195 17125
rect 10137 17116 10149 17119
rect 9824 17088 10149 17116
rect 9824 17076 9830 17088
rect 10137 17085 10149 17088
rect 10183 17085 10195 17119
rect 10137 17079 10195 17085
rect 10226 17076 10232 17128
rect 10284 17116 10290 17128
rect 10321 17119 10379 17125
rect 10321 17116 10333 17119
rect 10284 17088 10333 17116
rect 10284 17076 10290 17088
rect 10321 17085 10333 17088
rect 10367 17085 10379 17119
rect 10594 17116 10600 17128
rect 10555 17088 10600 17116
rect 10321 17079 10379 17085
rect 10594 17076 10600 17088
rect 10652 17076 10658 17128
rect 12158 17076 12164 17128
rect 12216 17116 12222 17128
rect 12216 17088 12261 17116
rect 12216 17076 12222 17088
rect 15378 17076 15384 17128
rect 15436 17116 15442 17128
rect 15841 17119 15899 17125
rect 15841 17116 15853 17119
rect 15436 17088 15853 17116
rect 15436 17076 15442 17088
rect 15841 17085 15853 17088
rect 15887 17085 15899 17119
rect 15841 17079 15899 17085
rect 16025 17119 16083 17125
rect 16025 17085 16037 17119
rect 16071 17085 16083 17119
rect 17126 17116 17132 17128
rect 17087 17088 17132 17116
rect 16025 17079 16083 17085
rect 10042 17048 10048 17060
rect 8036 17020 8248 17048
rect 6178 16980 6184 16992
rect 4448 16952 6184 16980
rect 3789 16943 3847 16949
rect 6178 16940 6184 16952
rect 6236 16940 6242 16992
rect 6546 16940 6552 16992
rect 6604 16980 6610 16992
rect 6822 16980 6828 16992
rect 6604 16952 6828 16980
rect 6604 16940 6610 16952
rect 6822 16940 6828 16952
rect 6880 16980 6886 16992
rect 7926 16980 7932 16992
rect 6880 16952 7932 16980
rect 6880 16940 6886 16952
rect 7926 16940 7932 16952
rect 7984 16980 7990 16992
rect 8021 16983 8079 16989
rect 8021 16980 8033 16983
rect 7984 16952 8033 16980
rect 7984 16940 7990 16952
rect 8021 16949 8033 16952
rect 8067 16949 8079 16983
rect 8220 16980 8248 17020
rect 9508 17020 10048 17048
rect 9508 16980 9536 17020
rect 10042 17008 10048 17020
rect 10100 17008 10106 17060
rect 13817 17051 13875 17057
rect 13817 17017 13829 17051
rect 13863 17048 13875 17051
rect 13998 17048 14004 17060
rect 13863 17020 14004 17048
rect 13863 17017 13875 17020
rect 13817 17011 13875 17017
rect 13998 17008 14004 17020
rect 14056 17048 14062 17060
rect 16040 17048 16068 17079
rect 17126 17076 17132 17088
rect 17184 17076 17190 17128
rect 17310 17116 17316 17128
rect 17271 17088 17316 17116
rect 17310 17076 17316 17088
rect 17368 17076 17374 17128
rect 17678 17076 17684 17128
rect 17736 17116 17742 17128
rect 18049 17119 18107 17125
rect 18049 17116 18061 17119
rect 17736 17088 18061 17116
rect 17736 17076 17742 17088
rect 18049 17085 18061 17088
rect 18095 17085 18107 17119
rect 18049 17079 18107 17085
rect 17497 17051 17555 17057
rect 17497 17048 17509 17051
rect 14056 17020 14412 17048
rect 16040 17020 17509 17048
rect 14056 17008 14062 17020
rect 8220 16952 9536 16980
rect 9585 16983 9643 16989
rect 8021 16943 8079 16949
rect 9585 16949 9597 16983
rect 9631 16980 9643 16983
rect 10134 16980 10140 16992
rect 9631 16952 10140 16980
rect 9631 16949 9643 16952
rect 9585 16943 9643 16949
rect 10134 16940 10140 16952
rect 10192 16940 10198 16992
rect 11146 16940 11152 16992
rect 11204 16980 11210 16992
rect 11609 16983 11667 16989
rect 11609 16980 11621 16983
rect 11204 16952 11621 16980
rect 11204 16940 11210 16952
rect 11609 16949 11621 16952
rect 11655 16949 11667 16983
rect 11609 16943 11667 16949
rect 13630 16940 13636 16992
rect 13688 16980 13694 16992
rect 13909 16983 13967 16989
rect 13909 16980 13921 16983
rect 13688 16952 13921 16980
rect 13688 16940 13694 16952
rect 13909 16949 13921 16952
rect 13955 16949 13967 16983
rect 14384 16980 14412 17020
rect 17497 17017 17509 17020
rect 17543 17017 17555 17051
rect 17497 17011 17555 17017
rect 14550 16980 14556 16992
rect 14384 16952 14556 16980
rect 13909 16943 13967 16949
rect 14550 16940 14556 16952
rect 14608 16940 14614 16992
rect 16485 16983 16543 16989
rect 16485 16949 16497 16983
rect 16531 16980 16543 16983
rect 19794 16980 19800 16992
rect 16531 16952 19800 16980
rect 16531 16949 16543 16952
rect 16485 16943 16543 16949
rect 19794 16940 19800 16952
rect 19852 16940 19858 16992
rect 21450 16980 21456 16992
rect 21411 16952 21456 16980
rect 21450 16940 21456 16952
rect 21508 16940 21514 16992
rect 1104 16890 21896 16912
rect 1104 16838 3549 16890
rect 3601 16838 3613 16890
rect 3665 16838 3677 16890
rect 3729 16838 3741 16890
rect 3793 16838 3805 16890
rect 3857 16838 8747 16890
rect 8799 16838 8811 16890
rect 8863 16838 8875 16890
rect 8927 16838 8939 16890
rect 8991 16838 9003 16890
rect 9055 16838 13945 16890
rect 13997 16838 14009 16890
rect 14061 16838 14073 16890
rect 14125 16838 14137 16890
rect 14189 16838 14201 16890
rect 14253 16838 19143 16890
rect 19195 16838 19207 16890
rect 19259 16838 19271 16890
rect 19323 16838 19335 16890
rect 19387 16838 19399 16890
rect 19451 16838 21896 16890
rect 1104 16816 21896 16838
rect 2225 16779 2283 16785
rect 2225 16745 2237 16779
rect 2271 16776 2283 16779
rect 2314 16776 2320 16788
rect 2271 16748 2320 16776
rect 2271 16745 2283 16748
rect 2225 16739 2283 16745
rect 2314 16736 2320 16748
rect 2372 16736 2378 16788
rect 4154 16736 4160 16788
rect 4212 16776 4218 16788
rect 4525 16779 4583 16785
rect 4525 16776 4537 16779
rect 4212 16748 4537 16776
rect 4212 16736 4218 16748
rect 4525 16745 4537 16748
rect 4571 16745 4583 16779
rect 4525 16739 4583 16745
rect 6365 16779 6423 16785
rect 6365 16745 6377 16779
rect 6411 16776 6423 16779
rect 6549 16779 6607 16785
rect 6549 16776 6561 16779
rect 6411 16748 6561 16776
rect 6411 16745 6423 16748
rect 6365 16739 6423 16745
rect 6549 16745 6561 16748
rect 6595 16776 6607 16779
rect 6638 16776 6644 16788
rect 6595 16748 6644 16776
rect 6595 16745 6607 16748
rect 6549 16739 6607 16745
rect 6638 16736 6644 16748
rect 6696 16736 6702 16788
rect 8202 16776 8208 16788
rect 8115 16748 8208 16776
rect 8202 16736 8208 16748
rect 8260 16776 8266 16788
rect 9309 16779 9367 16785
rect 9309 16776 9321 16779
rect 8260 16748 9321 16776
rect 8260 16736 8266 16748
rect 9309 16745 9321 16748
rect 9355 16776 9367 16779
rect 11793 16779 11851 16785
rect 9355 16748 10824 16776
rect 9355 16745 9367 16748
rect 9309 16739 9367 16745
rect 2958 16708 2964 16720
rect 2700 16680 2964 16708
rect 2700 16649 2728 16680
rect 2958 16668 2964 16680
rect 3016 16708 3022 16720
rect 3016 16680 6592 16708
rect 3016 16668 3022 16680
rect 6564 16652 6592 16680
rect 2685 16643 2743 16649
rect 2685 16609 2697 16643
rect 2731 16609 2743 16643
rect 2866 16640 2872 16652
rect 2827 16612 2872 16640
rect 2685 16603 2743 16609
rect 2866 16600 2872 16612
rect 2924 16600 2930 16652
rect 3973 16643 4031 16649
rect 3973 16609 3985 16643
rect 4019 16640 4031 16643
rect 5350 16640 5356 16652
rect 4019 16612 5356 16640
rect 4019 16609 4031 16612
rect 3973 16603 4031 16609
rect 5350 16600 5356 16612
rect 5408 16600 5414 16652
rect 6546 16600 6552 16652
rect 6604 16600 6610 16652
rect 6656 16649 6684 16736
rect 10796 16649 10824 16748
rect 11793 16745 11805 16779
rect 11839 16776 11851 16779
rect 11882 16776 11888 16788
rect 11839 16748 11888 16776
rect 11839 16745 11851 16748
rect 11793 16739 11851 16745
rect 11882 16736 11888 16748
rect 11940 16736 11946 16788
rect 13630 16776 13636 16788
rect 13188 16748 13636 16776
rect 11900 16649 11928 16736
rect 6641 16643 6699 16649
rect 6641 16609 6653 16643
rect 6687 16609 6699 16643
rect 6641 16603 6699 16609
rect 10781 16643 10839 16649
rect 10781 16609 10793 16643
rect 10827 16640 10839 16643
rect 11885 16643 11943 16649
rect 11885 16640 11897 16643
rect 10827 16612 11897 16640
rect 10827 16609 10839 16612
rect 10781 16603 10839 16609
rect 11885 16609 11897 16612
rect 11931 16609 11943 16643
rect 11885 16603 11943 16609
rect 1673 16575 1731 16581
rect 1673 16541 1685 16575
rect 1719 16541 1731 16575
rect 1673 16535 1731 16541
rect 2041 16575 2099 16581
rect 2041 16541 2053 16575
rect 2087 16572 2099 16575
rect 3234 16572 3240 16584
rect 2087 16544 3240 16572
rect 2087 16541 2099 16544
rect 2041 16535 2099 16541
rect 1688 16504 1716 16535
rect 3234 16532 3240 16544
rect 3292 16532 3298 16584
rect 4065 16575 4123 16581
rect 4065 16541 4077 16575
rect 4111 16572 4123 16575
rect 4154 16572 4160 16584
rect 4111 16544 4160 16572
rect 4111 16541 4123 16544
rect 4065 16535 4123 16541
rect 4154 16532 4160 16544
rect 4212 16532 4218 16584
rect 6178 16532 6184 16584
rect 6236 16572 6242 16584
rect 6897 16575 6955 16581
rect 6897 16572 6909 16575
rect 6236 16544 6909 16572
rect 6236 16532 6242 16544
rect 6897 16541 6909 16544
rect 6943 16541 6955 16575
rect 6897 16535 6955 16541
rect 10134 16532 10140 16584
rect 10192 16572 10198 16584
rect 10514 16575 10572 16581
rect 10514 16572 10526 16575
rect 10192 16544 10526 16572
rect 10192 16532 10198 16544
rect 10514 16541 10526 16544
rect 10560 16541 10572 16575
rect 10870 16572 10876 16584
rect 10831 16544 10876 16572
rect 10514 16535 10572 16541
rect 10870 16532 10876 16544
rect 10928 16532 10934 16584
rect 11238 16532 11244 16584
rect 11296 16532 11302 16584
rect 11790 16532 11796 16584
rect 11848 16572 11854 16584
rect 12141 16575 12199 16581
rect 12141 16572 12153 16575
rect 11848 16544 12153 16572
rect 11848 16532 11854 16544
rect 12141 16541 12153 16544
rect 12187 16572 12199 16575
rect 13188 16572 13216 16748
rect 13630 16736 13636 16748
rect 13688 16736 13694 16788
rect 13722 16736 13728 16788
rect 13780 16776 13786 16788
rect 13817 16779 13875 16785
rect 13817 16776 13829 16779
rect 13780 16748 13829 16776
rect 13780 16736 13786 16748
rect 13817 16745 13829 16748
rect 13863 16745 13875 16779
rect 13817 16739 13875 16745
rect 17221 16779 17279 16785
rect 17221 16745 17233 16779
rect 17267 16776 17279 16779
rect 17862 16776 17868 16788
rect 17267 16748 17868 16776
rect 17267 16745 17279 16748
rect 17221 16739 17279 16745
rect 13265 16711 13323 16717
rect 13265 16677 13277 16711
rect 13311 16677 13323 16711
rect 13538 16708 13544 16720
rect 13499 16680 13544 16708
rect 13265 16671 13323 16677
rect 13280 16640 13308 16671
rect 13538 16668 13544 16680
rect 13596 16668 13602 16720
rect 13832 16640 13860 16739
rect 17862 16736 17868 16748
rect 17920 16736 17926 16788
rect 18138 16736 18144 16788
rect 18196 16776 18202 16788
rect 18233 16779 18291 16785
rect 18233 16776 18245 16779
rect 18196 16748 18245 16776
rect 18196 16736 18202 16748
rect 18233 16745 18245 16748
rect 18279 16745 18291 16779
rect 20622 16776 20628 16788
rect 20583 16748 20628 16776
rect 18233 16739 18291 16745
rect 20622 16736 20628 16748
rect 20680 16736 20686 16788
rect 16117 16711 16175 16717
rect 16117 16677 16129 16711
rect 16163 16708 16175 16711
rect 16163 16680 16896 16708
rect 16163 16677 16175 16680
rect 16117 16671 16175 16677
rect 14093 16643 14151 16649
rect 14093 16640 14105 16643
rect 13280 16612 13492 16640
rect 13832 16612 14105 16640
rect 13354 16572 13360 16584
rect 12187 16544 13216 16572
rect 13315 16544 13360 16572
rect 12187 16541 12199 16544
rect 12141 16535 12199 16541
rect 13354 16532 13360 16544
rect 13412 16532 13418 16584
rect 2314 16504 2320 16516
rect 1688 16476 2320 16504
rect 2314 16464 2320 16476
rect 2372 16464 2378 16516
rect 2961 16507 3019 16513
rect 2961 16473 2973 16507
rect 3007 16504 3019 16507
rect 3421 16507 3479 16513
rect 3421 16504 3433 16507
rect 3007 16476 3433 16504
rect 3007 16473 3019 16476
rect 2961 16467 3019 16473
rect 3421 16473 3433 16476
rect 3467 16473 3479 16507
rect 3421 16467 3479 16473
rect 4890 16464 4896 16516
rect 4948 16504 4954 16516
rect 8386 16504 8392 16516
rect 4948 16476 8392 16504
rect 4948 16464 4954 16476
rect 8386 16464 8392 16476
rect 8444 16504 8450 16516
rect 10778 16504 10784 16516
rect 8444 16476 10784 16504
rect 8444 16464 8450 16476
rect 10778 16464 10784 16476
rect 10836 16464 10842 16516
rect 11256 16504 11284 16532
rect 12342 16504 12348 16516
rect 11256 16476 12348 16504
rect 12342 16464 12348 16476
rect 12400 16464 12406 16516
rect 13464 16504 13492 16612
rect 14093 16609 14105 16612
rect 14139 16609 14151 16643
rect 14093 16603 14151 16609
rect 16577 16643 16635 16649
rect 16577 16609 16589 16643
rect 16623 16609 16635 16643
rect 16868 16640 16896 16680
rect 16942 16668 16948 16720
rect 17000 16708 17006 16720
rect 17405 16711 17463 16717
rect 17405 16708 17417 16711
rect 17000 16680 17417 16708
rect 17000 16668 17006 16680
rect 17405 16677 17417 16680
rect 17451 16677 17463 16711
rect 17405 16671 17463 16677
rect 18782 16668 18788 16720
rect 18840 16708 18846 16720
rect 18840 16680 18920 16708
rect 18840 16668 18846 16680
rect 17957 16643 18015 16649
rect 16868 16612 17632 16640
rect 16577 16603 16635 16609
rect 13630 16532 13636 16584
rect 13688 16572 13694 16584
rect 16592 16572 16620 16603
rect 17494 16572 17500 16584
rect 13688 16544 17500 16572
rect 13688 16532 13694 16544
rect 17494 16532 17500 16544
rect 17552 16532 17558 16584
rect 17604 16572 17632 16612
rect 17957 16609 17969 16643
rect 18003 16609 18015 16643
rect 17957 16603 18015 16609
rect 17865 16575 17923 16581
rect 17865 16572 17877 16575
rect 17604 16544 17877 16572
rect 17865 16541 17877 16544
rect 17911 16541 17923 16575
rect 17972 16572 18000 16603
rect 18046 16600 18052 16652
rect 18104 16640 18110 16652
rect 18892 16649 18920 16680
rect 18693 16643 18751 16649
rect 18693 16640 18705 16643
rect 18104 16612 18705 16640
rect 18104 16600 18110 16612
rect 18693 16609 18705 16612
rect 18739 16609 18751 16643
rect 18693 16603 18751 16609
rect 18877 16643 18935 16649
rect 18877 16609 18889 16643
rect 18923 16609 18935 16643
rect 19610 16640 19616 16652
rect 18877 16603 18935 16609
rect 19306 16612 19616 16640
rect 18138 16572 18144 16584
rect 17972 16544 18144 16572
rect 17865 16535 17923 16541
rect 14338 16507 14396 16513
rect 14338 16504 14350 16507
rect 13464 16476 14350 16504
rect 14338 16473 14350 16476
rect 14384 16504 14396 16507
rect 17678 16504 17684 16516
rect 14384 16476 17684 16504
rect 14384 16473 14396 16476
rect 14338 16467 14396 16473
rect 17678 16464 17684 16476
rect 17736 16464 17742 16516
rect 17880 16504 17908 16535
rect 18138 16532 18144 16544
rect 18196 16532 18202 16584
rect 19306 16504 19334 16612
rect 19610 16600 19616 16612
rect 19668 16640 19674 16652
rect 20073 16643 20131 16649
rect 20073 16640 20085 16643
rect 19668 16612 20085 16640
rect 19668 16600 19674 16612
rect 20073 16609 20085 16612
rect 20119 16640 20131 16643
rect 20119 16612 20760 16640
rect 20119 16609 20131 16612
rect 20073 16603 20131 16609
rect 20732 16581 20760 16612
rect 20441 16575 20499 16581
rect 20441 16572 20453 16575
rect 17880 16476 19334 16504
rect 20272 16544 20453 16572
rect 1486 16436 1492 16448
rect 1447 16408 1492 16436
rect 1486 16396 1492 16408
rect 1544 16396 1550 16448
rect 2406 16436 2412 16448
rect 2367 16408 2412 16436
rect 2406 16396 2412 16408
rect 2464 16396 2470 16448
rect 3329 16439 3387 16445
rect 3329 16405 3341 16439
rect 3375 16436 3387 16439
rect 4157 16439 4215 16445
rect 4157 16436 4169 16439
rect 3375 16408 4169 16436
rect 3375 16405 3387 16408
rect 3329 16399 3387 16405
rect 4157 16405 4169 16408
rect 4203 16405 4215 16439
rect 8018 16436 8024 16448
rect 7979 16408 8024 16436
rect 4157 16399 4215 16405
rect 8018 16396 8024 16408
rect 8076 16396 8082 16448
rect 9214 16396 9220 16448
rect 9272 16436 9278 16448
rect 9401 16439 9459 16445
rect 9401 16436 9413 16439
rect 9272 16408 9413 16436
rect 9272 16396 9278 16408
rect 9401 16405 9413 16408
rect 9447 16405 9459 16439
rect 11054 16436 11060 16448
rect 11015 16408 11060 16436
rect 9401 16399 9459 16405
rect 11054 16396 11060 16408
rect 11112 16396 11118 16448
rect 11238 16396 11244 16448
rect 11296 16436 11302 16448
rect 15102 16436 15108 16448
rect 11296 16408 15108 16436
rect 11296 16396 11302 16408
rect 15102 16396 15108 16408
rect 15160 16396 15166 16448
rect 15378 16396 15384 16448
rect 15436 16436 15442 16448
rect 15473 16439 15531 16445
rect 15473 16436 15485 16439
rect 15436 16408 15485 16436
rect 15436 16396 15442 16408
rect 15473 16405 15485 16408
rect 15519 16405 15531 16439
rect 16390 16436 16396 16448
rect 16351 16408 16396 16436
rect 15473 16399 15531 16405
rect 16390 16396 16396 16408
rect 16448 16396 16454 16448
rect 16482 16396 16488 16448
rect 16540 16436 16546 16448
rect 16761 16439 16819 16445
rect 16761 16436 16773 16439
rect 16540 16408 16773 16436
rect 16540 16396 16546 16408
rect 16761 16405 16773 16408
rect 16807 16405 16819 16439
rect 16761 16399 16819 16405
rect 16853 16439 16911 16445
rect 16853 16405 16865 16439
rect 16899 16436 16911 16439
rect 17310 16436 17316 16448
rect 16899 16408 17316 16436
rect 16899 16405 16911 16408
rect 16853 16399 16911 16405
rect 17310 16396 17316 16408
rect 17368 16396 17374 16448
rect 17770 16436 17776 16448
rect 17731 16408 17776 16436
rect 17770 16396 17776 16408
rect 17828 16396 17834 16448
rect 18598 16436 18604 16448
rect 18559 16408 18604 16436
rect 18598 16396 18604 16408
rect 18656 16436 18662 16448
rect 20272 16445 20300 16544
rect 20441 16541 20453 16544
rect 20487 16541 20499 16575
rect 20441 16535 20499 16541
rect 20717 16575 20775 16581
rect 20717 16541 20729 16575
rect 20763 16541 20775 16575
rect 20717 16535 20775 16541
rect 20806 16532 20812 16584
rect 20864 16572 20870 16584
rect 21177 16575 21235 16581
rect 21177 16572 21189 16575
rect 20864 16544 21189 16572
rect 20864 16532 20870 16544
rect 21177 16541 21189 16544
rect 21223 16541 21235 16575
rect 21177 16535 21235 16541
rect 21269 16575 21327 16581
rect 21269 16541 21281 16575
rect 21315 16541 21327 16575
rect 21269 16535 21327 16541
rect 21284 16504 21312 16535
rect 20916 16476 21312 16504
rect 20916 16445 20944 16476
rect 20257 16439 20315 16445
rect 20257 16436 20269 16439
rect 18656 16408 20269 16436
rect 18656 16396 18662 16408
rect 20257 16405 20269 16408
rect 20303 16405 20315 16439
rect 20257 16399 20315 16405
rect 20901 16439 20959 16445
rect 20901 16405 20913 16439
rect 20947 16405 20959 16439
rect 20901 16399 20959 16405
rect 20990 16396 20996 16448
rect 21048 16436 21054 16448
rect 21450 16436 21456 16448
rect 21048 16408 21093 16436
rect 21411 16408 21456 16436
rect 21048 16396 21054 16408
rect 21450 16396 21456 16408
rect 21508 16396 21514 16448
rect 1104 16346 22056 16368
rect 1104 16294 6148 16346
rect 6200 16294 6212 16346
rect 6264 16294 6276 16346
rect 6328 16294 6340 16346
rect 6392 16294 6404 16346
rect 6456 16294 11346 16346
rect 11398 16294 11410 16346
rect 11462 16294 11474 16346
rect 11526 16294 11538 16346
rect 11590 16294 11602 16346
rect 11654 16294 16544 16346
rect 16596 16294 16608 16346
rect 16660 16294 16672 16346
rect 16724 16294 16736 16346
rect 16788 16294 16800 16346
rect 16852 16294 21742 16346
rect 21794 16294 21806 16346
rect 21858 16294 21870 16346
rect 21922 16294 21934 16346
rect 21986 16294 21998 16346
rect 22050 16294 22056 16346
rect 1104 16272 22056 16294
rect 2130 16232 2136 16244
rect 2091 16204 2136 16232
rect 2130 16192 2136 16204
rect 2188 16192 2194 16244
rect 2314 16192 2320 16244
rect 2372 16232 2378 16244
rect 2409 16235 2467 16241
rect 2409 16232 2421 16235
rect 2372 16204 2421 16232
rect 2372 16192 2378 16204
rect 2409 16201 2421 16204
rect 2455 16201 2467 16235
rect 2409 16195 2467 16201
rect 3605 16235 3663 16241
rect 3605 16201 3617 16235
rect 3651 16232 3663 16235
rect 4154 16232 4160 16244
rect 3651 16204 4160 16232
rect 3651 16201 3663 16204
rect 3605 16195 3663 16201
rect 4154 16192 4160 16204
rect 4212 16192 4218 16244
rect 4706 16192 4712 16244
rect 4764 16232 4770 16244
rect 4801 16235 4859 16241
rect 4801 16232 4813 16235
rect 4764 16204 4813 16232
rect 4764 16192 4770 16204
rect 4801 16201 4813 16204
rect 4847 16201 4859 16235
rect 4801 16195 4859 16201
rect 6181 16235 6239 16241
rect 6181 16201 6193 16235
rect 6227 16232 6239 16235
rect 6638 16232 6644 16244
rect 6227 16204 6644 16232
rect 6227 16201 6239 16204
rect 6181 16195 6239 16201
rect 3145 16167 3203 16173
rect 3145 16133 3157 16167
rect 3191 16164 3203 16167
rect 3789 16167 3847 16173
rect 3789 16164 3801 16167
rect 3191 16136 3801 16164
rect 3191 16133 3203 16136
rect 3145 16127 3203 16133
rect 3789 16133 3801 16136
rect 3835 16164 3847 16167
rect 3970 16164 3976 16176
rect 3835 16136 3976 16164
rect 3835 16133 3847 16136
rect 3789 16127 3847 16133
rect 3970 16124 3976 16136
rect 4028 16124 4034 16176
rect 1673 16099 1731 16105
rect 1673 16065 1685 16099
rect 1719 16065 1731 16099
rect 1673 16059 1731 16065
rect 1486 15892 1492 15904
rect 1447 15864 1492 15892
rect 1486 15852 1492 15864
rect 1544 15852 1550 15904
rect 1688 15892 1716 16059
rect 1946 16056 1952 16108
rect 2004 16096 2010 16108
rect 2041 16099 2099 16105
rect 2041 16096 2053 16099
rect 2004 16068 2053 16096
rect 2004 16056 2010 16068
rect 2041 16065 2053 16068
rect 2087 16065 2099 16099
rect 2314 16096 2320 16108
rect 2275 16068 2320 16096
rect 2041 16059 2099 16065
rect 2314 16056 2320 16068
rect 2372 16056 2378 16108
rect 2593 16099 2651 16105
rect 2593 16065 2605 16099
rect 2639 16096 2651 16099
rect 2774 16096 2780 16108
rect 2639 16068 2780 16096
rect 2639 16065 2651 16068
rect 2593 16059 2651 16065
rect 2774 16056 2780 16068
rect 2832 16096 2838 16108
rect 3237 16099 3295 16105
rect 2832 16068 2925 16096
rect 2832 16056 2838 16068
rect 3237 16065 3249 16099
rect 3283 16096 3295 16099
rect 4062 16096 4068 16108
rect 3283 16068 4068 16096
rect 3283 16065 3295 16068
rect 3237 16059 3295 16065
rect 4062 16056 4068 16068
rect 4120 16056 4126 16108
rect 5169 16099 5227 16105
rect 5169 16065 5181 16099
rect 5215 16096 5227 16099
rect 5442 16096 5448 16108
rect 5215 16068 5448 16096
rect 5215 16065 5227 16068
rect 5169 16059 5227 16065
rect 5442 16056 5448 16068
rect 5500 16056 5506 16108
rect 6380 16105 6408 16204
rect 6638 16192 6644 16204
rect 6696 16192 6702 16244
rect 9861 16235 9919 16241
rect 9861 16201 9873 16235
rect 9907 16201 9919 16235
rect 9861 16195 9919 16201
rect 10965 16235 11023 16241
rect 10965 16201 10977 16235
rect 11011 16232 11023 16235
rect 11146 16232 11152 16244
rect 11011 16204 11152 16232
rect 11011 16201 11023 16204
rect 10965 16195 11023 16201
rect 9876 16164 9904 16195
rect 11146 16192 11152 16204
rect 11204 16192 11210 16244
rect 11330 16232 11336 16244
rect 11291 16204 11336 16232
rect 11330 16192 11336 16204
rect 11388 16192 11394 16244
rect 11514 16192 11520 16244
rect 11572 16232 11578 16244
rect 12710 16232 12716 16244
rect 11572 16204 12716 16232
rect 11572 16192 11578 16204
rect 12710 16192 12716 16204
rect 12768 16192 12774 16244
rect 13722 16232 13728 16244
rect 13683 16204 13728 16232
rect 13722 16192 13728 16204
rect 13780 16192 13786 16244
rect 14642 16192 14648 16244
rect 14700 16232 14706 16244
rect 15102 16232 15108 16244
rect 14700 16204 15108 16232
rect 14700 16192 14706 16204
rect 15102 16192 15108 16204
rect 15160 16232 15166 16244
rect 16298 16232 16304 16244
rect 15160 16204 16304 16232
rect 15160 16192 15166 16204
rect 16298 16192 16304 16204
rect 16356 16192 16362 16244
rect 16390 16192 16396 16244
rect 16448 16232 16454 16244
rect 17129 16235 17187 16241
rect 17129 16232 17141 16235
rect 16448 16204 17141 16232
rect 16448 16192 16454 16204
rect 17129 16201 17141 16204
rect 17175 16201 17187 16235
rect 17129 16195 17187 16201
rect 17218 16192 17224 16244
rect 17276 16232 17282 16244
rect 17589 16235 17647 16241
rect 17589 16232 17601 16235
rect 17276 16204 17601 16232
rect 17276 16192 17282 16204
rect 17589 16201 17601 16204
rect 17635 16201 17647 16235
rect 17589 16195 17647 16201
rect 17954 16192 17960 16244
rect 18012 16232 18018 16244
rect 20530 16232 20536 16244
rect 18012 16204 18092 16232
rect 20491 16204 20536 16232
rect 18012 16192 18018 16204
rect 11238 16164 11244 16176
rect 9876 16136 11244 16164
rect 11238 16124 11244 16136
rect 11296 16124 11302 16176
rect 12728 16164 12756 16192
rect 16206 16164 16212 16176
rect 11992 16136 12296 16164
rect 12728 16136 16212 16164
rect 6365 16099 6423 16105
rect 6365 16065 6377 16099
rect 6411 16065 6423 16099
rect 6621 16099 6679 16105
rect 6621 16096 6633 16099
rect 6365 16059 6423 16065
rect 6472 16068 6633 16096
rect 2958 16028 2964 16040
rect 2919 16000 2964 16028
rect 2958 15988 2964 16000
rect 3016 15988 3022 16040
rect 5261 16031 5319 16037
rect 5261 15997 5273 16031
rect 5307 15997 5319 16031
rect 5261 15991 5319 15997
rect 1854 15960 1860 15972
rect 1815 15932 1860 15960
rect 1854 15920 1860 15932
rect 1912 15920 1918 15972
rect 5276 15960 5304 15991
rect 5350 15988 5356 16040
rect 5408 16028 5414 16040
rect 5408 16000 5453 16028
rect 5408 15988 5414 16000
rect 6270 15988 6276 16040
rect 6328 16028 6334 16040
rect 6472 16028 6500 16068
rect 6621 16065 6633 16068
rect 6667 16065 6679 16099
rect 6621 16059 6679 16065
rect 7190 16056 7196 16108
rect 7248 16096 7254 16108
rect 8202 16096 8208 16108
rect 7248 16068 8208 16096
rect 7248 16056 7254 16068
rect 8202 16056 8208 16068
rect 8260 16056 8266 16108
rect 9493 16099 9551 16105
rect 9493 16065 9505 16099
rect 9539 16096 9551 16099
rect 10042 16096 10048 16108
rect 9539 16068 10048 16096
rect 9539 16065 9551 16068
rect 9493 16059 9551 16065
rect 10042 16056 10048 16068
rect 10100 16056 10106 16108
rect 10134 16056 10140 16108
rect 10192 16096 10198 16108
rect 11992 16096 12020 16136
rect 10192 16068 12020 16096
rect 10192 16056 10198 16068
rect 12066 16056 12072 16108
rect 12124 16096 12130 16108
rect 12124 16068 12169 16096
rect 12124 16056 12130 16068
rect 9214 16028 9220 16040
rect 6328 16000 6500 16028
rect 9175 16000 9220 16028
rect 6328 15988 6334 16000
rect 9214 15988 9220 16000
rect 9272 15988 9278 16040
rect 9401 16031 9459 16037
rect 9401 15997 9413 16031
rect 9447 15997 9459 16031
rect 10686 16028 10692 16040
rect 10647 16000 10692 16028
rect 9401 15991 9459 15997
rect 6362 15960 6368 15972
rect 5276 15932 6368 15960
rect 6362 15920 6368 15932
rect 6420 15920 6426 15972
rect 9416 15960 9444 15991
rect 10686 15988 10692 16000
rect 10744 15988 10750 16040
rect 10873 16031 10931 16037
rect 10873 15997 10885 16031
rect 10919 16028 10931 16031
rect 11974 16028 11980 16040
rect 10919 16000 11980 16028
rect 10919 15997 10931 16000
rect 10873 15991 10931 15997
rect 11974 15988 11980 16000
rect 12032 15988 12038 16040
rect 12268 16037 12296 16136
rect 16206 16124 16212 16136
rect 16264 16124 16270 16176
rect 18064 16173 18092 16204
rect 20530 16192 20536 16204
rect 20588 16192 20594 16244
rect 20809 16235 20867 16241
rect 20809 16201 20821 16235
rect 20855 16232 20867 16235
rect 21174 16232 21180 16244
rect 20855 16204 21180 16232
rect 20855 16201 20867 16204
rect 20809 16195 20867 16201
rect 21174 16192 21180 16204
rect 21232 16192 21238 16244
rect 18049 16167 18107 16173
rect 18049 16133 18061 16167
rect 18095 16164 18107 16167
rect 18509 16167 18567 16173
rect 18509 16164 18521 16167
rect 18095 16136 18521 16164
rect 18095 16133 18107 16136
rect 18049 16127 18107 16133
rect 18509 16133 18521 16136
rect 18555 16164 18567 16167
rect 22370 16164 22376 16176
rect 18555 16136 22376 16164
rect 18555 16133 18567 16136
rect 18509 16127 18567 16133
rect 22370 16124 22376 16136
rect 22428 16124 22434 16176
rect 13722 16056 13728 16108
rect 13780 16096 13786 16108
rect 13817 16099 13875 16105
rect 13817 16096 13829 16099
rect 13780 16068 13829 16096
rect 13780 16056 13786 16068
rect 13817 16065 13829 16068
rect 13863 16065 13875 16099
rect 13817 16059 13875 16065
rect 13906 16056 13912 16108
rect 13964 16096 13970 16108
rect 14073 16099 14131 16105
rect 14073 16096 14085 16099
rect 13964 16068 14085 16096
rect 13964 16056 13970 16068
rect 14073 16065 14085 16068
rect 14119 16065 14131 16099
rect 14073 16059 14131 16065
rect 15470 16056 15476 16108
rect 15528 16096 15534 16108
rect 17957 16099 18015 16105
rect 15528 16068 17356 16096
rect 15528 16056 15534 16068
rect 17328 16037 17356 16068
rect 17957 16065 17969 16099
rect 18003 16096 18015 16099
rect 18782 16096 18788 16108
rect 18003 16068 18788 16096
rect 18003 16065 18015 16068
rect 17957 16059 18015 16065
rect 18782 16056 18788 16068
rect 18840 16056 18846 16108
rect 20254 16056 20260 16108
rect 20312 16096 20318 16108
rect 20349 16099 20407 16105
rect 20349 16096 20361 16099
rect 20312 16068 20361 16096
rect 20312 16056 20318 16068
rect 20349 16065 20361 16068
rect 20395 16065 20407 16099
rect 20349 16059 20407 16065
rect 20625 16099 20683 16105
rect 20625 16065 20637 16099
rect 20671 16065 20683 16099
rect 20898 16096 20904 16108
rect 20859 16068 20904 16096
rect 20625 16059 20683 16065
rect 12161 16031 12219 16037
rect 12161 15997 12173 16031
rect 12207 15997 12219 16031
rect 12161 15991 12219 15997
rect 12253 16031 12311 16037
rect 12253 15997 12265 16031
rect 12299 15997 12311 16031
rect 17221 16031 17279 16037
rect 17221 16028 17233 16031
rect 12253 15991 12311 15997
rect 16408 16000 17233 16028
rect 11701 15963 11759 15969
rect 11701 15960 11713 15963
rect 9416 15932 11713 15960
rect 11701 15929 11713 15932
rect 11747 15929 11759 15963
rect 12176 15960 12204 15991
rect 16408 15969 16436 16000
rect 17221 15997 17233 16000
rect 17267 15997 17279 16031
rect 17221 15991 17279 15997
rect 17313 16031 17371 16037
rect 17313 15997 17325 16031
rect 17359 16028 17371 16031
rect 17586 16028 17592 16040
rect 17359 16000 17592 16028
rect 17359 15997 17371 16000
rect 17313 15991 17371 15997
rect 16393 15963 16451 15969
rect 16393 15960 16405 15963
rect 11701 15923 11759 15929
rect 11992 15932 12204 15960
rect 15028 15932 16405 15960
rect 2314 15892 2320 15904
rect 1688 15864 2320 15892
rect 2314 15852 2320 15864
rect 2372 15852 2378 15904
rect 2958 15852 2964 15904
rect 3016 15892 3022 15904
rect 3326 15892 3332 15904
rect 3016 15864 3332 15892
rect 3016 15852 3022 15864
rect 3326 15852 3332 15864
rect 3384 15852 3390 15904
rect 7558 15852 7564 15904
rect 7616 15892 7622 15904
rect 7745 15895 7803 15901
rect 7745 15892 7757 15895
rect 7616 15864 7757 15892
rect 7616 15852 7622 15864
rect 7745 15861 7757 15864
rect 7791 15861 7803 15895
rect 7745 15855 7803 15861
rect 9858 15852 9864 15904
rect 9916 15892 9922 15904
rect 9953 15895 10011 15901
rect 9953 15892 9965 15895
rect 9916 15864 9965 15892
rect 9916 15852 9922 15864
rect 9953 15861 9965 15864
rect 9999 15861 10011 15895
rect 9953 15855 10011 15861
rect 10778 15852 10784 15904
rect 10836 15892 10842 15904
rect 11606 15892 11612 15904
rect 10836 15864 11612 15892
rect 10836 15852 10842 15864
rect 11606 15852 11612 15864
rect 11664 15892 11670 15904
rect 11992 15892 12020 15932
rect 11664 15864 12020 15892
rect 11664 15852 11670 15864
rect 12066 15852 12072 15904
rect 12124 15892 12130 15904
rect 12529 15895 12587 15901
rect 12529 15892 12541 15895
rect 12124 15864 12541 15892
rect 12124 15852 12130 15864
rect 12529 15861 12541 15864
rect 12575 15892 12587 15895
rect 12894 15892 12900 15904
rect 12575 15864 12900 15892
rect 12575 15861 12587 15864
rect 12529 15855 12587 15861
rect 12894 15852 12900 15864
rect 12952 15852 12958 15904
rect 13538 15852 13544 15904
rect 13596 15892 13602 15904
rect 15028 15892 15056 15932
rect 16393 15929 16405 15932
rect 16439 15929 16451 15963
rect 16393 15923 16451 15929
rect 16761 15963 16819 15969
rect 16761 15929 16773 15963
rect 16807 15960 16819 15963
rect 17034 15960 17040 15972
rect 16807 15932 17040 15960
rect 16807 15929 16819 15932
rect 16761 15923 16819 15929
rect 17034 15920 17040 15932
rect 17092 15920 17098 15972
rect 17236 15960 17264 15991
rect 17586 15988 17592 16000
rect 17644 15988 17650 16040
rect 18138 16028 18144 16040
rect 18099 16000 18144 16028
rect 18138 15988 18144 16000
rect 18196 15988 18202 16040
rect 20640 16028 20668 16059
rect 20898 16056 20904 16068
rect 20956 16056 20962 16108
rect 21269 16099 21327 16105
rect 21269 16065 21281 16099
rect 21315 16096 21327 16099
rect 21358 16096 21364 16108
rect 21315 16068 21364 16096
rect 21315 16065 21327 16068
rect 21269 16059 21327 16065
rect 21358 16056 21364 16068
rect 21416 16056 21422 16108
rect 20180 16000 20668 16028
rect 18598 15960 18604 15972
rect 17236 15932 18604 15960
rect 18598 15920 18604 15932
rect 18656 15920 18662 15972
rect 20180 15904 20208 16000
rect 21082 15960 21088 15972
rect 21043 15932 21088 15960
rect 21082 15920 21088 15932
rect 21140 15920 21146 15972
rect 15194 15892 15200 15904
rect 13596 15864 15056 15892
rect 15107 15864 15200 15892
rect 13596 15852 13602 15864
rect 15194 15852 15200 15864
rect 15252 15892 15258 15904
rect 15746 15892 15752 15904
rect 15252 15864 15752 15892
rect 15252 15852 15258 15864
rect 15746 15852 15752 15864
rect 15804 15852 15810 15904
rect 20162 15892 20168 15904
rect 20123 15864 20168 15892
rect 20162 15852 20168 15864
rect 20220 15852 20226 15904
rect 21450 15892 21456 15904
rect 21411 15864 21456 15892
rect 21450 15852 21456 15864
rect 21508 15852 21514 15904
rect 1104 15802 21896 15824
rect 1104 15750 3549 15802
rect 3601 15750 3613 15802
rect 3665 15750 3677 15802
rect 3729 15750 3741 15802
rect 3793 15750 3805 15802
rect 3857 15750 8747 15802
rect 8799 15750 8811 15802
rect 8863 15750 8875 15802
rect 8927 15750 8939 15802
rect 8991 15750 9003 15802
rect 9055 15750 13945 15802
rect 13997 15750 14009 15802
rect 14061 15750 14073 15802
rect 14125 15750 14137 15802
rect 14189 15750 14201 15802
rect 14253 15750 19143 15802
rect 19195 15750 19207 15802
rect 19259 15750 19271 15802
rect 19323 15750 19335 15802
rect 19387 15750 19399 15802
rect 19451 15750 21896 15802
rect 1104 15728 21896 15750
rect 1946 15688 1952 15700
rect 1907 15660 1952 15688
rect 1946 15648 1952 15660
rect 2004 15648 2010 15700
rect 2222 15688 2228 15700
rect 2183 15660 2228 15688
rect 2222 15648 2228 15660
rect 2280 15648 2286 15700
rect 5442 15688 5448 15700
rect 5403 15660 5448 15688
rect 5442 15648 5448 15660
rect 5500 15648 5506 15700
rect 6270 15688 6276 15700
rect 6231 15660 6276 15688
rect 6270 15648 6276 15660
rect 6328 15648 6334 15700
rect 6362 15648 6368 15700
rect 6420 15688 6426 15700
rect 8941 15691 8999 15697
rect 8941 15688 8953 15691
rect 6420 15660 8953 15688
rect 6420 15648 6426 15660
rect 8941 15657 8953 15660
rect 8987 15657 8999 15691
rect 10042 15688 10048 15700
rect 10003 15660 10048 15688
rect 8941 15651 8999 15657
rect 10042 15648 10048 15660
rect 10100 15648 10106 15700
rect 10870 15688 10876 15700
rect 10831 15660 10876 15688
rect 10870 15648 10876 15660
rect 10928 15648 10934 15700
rect 11054 15648 11060 15700
rect 11112 15688 11118 15700
rect 11793 15691 11851 15697
rect 11793 15688 11805 15691
rect 11112 15660 11805 15688
rect 11112 15648 11118 15660
rect 11793 15657 11805 15660
rect 11839 15657 11851 15691
rect 11974 15688 11980 15700
rect 11935 15660 11980 15688
rect 11793 15651 11851 15657
rect 2038 15580 2044 15632
rect 2096 15620 2102 15632
rect 2501 15623 2559 15629
rect 2501 15620 2513 15623
rect 2096 15592 2513 15620
rect 2096 15580 2102 15592
rect 2501 15589 2513 15592
rect 2547 15589 2559 15623
rect 6288 15620 6316 15648
rect 2501 15583 2559 15589
rect 5460 15592 6316 15620
rect 7837 15623 7895 15629
rect 5460 15564 5488 15592
rect 7837 15589 7849 15623
rect 7883 15620 7895 15623
rect 11514 15620 11520 15632
rect 7883 15592 11520 15620
rect 7883 15589 7895 15592
rect 7837 15583 7895 15589
rect 5442 15512 5448 15564
rect 5500 15512 5506 15564
rect 6089 15555 6147 15561
rect 6089 15521 6101 15555
rect 6135 15552 6147 15555
rect 6546 15552 6552 15564
rect 6135 15524 6552 15552
rect 6135 15521 6147 15524
rect 6089 15515 6147 15521
rect 6546 15512 6552 15524
rect 6604 15512 6610 15564
rect 1670 15484 1676 15496
rect 1631 15456 1676 15484
rect 1670 15444 1676 15456
rect 1728 15444 1734 15496
rect 2133 15487 2191 15493
rect 2133 15453 2145 15487
rect 2179 15453 2191 15487
rect 2406 15484 2412 15496
rect 2367 15456 2412 15484
rect 2133 15447 2191 15453
rect 2148 15416 2176 15447
rect 2406 15444 2412 15456
rect 2464 15444 2470 15496
rect 2685 15487 2743 15493
rect 2685 15453 2697 15487
rect 2731 15484 2743 15487
rect 2869 15487 2927 15493
rect 2869 15484 2881 15487
rect 2731 15456 2881 15484
rect 2731 15453 2743 15456
rect 2685 15447 2743 15453
rect 2869 15453 2881 15456
rect 2915 15484 2927 15487
rect 2915 15456 5856 15484
rect 2915 15453 2927 15456
rect 2869 15447 2927 15453
rect 3053 15419 3111 15425
rect 3053 15416 3065 15419
rect 2148 15388 3065 15416
rect 3053 15385 3065 15388
rect 3099 15416 3111 15419
rect 4614 15416 4620 15428
rect 3099 15388 4620 15416
rect 3099 15385 3111 15388
rect 3053 15379 3111 15385
rect 4614 15376 4620 15388
rect 4672 15376 4678 15428
rect 5828 15425 5856 15456
rect 6638 15444 6644 15496
rect 6696 15484 6702 15496
rect 7653 15487 7711 15493
rect 7653 15484 7665 15487
rect 6696 15456 7665 15484
rect 6696 15444 6702 15456
rect 7653 15453 7665 15456
rect 7699 15453 7711 15487
rect 7653 15447 7711 15453
rect 5813 15419 5871 15425
rect 5813 15385 5825 15419
rect 5859 15416 5871 15419
rect 6546 15416 6552 15428
rect 5859 15388 6552 15416
rect 5859 15385 5871 15388
rect 5813 15379 5871 15385
rect 6546 15376 6552 15388
rect 6604 15376 6610 15428
rect 7408 15419 7466 15425
rect 7408 15385 7420 15419
rect 7454 15416 7466 15419
rect 7742 15416 7748 15428
rect 7454 15388 7748 15416
rect 7454 15385 7466 15388
rect 7408 15379 7466 15385
rect 7742 15376 7748 15388
rect 7800 15376 7806 15428
rect 1486 15348 1492 15360
rect 1447 15320 1492 15348
rect 1486 15308 1492 15320
rect 1544 15308 1550 15360
rect 4522 15348 4528 15360
rect 4483 15320 4528 15348
rect 4522 15308 4528 15320
rect 4580 15308 4586 15360
rect 5905 15351 5963 15357
rect 5905 15317 5917 15351
rect 5951 15348 5963 15351
rect 7852 15348 7880 15583
rect 11514 15580 11520 15592
rect 11572 15580 11578 15632
rect 7926 15512 7932 15564
rect 7984 15552 7990 15564
rect 9493 15555 9551 15561
rect 9493 15552 9505 15555
rect 7984 15524 9505 15552
rect 7984 15512 7990 15524
rect 9493 15521 9505 15524
rect 9539 15521 9551 15555
rect 9493 15515 9551 15521
rect 10226 15512 10232 15564
rect 10284 15552 10290 15564
rect 10597 15555 10655 15561
rect 10597 15552 10609 15555
rect 10284 15524 10609 15552
rect 10284 15512 10290 15524
rect 10597 15521 10609 15524
rect 10643 15521 10655 15555
rect 11330 15552 11336 15564
rect 11291 15524 11336 15552
rect 10597 15515 10655 15521
rect 11330 15512 11336 15524
rect 11388 15512 11394 15564
rect 11425 15555 11483 15561
rect 11425 15521 11437 15555
rect 11471 15521 11483 15555
rect 11425 15515 11483 15521
rect 9306 15484 9312 15496
rect 9267 15456 9312 15484
rect 9306 15444 9312 15456
rect 9364 15444 9370 15496
rect 10134 15484 10140 15496
rect 9416 15456 10140 15484
rect 8202 15376 8208 15428
rect 8260 15416 8266 15428
rect 9416 15425 9444 15456
rect 10134 15444 10140 15456
rect 10192 15444 10198 15496
rect 11054 15444 11060 15496
rect 11112 15484 11118 15496
rect 11440 15484 11468 15515
rect 11112 15456 11468 15484
rect 11808 15484 11836 15651
rect 11974 15648 11980 15660
rect 12032 15648 12038 15700
rect 13722 15648 13728 15700
rect 13780 15688 13786 15700
rect 13817 15691 13875 15697
rect 13817 15688 13829 15691
rect 13780 15660 13829 15688
rect 13780 15648 13786 15660
rect 13817 15657 13829 15660
rect 13863 15657 13875 15691
rect 13817 15651 13875 15657
rect 12158 15512 12164 15564
rect 12216 15552 12222 15564
rect 12621 15555 12679 15561
rect 12621 15552 12633 15555
rect 12216 15524 12633 15552
rect 12216 15512 12222 15524
rect 12621 15521 12633 15524
rect 12667 15552 12679 15555
rect 13078 15552 13084 15564
rect 12667 15524 13084 15552
rect 12667 15521 12679 15524
rect 12621 15515 12679 15521
rect 13078 15512 13084 15524
rect 13136 15512 13142 15564
rect 13832 15552 13860 15651
rect 15470 15648 15476 15700
rect 15528 15688 15534 15700
rect 15565 15691 15623 15697
rect 15565 15688 15577 15691
rect 15528 15660 15577 15688
rect 15528 15648 15534 15660
rect 15565 15657 15577 15660
rect 15611 15657 15623 15691
rect 17037 15691 17095 15697
rect 15565 15651 15623 15657
rect 15948 15660 16988 15688
rect 14093 15555 14151 15561
rect 14093 15552 14105 15555
rect 13832 15524 14105 15552
rect 14093 15521 14105 15524
rect 14139 15521 14151 15555
rect 14093 15515 14151 15521
rect 12342 15484 12348 15496
rect 11808 15456 12204 15484
rect 12303 15456 12348 15484
rect 11112 15444 11118 15456
rect 9401 15419 9459 15425
rect 9401 15416 9413 15419
rect 8260 15388 9413 15416
rect 8260 15376 8266 15388
rect 9401 15385 9413 15388
rect 9447 15385 9459 15419
rect 9401 15379 9459 15385
rect 9953 15419 10011 15425
rect 9953 15385 9965 15419
rect 9999 15416 10011 15419
rect 10413 15419 10471 15425
rect 10413 15416 10425 15419
rect 9999 15388 10425 15416
rect 9999 15385 10011 15388
rect 9953 15379 10011 15385
rect 10413 15385 10425 15388
rect 10459 15385 10471 15419
rect 10413 15379 10471 15385
rect 11241 15419 11299 15425
rect 11241 15385 11253 15419
rect 11287 15416 11299 15419
rect 12066 15416 12072 15428
rect 11287 15388 12072 15416
rect 11287 15385 11299 15388
rect 11241 15379 11299 15385
rect 12066 15376 12072 15388
rect 12124 15376 12130 15428
rect 5951 15320 7880 15348
rect 5951 15317 5963 15320
rect 5905 15311 5963 15317
rect 9858 15308 9864 15360
rect 9916 15348 9922 15360
rect 10505 15351 10563 15357
rect 10505 15348 10517 15351
rect 9916 15320 10517 15348
rect 9916 15308 9922 15320
rect 10505 15317 10517 15320
rect 10551 15348 10563 15351
rect 10594 15348 10600 15360
rect 10551 15320 10600 15348
rect 10551 15317 10563 15320
rect 10505 15311 10563 15317
rect 10594 15308 10600 15320
rect 10652 15308 10658 15360
rect 11606 15308 11612 15360
rect 11664 15348 11670 15360
rect 11882 15348 11888 15360
rect 11664 15320 11888 15348
rect 11664 15308 11670 15320
rect 11882 15308 11888 15320
rect 11940 15308 11946 15360
rect 12176 15348 12204 15456
rect 12342 15444 12348 15456
rect 12400 15444 12406 15496
rect 12437 15487 12495 15493
rect 12437 15453 12449 15487
rect 12483 15484 12495 15487
rect 15948 15484 15976 15660
rect 16960 15620 16988 15660
rect 17037 15657 17049 15691
rect 17083 15688 17095 15691
rect 17126 15688 17132 15700
rect 17083 15660 17132 15688
rect 17083 15657 17095 15660
rect 17037 15651 17095 15657
rect 17126 15648 17132 15660
rect 17184 15648 17190 15700
rect 18138 15688 18144 15700
rect 17236 15660 18144 15688
rect 17236 15620 17264 15660
rect 18138 15648 18144 15660
rect 18196 15648 18202 15700
rect 20254 15688 20260 15700
rect 20215 15660 20260 15688
rect 20254 15648 20260 15660
rect 20312 15648 20318 15700
rect 20993 15691 21051 15697
rect 20993 15657 21005 15691
rect 21039 15688 21051 15691
rect 21266 15688 21272 15700
rect 21039 15660 21272 15688
rect 21039 15657 21051 15660
rect 20993 15651 21051 15657
rect 21266 15648 21272 15660
rect 21324 15648 21330 15700
rect 21453 15691 21511 15697
rect 21453 15657 21465 15691
rect 21499 15688 21511 15691
rect 21542 15688 21548 15700
rect 21499 15660 21548 15688
rect 21499 15657 21511 15660
rect 21453 15651 21511 15657
rect 21542 15648 21548 15660
rect 21600 15648 21606 15700
rect 21634 15620 21640 15632
rect 16960 15592 17264 15620
rect 17420 15592 21640 15620
rect 16942 15484 16948 15496
rect 12483 15456 15976 15484
rect 16903 15456 16948 15484
rect 12483 15453 12495 15456
rect 12437 15447 12495 15453
rect 12452 15348 12480 15447
rect 16942 15444 16948 15456
rect 17000 15444 17006 15496
rect 17420 15493 17448 15592
rect 21634 15580 21640 15592
rect 21692 15580 21698 15632
rect 17586 15552 17592 15564
rect 17547 15524 17592 15552
rect 17586 15512 17592 15524
rect 17644 15512 17650 15564
rect 18417 15555 18475 15561
rect 18417 15552 18429 15555
rect 17696 15524 18429 15552
rect 17405 15487 17463 15493
rect 17405 15453 17417 15487
rect 17451 15453 17463 15487
rect 17405 15447 17463 15453
rect 14366 15425 14372 15428
rect 14360 15379 14372 15425
rect 14424 15416 14430 15428
rect 16700 15419 16758 15425
rect 16700 15416 16712 15419
rect 14424 15388 14460 15416
rect 15488 15388 16712 15416
rect 14366 15376 14372 15379
rect 14424 15376 14430 15388
rect 15488 15357 15516 15388
rect 16700 15385 16712 15388
rect 16746 15416 16758 15419
rect 17696 15416 17724 15524
rect 18417 15521 18429 15524
rect 18463 15521 18475 15555
rect 18417 15515 18475 15521
rect 20717 15555 20775 15561
rect 20717 15521 20729 15555
rect 20763 15521 20775 15555
rect 20717 15515 20775 15521
rect 17954 15444 17960 15496
rect 18012 15484 18018 15496
rect 20073 15487 20131 15493
rect 20073 15484 20085 15487
rect 18012 15456 20085 15484
rect 18012 15444 18018 15456
rect 20073 15453 20085 15456
rect 20119 15453 20131 15487
rect 20732 15484 20760 15515
rect 20809 15487 20867 15493
rect 20809 15484 20821 15487
rect 20732 15456 20821 15484
rect 20073 15447 20131 15453
rect 20809 15453 20821 15456
rect 20855 15484 20867 15487
rect 20990 15484 20996 15496
rect 20855 15456 20996 15484
rect 20855 15453 20867 15456
rect 20809 15447 20867 15453
rect 20990 15444 20996 15456
rect 21048 15444 21054 15496
rect 21269 15487 21327 15493
rect 21269 15453 21281 15487
rect 21315 15453 21327 15487
rect 21269 15447 21327 15453
rect 16746 15388 17724 15416
rect 16746 15385 16758 15388
rect 16700 15379 16758 15385
rect 18138 15376 18144 15428
rect 18196 15416 18202 15428
rect 18325 15419 18383 15425
rect 18325 15416 18337 15419
rect 18196 15388 18337 15416
rect 18196 15376 18202 15388
rect 18325 15385 18337 15388
rect 18371 15416 18383 15419
rect 18874 15416 18880 15428
rect 18371 15388 18880 15416
rect 18371 15385 18383 15388
rect 18325 15379 18383 15385
rect 18874 15376 18880 15388
rect 18932 15376 18938 15428
rect 20714 15376 20720 15428
rect 20772 15416 20778 15428
rect 21284 15416 21312 15447
rect 22094 15416 22100 15428
rect 20772 15388 21312 15416
rect 21376 15388 22100 15416
rect 20772 15376 20778 15388
rect 12176 15320 12480 15348
rect 15473 15351 15531 15357
rect 15473 15317 15485 15351
rect 15519 15317 15531 15351
rect 15473 15311 15531 15317
rect 17497 15351 17555 15357
rect 17497 15317 17509 15351
rect 17543 15348 17555 15351
rect 17865 15351 17923 15357
rect 17865 15348 17877 15351
rect 17543 15320 17877 15348
rect 17543 15317 17555 15320
rect 17497 15311 17555 15317
rect 17865 15317 17877 15320
rect 17911 15317 17923 15351
rect 17865 15311 17923 15317
rect 18233 15351 18291 15357
rect 18233 15317 18245 15351
rect 18279 15348 18291 15351
rect 18414 15348 18420 15360
rect 18279 15320 18420 15348
rect 18279 15317 18291 15320
rect 18233 15311 18291 15317
rect 18414 15308 18420 15320
rect 18472 15348 18478 15360
rect 18693 15351 18751 15357
rect 18693 15348 18705 15351
rect 18472 15320 18705 15348
rect 18472 15308 18478 15320
rect 18693 15317 18705 15320
rect 18739 15348 18751 15351
rect 21376 15348 21404 15388
rect 22094 15376 22100 15388
rect 22152 15376 22158 15428
rect 18739 15320 21404 15348
rect 18739 15317 18751 15320
rect 18693 15311 18751 15317
rect 1104 15258 22056 15280
rect 1104 15206 6148 15258
rect 6200 15206 6212 15258
rect 6264 15206 6276 15258
rect 6328 15206 6340 15258
rect 6392 15206 6404 15258
rect 6456 15206 11346 15258
rect 11398 15206 11410 15258
rect 11462 15206 11474 15258
rect 11526 15206 11538 15258
rect 11590 15206 11602 15258
rect 11654 15206 16544 15258
rect 16596 15206 16608 15258
rect 16660 15206 16672 15258
rect 16724 15206 16736 15258
rect 16788 15206 16800 15258
rect 16852 15206 21742 15258
rect 21794 15206 21806 15258
rect 21858 15206 21870 15258
rect 21922 15206 21934 15258
rect 21986 15206 21998 15258
rect 22050 15206 22056 15258
rect 1104 15184 22056 15206
rect 1670 15104 1676 15156
rect 1728 15144 1734 15156
rect 1765 15147 1823 15153
rect 1765 15144 1777 15147
rect 1728 15116 1777 15144
rect 1728 15104 1734 15116
rect 1765 15113 1777 15116
rect 1811 15113 1823 15147
rect 1765 15107 1823 15113
rect 2041 15147 2099 15153
rect 2041 15113 2053 15147
rect 2087 15113 2099 15147
rect 2041 15107 2099 15113
rect 2056 15076 2084 15107
rect 2406 15104 2412 15156
rect 2464 15144 2470 15156
rect 2685 15147 2743 15153
rect 2685 15144 2697 15147
rect 2464 15116 2697 15144
rect 2464 15104 2470 15116
rect 2685 15113 2697 15116
rect 2731 15113 2743 15147
rect 3053 15147 3111 15153
rect 3053 15144 3065 15147
rect 2685 15107 2743 15113
rect 2792 15116 3065 15144
rect 2792 15076 2820 15116
rect 3053 15113 3065 15116
rect 3099 15144 3111 15147
rect 4430 15144 4436 15156
rect 3099 15116 4436 15144
rect 3099 15113 3111 15116
rect 3053 15107 3111 15113
rect 4430 15104 4436 15116
rect 4488 15104 4494 15156
rect 4522 15104 4528 15156
rect 4580 15144 4586 15156
rect 5169 15147 5227 15153
rect 5169 15144 5181 15147
rect 4580 15116 5181 15144
rect 4580 15104 4586 15116
rect 5169 15113 5181 15116
rect 5215 15113 5227 15147
rect 5169 15107 5227 15113
rect 6181 15147 6239 15153
rect 6181 15113 6193 15147
rect 6227 15144 6239 15147
rect 6638 15144 6644 15156
rect 6227 15116 6644 15144
rect 6227 15113 6239 15116
rect 6181 15107 6239 15113
rect 6638 15104 6644 15116
rect 6696 15144 6702 15156
rect 9122 15144 9128 15156
rect 6696 15116 9128 15144
rect 6696 15104 6702 15116
rect 1688 15048 2084 15076
rect 2240 15048 2820 15076
rect 1688 15017 1716 15048
rect 1673 15011 1731 15017
rect 1673 14977 1685 15011
rect 1719 14977 1731 15011
rect 1946 15008 1952 15020
rect 1907 14980 1952 15008
rect 1673 14971 1731 14977
rect 1946 14968 1952 14980
rect 2004 14968 2010 15020
rect 2240 15017 2268 15048
rect 5074 15036 5080 15088
rect 5132 15076 5138 15088
rect 5261 15079 5319 15085
rect 5261 15076 5273 15079
rect 5132 15048 5273 15076
rect 5132 15036 5138 15048
rect 5261 15045 5273 15048
rect 5307 15045 5319 15079
rect 5261 15039 5319 15045
rect 6457 15079 6515 15085
rect 6457 15045 6469 15079
rect 6503 15076 6515 15079
rect 6546 15076 6552 15088
rect 6503 15048 6552 15076
rect 6503 15045 6515 15048
rect 6457 15039 6515 15045
rect 6546 15036 6552 15048
rect 6604 15036 6610 15088
rect 2225 15011 2283 15017
rect 2225 14977 2237 15011
rect 2271 14977 2283 15011
rect 2225 14971 2283 14977
rect 2593 15011 2651 15017
rect 2593 14977 2605 15011
rect 2639 15008 2651 15011
rect 2774 15008 2780 15020
rect 2639 14980 2780 15008
rect 2639 14977 2651 14980
rect 2593 14971 2651 14977
rect 2774 14968 2780 14980
rect 2832 14968 2838 15020
rect 2869 15011 2927 15017
rect 2869 14977 2881 15011
rect 2915 15008 2927 15011
rect 4338 15008 4344 15020
rect 2915 14980 4016 15008
rect 4299 14980 4344 15008
rect 2915 14977 2927 14980
rect 2869 14971 2927 14977
rect 2409 14875 2467 14881
rect 2409 14841 2421 14875
rect 2455 14872 2467 14875
rect 2498 14872 2504 14884
rect 2455 14844 2504 14872
rect 2455 14841 2467 14844
rect 2409 14835 2467 14841
rect 2498 14832 2504 14844
rect 2556 14832 2562 14884
rect 3988 14881 4016 14980
rect 4338 14968 4344 14980
rect 4396 14968 4402 15020
rect 7558 15008 7564 15020
rect 4632 14980 7564 15008
rect 4632 14949 4660 14980
rect 7558 14968 7564 14980
rect 7616 14968 7622 15020
rect 7857 15011 7915 15017
rect 7857 14977 7869 15011
rect 7903 15008 7915 15011
rect 8018 15008 8024 15020
rect 7903 14980 8024 15008
rect 7903 14977 7915 14980
rect 7857 14971 7915 14977
rect 8018 14968 8024 14980
rect 8076 14968 8082 15020
rect 8128 15017 8156 15116
rect 9122 15104 9128 15116
rect 9180 15144 9186 15156
rect 9585 15147 9643 15153
rect 9585 15144 9597 15147
rect 9180 15116 9597 15144
rect 9180 15104 9186 15116
rect 9585 15113 9597 15116
rect 9631 15144 9643 15147
rect 11241 15147 11299 15153
rect 11241 15144 11253 15147
rect 9631 15116 11253 15144
rect 9631 15113 9643 15116
rect 9585 15107 9643 15113
rect 8570 15076 8576 15088
rect 8531 15048 8576 15076
rect 8570 15036 8576 15048
rect 8628 15036 8634 15088
rect 8113 15011 8171 15017
rect 8113 14977 8125 15011
rect 8159 14977 8171 15011
rect 8113 14971 8171 14977
rect 8202 14968 8208 15020
rect 8260 15008 8266 15020
rect 9784 15017 9812 15116
rect 11241 15113 11253 15116
rect 11287 15144 11299 15147
rect 11330 15144 11336 15156
rect 11287 15116 11336 15144
rect 11287 15113 11299 15116
rect 11241 15107 11299 15113
rect 11330 15104 11336 15116
rect 11388 15144 11394 15156
rect 13722 15144 13728 15156
rect 11388 15116 12434 15144
rect 13683 15116 13728 15144
rect 11388 15104 11394 15116
rect 12406 15076 12434 15116
rect 13722 15104 13728 15116
rect 13780 15144 13786 15156
rect 15381 15147 15439 15153
rect 15381 15144 15393 15147
rect 13780 15116 15393 15144
rect 13780 15104 13786 15116
rect 12406 15048 12940 15076
rect 8481 15011 8539 15017
rect 8481 15008 8493 15011
rect 8260 14980 8493 15008
rect 8260 14968 8266 14980
rect 8481 14977 8493 14980
rect 8527 14977 8539 15011
rect 8481 14971 8539 14977
rect 9769 15011 9827 15017
rect 9769 14977 9781 15011
rect 9815 14977 9827 15011
rect 9769 14971 9827 14977
rect 10036 15011 10094 15017
rect 10036 14977 10048 15011
rect 10082 15008 10094 15011
rect 10318 15008 10324 15020
rect 10082 14980 10324 15008
rect 10082 14977 10094 14980
rect 10036 14971 10094 14977
rect 10318 14968 10324 14980
rect 10376 14968 10382 15020
rect 12641 15011 12699 15017
rect 12641 14977 12653 15011
rect 12687 15008 12699 15011
rect 12802 15008 12808 15020
rect 12687 14980 12808 15008
rect 12687 14977 12699 14980
rect 12641 14971 12699 14977
rect 12802 14968 12808 14980
rect 12860 14968 12866 15020
rect 12912 15017 12940 15048
rect 12897 15011 12955 15017
rect 12897 14977 12909 15011
rect 12943 15008 12955 15011
rect 13722 15008 13728 15020
rect 12943 14980 13728 15008
rect 12943 14977 12955 14980
rect 12897 14971 12955 14977
rect 13722 14968 13728 14980
rect 13780 14968 13786 15020
rect 15212 15017 15240 15116
rect 15381 15113 15393 15116
rect 15427 15144 15439 15147
rect 15470 15144 15476 15156
rect 15427 15116 15476 15144
rect 15427 15113 15439 15116
rect 15381 15107 15439 15113
rect 15470 15104 15476 15116
rect 15528 15144 15534 15156
rect 16942 15144 16948 15156
rect 15528 15116 16948 15144
rect 15528 15104 15534 15116
rect 16942 15104 16948 15116
rect 17000 15104 17006 15156
rect 17313 15147 17371 15153
rect 17313 15113 17325 15147
rect 17359 15144 17371 15147
rect 18601 15147 18659 15153
rect 18601 15144 18613 15147
rect 17359 15116 18613 15144
rect 17359 15113 17371 15116
rect 17313 15107 17371 15113
rect 18601 15113 18613 15116
rect 18647 15113 18659 15147
rect 20714 15144 20720 15156
rect 20675 15116 20720 15144
rect 18601 15107 18659 15113
rect 20714 15104 20720 15116
rect 20772 15104 20778 15156
rect 20898 15104 20904 15156
rect 20956 15144 20962 15156
rect 20993 15147 21051 15153
rect 20993 15144 21005 15147
rect 20956 15116 21005 15144
rect 20956 15104 20962 15116
rect 20993 15113 21005 15116
rect 21039 15113 21051 15147
rect 20993 15107 21051 15113
rect 17865 15079 17923 15085
rect 17865 15045 17877 15079
rect 17911 15076 17923 15079
rect 18138 15076 18144 15088
rect 17911 15048 18144 15076
rect 17911 15045 17923 15048
rect 17865 15039 17923 15045
rect 18138 15036 18144 15048
rect 18196 15036 18202 15088
rect 14941 15011 14999 15017
rect 14941 14977 14953 15011
rect 14987 15008 14999 15011
rect 15197 15011 15255 15017
rect 14987 14980 15148 15008
rect 14987 14977 14999 14980
rect 14941 14971 14999 14977
rect 4433 14943 4491 14949
rect 4433 14909 4445 14943
rect 4479 14909 4491 14943
rect 4433 14903 4491 14909
rect 4617 14943 4675 14949
rect 4617 14909 4629 14943
rect 4663 14909 4675 14943
rect 5350 14940 5356 14952
rect 5311 14912 5356 14940
rect 4617 14903 4675 14909
rect 3973 14875 4031 14881
rect 3973 14841 3985 14875
rect 4019 14841 4031 14875
rect 4448 14872 4476 14903
rect 5350 14900 5356 14912
rect 5408 14900 5414 14952
rect 8297 14943 8355 14949
rect 8297 14909 8309 14943
rect 8343 14909 8355 14943
rect 15120 14940 15148 14980
rect 15197 14977 15209 15011
rect 15243 14977 15255 15011
rect 18966 15008 18972 15020
rect 18927 14980 18972 15008
rect 15197 14971 15255 14977
rect 18966 14968 18972 14980
rect 19024 14968 19030 15020
rect 19518 14968 19524 15020
rect 19576 15008 19582 15020
rect 20533 15011 20591 15017
rect 20533 15008 20545 15011
rect 19576 14980 20545 15008
rect 19576 14968 19582 14980
rect 20533 14977 20545 14980
rect 20579 14977 20591 15011
rect 20533 14971 20591 14977
rect 20809 15011 20867 15017
rect 20809 14977 20821 15011
rect 20855 14977 20867 15011
rect 20809 14971 20867 14977
rect 15378 14940 15384 14952
rect 15120 14912 15384 14940
rect 8297 14903 8355 14909
rect 4890 14872 4896 14884
rect 4448 14844 4896 14872
rect 3973 14835 4031 14841
rect 4890 14832 4896 14844
rect 4948 14832 4954 14884
rect 5534 14832 5540 14884
rect 5592 14872 5598 14884
rect 5592 14844 6868 14872
rect 5592 14832 5598 14844
rect 1486 14804 1492 14816
rect 1447 14776 1492 14804
rect 1486 14764 1492 14776
rect 1544 14764 1550 14816
rect 4154 14764 4160 14816
rect 4212 14804 4218 14816
rect 4801 14807 4859 14813
rect 4801 14804 4813 14807
rect 4212 14776 4813 14804
rect 4212 14764 4218 14776
rect 4801 14773 4813 14776
rect 4847 14773 4859 14807
rect 6730 14804 6736 14816
rect 6691 14776 6736 14804
rect 4801 14767 4859 14773
rect 6730 14764 6736 14776
rect 6788 14764 6794 14816
rect 6840 14804 6868 14844
rect 8110 14832 8116 14884
rect 8168 14872 8174 14884
rect 8312 14872 8340 14903
rect 15378 14900 15384 14912
rect 15436 14900 15442 14952
rect 15746 14900 15752 14952
rect 15804 14940 15810 14952
rect 17037 14943 17095 14949
rect 17037 14940 17049 14943
rect 15804 14912 17049 14940
rect 15804 14900 15810 14912
rect 17037 14909 17049 14912
rect 17083 14909 17095 14943
rect 17218 14940 17224 14952
rect 17179 14912 17224 14940
rect 17037 14903 17095 14909
rect 17218 14900 17224 14912
rect 17276 14900 17282 14952
rect 19058 14940 19064 14952
rect 19019 14912 19064 14940
rect 19058 14900 19064 14912
rect 19116 14900 19122 14952
rect 19153 14943 19211 14949
rect 19153 14909 19165 14943
rect 19199 14909 19211 14943
rect 20824 14940 20852 14971
rect 20898 14968 20904 15020
rect 20956 15008 20962 15020
rect 21269 15011 21327 15017
rect 21269 15008 21281 15011
rect 20956 14980 21281 15008
rect 20956 14968 20962 14980
rect 21269 14977 21281 14980
rect 21315 14977 21327 15011
rect 21269 14971 21327 14977
rect 20824 14912 21220 14940
rect 19153 14903 19211 14909
rect 8168 14844 8340 14872
rect 11149 14875 11207 14881
rect 8168 14832 8174 14844
rect 11149 14841 11161 14875
rect 11195 14872 11207 14875
rect 11698 14872 11704 14884
rect 11195 14844 11704 14872
rect 11195 14841 11207 14844
rect 11149 14835 11207 14841
rect 11698 14832 11704 14844
rect 11756 14832 11762 14884
rect 17681 14875 17739 14881
rect 17681 14841 17693 14875
rect 17727 14872 17739 14875
rect 17954 14872 17960 14884
rect 17727 14844 17960 14872
rect 17727 14841 17739 14844
rect 17681 14835 17739 14841
rect 17954 14832 17960 14844
rect 18012 14832 18018 14884
rect 18690 14832 18696 14884
rect 18748 14872 18754 14884
rect 19168 14872 19196 14903
rect 18748 14844 19196 14872
rect 18748 14832 18754 14844
rect 21192 14816 21220 14912
rect 8294 14804 8300 14816
rect 6840 14776 8300 14804
rect 8294 14764 8300 14776
rect 8352 14764 8358 14816
rect 8662 14764 8668 14816
rect 8720 14804 8726 14816
rect 8941 14807 8999 14813
rect 8941 14804 8953 14807
rect 8720 14776 8953 14804
rect 8720 14764 8726 14776
rect 8941 14773 8953 14776
rect 8987 14773 8999 14807
rect 11514 14804 11520 14816
rect 11475 14776 11520 14804
rect 8941 14767 8999 14773
rect 11514 14764 11520 14776
rect 11572 14764 11578 14816
rect 12986 14764 12992 14816
rect 13044 14804 13050 14816
rect 13817 14807 13875 14813
rect 13817 14804 13829 14807
rect 13044 14776 13829 14804
rect 13044 14764 13050 14776
rect 13817 14773 13829 14776
rect 13863 14773 13875 14807
rect 21174 14804 21180 14816
rect 21135 14776 21180 14804
rect 13817 14767 13875 14773
rect 21174 14764 21180 14776
rect 21232 14764 21238 14816
rect 21450 14804 21456 14816
rect 21411 14776 21456 14804
rect 21450 14764 21456 14776
rect 21508 14764 21514 14816
rect 1104 14714 21896 14736
rect 1104 14662 3549 14714
rect 3601 14662 3613 14714
rect 3665 14662 3677 14714
rect 3729 14662 3741 14714
rect 3793 14662 3805 14714
rect 3857 14662 8747 14714
rect 8799 14662 8811 14714
rect 8863 14662 8875 14714
rect 8927 14662 8939 14714
rect 8991 14662 9003 14714
rect 9055 14662 13945 14714
rect 13997 14662 14009 14714
rect 14061 14662 14073 14714
rect 14125 14662 14137 14714
rect 14189 14662 14201 14714
rect 14253 14662 19143 14714
rect 19195 14662 19207 14714
rect 19259 14662 19271 14714
rect 19323 14662 19335 14714
rect 19387 14662 19399 14714
rect 19451 14662 21896 14714
rect 1104 14640 21896 14662
rect 1946 14560 1952 14612
rect 2004 14600 2010 14612
rect 2869 14603 2927 14609
rect 2869 14600 2881 14603
rect 2004 14572 2881 14600
rect 2004 14560 2010 14572
rect 2869 14569 2881 14572
rect 2915 14569 2927 14603
rect 2869 14563 2927 14569
rect 4338 14560 4344 14612
rect 4396 14600 4402 14612
rect 4525 14603 4583 14609
rect 4525 14600 4537 14603
rect 4396 14572 4537 14600
rect 4396 14560 4402 14572
rect 4525 14569 4537 14572
rect 4571 14569 4583 14603
rect 7742 14600 7748 14612
rect 4525 14563 4583 14569
rect 6380 14572 7748 14600
rect 4706 14492 4712 14544
rect 4764 14532 4770 14544
rect 5350 14532 5356 14544
rect 4764 14504 5356 14532
rect 4764 14492 4770 14504
rect 5350 14492 5356 14504
rect 5408 14532 5414 14544
rect 5408 14504 5856 14532
rect 5408 14492 5414 14504
rect 3973 14467 4031 14473
rect 3973 14433 3985 14467
rect 4019 14464 4031 14467
rect 5442 14464 5448 14476
rect 4019 14436 5448 14464
rect 4019 14433 4031 14436
rect 3973 14427 4031 14433
rect 5442 14424 5448 14436
rect 5500 14424 5506 14476
rect 5828 14473 5856 14504
rect 5813 14467 5871 14473
rect 5813 14433 5825 14467
rect 5859 14464 5871 14467
rect 6380 14464 6408 14572
rect 7742 14560 7748 14572
rect 7800 14560 7806 14612
rect 9122 14600 9128 14612
rect 9083 14572 9128 14600
rect 9122 14560 9128 14572
rect 9180 14560 9186 14612
rect 10689 14603 10747 14609
rect 10689 14569 10701 14603
rect 10735 14600 10747 14603
rect 11054 14600 11060 14612
rect 10735 14572 11060 14600
rect 10735 14569 10747 14572
rect 10689 14563 10747 14569
rect 11054 14560 11060 14572
rect 11112 14560 11118 14612
rect 11330 14600 11336 14612
rect 11291 14572 11336 14600
rect 11330 14560 11336 14572
rect 11388 14560 11394 14612
rect 13722 14560 13728 14612
rect 13780 14600 13786 14612
rect 13817 14603 13875 14609
rect 13817 14600 13829 14603
rect 13780 14572 13829 14600
rect 13780 14560 13786 14572
rect 13817 14569 13829 14572
rect 13863 14569 13875 14603
rect 13817 14563 13875 14569
rect 14093 14603 14151 14609
rect 14093 14569 14105 14603
rect 14139 14600 14151 14603
rect 14366 14600 14372 14612
rect 14139 14572 14372 14600
rect 14139 14569 14151 14572
rect 14093 14563 14151 14569
rect 14366 14560 14372 14572
rect 14424 14560 14430 14612
rect 16853 14603 16911 14609
rect 14568 14572 15608 14600
rect 5859 14436 6408 14464
rect 7837 14467 7895 14473
rect 5859 14433 5871 14436
rect 5813 14427 5871 14433
rect 7837 14433 7849 14467
rect 7883 14464 7895 14467
rect 8570 14464 8576 14476
rect 7883 14436 8576 14464
rect 7883 14433 7895 14436
rect 7837 14427 7895 14433
rect 8570 14424 8576 14436
rect 8628 14424 8634 14476
rect 9140 14464 9168 14560
rect 9309 14467 9367 14473
rect 9309 14464 9321 14467
rect 9140 14436 9321 14464
rect 9309 14433 9321 14436
rect 9355 14433 9367 14467
rect 11348 14464 11376 14560
rect 12897 14535 12955 14541
rect 12897 14501 12909 14535
rect 12943 14501 12955 14535
rect 12897 14495 12955 14501
rect 11517 14467 11575 14473
rect 11517 14464 11529 14467
rect 11348 14436 11529 14464
rect 9309 14427 9367 14433
rect 11517 14433 11529 14436
rect 11563 14433 11575 14467
rect 12912 14464 12940 14495
rect 13906 14492 13912 14544
rect 13964 14532 13970 14544
rect 14568 14532 14596 14572
rect 13964 14504 14596 14532
rect 13964 14492 13970 14504
rect 15470 14464 15476 14476
rect 12912 14436 14504 14464
rect 15431 14436 15476 14464
rect 11517 14427 11575 14433
rect 1673 14399 1731 14405
rect 1673 14365 1685 14399
rect 1719 14396 1731 14399
rect 1762 14396 1768 14408
rect 1719 14368 1768 14396
rect 1719 14365 1731 14368
rect 1673 14359 1731 14365
rect 1762 14356 1768 14368
rect 1820 14356 1826 14408
rect 2038 14396 2044 14408
rect 1999 14368 2044 14396
rect 2038 14356 2044 14368
rect 2096 14356 2102 14408
rect 3053 14399 3111 14405
rect 3053 14365 3065 14399
rect 3099 14396 3111 14399
rect 3418 14396 3424 14408
rect 3099 14368 3424 14396
rect 3099 14365 3111 14368
rect 3053 14359 3111 14365
rect 3418 14356 3424 14368
rect 3476 14356 3482 14408
rect 4154 14396 4160 14408
rect 4115 14368 4160 14396
rect 4154 14356 4160 14368
rect 4212 14356 4218 14408
rect 5534 14396 5540 14408
rect 5495 14368 5540 14396
rect 5534 14356 5540 14368
rect 5592 14356 5598 14408
rect 6638 14356 6644 14408
rect 6696 14396 6702 14408
rect 7377 14399 7435 14405
rect 7377 14396 7389 14399
rect 6696 14368 7389 14396
rect 6696 14356 6702 14368
rect 7377 14365 7389 14368
rect 7423 14365 7435 14399
rect 7377 14359 7435 14365
rect 7466 14356 7472 14408
rect 7524 14396 7530 14408
rect 7929 14399 7987 14405
rect 7929 14396 7941 14399
rect 7524 14368 7941 14396
rect 7524 14356 7530 14368
rect 7929 14365 7941 14368
rect 7975 14365 7987 14399
rect 7929 14359 7987 14365
rect 8021 14399 8079 14405
rect 8021 14365 8033 14399
rect 8067 14396 8079 14399
rect 8294 14396 8300 14408
rect 8067 14368 8300 14396
rect 8067 14365 8079 14368
rect 8021 14359 8079 14365
rect 8294 14356 8300 14368
rect 8352 14356 8358 14408
rect 14476 14396 14504 14436
rect 15470 14424 15476 14436
rect 15528 14424 15534 14476
rect 15580 14464 15608 14572
rect 16853 14569 16865 14603
rect 16899 14600 16911 14603
rect 17218 14600 17224 14612
rect 16899 14572 17224 14600
rect 16899 14569 16911 14572
rect 16853 14563 16911 14569
rect 17218 14560 17224 14572
rect 17276 14560 17282 14612
rect 19058 14560 19064 14612
rect 19116 14600 19122 14612
rect 19245 14603 19303 14609
rect 19245 14600 19257 14603
rect 19116 14572 19257 14600
rect 19116 14560 19122 14572
rect 19245 14569 19257 14572
rect 19291 14569 19303 14603
rect 20990 14600 20996 14612
rect 19245 14563 19303 14569
rect 19628 14572 20996 14600
rect 16209 14467 16267 14473
rect 16209 14464 16221 14467
rect 15580 14436 16221 14464
rect 16209 14433 16221 14436
rect 16255 14464 16267 14467
rect 18690 14464 18696 14476
rect 16255 14436 18696 14464
rect 16255 14433 16267 14436
rect 16209 14427 16267 14433
rect 18690 14424 18696 14436
rect 18748 14424 18754 14476
rect 19628 14464 19656 14572
rect 20990 14560 20996 14572
rect 21048 14560 21054 14612
rect 20809 14535 20867 14541
rect 20809 14501 20821 14535
rect 20855 14501 20867 14535
rect 20809 14495 20867 14501
rect 19794 14464 19800 14476
rect 18800 14436 19656 14464
rect 19755 14436 19800 14464
rect 15206 14399 15264 14405
rect 15206 14396 15218 14399
rect 8404 14368 14412 14396
rect 14476 14368 15218 14396
rect 5629 14331 5687 14337
rect 5629 14297 5641 14331
rect 5675 14328 5687 14331
rect 5675 14300 6684 14328
rect 5675 14297 5687 14300
rect 5629 14291 5687 14297
rect 1486 14260 1492 14272
rect 1447 14232 1492 14260
rect 1486 14220 1492 14232
rect 1544 14220 1550 14272
rect 1854 14260 1860 14272
rect 1815 14232 1860 14260
rect 1854 14220 1860 14232
rect 1912 14220 1918 14272
rect 4065 14263 4123 14269
rect 4065 14229 4077 14263
rect 4111 14260 4123 14263
rect 4522 14260 4528 14272
rect 4111 14232 4528 14260
rect 4111 14229 4123 14232
rect 4065 14223 4123 14229
rect 4522 14220 4528 14232
rect 4580 14220 4586 14272
rect 5169 14263 5227 14269
rect 5169 14229 5181 14263
rect 5215 14260 5227 14263
rect 5350 14260 5356 14272
rect 5215 14232 5356 14260
rect 5215 14229 5227 14232
rect 5169 14223 5227 14229
rect 5350 14220 5356 14232
rect 5408 14220 5414 14272
rect 5994 14260 6000 14272
rect 5955 14232 6000 14260
rect 5994 14220 6000 14232
rect 6052 14220 6058 14272
rect 6656 14260 6684 14300
rect 6730 14288 6736 14340
rect 6788 14328 6794 14340
rect 7110 14331 7168 14337
rect 7110 14328 7122 14331
rect 6788 14300 7122 14328
rect 6788 14288 6794 14300
rect 7110 14297 7122 14300
rect 7156 14297 7168 14331
rect 7110 14291 7168 14297
rect 7484 14260 7512 14356
rect 8404 14269 8432 14368
rect 9576 14331 9634 14337
rect 9576 14297 9588 14331
rect 9622 14328 9634 14331
rect 10042 14328 10048 14340
rect 9622 14300 10048 14328
rect 9622 14297 9634 14300
rect 9576 14291 9634 14297
rect 10042 14288 10048 14300
rect 10100 14328 10106 14340
rect 10686 14328 10692 14340
rect 10100 14300 10692 14328
rect 10100 14288 10106 14300
rect 10686 14288 10692 14300
rect 10744 14288 10750 14340
rect 11514 14328 11520 14340
rect 10888 14300 11520 14328
rect 6656 14232 7512 14260
rect 8389 14263 8447 14269
rect 8389 14229 8401 14263
rect 8435 14229 8447 14263
rect 8389 14223 8447 14229
rect 9398 14220 9404 14272
rect 9456 14260 9462 14272
rect 10888 14260 10916 14300
rect 11514 14288 11520 14300
rect 11572 14328 11578 14340
rect 11762 14331 11820 14337
rect 11762 14328 11774 14331
rect 11572 14300 11774 14328
rect 11572 14288 11578 14300
rect 11762 14297 11774 14300
rect 11808 14297 11820 14331
rect 11762 14291 11820 14297
rect 9456 14232 10916 14260
rect 14384 14260 14412 14368
rect 15206 14365 15218 14368
rect 15252 14396 15264 14399
rect 15562 14396 15568 14408
rect 15252 14368 15568 14396
rect 15252 14365 15264 14368
rect 15206 14359 15264 14365
rect 15562 14356 15568 14368
rect 15620 14356 15626 14408
rect 16390 14356 16396 14408
rect 16448 14396 16454 14408
rect 16485 14399 16543 14405
rect 16485 14396 16497 14399
rect 16448 14368 16497 14396
rect 16448 14356 16454 14368
rect 16485 14365 16497 14368
rect 16531 14365 16543 14399
rect 18800 14396 18828 14436
rect 16485 14359 16543 14365
rect 18248 14368 18828 14396
rect 18877 14399 18935 14405
rect 16022 14288 16028 14340
rect 16080 14328 16086 14340
rect 18248 14328 18276 14368
rect 18877 14365 18889 14399
rect 18923 14396 18935 14399
rect 19058 14396 19064 14408
rect 18923 14368 19064 14396
rect 18923 14365 18935 14368
rect 18877 14359 18935 14365
rect 19058 14356 19064 14368
rect 19116 14356 19122 14408
rect 19628 14405 19656 14436
rect 19794 14424 19800 14436
rect 19852 14424 19858 14476
rect 19613 14399 19671 14405
rect 19613 14365 19625 14399
rect 19659 14365 19671 14399
rect 20622 14396 20628 14408
rect 20583 14368 20628 14396
rect 19613 14359 19671 14365
rect 20622 14356 20628 14368
rect 20680 14356 20686 14408
rect 20824 14396 20852 14495
rect 20901 14399 20959 14405
rect 20901 14396 20913 14399
rect 20824 14368 20913 14396
rect 20901 14365 20913 14368
rect 20947 14365 20959 14399
rect 20901 14359 20959 14365
rect 20990 14356 20996 14408
rect 21048 14396 21054 14408
rect 21269 14399 21327 14405
rect 21269 14396 21281 14399
rect 21048 14368 21281 14396
rect 21048 14356 21054 14368
rect 21269 14365 21281 14368
rect 21315 14365 21327 14399
rect 21269 14359 21327 14365
rect 16080 14300 18276 14328
rect 16080 14288 16086 14300
rect 16393 14263 16451 14269
rect 16393 14260 16405 14263
rect 14384 14232 16405 14260
rect 9456 14220 9462 14232
rect 16393 14229 16405 14232
rect 16439 14229 16451 14263
rect 16393 14223 16451 14229
rect 17589 14263 17647 14269
rect 17589 14229 17601 14263
rect 17635 14260 17647 14263
rect 17862 14260 17868 14272
rect 17635 14232 17868 14260
rect 17635 14229 17647 14232
rect 17589 14223 17647 14229
rect 17862 14220 17868 14232
rect 17920 14220 17926 14272
rect 18248 14260 18276 14300
rect 18506 14288 18512 14340
rect 18564 14328 18570 14340
rect 19705 14331 19763 14337
rect 19705 14328 19717 14331
rect 18564 14300 19717 14328
rect 18564 14288 18570 14300
rect 19705 14297 19717 14300
rect 19751 14297 19763 14331
rect 19705 14291 19763 14297
rect 18693 14263 18751 14269
rect 18693 14260 18705 14263
rect 18248 14232 18705 14260
rect 18693 14229 18705 14232
rect 18739 14229 18751 14263
rect 18693 14223 18751 14229
rect 19061 14263 19119 14269
rect 19061 14229 19073 14263
rect 19107 14260 19119 14263
rect 19518 14260 19524 14272
rect 19107 14232 19524 14260
rect 19107 14229 19119 14232
rect 19061 14223 19119 14229
rect 19518 14220 19524 14232
rect 19576 14220 19582 14272
rect 20070 14260 20076 14272
rect 20031 14232 20076 14260
rect 20070 14220 20076 14232
rect 20128 14220 20134 14272
rect 21082 14260 21088 14272
rect 21043 14232 21088 14260
rect 21082 14220 21088 14232
rect 21140 14220 21146 14272
rect 21450 14260 21456 14272
rect 21411 14232 21456 14260
rect 21450 14220 21456 14232
rect 21508 14220 21514 14272
rect 1104 14170 22056 14192
rect 1104 14118 6148 14170
rect 6200 14118 6212 14170
rect 6264 14118 6276 14170
rect 6328 14118 6340 14170
rect 6392 14118 6404 14170
rect 6456 14118 11346 14170
rect 11398 14118 11410 14170
rect 11462 14118 11474 14170
rect 11526 14118 11538 14170
rect 11590 14118 11602 14170
rect 11654 14118 16544 14170
rect 16596 14118 16608 14170
rect 16660 14118 16672 14170
rect 16724 14118 16736 14170
rect 16788 14118 16800 14170
rect 16852 14118 21742 14170
rect 21794 14118 21806 14170
rect 21858 14118 21870 14170
rect 21922 14118 21934 14170
rect 21986 14118 21998 14170
rect 22050 14118 22056 14170
rect 1104 14096 22056 14118
rect 1578 14016 1584 14068
rect 1636 14056 1642 14068
rect 1857 14059 1915 14065
rect 1857 14056 1869 14059
rect 1636 14028 1869 14056
rect 1636 14016 1642 14028
rect 1857 14025 1869 14028
rect 1903 14025 1915 14059
rect 4522 14056 4528 14068
rect 4483 14028 4528 14056
rect 1857 14019 1915 14025
rect 4522 14016 4528 14028
rect 4580 14016 4586 14068
rect 4890 14056 4896 14068
rect 4851 14028 4896 14056
rect 4890 14016 4896 14028
rect 4948 14016 4954 14068
rect 5350 14056 5356 14068
rect 5311 14028 5356 14056
rect 5350 14016 5356 14028
rect 5408 14016 5414 14068
rect 5905 14059 5963 14065
rect 5905 14025 5917 14059
rect 5951 14056 5963 14059
rect 6178 14056 6184 14068
rect 5951 14028 6184 14056
rect 5951 14025 5963 14028
rect 5905 14019 5963 14025
rect 6178 14016 6184 14028
rect 6236 14056 6242 14068
rect 6638 14056 6644 14068
rect 6236 14028 6644 14056
rect 6236 14016 6242 14028
rect 4065 13991 4123 13997
rect 4065 13957 4077 13991
rect 4111 13988 4123 13991
rect 4617 13991 4675 13997
rect 4617 13988 4629 13991
rect 4111 13960 4629 13988
rect 4111 13957 4123 13960
rect 4065 13951 4123 13957
rect 4617 13957 4629 13960
rect 4663 13988 4675 13991
rect 4982 13988 4988 14000
rect 4663 13960 4988 13988
rect 4663 13957 4675 13960
rect 4617 13951 4675 13957
rect 4982 13948 4988 13960
rect 5040 13948 5046 14000
rect 1670 13920 1676 13932
rect 1631 13892 1676 13920
rect 1670 13880 1676 13892
rect 1728 13880 1734 13932
rect 2041 13923 2099 13929
rect 2041 13889 2053 13923
rect 2087 13920 2099 13923
rect 2133 13923 2191 13929
rect 2133 13920 2145 13923
rect 2087 13892 2145 13920
rect 2087 13889 2099 13892
rect 2041 13883 2099 13889
rect 2133 13889 2145 13892
rect 2179 13889 2191 13923
rect 4154 13920 4160 13932
rect 4115 13892 4160 13920
rect 2133 13883 2191 13889
rect 1486 13716 1492 13728
rect 1447 13688 1492 13716
rect 1486 13676 1492 13688
rect 1544 13676 1550 13728
rect 2148 13716 2176 13883
rect 4154 13880 4160 13892
rect 4212 13880 4218 13932
rect 5261 13923 5319 13929
rect 5261 13889 5273 13923
rect 5307 13920 5319 13923
rect 6086 13920 6092 13932
rect 5307 13892 6092 13920
rect 5307 13889 5319 13892
rect 5261 13883 5319 13889
rect 6086 13880 6092 13892
rect 6144 13880 6150 13932
rect 6380 13929 6408 14028
rect 6638 14016 6644 14028
rect 6696 14056 6702 14068
rect 8297 14059 8355 14065
rect 8297 14056 8309 14059
rect 6696 14028 8309 14056
rect 6696 14016 6702 14028
rect 8297 14025 8309 14028
rect 8343 14025 8355 14059
rect 8297 14019 8355 14025
rect 9861 14059 9919 14065
rect 9861 14025 9873 14059
rect 9907 14056 9919 14059
rect 13173 14059 13231 14065
rect 9907 14028 13124 14056
rect 9907 14025 9919 14028
rect 9861 14019 9919 14025
rect 8312 13988 8340 14019
rect 10220 13991 10278 13997
rect 8312 13960 9996 13988
rect 6638 13929 6644 13932
rect 6365 13923 6423 13929
rect 6365 13889 6377 13923
rect 6411 13889 6423 13923
rect 6632 13920 6644 13929
rect 6599 13892 6644 13920
rect 6365 13883 6423 13889
rect 6632 13883 6644 13892
rect 6638 13880 6644 13883
rect 6696 13880 6702 13932
rect 8312 13920 8340 13960
rect 8478 13920 8484 13932
rect 8312 13892 8484 13920
rect 8478 13880 8484 13892
rect 8536 13880 8542 13932
rect 8570 13880 8576 13932
rect 8628 13920 8634 13932
rect 9968 13929 9996 13960
rect 10220 13957 10232 13991
rect 10266 13988 10278 13991
rect 11054 13988 11060 14000
rect 10266 13960 11060 13988
rect 10266 13957 10278 13960
rect 10220 13951 10278 13957
rect 11054 13948 11060 13960
rect 11112 13948 11118 14000
rect 13096 13988 13124 14028
rect 13173 14025 13185 14059
rect 13219 14056 13231 14059
rect 13354 14056 13360 14068
rect 13219 14028 13360 14056
rect 13219 14025 13231 14028
rect 13173 14019 13231 14025
rect 13354 14016 13360 14028
rect 13412 14016 13418 14068
rect 13722 14016 13728 14068
rect 13780 14056 13786 14068
rect 14001 14059 14059 14065
rect 14001 14056 14013 14059
rect 13780 14028 14013 14056
rect 13780 14016 13786 14028
rect 14001 14025 14013 14028
rect 14047 14025 14059 14059
rect 14001 14019 14059 14025
rect 13814 13988 13820 14000
rect 12406 13960 13032 13988
rect 13096 13960 13820 13988
rect 8748 13923 8806 13929
rect 8748 13920 8760 13923
rect 8628 13892 8760 13920
rect 8628 13880 8634 13892
rect 8748 13889 8760 13892
rect 8794 13920 8806 13923
rect 9953 13923 10011 13929
rect 8794 13892 9628 13920
rect 8794 13889 8806 13892
rect 8748 13883 8806 13889
rect 3973 13855 4031 13861
rect 3973 13821 3985 13855
rect 4019 13821 4031 13855
rect 5442 13852 5448 13864
rect 5403 13824 5448 13852
rect 3973 13815 4031 13821
rect 3988 13784 4016 13815
rect 5442 13812 5448 13824
rect 5500 13812 5506 13864
rect 9600 13852 9628 13892
rect 9953 13889 9965 13923
rect 9999 13889 10011 13923
rect 12406 13920 12434 13960
rect 9953 13883 10011 13889
rect 10060 13892 12434 13920
rect 12805 13923 12863 13929
rect 10060 13852 10088 13892
rect 12805 13889 12817 13923
rect 12851 13889 12863 13923
rect 13004 13920 13032 13960
rect 13814 13948 13820 13960
rect 13872 13948 13878 14000
rect 13906 13920 13912 13932
rect 13004 13892 13912 13920
rect 12805 13883 12863 13889
rect 9600 13824 10088 13852
rect 12529 13855 12587 13861
rect 12529 13821 12541 13855
rect 12575 13821 12587 13855
rect 12529 13815 12587 13821
rect 12713 13855 12771 13861
rect 12713 13821 12725 13855
rect 12759 13821 12771 13855
rect 12820 13852 12848 13883
rect 13906 13880 13912 13892
rect 13964 13880 13970 13932
rect 14016 13920 14044 14019
rect 14274 14016 14280 14068
rect 14332 14056 14338 14068
rect 15010 14056 15016 14068
rect 14332 14028 15016 14056
rect 14332 14016 14338 14028
rect 15010 14016 15016 14028
rect 15068 14016 15074 14068
rect 16390 14016 16396 14068
rect 16448 14056 16454 14068
rect 16669 14059 16727 14065
rect 16669 14056 16681 14059
rect 16448 14028 16681 14056
rect 16448 14016 16454 14028
rect 16669 14025 16681 14028
rect 16715 14025 16727 14059
rect 18230 14056 18236 14068
rect 18191 14028 18236 14056
rect 16669 14019 16727 14025
rect 18230 14016 18236 14028
rect 18288 14016 18294 14068
rect 18693 14059 18751 14065
rect 18693 14025 18705 14059
rect 18739 14056 18751 14059
rect 18874 14056 18880 14068
rect 18739 14028 18880 14056
rect 18739 14025 18751 14028
rect 18693 14019 18751 14025
rect 18874 14016 18880 14028
rect 18932 14016 18938 14068
rect 19058 14056 19064 14068
rect 19019 14028 19064 14056
rect 19058 14016 19064 14028
rect 19116 14016 19122 14068
rect 19153 14059 19211 14065
rect 19153 14025 19165 14059
rect 19199 14025 19211 14059
rect 19153 14019 19211 14025
rect 19521 14059 19579 14065
rect 19521 14025 19533 14059
rect 19567 14056 19579 14059
rect 20070 14056 20076 14068
rect 19567 14028 20076 14056
rect 19567 14025 19579 14028
rect 19521 14019 19579 14025
rect 16574 13988 16580 14000
rect 14292 13960 16580 13988
rect 14185 13923 14243 13929
rect 14185 13920 14197 13923
rect 14016 13892 14197 13920
rect 14185 13889 14197 13892
rect 14231 13889 14243 13923
rect 14185 13883 14243 13889
rect 14292 13852 14320 13960
rect 16574 13948 16580 13960
rect 16632 13948 16638 14000
rect 16868 13960 18920 13988
rect 14458 13929 14464 13932
rect 14452 13920 14464 13929
rect 14419 13892 14464 13920
rect 14452 13883 14464 13892
rect 14458 13880 14464 13883
rect 14516 13880 14522 13932
rect 15010 13880 15016 13932
rect 15068 13920 15074 13932
rect 16868 13920 16896 13960
rect 15068 13892 16896 13920
rect 15068 13880 15074 13892
rect 16942 13880 16948 13932
rect 17000 13920 17006 13932
rect 17037 13923 17095 13929
rect 17037 13920 17049 13923
rect 17000 13892 17049 13920
rect 17000 13880 17006 13892
rect 17037 13889 17049 13892
rect 17083 13889 17095 13923
rect 17144 13920 17172 13960
rect 17865 13923 17923 13929
rect 17144 13892 17264 13920
rect 17037 13883 17095 13889
rect 15838 13852 15844 13864
rect 12820 13824 14320 13852
rect 15799 13824 15844 13852
rect 12713 13815 12771 13821
rect 4706 13784 4712 13796
rect 3988 13756 4712 13784
rect 4706 13744 4712 13756
rect 4764 13744 4770 13796
rect 12544 13784 12572 13815
rect 10888 13756 12572 13784
rect 12728 13784 12756 13815
rect 15838 13812 15844 13824
rect 15896 13812 15902 13864
rect 17126 13852 17132 13864
rect 17087 13824 17132 13852
rect 17126 13812 17132 13824
rect 17184 13812 17190 13864
rect 17236 13861 17264 13892
rect 17865 13889 17877 13923
rect 17911 13920 17923 13923
rect 18230 13920 18236 13932
rect 17911 13892 18236 13920
rect 17911 13889 17923 13892
rect 17865 13883 17923 13889
rect 18230 13880 18236 13892
rect 18288 13880 18294 13932
rect 18892 13920 18920 13960
rect 18966 13948 18972 14000
rect 19024 13988 19030 14000
rect 19168 13988 19196 14019
rect 20070 14016 20076 14028
rect 20128 14016 20134 14068
rect 19024 13960 19196 13988
rect 19024 13948 19030 13960
rect 19794 13920 19800 13932
rect 18892 13892 19800 13920
rect 17221 13855 17279 13861
rect 17221 13821 17233 13855
rect 17267 13821 17279 13855
rect 17221 13815 17279 13821
rect 17589 13855 17647 13861
rect 17589 13821 17601 13855
rect 17635 13821 17647 13855
rect 17589 13815 17647 13821
rect 17773 13855 17831 13861
rect 17773 13821 17785 13855
rect 17819 13852 17831 13855
rect 18138 13852 18144 13864
rect 17819 13824 18144 13852
rect 17819 13821 17831 13824
rect 17773 13815 17831 13821
rect 13170 13784 13176 13796
rect 12728 13756 13176 13784
rect 7558 13716 7564 13728
rect 2148 13688 7564 13716
rect 7558 13676 7564 13688
rect 7616 13676 7622 13728
rect 7742 13716 7748 13728
rect 7655 13688 7748 13716
rect 7742 13676 7748 13688
rect 7800 13716 7806 13728
rect 7926 13716 7932 13728
rect 7800 13688 7932 13716
rect 7800 13676 7806 13688
rect 7926 13676 7932 13688
rect 7984 13676 7990 13728
rect 10318 13676 10324 13728
rect 10376 13716 10382 13728
rect 10888 13716 10916 13756
rect 13170 13744 13176 13756
rect 13228 13744 13234 13796
rect 15565 13787 15623 13793
rect 15565 13753 15577 13787
rect 15611 13784 15623 13787
rect 15746 13784 15752 13796
rect 15611 13756 15752 13784
rect 15611 13753 15623 13756
rect 15565 13747 15623 13753
rect 15746 13744 15752 13756
rect 15804 13784 15810 13796
rect 17604 13784 17632 13815
rect 18138 13812 18144 13824
rect 18196 13812 18202 13864
rect 18417 13855 18475 13861
rect 18417 13821 18429 13855
rect 18463 13821 18475 13855
rect 18598 13852 18604 13864
rect 18559 13824 18604 13852
rect 18417 13815 18475 13821
rect 15804 13756 17632 13784
rect 15804 13744 15810 13756
rect 17678 13744 17684 13796
rect 17736 13784 17742 13796
rect 18432 13784 18460 13815
rect 18598 13812 18604 13824
rect 18656 13812 18662 13864
rect 19720 13861 19748 13892
rect 19794 13880 19800 13892
rect 19852 13880 19858 13932
rect 21266 13920 21272 13932
rect 21227 13892 21272 13920
rect 21266 13880 21272 13892
rect 21324 13880 21330 13932
rect 19613 13855 19671 13861
rect 19613 13852 19625 13855
rect 19352 13824 19625 13852
rect 17736 13756 18460 13784
rect 17736 13744 17742 13756
rect 18966 13744 18972 13796
rect 19024 13784 19030 13796
rect 19352 13784 19380 13824
rect 19613 13821 19625 13824
rect 19659 13821 19671 13855
rect 19613 13815 19671 13821
rect 19705 13855 19763 13861
rect 19705 13821 19717 13855
rect 19751 13821 19763 13855
rect 19705 13815 19763 13821
rect 19024 13756 19380 13784
rect 19024 13744 19030 13756
rect 10376 13688 10916 13716
rect 11333 13719 11391 13725
rect 10376 13676 10382 13688
rect 11333 13685 11345 13719
rect 11379 13716 11391 13719
rect 11698 13716 11704 13728
rect 11379 13688 11704 13716
rect 11379 13685 11391 13688
rect 11333 13679 11391 13685
rect 11698 13676 11704 13688
rect 11756 13676 11762 13728
rect 12434 13676 12440 13728
rect 12492 13716 12498 13728
rect 15470 13716 15476 13728
rect 12492 13688 15476 13716
rect 12492 13676 12498 13688
rect 15470 13676 15476 13688
rect 15528 13676 15534 13728
rect 16022 13716 16028 13728
rect 15983 13688 16028 13716
rect 16022 13676 16028 13688
rect 16080 13676 16086 13728
rect 19628 13716 19656 13815
rect 21177 13787 21235 13793
rect 21177 13753 21189 13787
rect 21223 13784 21235 13787
rect 21542 13784 21548 13796
rect 21223 13756 21548 13784
rect 21223 13753 21235 13756
rect 21177 13747 21235 13753
rect 21542 13744 21548 13756
rect 21600 13744 21606 13796
rect 19702 13716 19708 13728
rect 19628 13688 19708 13716
rect 19702 13676 19708 13688
rect 19760 13676 19766 13728
rect 21450 13716 21456 13728
rect 21411 13688 21456 13716
rect 21450 13676 21456 13688
rect 21508 13676 21514 13728
rect 1104 13626 21896 13648
rect 1104 13574 3549 13626
rect 3601 13574 3613 13626
rect 3665 13574 3677 13626
rect 3729 13574 3741 13626
rect 3793 13574 3805 13626
rect 3857 13574 8747 13626
rect 8799 13574 8811 13626
rect 8863 13574 8875 13626
rect 8927 13574 8939 13626
rect 8991 13574 9003 13626
rect 9055 13574 13945 13626
rect 13997 13574 14009 13626
rect 14061 13574 14073 13626
rect 14125 13574 14137 13626
rect 14189 13574 14201 13626
rect 14253 13574 19143 13626
rect 19195 13574 19207 13626
rect 19259 13574 19271 13626
rect 19323 13574 19335 13626
rect 19387 13574 19399 13626
rect 19451 13574 21896 13626
rect 1104 13552 21896 13574
rect 1670 13472 1676 13524
rect 1728 13512 1734 13524
rect 1857 13515 1915 13521
rect 1857 13512 1869 13515
rect 1728 13484 1869 13512
rect 1728 13472 1734 13484
rect 1857 13481 1869 13484
rect 1903 13481 1915 13515
rect 1857 13475 1915 13481
rect 2774 13472 2780 13524
rect 2832 13512 2838 13524
rect 4065 13515 4123 13521
rect 4065 13512 4077 13515
rect 2832 13484 4077 13512
rect 2832 13472 2838 13484
rect 4065 13481 4077 13484
rect 4111 13481 4123 13515
rect 4065 13475 4123 13481
rect 5534 13472 5540 13524
rect 5592 13512 5598 13524
rect 6178 13512 6184 13524
rect 5592 13484 6184 13512
rect 5592 13472 5598 13484
rect 6178 13472 6184 13484
rect 6236 13472 6242 13524
rect 7837 13515 7895 13521
rect 7837 13512 7849 13515
rect 6564 13484 7849 13512
rect 1581 13447 1639 13453
rect 1581 13413 1593 13447
rect 1627 13444 1639 13447
rect 3050 13444 3056 13456
rect 1627 13416 3056 13444
rect 1627 13413 1639 13416
rect 1581 13407 1639 13413
rect 3050 13404 3056 13416
rect 3108 13404 3114 13456
rect 6086 13404 6092 13456
rect 6144 13444 6150 13456
rect 6564 13444 6592 13484
rect 7837 13481 7849 13484
rect 7883 13481 7895 13515
rect 7837 13475 7895 13481
rect 8478 13472 8484 13524
rect 8536 13512 8542 13524
rect 8665 13515 8723 13521
rect 8665 13512 8677 13515
rect 8536 13484 8677 13512
rect 8536 13472 8542 13484
rect 8665 13481 8677 13484
rect 8711 13512 8723 13515
rect 10413 13515 10471 13521
rect 10413 13512 10425 13515
rect 8711 13484 10425 13512
rect 8711 13481 8723 13484
rect 8665 13475 8723 13481
rect 8496 13444 8524 13472
rect 6144 13416 6592 13444
rect 7760 13416 8524 13444
rect 6144 13404 6150 13416
rect 7760 13388 7788 13416
rect 4709 13379 4767 13385
rect 4709 13345 4721 13379
rect 4755 13376 4767 13379
rect 5626 13376 5632 13388
rect 4755 13348 5632 13376
rect 4755 13345 4767 13348
rect 4709 13339 4767 13345
rect 5626 13336 5632 13348
rect 5684 13376 5690 13388
rect 5994 13376 6000 13388
rect 5684 13348 6000 13376
rect 5684 13336 5690 13348
rect 5994 13336 6000 13348
rect 6052 13336 6058 13388
rect 7742 13336 7748 13388
rect 7800 13376 7806 13388
rect 7800 13348 7893 13376
rect 7800 13336 7806 13348
rect 7926 13336 7932 13388
rect 7984 13376 7990 13388
rect 8956 13385 8984 13484
rect 10413 13481 10425 13484
rect 10459 13512 10471 13515
rect 11149 13515 11207 13521
rect 11149 13512 11161 13515
rect 10459 13484 11161 13512
rect 10459 13481 10471 13484
rect 10413 13475 10471 13481
rect 11149 13481 11161 13484
rect 11195 13481 11207 13515
rect 12805 13515 12863 13521
rect 11149 13475 11207 13481
rect 11348 13484 12756 13512
rect 10318 13444 10324 13456
rect 10279 13416 10324 13444
rect 10318 13404 10324 13416
rect 10376 13404 10382 13456
rect 8389 13379 8447 13385
rect 8389 13376 8401 13379
rect 7984 13348 8401 13376
rect 7984 13336 7990 13348
rect 8389 13345 8401 13348
rect 8435 13345 8447 13379
rect 8389 13339 8447 13345
rect 8941 13379 8999 13385
rect 8941 13345 8953 13379
rect 8987 13345 8999 13379
rect 8941 13339 8999 13345
rect 1394 13308 1400 13320
rect 1355 13280 1400 13308
rect 1394 13268 1400 13280
rect 1452 13308 1458 13320
rect 1673 13311 1731 13317
rect 1673 13308 1685 13311
rect 1452 13280 1685 13308
rect 1452 13268 1458 13280
rect 1673 13277 1685 13280
rect 1719 13277 1731 13311
rect 1673 13271 1731 13277
rect 2041 13311 2099 13317
rect 2041 13277 2053 13311
rect 2087 13308 2099 13311
rect 2314 13308 2320 13320
rect 2087 13280 2320 13308
rect 2087 13277 2099 13280
rect 2041 13271 2099 13277
rect 2314 13268 2320 13280
rect 2372 13268 2378 13320
rect 3970 13268 3976 13320
rect 4028 13308 4034 13320
rect 7489 13311 7547 13317
rect 7489 13308 7501 13311
rect 4028 13280 7236 13308
rect 4028 13268 4034 13280
rect 5350 13200 5356 13252
rect 5408 13240 5414 13252
rect 7098 13240 7104 13252
rect 5408 13212 7104 13240
rect 5408 13200 5414 13212
rect 7098 13200 7104 13212
rect 7156 13200 7162 13252
rect 2222 13172 2228 13184
rect 2183 13144 2228 13172
rect 2222 13132 2228 13144
rect 2280 13132 2286 13184
rect 4430 13172 4436 13184
rect 4391 13144 4436 13172
rect 4430 13132 4436 13144
rect 4488 13132 4494 13184
rect 4525 13175 4583 13181
rect 4525 13141 4537 13175
rect 4571 13172 4583 13175
rect 5442 13172 5448 13184
rect 4571 13144 5448 13172
rect 4571 13141 4583 13144
rect 4525 13135 4583 13141
rect 5442 13132 5448 13144
rect 5500 13132 5506 13184
rect 6365 13175 6423 13181
rect 6365 13141 6377 13175
rect 6411 13172 6423 13175
rect 6822 13172 6828 13184
rect 6411 13144 6828 13172
rect 6411 13141 6423 13144
rect 6365 13135 6423 13141
rect 6822 13132 6828 13144
rect 6880 13132 6886 13184
rect 7208 13172 7236 13280
rect 7300 13280 7501 13308
rect 7300 13252 7328 13280
rect 7489 13277 7501 13280
rect 7535 13308 7547 13311
rect 8110 13308 8116 13320
rect 7535 13280 8116 13308
rect 7535 13277 7547 13280
rect 7489 13271 7547 13277
rect 8110 13268 8116 13280
rect 8168 13268 8174 13320
rect 8202 13268 8208 13320
rect 8260 13308 8266 13320
rect 8297 13311 8355 13317
rect 8297 13308 8309 13311
rect 8260 13280 8309 13308
rect 8260 13268 8266 13280
rect 8297 13277 8309 13280
rect 8343 13277 8355 13311
rect 9766 13308 9772 13320
rect 8297 13271 8355 13277
rect 9140 13280 9772 13308
rect 7282 13200 7288 13252
rect 7340 13200 7346 13252
rect 9140 13240 9168 13280
rect 9766 13268 9772 13280
rect 9824 13268 9830 13320
rect 7484 13212 9168 13240
rect 9208 13243 9266 13249
rect 7484 13172 7512 13212
rect 9208 13209 9220 13243
rect 9254 13240 9266 13243
rect 11348 13240 11376 13484
rect 12728 13444 12756 13484
rect 12805 13481 12817 13515
rect 12851 13512 12863 13515
rect 13170 13512 13176 13524
rect 12851 13484 13176 13512
rect 12851 13481 12863 13484
rect 12805 13475 12863 13481
rect 13170 13472 13176 13484
rect 13228 13472 13234 13524
rect 18230 13512 18236 13524
rect 14200 13484 17264 13512
rect 18191 13484 18236 13512
rect 12728 13416 13492 13444
rect 13464 13385 13492 13416
rect 13449 13379 13507 13385
rect 13449 13345 13461 13379
rect 13495 13376 13507 13379
rect 14200 13376 14228 13484
rect 15841 13447 15899 13453
rect 15841 13444 15853 13447
rect 14568 13416 15853 13444
rect 14366 13376 14372 13388
rect 13495 13348 14228 13376
rect 14327 13348 14372 13376
rect 13495 13345 13507 13348
rect 13449 13339 13507 13345
rect 14366 13336 14372 13348
rect 14424 13336 14430 13388
rect 12710 13308 12716 13320
rect 12671 13280 12716 13308
rect 12710 13268 12716 13280
rect 12768 13268 12774 13320
rect 14568 13317 14596 13416
rect 15841 13413 15853 13416
rect 15887 13413 15899 13447
rect 15841 13407 15899 13413
rect 16574 13404 16580 13456
rect 16632 13444 16638 13456
rect 16669 13447 16727 13453
rect 16669 13444 16681 13447
rect 16632 13416 16681 13444
rect 16632 13404 16638 13416
rect 16669 13413 16681 13416
rect 16715 13413 16727 13447
rect 16669 13407 16727 13413
rect 15470 13376 15476 13388
rect 15431 13348 15476 13376
rect 15470 13336 15476 13348
rect 15528 13336 15534 13388
rect 15562 13336 15568 13388
rect 15620 13376 15626 13388
rect 17236 13385 17264 13484
rect 18230 13472 18236 13484
rect 18288 13472 18294 13524
rect 20990 13512 20996 13524
rect 20951 13484 20996 13512
rect 20990 13472 20996 13484
rect 21048 13472 21054 13524
rect 21269 13515 21327 13521
rect 21269 13481 21281 13515
rect 21315 13512 21327 13515
rect 21358 13512 21364 13524
rect 21315 13484 21364 13512
rect 21315 13481 21327 13484
rect 21269 13475 21327 13481
rect 21358 13472 21364 13484
rect 21416 13472 21422 13524
rect 16393 13379 16451 13385
rect 16393 13376 16405 13379
rect 15620 13348 16405 13376
rect 15620 13336 15626 13348
rect 16393 13345 16405 13348
rect 16439 13345 16451 13379
rect 16393 13339 16451 13345
rect 17221 13379 17279 13385
rect 17221 13345 17233 13379
rect 17267 13345 17279 13379
rect 17586 13376 17592 13388
rect 17547 13348 17592 13376
rect 17221 13339 17279 13345
rect 17586 13336 17592 13348
rect 17644 13336 17650 13388
rect 18966 13376 18972 13388
rect 18927 13348 18972 13376
rect 18966 13336 18972 13348
rect 19024 13336 19030 13388
rect 21358 13376 21364 13388
rect 19352 13348 21364 13376
rect 14553 13311 14611 13317
rect 14553 13277 14565 13311
rect 14599 13277 14611 13311
rect 14553 13271 14611 13277
rect 15838 13268 15844 13320
rect 15896 13308 15902 13320
rect 16209 13311 16267 13317
rect 16209 13308 16221 13311
rect 15896 13280 16221 13308
rect 15896 13268 15902 13280
rect 16209 13277 16221 13280
rect 16255 13277 16267 13311
rect 17862 13308 17868 13320
rect 17823 13280 17868 13308
rect 16209 13271 16267 13277
rect 17862 13268 17868 13280
rect 17920 13268 17926 13320
rect 18690 13268 18696 13320
rect 18748 13308 18754 13320
rect 19245 13311 19303 13317
rect 19245 13308 19257 13311
rect 18748 13280 19257 13308
rect 18748 13268 18754 13280
rect 19245 13277 19257 13280
rect 19291 13277 19303 13311
rect 19245 13271 19303 13277
rect 9254 13212 11376 13240
rect 9254 13209 9266 13212
rect 9208 13203 9266 13209
rect 7208 13144 7512 13172
rect 7558 13132 7564 13184
rect 7616 13172 7622 13184
rect 8205 13175 8263 13181
rect 8205 13172 8217 13175
rect 7616 13144 8217 13172
rect 7616 13132 7622 13144
rect 8205 13141 8217 13144
rect 8251 13172 8263 13175
rect 8294 13172 8300 13184
rect 8251 13144 8300 13172
rect 8251 13141 8263 13144
rect 8205 13135 8263 13141
rect 8294 13132 8300 13144
rect 8352 13172 8358 13184
rect 9674 13172 9680 13184
rect 8352 13144 9680 13172
rect 8352 13132 8358 13144
rect 9674 13132 9680 13144
rect 9732 13132 9738 13184
rect 9766 13132 9772 13184
rect 9824 13172 9830 13184
rect 11238 13172 11244 13184
rect 9824 13144 11244 13172
rect 9824 13132 9830 13144
rect 11238 13132 11244 13144
rect 11296 13132 11302 13184
rect 11348 13181 11376 13212
rect 11698 13200 11704 13252
rect 11756 13240 11762 13252
rect 12342 13240 12348 13252
rect 11756 13212 12348 13240
rect 11756 13200 11762 13212
rect 12342 13200 12348 13212
rect 12400 13240 12406 13252
rect 12446 13243 12504 13249
rect 12446 13240 12458 13243
rect 12400 13212 12458 13240
rect 12400 13200 12406 13212
rect 12446 13209 12458 13212
rect 12492 13209 12504 13243
rect 13265 13243 13323 13249
rect 13265 13240 13277 13243
rect 12446 13203 12504 13209
rect 12820 13212 13277 13240
rect 11333 13175 11391 13181
rect 11333 13141 11345 13175
rect 11379 13141 11391 13175
rect 11333 13135 11391 13141
rect 12250 13132 12256 13184
rect 12308 13172 12314 13184
rect 12820 13172 12848 13212
rect 13265 13209 13277 13212
rect 13311 13209 13323 13243
rect 13265 13203 13323 13209
rect 14461 13243 14519 13249
rect 14461 13209 14473 13243
rect 14507 13240 14519 13243
rect 15381 13243 15439 13249
rect 14507 13212 15056 13240
rect 14507 13209 14519 13212
rect 14461 13203 14519 13209
rect 13170 13172 13176 13184
rect 12308 13144 12848 13172
rect 13131 13144 13176 13172
rect 12308 13132 12314 13144
rect 13170 13132 13176 13144
rect 13228 13132 13234 13184
rect 14918 13172 14924 13184
rect 14879 13144 14924 13172
rect 14918 13132 14924 13144
rect 14976 13132 14982 13184
rect 15028 13181 15056 13212
rect 15381 13209 15393 13243
rect 15427 13240 15439 13243
rect 19352 13240 19380 13348
rect 21358 13336 21364 13348
rect 21416 13336 21422 13388
rect 20809 13311 20867 13317
rect 20809 13308 20821 13311
rect 15427 13212 19380 13240
rect 19444 13280 20821 13308
rect 15427 13209 15439 13212
rect 15381 13203 15439 13209
rect 15013 13175 15071 13181
rect 15013 13141 15025 13175
rect 15059 13141 15071 13175
rect 15013 13135 15071 13141
rect 15562 13132 15568 13184
rect 15620 13172 15626 13184
rect 16022 13172 16028 13184
rect 15620 13144 16028 13172
rect 15620 13132 15626 13144
rect 16022 13132 16028 13144
rect 16080 13172 16086 13184
rect 16301 13175 16359 13181
rect 16301 13172 16313 13175
rect 16080 13144 16313 13172
rect 16080 13132 16086 13144
rect 16301 13141 16313 13144
rect 16347 13141 16359 13175
rect 17034 13172 17040 13184
rect 16995 13144 17040 13172
rect 16301 13135 16359 13141
rect 17034 13132 17040 13144
rect 17092 13132 17098 13184
rect 17126 13132 17132 13184
rect 17184 13172 17190 13184
rect 17770 13172 17776 13184
rect 17184 13144 17229 13172
rect 17731 13144 17776 13172
rect 17184 13132 17190 13144
rect 17770 13132 17776 13144
rect 17828 13132 17834 13184
rect 19444 13181 19472 13280
rect 20809 13277 20821 13280
rect 20855 13277 20867 13311
rect 20809 13271 20867 13277
rect 21085 13311 21143 13317
rect 21085 13277 21097 13311
rect 21131 13277 21143 13311
rect 21542 13308 21548 13320
rect 21503 13280 21548 13308
rect 21085 13271 21143 13277
rect 21100 13240 21128 13271
rect 21542 13268 21548 13280
rect 21600 13268 21606 13320
rect 20824 13212 21128 13240
rect 20824 13184 20852 13212
rect 19429 13175 19487 13181
rect 19429 13141 19441 13175
rect 19475 13141 19487 13175
rect 19429 13135 19487 13141
rect 20717 13175 20775 13181
rect 20717 13141 20729 13175
rect 20763 13172 20775 13175
rect 20806 13172 20812 13184
rect 20763 13144 20812 13172
rect 20763 13141 20775 13144
rect 20717 13135 20775 13141
rect 20806 13132 20812 13144
rect 20864 13132 20870 13184
rect 21361 13175 21419 13181
rect 21361 13141 21373 13175
rect 21407 13172 21419 13175
rect 21634 13172 21640 13184
rect 21407 13144 21640 13172
rect 21407 13141 21419 13144
rect 21361 13135 21419 13141
rect 21634 13132 21640 13144
rect 21692 13132 21698 13184
rect 1104 13082 22056 13104
rect 1104 13030 6148 13082
rect 6200 13030 6212 13082
rect 6264 13030 6276 13082
rect 6328 13030 6340 13082
rect 6392 13030 6404 13082
rect 6456 13030 11346 13082
rect 11398 13030 11410 13082
rect 11462 13030 11474 13082
rect 11526 13030 11538 13082
rect 11590 13030 11602 13082
rect 11654 13030 16544 13082
rect 16596 13030 16608 13082
rect 16660 13030 16672 13082
rect 16724 13030 16736 13082
rect 16788 13030 16800 13082
rect 16852 13030 21742 13082
rect 21794 13030 21806 13082
rect 21858 13030 21870 13082
rect 21922 13030 21934 13082
rect 21986 13030 21998 13082
rect 22050 13030 22056 13082
rect 1104 13008 22056 13030
rect 2314 12968 2320 12980
rect 2275 12940 2320 12968
rect 2314 12928 2320 12940
rect 2372 12928 2378 12980
rect 3421 12971 3479 12977
rect 3421 12937 3433 12971
rect 3467 12968 3479 12971
rect 3973 12971 4031 12977
rect 3973 12968 3985 12971
rect 3467 12940 3985 12968
rect 3467 12937 3479 12940
rect 3421 12931 3479 12937
rect 3973 12937 3985 12940
rect 4019 12937 4031 12971
rect 3973 12931 4031 12937
rect 5353 12971 5411 12977
rect 5353 12937 5365 12971
rect 5399 12968 5411 12971
rect 5534 12968 5540 12980
rect 5399 12940 5540 12968
rect 5399 12937 5411 12940
rect 5353 12931 5411 12937
rect 5534 12928 5540 12940
rect 5592 12968 5598 12980
rect 5994 12968 6000 12980
rect 5592 12940 6000 12968
rect 5592 12928 5598 12940
rect 5994 12928 6000 12940
rect 6052 12928 6058 12980
rect 6822 12928 6828 12980
rect 6880 12968 6886 12980
rect 8294 12968 8300 12980
rect 6880 12940 7880 12968
rect 8255 12940 8300 12968
rect 6880 12928 6886 12940
rect 2961 12903 3019 12909
rect 2961 12869 2973 12903
rect 3007 12900 3019 12903
rect 5905 12903 5963 12909
rect 3007 12872 5764 12900
rect 3007 12869 3019 12872
rect 2961 12863 3019 12869
rect 2498 12832 2504 12844
rect 2459 12804 2504 12832
rect 2498 12792 2504 12804
rect 2556 12792 2562 12844
rect 3050 12832 3056 12844
rect 3011 12804 3056 12832
rect 3050 12792 3056 12804
rect 3108 12792 3114 12844
rect 3142 12792 3148 12844
rect 3200 12832 3206 12844
rect 3881 12835 3939 12841
rect 3881 12832 3893 12835
rect 3200 12804 3893 12832
rect 3200 12792 3206 12804
rect 3881 12801 3893 12804
rect 3927 12801 3939 12835
rect 5350 12832 5356 12844
rect 3881 12795 3939 12801
rect 4080 12804 5356 12832
rect 1949 12767 2007 12773
rect 1949 12733 1961 12767
rect 1995 12733 2007 12767
rect 2222 12764 2228 12776
rect 2183 12736 2228 12764
rect 1949 12727 2007 12733
rect 1964 12628 1992 12727
rect 2222 12724 2228 12736
rect 2280 12724 2286 12776
rect 2869 12767 2927 12773
rect 2869 12733 2881 12767
rect 2915 12764 2927 12767
rect 4080 12764 4108 12804
rect 5350 12792 5356 12804
rect 5408 12792 5414 12844
rect 2915 12736 4108 12764
rect 4157 12767 4215 12773
rect 2915 12733 2927 12736
rect 2869 12727 2927 12733
rect 4157 12733 4169 12767
rect 4203 12733 4215 12767
rect 4890 12764 4896 12776
rect 4851 12736 4896 12764
rect 4157 12727 4215 12733
rect 3418 12656 3424 12708
rect 3476 12696 3482 12708
rect 3513 12699 3571 12705
rect 3513 12696 3525 12699
rect 3476 12668 3525 12696
rect 3476 12656 3482 12668
rect 3513 12665 3525 12668
rect 3559 12665 3571 12699
rect 3513 12659 3571 12665
rect 3970 12628 3976 12640
rect 1964 12600 3976 12628
rect 3970 12588 3976 12600
rect 4028 12588 4034 12640
rect 4172 12628 4200 12727
rect 4890 12724 4896 12736
rect 4948 12724 4954 12776
rect 5442 12696 5448 12708
rect 5403 12668 5448 12696
rect 5442 12656 5448 12668
rect 5500 12656 5506 12708
rect 5736 12696 5764 12872
rect 5905 12869 5917 12903
rect 5951 12900 5963 12903
rect 7006 12900 7012 12912
rect 5951 12872 7012 12900
rect 5951 12869 5963 12872
rect 5905 12863 5963 12869
rect 7006 12860 7012 12872
rect 7064 12860 7070 12912
rect 7190 12860 7196 12912
rect 7248 12900 7254 12912
rect 7478 12903 7536 12909
rect 7478 12900 7490 12903
rect 7248 12872 7490 12900
rect 7248 12860 7254 12872
rect 7478 12869 7490 12872
rect 7524 12869 7536 12903
rect 7478 12863 7536 12869
rect 5813 12835 5871 12841
rect 5813 12801 5825 12835
rect 5859 12832 5871 12835
rect 6362 12832 6368 12844
rect 5859 12804 6368 12832
rect 5859 12801 5871 12804
rect 5813 12795 5871 12801
rect 6362 12792 6368 12804
rect 6420 12792 6426 12844
rect 7742 12832 7748 12844
rect 7703 12804 7748 12832
rect 7742 12792 7748 12804
rect 7800 12792 7806 12844
rect 7852 12832 7880 12940
rect 8294 12928 8300 12940
rect 8352 12928 8358 12980
rect 8662 12928 8668 12980
rect 8720 12968 8726 12980
rect 8849 12971 8907 12977
rect 8849 12968 8861 12971
rect 8720 12940 8861 12968
rect 8720 12928 8726 12940
rect 8849 12937 8861 12940
rect 8895 12937 8907 12971
rect 9490 12968 9496 12980
rect 9451 12940 9496 12968
rect 8849 12931 8907 12937
rect 9490 12928 9496 12940
rect 9548 12928 9554 12980
rect 9585 12971 9643 12977
rect 9585 12937 9597 12971
rect 9631 12968 9643 12971
rect 9674 12968 9680 12980
rect 9631 12940 9680 12968
rect 9631 12937 9643 12940
rect 9585 12931 9643 12937
rect 9674 12928 9680 12940
rect 9732 12928 9738 12980
rect 9766 12928 9772 12980
rect 9824 12928 9830 12980
rect 9953 12971 10011 12977
rect 9953 12937 9965 12971
rect 9999 12937 10011 12971
rect 9953 12931 10011 12937
rect 8754 12900 8760 12912
rect 8715 12872 8760 12900
rect 8754 12860 8760 12872
rect 8812 12860 8818 12912
rect 9508 12900 9536 12928
rect 9784 12900 9812 12928
rect 9508 12872 9812 12900
rect 9968 12900 9996 12931
rect 10134 12928 10140 12980
rect 10192 12968 10198 12980
rect 10321 12971 10379 12977
rect 10321 12968 10333 12971
rect 10192 12940 10333 12968
rect 10192 12928 10198 12940
rect 10321 12937 10333 12940
rect 10367 12937 10379 12971
rect 10321 12931 10379 12937
rect 11238 12928 11244 12980
rect 11296 12968 11302 12980
rect 11793 12971 11851 12977
rect 11793 12968 11805 12971
rect 11296 12940 11805 12968
rect 11296 12928 11302 12940
rect 11793 12937 11805 12940
rect 11839 12937 11851 12971
rect 11793 12931 11851 12937
rect 11882 12928 11888 12980
rect 11940 12968 11946 12980
rect 12250 12968 12256 12980
rect 11940 12940 11985 12968
rect 12211 12940 12256 12968
rect 11940 12928 11946 12940
rect 12250 12928 12256 12940
rect 12308 12928 12314 12980
rect 12618 12928 12624 12980
rect 12676 12968 12682 12980
rect 16945 12971 17003 12977
rect 16945 12968 16957 12971
rect 12676 12940 16957 12968
rect 12676 12928 12682 12940
rect 16945 12937 16957 12940
rect 16991 12937 17003 12971
rect 16945 12931 17003 12937
rect 17034 12928 17040 12980
rect 17092 12968 17098 12980
rect 17497 12971 17555 12977
rect 17497 12968 17509 12971
rect 17092 12940 17509 12968
rect 17092 12928 17098 12940
rect 17497 12937 17509 12940
rect 17543 12937 17555 12971
rect 17497 12931 17555 12937
rect 18598 12928 18604 12980
rect 18656 12968 18662 12980
rect 19061 12971 19119 12977
rect 19061 12968 19073 12971
rect 18656 12940 19073 12968
rect 18656 12928 18662 12940
rect 19061 12937 19073 12940
rect 19107 12937 19119 12971
rect 19061 12931 19119 12937
rect 19981 12971 20039 12977
rect 19981 12937 19993 12971
rect 20027 12968 20039 12971
rect 20714 12968 20720 12980
rect 20027 12940 20720 12968
rect 20027 12937 20039 12940
rect 19981 12931 20039 12937
rect 20714 12928 20720 12940
rect 20772 12928 20778 12980
rect 20990 12968 20996 12980
rect 20951 12940 20996 12968
rect 20990 12928 20996 12940
rect 21048 12928 21054 12980
rect 12434 12900 12440 12912
rect 9968 12872 12440 12900
rect 12434 12860 12440 12872
rect 12492 12860 12498 12912
rect 14553 12903 14611 12909
rect 14553 12900 14565 12903
rect 12820 12872 14565 12900
rect 7852 12804 8984 12832
rect 6086 12764 6092 12776
rect 6047 12736 6092 12764
rect 6086 12724 6092 12736
rect 6144 12724 6150 12776
rect 7834 12724 7840 12776
rect 7892 12764 7898 12776
rect 8956 12773 8984 12804
rect 9306 12792 9312 12844
rect 9364 12832 9370 12844
rect 10413 12835 10471 12841
rect 10413 12832 10425 12835
rect 9364 12804 10425 12832
rect 9364 12792 9370 12804
rect 10413 12801 10425 12804
rect 10459 12801 10471 12835
rect 12158 12832 12164 12844
rect 10413 12795 10471 12801
rect 10520 12804 12164 12832
rect 8021 12767 8079 12773
rect 8021 12764 8033 12767
rect 7892 12736 8033 12764
rect 7892 12724 7898 12736
rect 8021 12733 8033 12736
rect 8067 12764 8079 12767
rect 8941 12767 8999 12773
rect 8067 12736 8892 12764
rect 8067 12733 8079 12736
rect 8021 12727 8079 12733
rect 8389 12699 8447 12705
rect 8389 12696 8401 12699
rect 5736 12668 6500 12696
rect 6270 12628 6276 12640
rect 4172 12600 6276 12628
rect 6270 12588 6276 12600
rect 6328 12628 6334 12640
rect 6365 12631 6423 12637
rect 6365 12628 6377 12631
rect 6328 12600 6377 12628
rect 6328 12588 6334 12600
rect 6365 12597 6377 12600
rect 6411 12597 6423 12631
rect 6472 12628 6500 12668
rect 7760 12668 8401 12696
rect 7760 12628 7788 12668
rect 8389 12665 8401 12668
rect 8435 12665 8447 12699
rect 8864 12696 8892 12736
rect 8941 12733 8953 12767
rect 8987 12733 8999 12767
rect 9398 12764 9404 12776
rect 9359 12736 9404 12764
rect 8941 12727 8999 12733
rect 9398 12724 9404 12736
rect 9456 12724 9462 12776
rect 10134 12764 10140 12776
rect 10095 12736 10140 12764
rect 10134 12724 10140 12736
rect 10192 12724 10198 12776
rect 10520 12696 10548 12804
rect 12158 12792 12164 12804
rect 12216 12792 12222 12844
rect 12621 12835 12679 12841
rect 12621 12832 12633 12835
rect 12452 12804 12633 12832
rect 11698 12764 11704 12776
rect 11659 12736 11704 12764
rect 11698 12724 11704 12736
rect 11756 12724 11762 12776
rect 11882 12724 11888 12776
rect 11940 12764 11946 12776
rect 12452 12764 12480 12804
rect 12621 12801 12633 12804
rect 12667 12832 12679 12835
rect 12710 12832 12716 12844
rect 12667 12804 12716 12832
rect 12667 12801 12679 12804
rect 12621 12795 12679 12801
rect 12710 12792 12716 12804
rect 12768 12832 12774 12844
rect 12820 12832 12848 12872
rect 14553 12869 14565 12872
rect 14599 12900 14611 12903
rect 16206 12900 16212 12912
rect 14599 12872 16068 12900
rect 16167 12872 16212 12900
rect 14599 12869 14611 12872
rect 14553 12863 14611 12869
rect 12986 12841 12992 12844
rect 12768 12804 12848 12832
rect 12768 12792 12774 12804
rect 12980 12795 12992 12841
rect 13044 12832 13050 12844
rect 13354 12832 13360 12844
rect 13044 12804 13360 12832
rect 12986 12792 12992 12795
rect 13044 12792 13050 12804
rect 13354 12792 13360 12804
rect 13412 12792 13418 12844
rect 15746 12792 15752 12844
rect 15804 12841 15810 12844
rect 16040 12841 16068 12872
rect 16206 12860 16212 12872
rect 16264 12860 16270 12912
rect 16485 12903 16543 12909
rect 16485 12869 16497 12903
rect 16531 12900 16543 12903
rect 17865 12903 17923 12909
rect 17865 12900 17877 12903
rect 16531 12872 17877 12900
rect 16531 12869 16543 12872
rect 16485 12863 16543 12869
rect 17865 12869 17877 12872
rect 17911 12869 17923 12903
rect 17865 12863 17923 12869
rect 15804 12832 15816 12841
rect 16025 12835 16083 12841
rect 15804 12804 15849 12832
rect 15804 12795 15816 12804
rect 16025 12801 16037 12835
rect 16071 12801 16083 12835
rect 16224 12832 16252 12860
rect 17037 12835 17095 12841
rect 17037 12832 17049 12835
rect 16224 12804 17049 12832
rect 16025 12795 16083 12801
rect 17037 12801 17049 12804
rect 17083 12801 17095 12835
rect 17037 12795 17095 12801
rect 15804 12792 15810 12795
rect 17494 12792 17500 12844
rect 17552 12832 17558 12844
rect 18693 12835 18751 12841
rect 17552 12804 18092 12832
rect 17552 12792 17558 12804
rect 16758 12764 16764 12776
rect 11940 12736 12480 12764
rect 16719 12736 16764 12764
rect 11940 12724 11946 12736
rect 16758 12724 16764 12736
rect 16816 12724 16822 12776
rect 18064 12773 18092 12804
rect 18693 12801 18705 12835
rect 18739 12832 18751 12835
rect 18966 12832 18972 12844
rect 18739 12804 18972 12832
rect 18739 12801 18751 12804
rect 18693 12795 18751 12801
rect 18966 12792 18972 12804
rect 19024 12792 19030 12844
rect 19518 12792 19524 12844
rect 19576 12832 19582 12844
rect 19797 12835 19855 12841
rect 19797 12832 19809 12835
rect 19576 12804 19809 12832
rect 19576 12792 19582 12804
rect 19797 12801 19809 12804
rect 19843 12801 19855 12835
rect 19797 12795 19855 12801
rect 20809 12835 20867 12841
rect 20809 12801 20821 12835
rect 20855 12832 20867 12835
rect 21082 12832 21088 12844
rect 20855 12804 21088 12832
rect 20855 12801 20867 12804
rect 20809 12795 20867 12801
rect 21082 12792 21088 12804
rect 21140 12792 21146 12844
rect 21450 12832 21456 12844
rect 21411 12804 21456 12832
rect 21450 12792 21456 12804
rect 21508 12792 21514 12844
rect 17957 12767 18015 12773
rect 17957 12764 17969 12767
rect 17052 12736 17969 12764
rect 17052 12708 17080 12736
rect 17957 12733 17969 12736
rect 18003 12733 18015 12767
rect 17957 12727 18015 12733
rect 18049 12767 18107 12773
rect 18049 12733 18061 12767
rect 18095 12733 18107 12767
rect 18414 12764 18420 12776
rect 18375 12736 18420 12764
rect 18049 12727 18107 12733
rect 18414 12724 18420 12736
rect 18472 12724 18478 12776
rect 18601 12767 18659 12773
rect 18601 12733 18613 12767
rect 18647 12733 18659 12767
rect 20254 12764 20260 12776
rect 20215 12736 20260 12764
rect 18601 12727 18659 12733
rect 8864 12668 10548 12696
rect 10781 12699 10839 12705
rect 8389 12659 8447 12665
rect 10781 12665 10793 12699
rect 10827 12696 10839 12699
rect 12618 12696 12624 12708
rect 10827 12668 11836 12696
rect 10827 12665 10839 12668
rect 10781 12659 10839 12665
rect 6472 12600 7788 12628
rect 6365 12591 6423 12597
rect 8294 12588 8300 12640
rect 8352 12628 8358 12640
rect 9490 12628 9496 12640
rect 8352 12600 9496 12628
rect 8352 12588 8358 12600
rect 9490 12588 9496 12600
rect 9548 12588 9554 12640
rect 9674 12588 9680 12640
rect 9732 12628 9738 12640
rect 10873 12631 10931 12637
rect 10873 12628 10885 12631
rect 9732 12600 10885 12628
rect 9732 12588 9738 12600
rect 10873 12597 10885 12600
rect 10919 12628 10931 12631
rect 10962 12628 10968 12640
rect 10919 12600 10968 12628
rect 10919 12597 10931 12600
rect 10873 12591 10931 12597
rect 10962 12588 10968 12600
rect 11020 12588 11026 12640
rect 11808 12628 11836 12668
rect 11992 12668 12624 12696
rect 11992 12628 12020 12668
rect 12618 12656 12624 12668
rect 12676 12656 12682 12708
rect 14645 12699 14703 12705
rect 14645 12696 14657 12699
rect 13648 12668 14657 12696
rect 13648 12640 13676 12668
rect 14645 12665 14657 12668
rect 14691 12665 14703 12699
rect 14645 12659 14703 12665
rect 16040 12668 16252 12696
rect 11808 12600 12020 12628
rect 12158 12588 12164 12640
rect 12216 12628 12222 12640
rect 12894 12628 12900 12640
rect 12216 12600 12900 12628
rect 12216 12588 12222 12600
rect 12894 12588 12900 12600
rect 12952 12588 12958 12640
rect 13630 12588 13636 12640
rect 13688 12588 13694 12640
rect 14093 12631 14151 12637
rect 14093 12597 14105 12631
rect 14139 12628 14151 12631
rect 14458 12628 14464 12640
rect 14139 12600 14464 12628
rect 14139 12597 14151 12600
rect 14093 12591 14151 12597
rect 14458 12588 14464 12600
rect 14516 12628 14522 12640
rect 16040 12628 16068 12668
rect 14516 12600 16068 12628
rect 16224 12628 16252 12668
rect 17034 12656 17040 12708
rect 17092 12656 17098 12708
rect 17405 12699 17463 12705
rect 17405 12665 17417 12699
rect 17451 12696 17463 12699
rect 18616 12696 18644 12727
rect 20254 12724 20260 12736
rect 20312 12724 20318 12776
rect 17451 12668 18644 12696
rect 17451 12665 17463 12668
rect 17405 12659 17463 12665
rect 20714 12656 20720 12708
rect 20772 12696 20778 12708
rect 21269 12699 21327 12705
rect 21269 12696 21281 12699
rect 20772 12668 21281 12696
rect 20772 12656 20778 12668
rect 21269 12665 21281 12668
rect 21315 12665 21327 12699
rect 21269 12659 21327 12665
rect 17586 12628 17592 12640
rect 16224 12600 17592 12628
rect 14516 12588 14522 12600
rect 17586 12588 17592 12600
rect 17644 12588 17650 12640
rect 1104 12538 21896 12560
rect 1104 12486 3549 12538
rect 3601 12486 3613 12538
rect 3665 12486 3677 12538
rect 3729 12486 3741 12538
rect 3793 12486 3805 12538
rect 3857 12486 8747 12538
rect 8799 12486 8811 12538
rect 8863 12486 8875 12538
rect 8927 12486 8939 12538
rect 8991 12486 9003 12538
rect 9055 12486 13945 12538
rect 13997 12486 14009 12538
rect 14061 12486 14073 12538
rect 14125 12486 14137 12538
rect 14189 12486 14201 12538
rect 14253 12486 19143 12538
rect 19195 12486 19207 12538
rect 19259 12486 19271 12538
rect 19323 12486 19335 12538
rect 19387 12486 19399 12538
rect 19451 12486 21896 12538
rect 1104 12464 21896 12486
rect 2038 12384 2044 12436
rect 2096 12424 2102 12436
rect 2133 12427 2191 12433
rect 2133 12424 2145 12427
rect 2096 12396 2145 12424
rect 2096 12384 2102 12396
rect 2133 12393 2145 12396
rect 2179 12393 2191 12427
rect 2133 12387 2191 12393
rect 2777 12427 2835 12433
rect 2777 12393 2789 12427
rect 2823 12424 2835 12427
rect 3050 12424 3056 12436
rect 2823 12396 3056 12424
rect 2823 12393 2835 12396
rect 2777 12387 2835 12393
rect 3050 12384 3056 12396
rect 3108 12384 3114 12436
rect 3878 12424 3884 12436
rect 3252 12396 3884 12424
rect 1670 12356 1676 12368
rect 1631 12328 1676 12356
rect 1670 12316 1676 12328
rect 1728 12316 1734 12368
rect 3252 12297 3280 12396
rect 3878 12384 3884 12396
rect 3936 12384 3942 12436
rect 4430 12424 4436 12436
rect 4391 12396 4436 12424
rect 4430 12384 4436 12396
rect 4488 12384 4494 12436
rect 6362 12384 6368 12436
rect 6420 12424 6426 12436
rect 7101 12427 7159 12433
rect 7101 12424 7113 12427
rect 6420 12396 7113 12424
rect 6420 12384 6426 12396
rect 7101 12393 7113 12396
rect 7147 12393 7159 12427
rect 9490 12424 9496 12436
rect 7101 12387 7159 12393
rect 7208 12396 9496 12424
rect 5718 12316 5724 12368
rect 5776 12356 5782 12368
rect 7208 12356 7236 12396
rect 9490 12384 9496 12396
rect 9548 12384 9554 12436
rect 9766 12424 9772 12436
rect 9727 12396 9772 12424
rect 9766 12384 9772 12396
rect 9824 12384 9830 12436
rect 10060 12396 10272 12424
rect 8018 12356 8024 12368
rect 5776 12328 7236 12356
rect 7668 12328 8024 12356
rect 5776 12316 5782 12328
rect 2593 12291 2651 12297
rect 2593 12288 2605 12291
rect 1504 12260 2605 12288
rect 1504 12232 1532 12260
rect 2593 12257 2605 12260
rect 2639 12257 2651 12291
rect 2593 12251 2651 12257
rect 3237 12291 3295 12297
rect 3237 12257 3249 12291
rect 3283 12257 3295 12291
rect 3237 12251 3295 12257
rect 3421 12291 3479 12297
rect 3421 12257 3433 12291
rect 3467 12288 3479 12291
rect 5077 12291 5135 12297
rect 3467 12260 5028 12288
rect 3467 12257 3479 12260
rect 3421 12251 3479 12257
rect 1486 12220 1492 12232
rect 1447 12192 1492 12220
rect 1486 12180 1492 12192
rect 1544 12180 1550 12232
rect 1946 12180 1952 12232
rect 2004 12220 2010 12232
rect 2317 12223 2375 12229
rect 2317 12220 2329 12223
rect 2004 12192 2329 12220
rect 2004 12180 2010 12192
rect 2317 12189 2329 12192
rect 2363 12189 2375 12223
rect 2317 12183 2375 12189
rect 2958 12180 2964 12232
rect 3016 12220 3022 12232
rect 3145 12223 3203 12229
rect 3145 12220 3157 12223
rect 3016 12192 3157 12220
rect 3016 12180 3022 12192
rect 3145 12189 3157 12192
rect 3191 12220 3203 12223
rect 3973 12223 4031 12229
rect 3973 12220 3985 12223
rect 3191 12192 3985 12220
rect 3191 12189 3203 12192
rect 3145 12183 3203 12189
rect 3973 12189 3985 12192
rect 4019 12189 4031 12223
rect 3973 12183 4031 12189
rect 4801 12223 4859 12229
rect 4801 12189 4813 12223
rect 4847 12220 4859 12223
rect 4890 12220 4896 12232
rect 4847 12192 4896 12220
rect 4847 12189 4859 12192
rect 4801 12183 4859 12189
rect 4890 12180 4896 12192
rect 4948 12180 4954 12232
rect 5000 12220 5028 12260
rect 5077 12257 5089 12291
rect 5123 12288 5135 12291
rect 6086 12288 6092 12300
rect 5123 12260 6092 12288
rect 5123 12257 5135 12260
rect 5077 12251 5135 12257
rect 6086 12248 6092 12260
rect 6144 12288 6150 12300
rect 6730 12288 6736 12300
rect 6144 12260 6736 12288
rect 6144 12248 6150 12260
rect 6730 12248 6736 12260
rect 6788 12248 6794 12300
rect 7098 12248 7104 12300
rect 7156 12288 7162 12300
rect 7668 12297 7696 12328
rect 8018 12316 8024 12328
rect 8076 12316 8082 12368
rect 8757 12359 8815 12365
rect 8757 12325 8769 12359
rect 8803 12356 8815 12359
rect 10060 12356 10088 12396
rect 8803 12328 9352 12356
rect 8803 12325 8815 12328
rect 8757 12319 8815 12325
rect 7653 12291 7711 12297
rect 7653 12288 7665 12291
rect 7156 12260 7665 12288
rect 7156 12248 7162 12260
rect 7653 12257 7665 12260
rect 7699 12257 7711 12291
rect 8110 12288 8116 12300
rect 8071 12260 8116 12288
rect 7653 12251 7711 12257
rect 8110 12248 8116 12260
rect 8168 12248 8174 12300
rect 8294 12288 8300 12300
rect 8255 12260 8300 12288
rect 8294 12248 8300 12260
rect 8352 12248 8358 12300
rect 9214 12288 9220 12300
rect 9175 12260 9220 12288
rect 9214 12248 9220 12260
rect 9272 12248 9278 12300
rect 9324 12297 9352 12328
rect 9646 12328 10088 12356
rect 10244 12356 10272 12396
rect 10318 12384 10324 12436
rect 10376 12424 10382 12436
rect 12986 12424 12992 12436
rect 10376 12396 12992 12424
rect 10376 12384 10382 12396
rect 12986 12384 12992 12396
rect 13044 12384 13050 12436
rect 13170 12424 13176 12436
rect 13131 12396 13176 12424
rect 13170 12384 13176 12396
rect 13228 12384 13234 12436
rect 16758 12424 16764 12436
rect 14108 12396 16764 12424
rect 10244 12328 12756 12356
rect 9309 12291 9367 12297
rect 9309 12257 9321 12291
rect 9355 12257 9367 12291
rect 9646 12288 9674 12328
rect 9309 12251 9367 12257
rect 9416 12260 9674 12288
rect 10045 12291 10103 12297
rect 6181 12223 6239 12229
rect 5000 12192 6132 12220
rect 1854 12152 1860 12164
rect 1815 12124 1860 12152
rect 1854 12112 1860 12124
rect 1912 12152 1918 12164
rect 2409 12155 2467 12161
rect 2409 12152 2421 12155
rect 1912 12124 2421 12152
rect 1912 12112 1918 12124
rect 2409 12121 2421 12124
rect 2455 12121 2467 12155
rect 2409 12115 2467 12121
rect 1949 12087 2007 12093
rect 1949 12053 1961 12087
rect 1995 12084 2007 12087
rect 2682 12084 2688 12096
rect 1995 12056 2688 12084
rect 1995 12053 2007 12056
rect 1949 12047 2007 12053
rect 2682 12044 2688 12056
rect 2740 12044 2746 12096
rect 4890 12084 4896 12096
rect 4851 12056 4896 12084
rect 4890 12044 4896 12056
rect 4948 12044 4954 12096
rect 5074 12044 5080 12096
rect 5132 12084 5138 12096
rect 5350 12084 5356 12096
rect 5132 12056 5356 12084
rect 5132 12044 5138 12056
rect 5350 12044 5356 12056
rect 5408 12044 5414 12096
rect 5994 12084 6000 12096
rect 5955 12056 6000 12084
rect 5994 12044 6000 12056
rect 6052 12044 6058 12096
rect 6104 12084 6132 12192
rect 6181 12189 6193 12223
rect 6227 12189 6239 12223
rect 6181 12183 6239 12189
rect 6457 12223 6515 12229
rect 6457 12189 6469 12223
rect 6503 12220 6515 12223
rect 6638 12220 6644 12232
rect 6503 12192 6644 12220
rect 6503 12189 6515 12192
rect 6457 12183 6515 12189
rect 6196 12152 6224 12183
rect 6638 12180 6644 12192
rect 6696 12180 6702 12232
rect 7469 12223 7527 12229
rect 7469 12189 7481 12223
rect 7515 12220 7527 12223
rect 7834 12220 7840 12232
rect 7515 12192 7840 12220
rect 7515 12189 7527 12192
rect 7469 12183 7527 12189
rect 7834 12180 7840 12192
rect 7892 12180 7898 12232
rect 8386 12220 8392 12232
rect 8347 12192 8392 12220
rect 8386 12180 8392 12192
rect 8444 12180 8450 12232
rect 7374 12152 7380 12164
rect 6196 12124 7380 12152
rect 7374 12112 7380 12124
rect 7432 12112 7438 12164
rect 7650 12112 7656 12164
rect 7708 12152 7714 12164
rect 7708 12124 8791 12152
rect 7708 12112 7714 12124
rect 6730 12084 6736 12096
rect 6104 12056 6736 12084
rect 6730 12044 6736 12056
rect 6788 12044 6794 12096
rect 7561 12087 7619 12093
rect 7561 12053 7573 12087
rect 7607 12084 7619 12087
rect 8662 12084 8668 12096
rect 7607 12056 8668 12084
rect 7607 12053 7619 12056
rect 7561 12047 7619 12053
rect 8662 12044 8668 12056
rect 8720 12044 8726 12096
rect 8763 12084 8791 12124
rect 9306 12112 9312 12164
rect 9364 12152 9370 12164
rect 9416 12161 9444 12260
rect 10045 12257 10057 12291
rect 10091 12288 10103 12291
rect 10318 12288 10324 12300
rect 10091 12260 10324 12288
rect 10091 12257 10103 12260
rect 10045 12251 10103 12257
rect 10318 12248 10324 12260
rect 10376 12248 10382 12300
rect 10502 12248 10508 12300
rect 10560 12288 10566 12300
rect 11241 12291 11299 12297
rect 11241 12288 11253 12291
rect 10560 12260 11253 12288
rect 10560 12248 10566 12260
rect 11241 12257 11253 12260
rect 11287 12257 11299 12291
rect 11241 12251 11299 12257
rect 12342 12248 12348 12300
rect 12400 12288 12406 12300
rect 12728 12297 12756 12328
rect 12802 12316 12808 12368
rect 12860 12356 12866 12368
rect 14108 12356 14136 12396
rect 16758 12384 16764 12396
rect 16816 12424 16822 12436
rect 18601 12427 18659 12433
rect 16816 12396 18552 12424
rect 16816 12384 16822 12396
rect 12860 12328 14136 12356
rect 12860 12316 12866 12328
rect 15378 12316 15384 12368
rect 15436 12356 15442 12368
rect 15473 12359 15531 12365
rect 15473 12356 15485 12359
rect 15436 12328 15485 12356
rect 15436 12316 15442 12328
rect 15473 12325 15485 12328
rect 15519 12356 15531 12359
rect 18524 12356 18552 12396
rect 18601 12393 18613 12427
rect 18647 12424 18659 12427
rect 18690 12424 18696 12436
rect 18647 12396 18696 12424
rect 18647 12393 18659 12396
rect 18601 12387 18659 12393
rect 18690 12384 18696 12396
rect 18748 12384 18754 12436
rect 18874 12384 18880 12436
rect 18932 12424 18938 12436
rect 19245 12427 19303 12433
rect 19245 12424 19257 12427
rect 18932 12396 19257 12424
rect 18932 12384 18938 12396
rect 19245 12393 19257 12396
rect 19291 12393 19303 12427
rect 19245 12387 19303 12393
rect 21361 12427 21419 12433
rect 21361 12393 21373 12427
rect 21407 12424 21419 12427
rect 22094 12424 22100 12436
rect 21407 12396 22100 12424
rect 21407 12393 21419 12396
rect 21361 12387 21419 12393
rect 22094 12384 22100 12396
rect 22152 12384 22158 12436
rect 19610 12356 19616 12368
rect 15519 12328 18000 12356
rect 18524 12328 19616 12356
rect 15519 12325 15531 12328
rect 15473 12319 15531 12325
rect 12621 12291 12679 12297
rect 12621 12288 12633 12291
rect 12400 12260 12633 12288
rect 12400 12248 12406 12260
rect 12621 12257 12633 12260
rect 12667 12257 12679 12291
rect 12621 12251 12679 12257
rect 12713 12291 12771 12297
rect 12713 12257 12725 12291
rect 12759 12257 12771 12291
rect 16853 12291 16911 12297
rect 12713 12251 12771 12257
rect 12820 12260 14228 12288
rect 9490 12180 9496 12232
rect 9548 12220 9554 12232
rect 9950 12220 9956 12232
rect 9548 12192 9956 12220
rect 9548 12180 9554 12192
rect 9950 12180 9956 12192
rect 10008 12220 10014 12232
rect 10229 12223 10287 12229
rect 10229 12220 10241 12223
rect 10008 12192 10241 12220
rect 10008 12180 10014 12192
rect 10229 12189 10241 12192
rect 10275 12189 10287 12223
rect 10229 12183 10287 12189
rect 10778 12180 10784 12232
rect 10836 12220 10842 12232
rect 11517 12223 11575 12229
rect 11517 12220 11529 12223
rect 10836 12192 11529 12220
rect 10836 12180 10842 12192
rect 11517 12189 11529 12192
rect 11563 12189 11575 12223
rect 12636 12220 12664 12251
rect 12820 12220 12848 12260
rect 14093 12223 14151 12229
rect 14093 12220 14105 12223
rect 12636 12192 12848 12220
rect 13924 12192 14105 12220
rect 11517 12183 11575 12189
rect 9401 12155 9459 12161
rect 9401 12152 9413 12155
rect 9364 12124 9413 12152
rect 9364 12112 9370 12124
rect 9401 12121 9413 12124
rect 9447 12121 9459 12155
rect 9401 12115 9459 12121
rect 9766 12112 9772 12164
rect 9824 12152 9830 12164
rect 11149 12155 11207 12161
rect 11149 12152 11161 12155
rect 9824 12124 11161 12152
rect 9824 12112 9830 12124
rect 11149 12121 11161 12124
rect 11195 12121 11207 12155
rect 11149 12115 11207 12121
rect 11698 12112 11704 12164
rect 11756 12152 11762 12164
rect 12526 12152 12532 12164
rect 11756 12124 12532 12152
rect 11756 12112 11762 12124
rect 12526 12112 12532 12124
rect 12584 12112 12590 12164
rect 12805 12155 12863 12161
rect 12805 12152 12817 12155
rect 12636 12124 12817 12152
rect 10137 12087 10195 12093
rect 10137 12084 10149 12087
rect 8763 12056 10149 12084
rect 10137 12053 10149 12056
rect 10183 12053 10195 12087
rect 10594 12084 10600 12096
rect 10555 12056 10600 12084
rect 10137 12047 10195 12053
rect 10594 12044 10600 12056
rect 10652 12044 10658 12096
rect 10689 12087 10747 12093
rect 10689 12053 10701 12087
rect 10735 12084 10747 12087
rect 10870 12084 10876 12096
rect 10735 12056 10876 12084
rect 10735 12053 10747 12056
rect 10689 12047 10747 12053
rect 10870 12044 10876 12056
rect 10928 12044 10934 12096
rect 11054 12084 11060 12096
rect 11015 12056 11060 12084
rect 11054 12044 11060 12056
rect 11112 12044 11118 12096
rect 12158 12084 12164 12096
rect 12119 12056 12164 12084
rect 12158 12044 12164 12056
rect 12216 12044 12222 12096
rect 12250 12044 12256 12096
rect 12308 12084 12314 12096
rect 12636 12084 12664 12124
rect 12805 12121 12817 12124
rect 12851 12121 12863 12155
rect 12805 12115 12863 12121
rect 13924 12093 13952 12192
rect 14093 12189 14105 12192
rect 14139 12189 14151 12223
rect 14200 12220 14228 12260
rect 16853 12257 16865 12291
rect 16899 12288 16911 12291
rect 17034 12288 17040 12300
rect 16899 12260 17040 12288
rect 16899 12257 16911 12260
rect 16853 12251 16911 12257
rect 17034 12248 17040 12260
rect 17092 12248 17098 12300
rect 17494 12288 17500 12300
rect 17455 12260 17500 12288
rect 17494 12248 17500 12260
rect 17552 12248 17558 12300
rect 17972 12297 18000 12328
rect 19610 12316 19616 12328
rect 19668 12356 19674 12368
rect 21177 12359 21235 12365
rect 19668 12328 20668 12356
rect 19668 12316 19674 12328
rect 17957 12291 18015 12297
rect 17957 12257 17969 12291
rect 18003 12257 18015 12291
rect 17957 12251 18015 12257
rect 18414 12248 18420 12300
rect 18472 12288 18478 12300
rect 20640 12297 20668 12328
rect 21177 12325 21189 12359
rect 21223 12356 21235 12359
rect 21450 12356 21456 12368
rect 21223 12328 21456 12356
rect 21223 12325 21235 12328
rect 21177 12319 21235 12325
rect 21450 12316 21456 12328
rect 21508 12316 21514 12368
rect 19797 12291 19855 12297
rect 19797 12288 19809 12291
rect 18472 12260 19809 12288
rect 18472 12248 18478 12260
rect 19797 12257 19809 12260
rect 19843 12257 19855 12291
rect 19797 12251 19855 12257
rect 20625 12291 20683 12297
rect 20625 12257 20637 12291
rect 20671 12257 20683 12291
rect 20625 12251 20683 12257
rect 17512 12220 17540 12248
rect 14200 12192 17540 12220
rect 14093 12183 14151 12189
rect 17862 12180 17868 12232
rect 17920 12220 17926 12232
rect 18693 12223 18751 12229
rect 18693 12220 18705 12223
rect 17920 12192 18705 12220
rect 17920 12180 17926 12192
rect 18693 12189 18705 12192
rect 18739 12189 18751 12223
rect 18693 12183 18751 12189
rect 20254 12180 20260 12232
rect 20312 12220 20318 12232
rect 20441 12223 20499 12229
rect 20441 12220 20453 12223
rect 20312 12192 20453 12220
rect 20312 12180 20318 12192
rect 20441 12189 20453 12192
rect 20487 12189 20499 12223
rect 20441 12183 20499 12189
rect 13998 12112 14004 12164
rect 14056 12152 14062 12164
rect 14360 12155 14418 12161
rect 14360 12152 14372 12155
rect 14056 12124 14372 12152
rect 14056 12112 14062 12124
rect 14360 12121 14372 12124
rect 14406 12152 14418 12155
rect 18874 12152 18880 12164
rect 14406 12124 18880 12152
rect 14406 12121 14418 12124
rect 14360 12115 14418 12121
rect 18874 12112 18880 12124
rect 18932 12112 18938 12164
rect 19613 12155 19671 12161
rect 19613 12121 19625 12155
rect 19659 12152 19671 12155
rect 20530 12152 20536 12164
rect 19659 12124 20116 12152
rect 20491 12124 20536 12152
rect 19659 12121 19671 12124
rect 19613 12115 19671 12121
rect 12308 12056 12664 12084
rect 13909 12087 13967 12093
rect 12308 12044 12314 12056
rect 13909 12053 13921 12087
rect 13955 12084 13967 12087
rect 14182 12084 14188 12096
rect 13955 12056 14188 12084
rect 13955 12053 13967 12056
rect 13909 12047 13967 12053
rect 14182 12044 14188 12056
rect 14240 12044 14246 12096
rect 16945 12087 17003 12093
rect 16945 12053 16957 12087
rect 16991 12084 17003 12087
rect 17126 12084 17132 12096
rect 16991 12056 17132 12084
rect 16991 12053 17003 12056
rect 16945 12047 17003 12053
rect 17126 12044 17132 12056
rect 17184 12044 17190 12096
rect 17218 12044 17224 12096
rect 17276 12084 17282 12096
rect 17313 12087 17371 12093
rect 17313 12084 17325 12087
rect 17276 12056 17325 12084
rect 17276 12044 17282 12056
rect 17313 12053 17325 12056
rect 17359 12053 17371 12087
rect 17313 12047 17371 12053
rect 17405 12087 17463 12093
rect 17405 12053 17417 12087
rect 17451 12084 17463 12087
rect 17862 12084 17868 12096
rect 17451 12056 17868 12084
rect 17451 12053 17463 12056
rect 17405 12047 17463 12053
rect 17862 12044 17868 12056
rect 17920 12044 17926 12096
rect 18138 12084 18144 12096
rect 18099 12056 18144 12084
rect 18138 12044 18144 12056
rect 18196 12044 18202 12096
rect 18233 12087 18291 12093
rect 18233 12053 18245 12087
rect 18279 12084 18291 12087
rect 18322 12084 18328 12096
rect 18279 12056 18328 12084
rect 18279 12053 18291 12056
rect 18233 12047 18291 12053
rect 18322 12044 18328 12056
rect 18380 12044 18386 12096
rect 19702 12084 19708 12096
rect 19663 12056 19708 12084
rect 19702 12044 19708 12056
rect 19760 12044 19766 12096
rect 20088 12093 20116 12124
rect 20530 12112 20536 12124
rect 20588 12112 20594 12164
rect 20993 12155 21051 12161
rect 20993 12121 21005 12155
rect 21039 12152 21051 12155
rect 21450 12152 21456 12164
rect 21039 12124 21456 12152
rect 21039 12121 21051 12124
rect 20993 12115 21051 12121
rect 21450 12112 21456 12124
rect 21508 12112 21514 12164
rect 20073 12087 20131 12093
rect 20073 12053 20085 12087
rect 20119 12053 20131 12087
rect 20073 12047 20131 12053
rect 1104 11994 22056 12016
rect 1104 11942 6148 11994
rect 6200 11942 6212 11994
rect 6264 11942 6276 11994
rect 6328 11942 6340 11994
rect 6392 11942 6404 11994
rect 6456 11942 11346 11994
rect 11398 11942 11410 11994
rect 11462 11942 11474 11994
rect 11526 11942 11538 11994
rect 11590 11942 11602 11994
rect 11654 11942 16544 11994
rect 16596 11942 16608 11994
rect 16660 11942 16672 11994
rect 16724 11942 16736 11994
rect 16788 11942 16800 11994
rect 16852 11942 21742 11994
rect 21794 11942 21806 11994
rect 21858 11942 21870 11994
rect 21922 11942 21934 11994
rect 21986 11942 21998 11994
rect 22050 11942 22056 11994
rect 1104 11920 22056 11942
rect 1762 11840 1768 11892
rect 1820 11880 1826 11892
rect 1857 11883 1915 11889
rect 1857 11880 1869 11883
rect 1820 11852 1869 11880
rect 1820 11840 1826 11852
rect 1857 11849 1869 11852
rect 1903 11849 1915 11883
rect 1857 11843 1915 11849
rect 2317 11883 2375 11889
rect 2317 11849 2329 11883
rect 2363 11880 2375 11883
rect 4246 11880 4252 11892
rect 2363 11852 4252 11880
rect 2363 11849 2375 11852
rect 2317 11843 2375 11849
rect 4246 11840 4252 11852
rect 4304 11840 4310 11892
rect 5718 11880 5724 11892
rect 5679 11852 5724 11880
rect 5718 11840 5724 11852
rect 5776 11840 5782 11892
rect 6638 11880 6644 11892
rect 6104 11852 6644 11880
rect 2593 11815 2651 11821
rect 2593 11812 2605 11815
rect 1504 11784 2605 11812
rect 1394 11704 1400 11756
rect 1452 11744 1458 11756
rect 1504 11753 1532 11784
rect 2593 11781 2605 11784
rect 2639 11781 2651 11815
rect 2593 11775 2651 11781
rect 4798 11772 4804 11824
rect 4856 11812 4862 11824
rect 6104 11812 6132 11852
rect 6638 11840 6644 11852
rect 6696 11840 6702 11892
rect 7742 11840 7748 11892
rect 7800 11880 7806 11892
rect 8941 11883 8999 11889
rect 8941 11880 8953 11883
rect 7800 11852 8953 11880
rect 7800 11840 7806 11852
rect 8941 11849 8953 11852
rect 8987 11880 8999 11883
rect 10870 11880 10876 11892
rect 8987 11852 9168 11880
rect 10831 11852 10876 11880
rect 8987 11849 8999 11852
rect 8941 11843 8999 11849
rect 4856 11784 6132 11812
rect 6564 11784 7604 11812
rect 4856 11772 4862 11784
rect 1489 11747 1547 11753
rect 1489 11744 1501 11747
rect 1452 11716 1501 11744
rect 1452 11704 1458 11716
rect 1489 11713 1501 11716
rect 1535 11713 1547 11747
rect 1489 11707 1547 11713
rect 2041 11747 2099 11753
rect 2041 11713 2053 11747
rect 2087 11713 2099 11747
rect 2041 11707 2099 11713
rect 1302 11636 1308 11688
rect 1360 11676 1366 11688
rect 1670 11676 1676 11688
rect 1360 11648 1676 11676
rect 1360 11636 1366 11648
rect 1670 11636 1676 11648
rect 1728 11636 1734 11688
rect 2056 11676 2084 11707
rect 2130 11704 2136 11756
rect 2188 11744 2194 11756
rect 2409 11747 2467 11753
rect 2409 11744 2421 11747
rect 2188 11716 2421 11744
rect 2188 11704 2194 11716
rect 2409 11713 2421 11716
rect 2455 11713 2467 11747
rect 2409 11707 2467 11713
rect 5258 11704 5264 11756
rect 5316 11744 5322 11756
rect 5316 11716 5948 11744
rect 5316 11704 5322 11716
rect 2590 11676 2596 11688
rect 2056 11648 2596 11676
rect 2590 11636 2596 11648
rect 2648 11636 2654 11688
rect 5626 11636 5632 11688
rect 5684 11676 5690 11688
rect 5813 11679 5871 11685
rect 5813 11676 5825 11679
rect 5684 11648 5825 11676
rect 5684 11636 5690 11648
rect 5813 11645 5825 11648
rect 5859 11645 5871 11679
rect 5813 11639 5871 11645
rect 5920 11608 5948 11716
rect 6012 11685 6040 11784
rect 6086 11704 6092 11756
rect 6144 11744 6150 11756
rect 6270 11744 6276 11756
rect 6144 11716 6276 11744
rect 6144 11704 6150 11716
rect 6270 11704 6276 11716
rect 6328 11744 6334 11756
rect 6365 11747 6423 11753
rect 6365 11744 6377 11747
rect 6328 11716 6377 11744
rect 6328 11704 6334 11716
rect 6365 11713 6377 11716
rect 6411 11713 6423 11747
rect 6564 11744 6592 11784
rect 6638 11753 6644 11756
rect 6365 11707 6423 11713
rect 6472 11716 6592 11744
rect 5997 11679 6055 11685
rect 5997 11645 6009 11679
rect 6043 11645 6055 11679
rect 6472 11676 6500 11716
rect 6632 11707 6644 11753
rect 6696 11744 6702 11756
rect 6696 11716 6732 11744
rect 6638 11704 6644 11707
rect 6696 11704 6702 11716
rect 5997 11639 6055 11645
rect 6380 11648 6500 11676
rect 7576 11676 7604 11784
rect 9140 11756 9168 11852
rect 10870 11840 10876 11852
rect 10928 11840 10934 11892
rect 14274 11880 14280 11892
rect 11532 11852 13860 11880
rect 14235 11852 14280 11880
rect 10502 11812 10508 11824
rect 9416 11784 10508 11812
rect 9416 11756 9444 11784
rect 10502 11772 10508 11784
rect 10560 11772 10566 11824
rect 10594 11772 10600 11824
rect 10652 11812 10658 11824
rect 11532 11812 11560 11852
rect 12158 11821 12164 11824
rect 12152 11812 12164 11821
rect 10652 11784 11560 11812
rect 12119 11784 12164 11812
rect 10652 11772 10658 11784
rect 12152 11775 12164 11784
rect 12158 11772 12164 11775
rect 12216 11772 12222 11824
rect 8205 11747 8263 11753
rect 8205 11713 8217 11747
rect 8251 11744 8263 11747
rect 9122 11744 9128 11756
rect 8251 11716 8892 11744
rect 9035 11716 9128 11744
rect 8251 11713 8263 11716
rect 8205 11707 8263 11713
rect 8294 11676 8300 11688
rect 7576 11648 8300 11676
rect 6380 11608 6408 11648
rect 8294 11636 8300 11648
rect 8352 11636 8358 11688
rect 8389 11679 8447 11685
rect 8389 11645 8401 11679
rect 8435 11645 8447 11679
rect 8389 11639 8447 11645
rect 5920 11580 6408 11608
rect 7745 11611 7803 11617
rect 7745 11577 7757 11611
rect 7791 11608 7803 11611
rect 8110 11608 8116 11620
rect 7791 11580 8116 11608
rect 7791 11577 7803 11580
rect 7745 11571 7803 11577
rect 8110 11568 8116 11580
rect 8168 11568 8174 11620
rect 8404 11608 8432 11639
rect 8220 11580 8432 11608
rect 4062 11500 4068 11552
rect 4120 11540 4126 11552
rect 5353 11543 5411 11549
rect 5353 11540 5365 11543
rect 4120 11512 5365 11540
rect 4120 11500 4126 11512
rect 5353 11509 5365 11512
rect 5399 11509 5411 11543
rect 5353 11503 5411 11509
rect 5442 11500 5448 11552
rect 5500 11540 5506 11552
rect 5626 11540 5632 11552
rect 5500 11512 5632 11540
rect 5500 11500 5506 11512
rect 5626 11500 5632 11512
rect 5684 11500 5690 11552
rect 7006 11500 7012 11552
rect 7064 11540 7070 11552
rect 7837 11543 7895 11549
rect 7837 11540 7849 11543
rect 7064 11512 7849 11540
rect 7064 11500 7070 11512
rect 7837 11509 7849 11512
rect 7883 11509 7895 11543
rect 7837 11503 7895 11509
rect 8018 11500 8024 11552
rect 8076 11540 8082 11552
rect 8220 11540 8248 11580
rect 8662 11540 8668 11552
rect 8076 11512 8248 11540
rect 8623 11512 8668 11540
rect 8076 11500 8082 11512
rect 8662 11500 8668 11512
rect 8720 11500 8726 11552
rect 8864 11540 8892 11716
rect 9122 11704 9128 11716
rect 9180 11704 9186 11756
rect 9398 11753 9404 11756
rect 9392 11744 9404 11753
rect 9359 11716 9404 11744
rect 9392 11707 9404 11716
rect 9398 11704 9404 11707
rect 9456 11704 9462 11756
rect 9674 11704 9680 11756
rect 9732 11744 9738 11756
rect 10965 11747 11023 11753
rect 10965 11744 10977 11747
rect 9732 11716 10977 11744
rect 9732 11704 9738 11716
rect 10965 11713 10977 11716
rect 11011 11713 11023 11747
rect 13262 11744 13268 11756
rect 10965 11707 11023 11713
rect 11348 11716 13268 11744
rect 10778 11676 10784 11688
rect 10520 11648 10784 11676
rect 10520 11617 10548 11648
rect 10778 11636 10784 11648
rect 10836 11636 10842 11688
rect 11348 11617 11376 11716
rect 13262 11704 13268 11716
rect 13320 11704 13326 11756
rect 13832 11744 13860 11852
rect 14274 11840 14280 11852
rect 14332 11840 14338 11892
rect 16945 11883 17003 11889
rect 16945 11880 16957 11883
rect 14660 11852 16957 11880
rect 14660 11744 14688 11852
rect 16945 11849 16957 11852
rect 16991 11849 17003 11883
rect 16945 11843 17003 11849
rect 17497 11883 17555 11889
rect 17497 11849 17509 11883
rect 17543 11880 17555 11883
rect 17770 11880 17776 11892
rect 17543 11852 17776 11880
rect 17543 11849 17555 11852
rect 17497 11843 17555 11849
rect 17770 11840 17776 11852
rect 17828 11840 17834 11892
rect 18322 11880 18328 11892
rect 18283 11852 18328 11880
rect 18322 11840 18328 11852
rect 18380 11840 18386 11892
rect 18785 11883 18843 11889
rect 18785 11849 18797 11883
rect 18831 11880 18843 11883
rect 19153 11883 19211 11889
rect 19153 11880 19165 11883
rect 18831 11852 19165 11880
rect 18831 11849 18843 11852
rect 18785 11843 18843 11849
rect 19153 11849 19165 11852
rect 19199 11849 19211 11883
rect 19153 11843 19211 11849
rect 20349 11883 20407 11889
rect 20349 11849 20361 11883
rect 20395 11880 20407 11883
rect 20530 11880 20536 11892
rect 20395 11852 20536 11880
rect 20395 11849 20407 11852
rect 20349 11843 20407 11849
rect 20530 11840 20536 11852
rect 20588 11840 20594 11892
rect 21358 11880 21364 11892
rect 21319 11852 21364 11880
rect 21358 11840 21364 11852
rect 21416 11840 21422 11892
rect 16114 11772 16120 11824
rect 16172 11812 16178 11824
rect 17310 11812 17316 11824
rect 16172 11784 17316 11812
rect 16172 11772 16178 11784
rect 17310 11772 17316 11784
rect 17368 11812 17374 11824
rect 17957 11815 18015 11821
rect 17368 11784 17908 11812
rect 17368 11772 17374 11784
rect 13832 11716 14688 11744
rect 15401 11747 15459 11753
rect 15401 11713 15413 11747
rect 15447 11744 15459 11747
rect 15562 11744 15568 11756
rect 15447 11716 15568 11744
rect 15447 11713 15459 11716
rect 15401 11707 15459 11713
rect 15562 11704 15568 11716
rect 15620 11704 15626 11756
rect 17037 11747 17095 11753
rect 17037 11713 17049 11747
rect 17083 11744 17095 11747
rect 17126 11744 17132 11756
rect 17083 11716 17132 11744
rect 17083 11713 17095 11716
rect 17037 11707 17095 11713
rect 17126 11704 17132 11716
rect 17184 11704 17190 11756
rect 17880 11753 17908 11784
rect 17957 11781 17969 11815
rect 18003 11812 18015 11815
rect 18003 11784 19104 11812
rect 18003 11781 18015 11784
rect 17957 11775 18015 11781
rect 17865 11747 17923 11753
rect 17865 11713 17877 11747
rect 17911 11713 17923 11747
rect 18690 11744 18696 11756
rect 18651 11716 18696 11744
rect 17865 11707 17923 11713
rect 18690 11704 18696 11716
rect 18748 11704 18754 11756
rect 19076 11688 19104 11784
rect 19242 11772 19248 11824
rect 19300 11812 19306 11824
rect 19521 11815 19579 11821
rect 19521 11812 19533 11815
rect 19300 11784 19533 11812
rect 19300 11772 19306 11784
rect 19521 11781 19533 11784
rect 19567 11812 19579 11815
rect 20806 11812 20812 11824
rect 19567 11784 20812 11812
rect 19567 11781 19579 11784
rect 19521 11775 19579 11781
rect 20806 11772 20812 11784
rect 20864 11772 20870 11824
rect 21269 11747 21327 11753
rect 21269 11713 21281 11747
rect 21315 11744 21327 11747
rect 21542 11744 21548 11756
rect 21315 11716 21548 11744
rect 21315 11713 21327 11716
rect 21269 11707 21327 11713
rect 21542 11704 21548 11716
rect 21600 11704 21606 11756
rect 11882 11676 11888 11688
rect 11716 11648 11888 11676
rect 10505 11611 10563 11617
rect 10505 11577 10517 11611
rect 10551 11577 10563 11611
rect 10505 11571 10563 11577
rect 11333 11611 11391 11617
rect 11333 11577 11345 11611
rect 11379 11577 11391 11611
rect 11333 11571 11391 11577
rect 10410 11540 10416 11552
rect 8864 11512 10416 11540
rect 10410 11500 10416 11512
rect 10468 11500 10474 11552
rect 11606 11500 11612 11552
rect 11664 11540 11670 11552
rect 11716 11549 11744 11648
rect 11882 11636 11888 11648
rect 11940 11636 11946 11688
rect 15654 11676 15660 11688
rect 15615 11648 15660 11676
rect 15654 11636 15660 11648
rect 15712 11636 15718 11688
rect 16853 11679 16911 11685
rect 16853 11645 16865 11679
rect 16899 11676 16911 11679
rect 17586 11676 17592 11688
rect 16899 11648 17592 11676
rect 16899 11645 16911 11648
rect 16853 11639 16911 11645
rect 17586 11636 17592 11648
rect 17644 11636 17650 11688
rect 17954 11636 17960 11688
rect 18012 11676 18018 11688
rect 18049 11679 18107 11685
rect 18049 11676 18061 11679
rect 18012 11648 18061 11676
rect 18012 11636 18018 11648
rect 18049 11645 18061 11648
rect 18095 11645 18107 11679
rect 18874 11676 18880 11688
rect 18835 11648 18880 11676
rect 18049 11639 18107 11645
rect 18874 11636 18880 11648
rect 18932 11636 18938 11688
rect 19058 11636 19064 11688
rect 19116 11676 19122 11688
rect 19613 11679 19671 11685
rect 19613 11676 19625 11679
rect 19116 11648 19625 11676
rect 19116 11636 19122 11648
rect 19613 11645 19625 11648
rect 19659 11645 19671 11679
rect 19794 11676 19800 11688
rect 19755 11648 19800 11676
rect 19613 11639 19671 11645
rect 19794 11636 19800 11648
rect 19852 11636 19858 11688
rect 19978 11676 19984 11688
rect 19939 11648 19984 11676
rect 19978 11636 19984 11648
rect 20036 11636 20042 11688
rect 20717 11679 20775 11685
rect 20717 11645 20729 11679
rect 20763 11676 20775 11679
rect 21358 11676 21364 11688
rect 20763 11648 21364 11676
rect 20763 11645 20775 11648
rect 20717 11639 20775 11645
rect 21358 11636 21364 11648
rect 21416 11636 21422 11688
rect 14093 11611 14151 11617
rect 14093 11577 14105 11611
rect 14139 11608 14151 11611
rect 14274 11608 14280 11620
rect 14139 11580 14280 11608
rect 14139 11577 14151 11580
rect 14093 11571 14151 11577
rect 14274 11568 14280 11580
rect 14332 11568 14338 11620
rect 17405 11611 17463 11617
rect 17405 11577 17417 11611
rect 17451 11608 17463 11611
rect 18230 11608 18236 11620
rect 17451 11580 18236 11608
rect 17451 11577 17463 11580
rect 17405 11571 17463 11577
rect 18230 11568 18236 11580
rect 18288 11568 18294 11620
rect 18322 11568 18328 11620
rect 18380 11608 18386 11620
rect 19242 11608 19248 11620
rect 18380 11580 19248 11608
rect 18380 11568 18386 11580
rect 19242 11568 19248 11580
rect 19300 11568 19306 11620
rect 20901 11611 20959 11617
rect 20901 11577 20913 11611
rect 20947 11608 20959 11611
rect 21450 11608 21456 11620
rect 20947 11580 21456 11608
rect 20947 11577 20959 11580
rect 20901 11571 20959 11577
rect 21450 11568 21456 11580
rect 21508 11568 21514 11620
rect 11701 11543 11759 11549
rect 11701 11540 11713 11543
rect 11664 11512 11713 11540
rect 11664 11500 11670 11512
rect 11701 11509 11713 11512
rect 11747 11509 11759 11543
rect 11701 11503 11759 11509
rect 12986 11500 12992 11552
rect 13044 11540 13050 11552
rect 13265 11543 13323 11549
rect 13265 11540 13277 11543
rect 13044 11512 13277 11540
rect 13044 11500 13050 11512
rect 13265 11509 13277 11512
rect 13311 11509 13323 11543
rect 13265 11503 13323 11509
rect 13354 11500 13360 11552
rect 13412 11540 13418 11552
rect 16574 11540 16580 11552
rect 13412 11512 16580 11540
rect 13412 11500 13418 11512
rect 16574 11500 16580 11512
rect 16632 11500 16638 11552
rect 17770 11500 17776 11552
rect 17828 11540 17834 11552
rect 20162 11540 20168 11552
rect 17828 11512 20168 11540
rect 17828 11500 17834 11512
rect 20162 11500 20168 11512
rect 20220 11500 20226 11552
rect 21082 11540 21088 11552
rect 21043 11512 21088 11540
rect 21082 11500 21088 11512
rect 21140 11500 21146 11552
rect 1104 11450 21896 11472
rect 1104 11398 3549 11450
rect 3601 11398 3613 11450
rect 3665 11398 3677 11450
rect 3729 11398 3741 11450
rect 3793 11398 3805 11450
rect 3857 11398 8747 11450
rect 8799 11398 8811 11450
rect 8863 11398 8875 11450
rect 8927 11398 8939 11450
rect 8991 11398 9003 11450
rect 9055 11398 13945 11450
rect 13997 11398 14009 11450
rect 14061 11398 14073 11450
rect 14125 11398 14137 11450
rect 14189 11398 14201 11450
rect 14253 11398 19143 11450
rect 19195 11398 19207 11450
rect 19259 11398 19271 11450
rect 19323 11398 19335 11450
rect 19387 11398 19399 11450
rect 19451 11398 21896 11450
rect 1104 11376 21896 11398
rect 1946 11336 1952 11348
rect 1907 11308 1952 11336
rect 1946 11296 1952 11308
rect 2004 11296 2010 11348
rect 6914 11336 6920 11348
rect 2746 11308 6920 11336
rect 1673 11271 1731 11277
rect 1673 11237 1685 11271
rect 1719 11268 1731 11271
rect 2746 11268 2774 11308
rect 6914 11296 6920 11308
rect 6972 11296 6978 11348
rect 7282 11336 7288 11348
rect 7243 11308 7288 11336
rect 7282 11296 7288 11308
rect 7340 11296 7346 11348
rect 9122 11296 9128 11348
rect 9180 11336 9186 11348
rect 10689 11339 10747 11345
rect 10689 11336 10701 11339
rect 9180 11308 10701 11336
rect 9180 11296 9186 11308
rect 10689 11305 10701 11308
rect 10735 11336 10747 11339
rect 11606 11336 11612 11348
rect 10735 11308 11612 11336
rect 10735 11305 10747 11308
rect 10689 11299 10747 11305
rect 5902 11268 5908 11280
rect 1719 11240 2774 11268
rect 4356 11240 5908 11268
rect 1719 11237 1731 11240
rect 1673 11231 1731 11237
rect 2685 11203 2743 11209
rect 2685 11169 2697 11203
rect 2731 11200 2743 11203
rect 4356 11200 4384 11240
rect 5902 11228 5908 11240
rect 5960 11228 5966 11280
rect 8757 11271 8815 11277
rect 8757 11237 8769 11271
rect 8803 11237 8815 11271
rect 8757 11231 8815 11237
rect 2731 11172 4384 11200
rect 4433 11203 4491 11209
rect 2731 11169 2743 11172
rect 2685 11163 2743 11169
rect 4433 11169 4445 11203
rect 4479 11169 4491 11203
rect 4433 11163 4491 11169
rect 5077 11203 5135 11209
rect 5077 11169 5089 11203
rect 5123 11200 5135 11203
rect 5166 11200 5172 11212
rect 5123 11172 5172 11200
rect 5123 11169 5135 11172
rect 5077 11163 5135 11169
rect 1765 11135 1823 11141
rect 1765 11101 1777 11135
rect 1811 11132 1823 11135
rect 2222 11132 2228 11144
rect 1811 11104 2228 11132
rect 1811 11101 1823 11104
rect 1765 11095 1823 11101
rect 2222 11092 2228 11104
rect 2280 11092 2286 11144
rect 2501 11135 2559 11141
rect 2501 11101 2513 11135
rect 2547 11132 2559 11135
rect 3234 11132 3240 11144
rect 2547 11104 3240 11132
rect 2547 11101 2559 11104
rect 2501 11095 2559 11101
rect 3234 11092 3240 11104
rect 3292 11092 3298 11144
rect 4157 11135 4215 11141
rect 4157 11101 4169 11135
rect 4203 11132 4215 11135
rect 4338 11132 4344 11144
rect 4203 11104 4344 11132
rect 4203 11101 4215 11104
rect 4157 11095 4215 11101
rect 4338 11092 4344 11104
rect 4396 11092 4402 11144
rect 4448 11132 4476 11163
rect 5166 11160 5172 11172
rect 5224 11160 5230 11212
rect 8478 11160 8484 11212
rect 8536 11200 8542 11212
rect 8772 11200 8800 11231
rect 10704 11200 10732 11299
rect 11606 11296 11612 11308
rect 11664 11336 11670 11348
rect 11664 11308 13952 11336
rect 11664 11296 11670 11308
rect 10873 11203 10931 11209
rect 10873 11200 10885 11203
rect 8536 11172 9076 11200
rect 10704 11172 10885 11200
rect 8536 11160 8542 11172
rect 4798 11132 4804 11144
rect 4448 11104 4804 11132
rect 4798 11092 4804 11104
rect 4856 11092 4862 11144
rect 5813 11135 5871 11141
rect 5813 11101 5825 11135
rect 5859 11132 5871 11135
rect 5905 11135 5963 11141
rect 5905 11132 5917 11135
rect 5859 11104 5917 11132
rect 5859 11101 5871 11104
rect 5813 11095 5871 11101
rect 5905 11101 5917 11104
rect 5951 11132 5963 11135
rect 6546 11132 6552 11144
rect 5951 11104 6552 11132
rect 5951 11101 5963 11104
rect 5905 11095 5963 11101
rect 6288 11076 6316 11104
rect 6546 11092 6552 11104
rect 6604 11132 6610 11144
rect 7377 11135 7435 11141
rect 7377 11132 7389 11135
rect 6604 11104 7389 11132
rect 6604 11092 6610 11104
rect 7377 11101 7389 11104
rect 7423 11132 7435 11135
rect 8941 11135 8999 11141
rect 8941 11132 8953 11135
rect 7423 11104 8953 11132
rect 7423 11101 7435 11104
rect 7377 11095 7435 11101
rect 8941 11101 8953 11104
rect 8987 11101 8999 11135
rect 9048 11132 9076 11172
rect 10873 11169 10885 11172
rect 10919 11169 10931 11203
rect 10873 11163 10931 11169
rect 12250 11160 12256 11212
rect 12308 11200 12314 11212
rect 12360 11209 12388 11308
rect 13725 11271 13783 11277
rect 13725 11237 13737 11271
rect 13771 11268 13783 11271
rect 13814 11268 13820 11280
rect 13771 11240 13820 11268
rect 13771 11237 13783 11240
rect 13725 11231 13783 11237
rect 13814 11228 13820 11240
rect 13872 11228 13878 11280
rect 12345 11203 12403 11209
rect 12345 11200 12357 11203
rect 12308 11172 12357 11200
rect 12308 11160 12314 11172
rect 12345 11169 12357 11172
rect 12391 11169 12403 11203
rect 12345 11163 12403 11169
rect 9214 11141 9220 11144
rect 9208 11132 9220 11141
rect 9048 11104 9220 11132
rect 8941 11095 8999 11101
rect 9208 11095 9220 11104
rect 9214 11092 9220 11095
rect 9272 11092 9278 11144
rect 10778 11132 10784 11144
rect 9324 11104 10784 11132
rect 1486 11064 1492 11076
rect 1447 11036 1492 11064
rect 1486 11024 1492 11036
rect 1544 11064 1550 11076
rect 2869 11067 2927 11073
rect 2869 11064 2881 11067
rect 1544 11036 2881 11064
rect 1544 11024 1550 11036
rect 2869 11033 2881 11036
rect 2915 11033 2927 11067
rect 2869 11027 2927 11033
rect 3326 11024 3332 11076
rect 3384 11064 3390 11076
rect 4617 11067 4675 11073
rect 4617 11064 4629 11067
rect 3384 11036 4629 11064
rect 3384 11024 3390 11036
rect 4617 11033 4629 11036
rect 4663 11033 4675 11067
rect 4617 11027 4675 11033
rect 5074 11024 5080 11076
rect 5132 11064 5138 11076
rect 6150 11067 6208 11073
rect 6150 11064 6162 11067
rect 5132 11036 6162 11064
rect 5132 11024 5138 11036
rect 6150 11033 6162 11036
rect 6196 11033 6208 11067
rect 6150 11027 6208 11033
rect 6270 11024 6276 11076
rect 6328 11024 6334 11076
rect 7644 11067 7702 11073
rect 7644 11033 7656 11067
rect 7690 11064 7702 11067
rect 8110 11064 8116 11076
rect 7690 11036 8116 11064
rect 7690 11033 7702 11036
rect 7644 11027 7702 11033
rect 8110 11024 8116 11036
rect 8168 11024 8174 11076
rect 8294 11024 8300 11076
rect 8352 11064 8358 11076
rect 9324 11064 9352 11104
rect 10778 11092 10784 11104
rect 10836 11092 10842 11144
rect 11140 11135 11198 11141
rect 11140 11101 11152 11135
rect 11186 11132 11198 11135
rect 11698 11132 11704 11144
rect 11186 11104 11704 11132
rect 11186 11101 11198 11104
rect 11140 11095 11198 11101
rect 11698 11092 11704 11104
rect 11756 11092 11762 11144
rect 13924 11141 13952 11308
rect 14734 11296 14740 11348
rect 14792 11336 14798 11348
rect 15841 11339 15899 11345
rect 14792 11308 15056 11336
rect 14792 11296 14798 11308
rect 15028 11268 15056 11308
rect 15841 11305 15853 11339
rect 15887 11336 15899 11339
rect 16942 11336 16948 11348
rect 15887 11308 16948 11336
rect 15887 11305 15899 11308
rect 15841 11299 15899 11305
rect 16942 11296 16948 11308
rect 17000 11296 17006 11348
rect 17126 11336 17132 11348
rect 17087 11308 17132 11336
rect 17126 11296 17132 11308
rect 17184 11296 17190 11348
rect 17310 11336 17316 11348
rect 17271 11308 17316 11336
rect 17310 11296 17316 11308
rect 17368 11296 17374 11348
rect 18690 11296 18696 11348
rect 18748 11336 18754 11348
rect 19245 11339 19303 11345
rect 19245 11336 19257 11339
rect 18748 11308 19257 11336
rect 18748 11296 18754 11308
rect 19245 11305 19257 11308
rect 19291 11305 19303 11339
rect 20162 11336 20168 11348
rect 20123 11308 20168 11336
rect 19245 11299 19303 11305
rect 20162 11296 20168 11308
rect 20220 11336 20226 11348
rect 20806 11336 20812 11348
rect 20220 11308 20812 11336
rect 20220 11296 20226 11308
rect 20806 11296 20812 11308
rect 20864 11336 20870 11348
rect 21174 11336 21180 11348
rect 20864 11308 21180 11336
rect 20864 11296 20870 11308
rect 21174 11296 21180 11308
rect 21232 11296 21238 11348
rect 15473 11271 15531 11277
rect 15028 11240 15148 11268
rect 15120 11200 15148 11240
rect 15473 11237 15485 11271
rect 15519 11268 15531 11271
rect 15562 11268 15568 11280
rect 15519 11240 15568 11268
rect 15519 11237 15531 11240
rect 15473 11231 15531 11237
rect 15562 11228 15568 11240
rect 15620 11268 15626 11280
rect 17678 11268 17684 11280
rect 15620 11240 17684 11268
rect 15620 11228 15626 11240
rect 17678 11228 17684 11240
rect 17736 11228 17742 11280
rect 18782 11228 18788 11280
rect 18840 11268 18846 11280
rect 20625 11271 20683 11277
rect 20625 11268 20637 11271
rect 18840 11240 20637 11268
rect 18840 11228 18846 11240
rect 20625 11237 20637 11240
rect 20671 11237 20683 11271
rect 20625 11231 20683 11237
rect 16206 11200 16212 11212
rect 15120 11172 16212 11200
rect 16206 11160 16212 11172
rect 16264 11160 16270 11212
rect 16574 11200 16580 11212
rect 16487 11172 16580 11200
rect 16574 11160 16580 11172
rect 16632 11200 16638 11212
rect 17954 11200 17960 11212
rect 16632 11172 17960 11200
rect 16632 11160 16638 11172
rect 17954 11160 17960 11172
rect 18012 11160 18018 11212
rect 18690 11160 18696 11212
rect 18748 11200 18754 11212
rect 19058 11200 19064 11212
rect 18748 11172 19064 11200
rect 18748 11160 18754 11172
rect 19058 11160 19064 11172
rect 19116 11160 19122 11212
rect 19794 11200 19800 11212
rect 19755 11172 19800 11200
rect 19794 11160 19800 11172
rect 19852 11160 19858 11212
rect 20901 11203 20959 11209
rect 20901 11169 20913 11203
rect 20947 11200 20959 11203
rect 21174 11200 21180 11212
rect 20947 11172 21180 11200
rect 20947 11169 20959 11172
rect 20901 11163 20959 11169
rect 21174 11160 21180 11172
rect 21232 11160 21238 11212
rect 13909 11135 13967 11141
rect 12268 11104 13860 11132
rect 8352 11036 9352 11064
rect 8352 11024 8358 11036
rect 9398 11024 9404 11076
rect 9456 11064 9462 11076
rect 9456 11036 10364 11064
rect 9456 11024 9462 11036
rect 2038 10956 2044 11008
rect 2096 10996 2102 11008
rect 2406 10996 2412 11008
rect 2096 10968 2141 10996
rect 2367 10968 2412 10996
rect 2096 10956 2102 10968
rect 2406 10956 2412 10968
rect 2464 10956 2470 11008
rect 2774 10956 2780 11008
rect 2832 10996 2838 11008
rect 3789 10999 3847 11005
rect 3789 10996 3801 10999
rect 2832 10968 3801 10996
rect 2832 10956 2838 10968
rect 3789 10965 3801 10968
rect 3835 10965 3847 10999
rect 4246 10996 4252 11008
rect 4207 10968 4252 10996
rect 3789 10959 3847 10965
rect 4246 10956 4252 10968
rect 4304 10956 4310 11008
rect 10336 11005 10364 11036
rect 12268 11005 12296 11104
rect 12612 11067 12670 11073
rect 12612 11033 12624 11067
rect 12658 11064 12670 11067
rect 13078 11064 13084 11076
rect 12658 11036 13084 11064
rect 12658 11033 12670 11036
rect 12612 11027 12670 11033
rect 13078 11024 13084 11036
rect 13136 11024 13142 11076
rect 13832 11064 13860 11104
rect 13909 11101 13921 11135
rect 13955 11132 13967 11135
rect 14090 11132 14096 11144
rect 13955 11104 14096 11132
rect 13955 11101 13967 11104
rect 13909 11095 13967 11101
rect 14090 11092 14096 11104
rect 14148 11092 14154 11144
rect 18414 11132 18420 11144
rect 14384 11104 18420 11132
rect 14384 11073 14412 11104
rect 18414 11092 18420 11104
rect 18472 11092 18478 11144
rect 18598 11092 18604 11144
rect 18656 11132 18662 11144
rect 18785 11135 18843 11141
rect 18785 11132 18797 11135
rect 18656 11104 18797 11132
rect 18656 11092 18662 11104
rect 18785 11101 18797 11104
rect 18831 11101 18843 11135
rect 18969 11135 19027 11141
rect 18969 11132 18981 11135
rect 18785 11095 18843 11101
rect 18892 11104 18981 11132
rect 14338 11067 14412 11073
rect 14338 11064 14350 11067
rect 13832 11036 14350 11064
rect 14338 11033 14350 11036
rect 14384 11036 14412 11067
rect 14384 11033 14396 11036
rect 14338 11027 14396 11033
rect 14458 11024 14464 11076
rect 14516 11064 14522 11076
rect 15749 11067 15807 11073
rect 15749 11064 15761 11067
rect 14516 11036 15761 11064
rect 14516 11024 14522 11036
rect 15749 11033 15761 11036
rect 15795 11033 15807 11067
rect 15749 11027 15807 11033
rect 16206 11024 16212 11076
rect 16264 11064 16270 11076
rect 16669 11067 16727 11073
rect 16669 11064 16681 11067
rect 16264 11036 16681 11064
rect 16264 11024 16270 11036
rect 16669 11033 16681 11036
rect 16715 11033 16727 11067
rect 16669 11027 16727 11033
rect 16761 11067 16819 11073
rect 16761 11033 16773 11067
rect 16807 11064 16819 11067
rect 17954 11064 17960 11076
rect 16807 11036 17960 11064
rect 16807 11033 16819 11036
rect 16761 11027 16819 11033
rect 17954 11024 17960 11036
rect 18012 11024 18018 11076
rect 18322 11024 18328 11076
rect 18380 11064 18386 11076
rect 18892 11064 18920 11104
rect 18969 11101 18981 11104
rect 19015 11101 19027 11135
rect 18969 11095 19027 11101
rect 19613 11135 19671 11141
rect 19613 11101 19625 11135
rect 19659 11132 19671 11135
rect 19978 11132 19984 11144
rect 19659 11104 19984 11132
rect 19659 11101 19671 11104
rect 19613 11095 19671 11101
rect 19978 11092 19984 11104
rect 20036 11092 20042 11144
rect 20809 11135 20867 11141
rect 20809 11101 20821 11135
rect 20855 11101 20867 11135
rect 20809 11095 20867 11101
rect 18380 11036 18920 11064
rect 18380 11024 18386 11036
rect 19242 11024 19248 11076
rect 19300 11064 19306 11076
rect 19705 11067 19763 11073
rect 19705 11064 19717 11067
rect 19300 11036 19717 11064
rect 19300 11024 19306 11036
rect 19705 11033 19717 11036
rect 19751 11064 19763 11067
rect 20346 11064 20352 11076
rect 19751 11036 20352 11064
rect 19751 11033 19763 11036
rect 19705 11027 19763 11033
rect 20346 11024 20352 11036
rect 20404 11024 20410 11076
rect 20530 11064 20536 11076
rect 20491 11036 20536 11064
rect 20530 11024 20536 11036
rect 20588 11064 20594 11076
rect 20824 11064 20852 11095
rect 20990 11092 20996 11144
rect 21048 11132 21054 11144
rect 21269 11135 21327 11141
rect 21269 11132 21281 11135
rect 21048 11104 21281 11132
rect 21048 11092 21054 11104
rect 21269 11101 21281 11104
rect 21315 11101 21327 11135
rect 21450 11132 21456 11144
rect 21411 11104 21456 11132
rect 21269 11095 21327 11101
rect 21450 11092 21456 11104
rect 21508 11092 21514 11144
rect 21082 11064 21088 11076
rect 20588 11036 20852 11064
rect 21043 11036 21088 11064
rect 20588 11024 20594 11036
rect 21082 11024 21088 11036
rect 21140 11024 21146 11076
rect 10321 10999 10379 11005
rect 10321 10965 10333 10999
rect 10367 10965 10379 10999
rect 10321 10959 10379 10965
rect 12253 10999 12311 11005
rect 12253 10965 12265 10999
rect 12299 10965 12311 10999
rect 13096 10996 13124 11024
rect 16390 10996 16396 11008
rect 13096 10968 16396 10996
rect 12253 10959 12311 10965
rect 16390 10956 16396 10968
rect 16448 10956 16454 11008
rect 19426 10956 19432 11008
rect 19484 10996 19490 11008
rect 19886 10996 19892 11008
rect 19484 10968 19892 10996
rect 19484 10956 19490 10968
rect 19886 10956 19892 10968
rect 19944 10956 19950 11008
rect 1104 10906 22056 10928
rect 1104 10854 6148 10906
rect 6200 10854 6212 10906
rect 6264 10854 6276 10906
rect 6328 10854 6340 10906
rect 6392 10854 6404 10906
rect 6456 10854 11346 10906
rect 11398 10854 11410 10906
rect 11462 10854 11474 10906
rect 11526 10854 11538 10906
rect 11590 10854 11602 10906
rect 11654 10854 16544 10906
rect 16596 10854 16608 10906
rect 16660 10854 16672 10906
rect 16724 10854 16736 10906
rect 16788 10854 16800 10906
rect 16852 10854 21742 10906
rect 21794 10854 21806 10906
rect 21858 10854 21870 10906
rect 21922 10854 21934 10906
rect 21986 10854 21998 10906
rect 22050 10854 22056 10906
rect 1104 10832 22056 10854
rect 1765 10795 1823 10801
rect 1765 10761 1777 10795
rect 1811 10792 1823 10795
rect 2038 10792 2044 10804
rect 1811 10764 2044 10792
rect 1811 10761 1823 10764
rect 1765 10755 1823 10761
rect 2038 10752 2044 10764
rect 2096 10752 2102 10804
rect 2222 10792 2228 10804
rect 2183 10764 2228 10792
rect 2222 10752 2228 10764
rect 2280 10752 2286 10804
rect 2317 10795 2375 10801
rect 2317 10761 2329 10795
rect 2363 10792 2375 10795
rect 2406 10792 2412 10804
rect 2363 10764 2412 10792
rect 2363 10761 2375 10764
rect 2317 10755 2375 10761
rect 2406 10752 2412 10764
rect 2464 10752 2470 10804
rect 2774 10752 2780 10804
rect 2832 10792 2838 10804
rect 3789 10795 3847 10801
rect 2832 10764 2877 10792
rect 2832 10752 2838 10764
rect 3789 10761 3801 10795
rect 3835 10792 3847 10795
rect 3970 10792 3976 10804
rect 3835 10764 3976 10792
rect 3835 10761 3847 10764
rect 3789 10755 3847 10761
rect 3970 10752 3976 10764
rect 4028 10752 4034 10804
rect 4154 10752 4160 10804
rect 4212 10792 4218 10804
rect 4614 10792 4620 10804
rect 4212 10764 4620 10792
rect 4212 10752 4218 10764
rect 4614 10752 4620 10764
rect 4672 10752 4678 10804
rect 4706 10752 4712 10804
rect 4764 10752 4770 10804
rect 10134 10752 10140 10804
rect 10192 10792 10198 10804
rect 10321 10795 10379 10801
rect 10321 10792 10333 10795
rect 10192 10764 10333 10792
rect 10192 10752 10198 10764
rect 10321 10761 10333 10764
rect 10367 10761 10379 10795
rect 10321 10755 10379 10761
rect 10410 10752 10416 10804
rect 10468 10792 10474 10804
rect 10781 10795 10839 10801
rect 10781 10792 10793 10795
rect 10468 10764 10793 10792
rect 10468 10752 10474 10764
rect 10781 10761 10793 10764
rect 10827 10761 10839 10795
rect 12250 10792 12256 10804
rect 12211 10764 12256 10792
rect 10781 10755 10839 10761
rect 12250 10752 12256 10764
rect 12308 10752 12314 10804
rect 14090 10752 14096 10804
rect 14148 10792 14154 10804
rect 14185 10795 14243 10801
rect 14185 10792 14197 10795
rect 14148 10764 14197 10792
rect 14148 10752 14154 10764
rect 14185 10761 14197 10764
rect 14231 10792 14243 10795
rect 15654 10792 15660 10804
rect 14231 10764 15660 10792
rect 14231 10761 14243 10764
rect 14185 10755 14243 10761
rect 15654 10752 15660 10764
rect 15712 10752 15718 10804
rect 16758 10752 16764 10804
rect 16816 10792 16822 10804
rect 17034 10792 17040 10804
rect 16816 10764 17040 10792
rect 16816 10752 16822 10764
rect 17034 10752 17040 10764
rect 17092 10752 17098 10804
rect 17681 10795 17739 10801
rect 17681 10761 17693 10795
rect 17727 10792 17739 10795
rect 18049 10795 18107 10801
rect 18049 10792 18061 10795
rect 17727 10764 18061 10792
rect 17727 10761 17739 10764
rect 17681 10755 17739 10761
rect 18049 10761 18061 10764
rect 18095 10761 18107 10795
rect 18049 10755 18107 10761
rect 18138 10752 18144 10804
rect 18196 10792 18202 10804
rect 18509 10795 18567 10801
rect 18509 10792 18521 10795
rect 18196 10764 18521 10792
rect 18196 10752 18202 10764
rect 18509 10761 18521 10764
rect 18555 10761 18567 10795
rect 18509 10755 18567 10761
rect 19702 10752 19708 10804
rect 19760 10792 19766 10804
rect 19797 10795 19855 10801
rect 19797 10792 19809 10795
rect 19760 10764 19809 10792
rect 19760 10752 19766 10764
rect 19797 10761 19809 10764
rect 19843 10761 19855 10795
rect 19797 10755 19855 10761
rect 19886 10752 19892 10804
rect 19944 10752 19950 10804
rect 20073 10795 20131 10801
rect 20073 10761 20085 10795
rect 20119 10792 20131 10795
rect 20622 10792 20628 10804
rect 20119 10764 20628 10792
rect 20119 10761 20131 10764
rect 20073 10755 20131 10761
rect 20622 10752 20628 10764
rect 20680 10752 20686 10804
rect 20806 10792 20812 10804
rect 20767 10764 20812 10792
rect 20806 10752 20812 10764
rect 20864 10752 20870 10804
rect 4724 10724 4752 10752
rect 5166 10724 5172 10736
rect 4632 10696 5172 10724
rect 1762 10616 1768 10668
rect 1820 10656 1826 10668
rect 1857 10659 1915 10665
rect 1857 10656 1869 10659
rect 1820 10628 1869 10656
rect 1820 10616 1826 10628
rect 1857 10625 1869 10628
rect 1903 10625 1915 10659
rect 2682 10656 2688 10668
rect 2643 10628 2688 10656
rect 1857 10619 1915 10625
rect 2682 10616 2688 10628
rect 2740 10616 2746 10668
rect 4632 10665 4660 10696
rect 5166 10684 5172 10696
rect 5224 10684 5230 10736
rect 7374 10684 7380 10736
rect 7432 10724 7438 10736
rect 7478 10727 7536 10733
rect 7478 10724 7490 10727
rect 7432 10696 7490 10724
rect 7432 10684 7438 10696
rect 7478 10693 7490 10696
rect 7524 10693 7536 10727
rect 7478 10687 7536 10693
rect 9208 10727 9266 10733
rect 9208 10693 9220 10727
rect 9254 10724 9266 10727
rect 12158 10724 12164 10736
rect 9254 10696 12164 10724
rect 9254 10693 9266 10696
rect 9208 10687 9266 10693
rect 12158 10684 12164 10696
rect 12216 10684 12222 10736
rect 15378 10684 15384 10736
rect 15436 10733 15442 10736
rect 15436 10724 15448 10733
rect 19610 10724 19616 10736
rect 15436 10696 15481 10724
rect 19352 10696 19616 10724
rect 15436 10687 15448 10696
rect 15436 10684 15442 10687
rect 4617 10659 4675 10665
rect 4617 10625 4629 10659
rect 4663 10625 4675 10659
rect 4617 10619 4675 10625
rect 4709 10659 4767 10665
rect 4709 10625 4721 10659
rect 4755 10656 4767 10659
rect 5353 10659 5411 10665
rect 5353 10656 5365 10659
rect 4755 10628 5365 10656
rect 4755 10625 4767 10628
rect 4709 10619 4767 10625
rect 5353 10625 5365 10628
rect 5399 10656 5411 10659
rect 10689 10659 10747 10665
rect 5399 10628 10640 10656
rect 5399 10625 5411 10628
rect 5353 10619 5411 10625
rect 1673 10591 1731 10597
rect 1673 10557 1685 10591
rect 1719 10557 1731 10591
rect 2958 10588 2964 10600
rect 2919 10560 2964 10588
rect 1673 10551 1731 10557
rect 1688 10520 1716 10551
rect 2958 10548 2964 10560
rect 3016 10548 3022 10600
rect 3878 10588 3884 10600
rect 3839 10560 3884 10588
rect 3878 10548 3884 10560
rect 3936 10548 3942 10600
rect 4065 10591 4123 10597
rect 4065 10557 4077 10591
rect 4111 10588 4123 10591
rect 4154 10588 4160 10600
rect 4111 10560 4160 10588
rect 4111 10557 4123 10560
rect 4065 10551 4123 10557
rect 4154 10548 4160 10560
rect 4212 10548 4218 10600
rect 4798 10588 4804 10600
rect 4759 10560 4804 10588
rect 4798 10548 4804 10560
rect 4856 10548 4862 10600
rect 5074 10548 5080 10600
rect 5132 10548 5138 10600
rect 7745 10591 7803 10597
rect 7745 10557 7757 10591
rect 7791 10557 7803 10591
rect 8941 10591 8999 10597
rect 8941 10588 8953 10591
rect 7745 10551 7803 10557
rect 8772 10560 8953 10588
rect 5092 10520 5120 10548
rect 1688 10492 5120 10520
rect 6181 10523 6239 10529
rect 6181 10489 6193 10523
rect 6227 10520 6239 10523
rect 6546 10520 6552 10532
rect 6227 10492 6552 10520
rect 6227 10489 6239 10492
rect 6181 10483 6239 10489
rect 6546 10480 6552 10492
rect 6604 10480 6610 10532
rect 3418 10452 3424 10464
rect 3379 10424 3424 10452
rect 3418 10412 3424 10424
rect 3476 10412 3482 10464
rect 4246 10452 4252 10464
rect 4207 10424 4252 10452
rect 4246 10412 4252 10424
rect 4304 10412 4310 10464
rect 5166 10452 5172 10464
rect 5127 10424 5172 10452
rect 5166 10412 5172 10424
rect 5224 10412 5230 10464
rect 6362 10452 6368 10464
rect 6323 10424 6368 10452
rect 6362 10412 6368 10424
rect 6420 10412 6426 10464
rect 6564 10452 6592 10480
rect 7760 10452 7788 10551
rect 8772 10461 8800 10560
rect 8941 10557 8953 10560
rect 8987 10557 8999 10591
rect 8941 10551 8999 10557
rect 10505 10591 10563 10597
rect 10505 10557 10517 10591
rect 10551 10557 10563 10591
rect 10612 10588 10640 10628
rect 10689 10625 10701 10659
rect 10735 10656 10747 10659
rect 10778 10656 10784 10668
rect 10735 10628 10784 10656
rect 10735 10625 10747 10628
rect 10689 10619 10747 10625
rect 10778 10616 10784 10628
rect 10836 10616 10842 10668
rect 17313 10659 17371 10665
rect 17313 10625 17325 10659
rect 17359 10656 17371 10659
rect 17402 10656 17408 10668
rect 17359 10628 17408 10656
rect 17359 10625 17371 10628
rect 17313 10619 17371 10625
rect 17402 10616 17408 10628
rect 17460 10616 17466 10668
rect 18141 10659 18199 10665
rect 18141 10625 18153 10659
rect 18187 10656 18199 10659
rect 18322 10656 18328 10668
rect 18187 10628 18328 10656
rect 18187 10625 18199 10628
rect 18141 10619 18199 10625
rect 18322 10616 18328 10628
rect 18380 10616 18386 10668
rect 19352 10656 19380 10696
rect 19610 10684 19616 10696
rect 19668 10724 19674 10736
rect 19904 10724 19932 10752
rect 19668 10696 19932 10724
rect 19668 10684 19674 10696
rect 19260 10628 19380 10656
rect 14642 10588 14648 10600
rect 10612 10560 14648 10588
rect 10505 10551 10563 10557
rect 7837 10455 7895 10461
rect 7837 10452 7849 10455
rect 6564 10424 7849 10452
rect 7837 10421 7849 10424
rect 7883 10452 7895 10455
rect 8573 10455 8631 10461
rect 8573 10452 8585 10455
rect 7883 10424 8585 10452
rect 7883 10421 7895 10424
rect 7837 10415 7895 10421
rect 8573 10421 8585 10424
rect 8619 10452 8631 10455
rect 8757 10455 8815 10461
rect 8757 10452 8769 10455
rect 8619 10424 8769 10452
rect 8619 10421 8631 10424
rect 8573 10415 8631 10421
rect 8757 10421 8769 10424
rect 8803 10421 8815 10455
rect 10520 10452 10548 10551
rect 14642 10548 14648 10560
rect 14700 10548 14706 10600
rect 15654 10588 15660 10600
rect 15615 10560 15660 10588
rect 15654 10548 15660 10560
rect 15712 10548 15718 10600
rect 16390 10548 16396 10600
rect 16448 10588 16454 10600
rect 17034 10588 17040 10600
rect 16448 10560 17040 10588
rect 16448 10548 16454 10560
rect 17034 10548 17040 10560
rect 17092 10548 17098 10600
rect 17218 10588 17224 10600
rect 17179 10560 17224 10588
rect 17218 10548 17224 10560
rect 17276 10548 17282 10600
rect 17957 10591 18015 10597
rect 17957 10557 17969 10591
rect 18003 10588 18015 10591
rect 18874 10588 18880 10600
rect 18003 10560 18880 10588
rect 18003 10557 18015 10560
rect 17957 10551 18015 10557
rect 18874 10548 18880 10560
rect 18932 10548 18938 10600
rect 19260 10597 19288 10628
rect 19426 10616 19432 10668
rect 19484 10656 19490 10668
rect 19889 10659 19947 10665
rect 19484 10628 19577 10656
rect 19484 10616 19490 10628
rect 19889 10625 19901 10659
rect 19935 10656 19947 10659
rect 19978 10656 19984 10668
rect 19935 10628 19984 10656
rect 19935 10625 19947 10628
rect 19889 10619 19947 10625
rect 19978 10616 19984 10628
rect 20036 10616 20042 10668
rect 20070 10616 20076 10668
rect 20128 10656 20134 10668
rect 20165 10659 20223 10665
rect 20165 10656 20177 10659
rect 20128 10628 20177 10656
rect 20128 10616 20134 10628
rect 20165 10625 20177 10628
rect 20211 10656 20223 10659
rect 20717 10659 20775 10665
rect 20717 10656 20729 10659
rect 20211 10628 20729 10656
rect 20211 10625 20223 10628
rect 20165 10619 20223 10625
rect 20717 10625 20729 10628
rect 20763 10625 20775 10659
rect 21450 10656 21456 10668
rect 21411 10628 21456 10656
rect 20717 10619 20775 10625
rect 21450 10616 21456 10628
rect 21508 10616 21514 10668
rect 19245 10591 19303 10597
rect 19245 10557 19257 10591
rect 19291 10557 19303 10591
rect 19245 10551 19303 10557
rect 19337 10591 19395 10597
rect 19337 10557 19349 10591
rect 19383 10557 19395 10591
rect 19337 10551 19395 10557
rect 11149 10523 11207 10529
rect 11149 10489 11161 10523
rect 11195 10520 11207 10523
rect 11195 10492 14780 10520
rect 11195 10489 11207 10492
rect 11149 10483 11207 10489
rect 14277 10455 14335 10461
rect 14277 10452 14289 10455
rect 10520 10424 14289 10452
rect 8757 10415 8815 10421
rect 14277 10421 14289 10424
rect 14323 10452 14335 10455
rect 14458 10452 14464 10464
rect 14323 10424 14464 10452
rect 14323 10421 14335 10424
rect 14277 10415 14335 10421
rect 14458 10412 14464 10424
rect 14516 10412 14522 10464
rect 14752 10452 14780 10492
rect 18690 10480 18696 10532
rect 18748 10520 18754 10532
rect 19352 10520 19380 10551
rect 18748 10492 19380 10520
rect 18748 10480 18754 10492
rect 16390 10452 16396 10464
rect 14752 10424 16396 10452
rect 16390 10412 16396 10424
rect 16448 10412 16454 10464
rect 18874 10412 18880 10464
rect 18932 10452 18938 10464
rect 18969 10455 19027 10461
rect 18969 10452 18981 10455
rect 18932 10424 18981 10452
rect 18932 10412 18938 10424
rect 18969 10421 18981 10424
rect 19015 10452 19027 10455
rect 19444 10452 19472 10616
rect 20806 10548 20812 10600
rect 20864 10588 20870 10600
rect 20901 10591 20959 10597
rect 20901 10588 20913 10591
rect 20864 10560 20913 10588
rect 20864 10548 20870 10560
rect 20901 10557 20913 10560
rect 20947 10557 20959 10591
rect 20901 10551 20959 10557
rect 20714 10480 20720 10532
rect 20772 10520 20778 10532
rect 21269 10523 21327 10529
rect 21269 10520 21281 10523
rect 20772 10492 21281 10520
rect 20772 10480 20778 10492
rect 21269 10489 21281 10492
rect 21315 10489 21327 10523
rect 21269 10483 21327 10489
rect 19015 10424 19472 10452
rect 20349 10455 20407 10461
rect 19015 10421 19027 10424
rect 18969 10415 19027 10421
rect 20349 10421 20361 10455
rect 20395 10452 20407 10455
rect 20622 10452 20628 10464
rect 20395 10424 20628 10452
rect 20395 10421 20407 10424
rect 20349 10415 20407 10421
rect 20622 10412 20628 10424
rect 20680 10412 20686 10464
rect 1104 10362 21896 10384
rect 1104 10310 3549 10362
rect 3601 10310 3613 10362
rect 3665 10310 3677 10362
rect 3729 10310 3741 10362
rect 3793 10310 3805 10362
rect 3857 10310 8747 10362
rect 8799 10310 8811 10362
rect 8863 10310 8875 10362
rect 8927 10310 8939 10362
rect 8991 10310 9003 10362
rect 9055 10310 13945 10362
rect 13997 10310 14009 10362
rect 14061 10310 14073 10362
rect 14125 10310 14137 10362
rect 14189 10310 14201 10362
rect 14253 10310 19143 10362
rect 19195 10310 19207 10362
rect 19259 10310 19271 10362
rect 19323 10310 19335 10362
rect 19387 10310 19399 10362
rect 19451 10310 21896 10362
rect 1104 10288 21896 10310
rect 2314 10248 2320 10260
rect 2275 10220 2320 10248
rect 2314 10208 2320 10220
rect 2372 10208 2378 10260
rect 2682 10208 2688 10260
rect 2740 10248 2746 10260
rect 2777 10251 2835 10257
rect 2777 10248 2789 10251
rect 2740 10220 2789 10248
rect 2740 10208 2746 10220
rect 2777 10217 2789 10220
rect 2823 10217 2835 10251
rect 2777 10211 2835 10217
rect 3878 10208 3884 10260
rect 3936 10248 3942 10260
rect 3973 10251 4031 10257
rect 3973 10248 3985 10251
rect 3936 10220 3985 10248
rect 3936 10208 3942 10220
rect 3973 10217 3985 10220
rect 4019 10217 4031 10251
rect 3973 10211 4031 10217
rect 5166 10208 5172 10260
rect 5224 10248 5230 10260
rect 10226 10248 10232 10260
rect 5224 10220 10232 10248
rect 5224 10208 5230 10220
rect 10226 10208 10232 10220
rect 10284 10208 10290 10260
rect 10321 10251 10379 10257
rect 10321 10217 10333 10251
rect 10367 10248 10379 10251
rect 17218 10248 17224 10260
rect 10367 10220 17224 10248
rect 10367 10217 10379 10220
rect 10321 10211 10379 10217
rect 17218 10208 17224 10220
rect 17276 10208 17282 10260
rect 17402 10248 17408 10260
rect 17363 10220 17408 10248
rect 17402 10208 17408 10220
rect 17460 10208 17466 10260
rect 18322 10248 18328 10260
rect 18283 10220 18328 10248
rect 18322 10208 18328 10220
rect 18380 10208 18386 10260
rect 19150 10248 19156 10260
rect 18800 10220 19156 10248
rect 1673 10183 1731 10189
rect 1673 10149 1685 10183
rect 1719 10180 1731 10183
rect 2222 10180 2228 10192
rect 1719 10152 2228 10180
rect 1719 10149 1731 10152
rect 1673 10143 1731 10149
rect 2222 10140 2228 10152
rect 2280 10140 2286 10192
rect 4154 10140 4160 10192
rect 4212 10180 4218 10192
rect 5718 10180 5724 10192
rect 4212 10152 5724 10180
rect 4212 10140 4218 10152
rect 5718 10140 5724 10152
rect 5776 10140 5782 10192
rect 13078 10180 13084 10192
rect 13039 10152 13084 10180
rect 13078 10140 13084 10152
rect 13136 10140 13142 10192
rect 18233 10183 18291 10189
rect 18233 10149 18245 10183
rect 18279 10180 18291 10183
rect 18800 10180 18828 10220
rect 19150 10208 19156 10220
rect 19208 10208 19214 10260
rect 19794 10248 19800 10260
rect 19260 10220 19800 10248
rect 18279 10152 18828 10180
rect 18279 10149 18291 10152
rect 18233 10143 18291 10149
rect 2038 10112 2044 10124
rect 1999 10084 2044 10112
rect 2038 10072 2044 10084
rect 2096 10072 2102 10124
rect 3050 10072 3056 10124
rect 3108 10112 3114 10124
rect 3326 10112 3332 10124
rect 3108 10084 3332 10112
rect 3108 10072 3114 10084
rect 3326 10072 3332 10084
rect 3384 10072 3390 10124
rect 4617 10115 4675 10121
rect 4617 10081 4629 10115
rect 4663 10112 4675 10115
rect 4798 10112 4804 10124
rect 4663 10084 4804 10112
rect 4663 10081 4675 10084
rect 4617 10075 4675 10081
rect 4798 10072 4804 10084
rect 4856 10112 4862 10124
rect 9769 10115 9827 10121
rect 4856 10084 5396 10112
rect 4856 10072 4862 10084
rect 1486 10044 1492 10056
rect 1447 10016 1492 10044
rect 1486 10004 1492 10016
rect 1544 10004 1550 10056
rect 2130 10044 2136 10056
rect 2091 10016 2136 10044
rect 2130 10004 2136 10016
rect 2188 10044 2194 10056
rect 2409 10047 2467 10053
rect 2409 10044 2421 10047
rect 2188 10016 2421 10044
rect 2188 10004 2194 10016
rect 2409 10013 2421 10016
rect 2455 10013 2467 10047
rect 3145 10047 3203 10053
rect 3145 10044 3157 10047
rect 2409 10007 2467 10013
rect 2746 10016 3157 10044
rect 1854 9976 1860 9988
rect 1815 9948 1860 9976
rect 1854 9936 1860 9948
rect 1912 9976 1918 9988
rect 2593 9979 2651 9985
rect 2593 9976 2605 9979
rect 1912 9948 2605 9976
rect 1912 9936 1918 9948
rect 2593 9945 2605 9948
rect 2639 9945 2651 9979
rect 2593 9939 2651 9945
rect 1946 9868 1952 9920
rect 2004 9908 2010 9920
rect 2746 9908 2774 10016
rect 3145 10013 3157 10016
rect 3191 10044 3203 10047
rect 3970 10044 3976 10056
rect 3191 10016 3976 10044
rect 3191 10013 3203 10016
rect 3145 10007 3203 10013
rect 3970 10004 3976 10016
rect 4028 10004 4034 10056
rect 4430 10044 4436 10056
rect 4343 10016 4436 10044
rect 4430 10004 4436 10016
rect 4488 10044 4494 10056
rect 4893 10047 4951 10053
rect 4893 10044 4905 10047
rect 4488 10016 4905 10044
rect 4488 10004 4494 10016
rect 4893 10013 4905 10016
rect 4939 10044 4951 10047
rect 5166 10044 5172 10056
rect 4939 10016 5172 10044
rect 4939 10013 4951 10016
rect 4893 10007 4951 10013
rect 5166 10004 5172 10016
rect 5224 10004 5230 10056
rect 3237 9979 3295 9985
rect 3237 9945 3249 9979
rect 3283 9976 3295 9979
rect 4614 9976 4620 9988
rect 3283 9948 4620 9976
rect 3283 9945 3295 9948
rect 3237 9939 3295 9945
rect 4614 9936 4620 9948
rect 4672 9936 4678 9988
rect 5368 9976 5396 10084
rect 9769 10081 9781 10115
rect 9815 10081 9827 10115
rect 15654 10112 15660 10124
rect 15615 10084 15660 10112
rect 9769 10075 9827 10081
rect 5445 10047 5503 10053
rect 5445 10013 5457 10047
rect 5491 10044 5503 10047
rect 5629 10047 5687 10053
rect 5629 10044 5641 10047
rect 5491 10016 5641 10044
rect 5491 10013 5503 10016
rect 5445 10007 5503 10013
rect 5629 10013 5641 10016
rect 5675 10044 5687 10047
rect 6546 10044 6552 10056
rect 5675 10016 6552 10044
rect 5675 10013 5687 10016
rect 5629 10007 5687 10013
rect 6546 10004 6552 10016
rect 6604 10044 6610 10056
rect 7101 10047 7159 10053
rect 7101 10044 7113 10047
rect 6604 10016 7113 10044
rect 6604 10004 6610 10016
rect 7101 10013 7113 10016
rect 7147 10013 7159 10047
rect 7101 10007 7159 10013
rect 6856 9979 6914 9985
rect 6856 9976 6868 9979
rect 5368 9948 6868 9976
rect 6856 9945 6868 9948
rect 6902 9976 6914 9979
rect 8018 9976 8024 9988
rect 6902 9948 8024 9976
rect 6902 9945 6914 9948
rect 6856 9939 6914 9945
rect 8018 9936 8024 9948
rect 8076 9936 8082 9988
rect 9784 9976 9812 10075
rect 15654 10072 15660 10084
rect 15712 10072 15718 10124
rect 16574 10112 16580 10124
rect 16535 10084 16580 10112
rect 16574 10072 16580 10084
rect 16632 10072 16638 10124
rect 16850 10112 16856 10124
rect 16811 10084 16856 10112
rect 16850 10072 16856 10084
rect 16908 10072 16914 10124
rect 17034 10072 17040 10124
rect 17092 10112 17098 10124
rect 18877 10115 18935 10121
rect 18877 10112 18889 10115
rect 17092 10084 18889 10112
rect 17092 10072 17098 10084
rect 18877 10081 18889 10084
rect 18923 10112 18935 10115
rect 19260 10112 19288 10220
rect 19794 10208 19800 10220
rect 19852 10208 19858 10260
rect 19978 10248 19984 10260
rect 19939 10220 19984 10248
rect 19978 10208 19984 10220
rect 20036 10208 20042 10260
rect 21177 10251 21235 10257
rect 21177 10217 21189 10251
rect 21223 10248 21235 10251
rect 21266 10248 21272 10260
rect 21223 10220 21272 10248
rect 21223 10217 21235 10220
rect 21177 10211 21235 10217
rect 21266 10208 21272 10220
rect 21324 10208 21330 10260
rect 21358 10208 21364 10260
rect 21416 10248 21422 10260
rect 21416 10220 21461 10248
rect 21416 10208 21422 10220
rect 19426 10140 19432 10192
rect 19484 10180 19490 10192
rect 19484 10152 21496 10180
rect 19484 10140 19490 10152
rect 18923 10084 19288 10112
rect 19337 10115 19395 10121
rect 18923 10081 18935 10084
rect 18877 10075 18935 10081
rect 19337 10081 19349 10115
rect 19383 10081 19395 10115
rect 20622 10112 20628 10124
rect 20583 10084 20628 10112
rect 19337 10075 19395 10081
rect 11609 10047 11667 10053
rect 11609 10013 11621 10047
rect 11655 10044 11667 10047
rect 11701 10047 11759 10053
rect 11701 10044 11713 10047
rect 11655 10016 11713 10044
rect 11655 10013 11667 10016
rect 11609 10007 11667 10013
rect 11701 10013 11713 10016
rect 11747 10044 11759 10047
rect 12250 10044 12256 10056
rect 11747 10016 12256 10044
rect 11747 10013 11759 10016
rect 11701 10007 11759 10013
rect 12250 10004 12256 10016
rect 12308 10004 12314 10056
rect 14185 10047 14243 10053
rect 14185 10013 14197 10047
rect 14231 10044 14243 10047
rect 15672 10044 15700 10072
rect 14231 10016 15700 10044
rect 16592 10044 16620 10072
rect 16945 10047 17003 10053
rect 16945 10044 16957 10047
rect 16592 10016 16957 10044
rect 14231 10013 14243 10016
rect 14185 10007 14243 10013
rect 16945 10013 16957 10016
rect 16991 10013 17003 10047
rect 16945 10007 17003 10013
rect 18506 10004 18512 10056
rect 18564 10044 18570 10056
rect 18693 10047 18751 10053
rect 18693 10044 18705 10047
rect 18564 10016 18705 10044
rect 18564 10004 18570 10016
rect 18693 10013 18705 10016
rect 18739 10044 18751 10047
rect 18782 10044 18788 10056
rect 18739 10016 18788 10044
rect 18739 10013 18751 10016
rect 18693 10007 18751 10013
rect 18782 10004 18788 10016
rect 18840 10004 18846 10056
rect 11974 9985 11980 9988
rect 11946 9979 11980 9985
rect 11946 9976 11958 9979
rect 9784 9948 11958 9976
rect 11946 9945 11958 9948
rect 12032 9976 12038 9988
rect 12032 9948 12094 9976
rect 11946 9939 11980 9945
rect 11974 9936 11980 9939
rect 12032 9936 12038 9948
rect 12158 9936 12164 9988
rect 12216 9976 12222 9988
rect 15378 9976 15384 9988
rect 15436 9985 15442 9988
rect 12216 9948 14320 9976
rect 15348 9948 15384 9976
rect 12216 9936 12222 9948
rect 4338 9908 4344 9920
rect 2004 9880 2774 9908
rect 4299 9880 4344 9908
rect 2004 9868 2010 9880
rect 4338 9868 4344 9880
rect 4396 9868 4402 9920
rect 4706 9868 4712 9920
rect 4764 9908 4770 9920
rect 6362 9908 6368 9920
rect 4764 9880 6368 9908
rect 4764 9868 4770 9880
rect 6362 9868 6368 9880
rect 6420 9908 6426 9920
rect 6730 9908 6736 9920
rect 6420 9880 6736 9908
rect 6420 9868 6426 9880
rect 6730 9868 6736 9880
rect 6788 9868 6794 9920
rect 9766 9868 9772 9920
rect 9824 9908 9830 9920
rect 9861 9911 9919 9917
rect 9861 9908 9873 9911
rect 9824 9880 9873 9908
rect 9824 9868 9830 9880
rect 9861 9877 9873 9880
rect 9907 9877 9919 9911
rect 9861 9871 9919 9877
rect 9950 9868 9956 9920
rect 10008 9908 10014 9920
rect 14292 9917 14320 9948
rect 15378 9936 15384 9948
rect 15436 9939 15448 9985
rect 19352 9976 19380 10075
rect 20622 10072 20628 10084
rect 20680 10072 20686 10124
rect 20717 10115 20775 10121
rect 20717 10081 20729 10115
rect 20763 10081 20775 10115
rect 20717 10075 20775 10081
rect 19518 10044 19524 10056
rect 19479 10016 19524 10044
rect 19518 10004 19524 10016
rect 19576 10004 19582 10056
rect 19702 10004 19708 10056
rect 19760 10044 19766 10056
rect 20732 10044 20760 10075
rect 21468 10056 21496 10152
rect 19760 10016 20760 10044
rect 20993 10047 21051 10053
rect 19760 10004 19766 10016
rect 20993 10013 21005 10047
rect 21039 10013 21051 10047
rect 21450 10044 21456 10056
rect 21363 10016 21456 10044
rect 20993 10007 21051 10013
rect 20438 9976 20444 9988
rect 15488 9948 19380 9976
rect 19444 9948 20444 9976
rect 15436 9936 15442 9939
rect 14277 9911 14335 9917
rect 10008 9880 10053 9908
rect 10008 9868 10014 9880
rect 14277 9877 14289 9911
rect 14323 9908 14335 9911
rect 15488 9908 15516 9948
rect 14323 9880 15516 9908
rect 14323 9877 14335 9880
rect 14277 9871 14335 9877
rect 16758 9868 16764 9920
rect 16816 9908 16822 9920
rect 17037 9911 17095 9917
rect 17037 9908 17049 9911
rect 16816 9880 17049 9908
rect 16816 9868 16822 9880
rect 17037 9877 17049 9880
rect 17083 9908 17095 9911
rect 17218 9908 17224 9920
rect 17083 9880 17224 9908
rect 17083 9877 17095 9880
rect 17037 9871 17095 9877
rect 17218 9868 17224 9880
rect 17276 9868 17282 9920
rect 17954 9868 17960 9920
rect 18012 9908 18018 9920
rect 18785 9911 18843 9917
rect 18785 9908 18797 9911
rect 18012 9880 18797 9908
rect 18012 9868 18018 9880
rect 18785 9877 18797 9880
rect 18831 9908 18843 9911
rect 19444 9908 19472 9948
rect 20438 9936 20444 9948
rect 20496 9936 20502 9988
rect 20622 9936 20628 9988
rect 20680 9976 20686 9988
rect 21008 9976 21036 10007
rect 21450 10004 21456 10016
rect 21508 10004 21514 10056
rect 20680 9948 21036 9976
rect 20680 9936 20686 9948
rect 18831 9880 19472 9908
rect 18831 9877 18843 9880
rect 18785 9871 18843 9877
rect 19610 9868 19616 9920
rect 19668 9908 19674 9920
rect 20162 9908 20168 9920
rect 19668 9880 19713 9908
rect 20123 9880 20168 9908
rect 19668 9868 19674 9880
rect 20162 9868 20168 9880
rect 20220 9868 20226 9920
rect 20530 9908 20536 9920
rect 20491 9880 20536 9908
rect 20530 9868 20536 9880
rect 20588 9868 20594 9920
rect 1104 9818 22056 9840
rect 1104 9766 6148 9818
rect 6200 9766 6212 9818
rect 6264 9766 6276 9818
rect 6328 9766 6340 9818
rect 6392 9766 6404 9818
rect 6456 9766 11346 9818
rect 11398 9766 11410 9818
rect 11462 9766 11474 9818
rect 11526 9766 11538 9818
rect 11590 9766 11602 9818
rect 11654 9766 16544 9818
rect 16596 9766 16608 9818
rect 16660 9766 16672 9818
rect 16724 9766 16736 9818
rect 16788 9766 16800 9818
rect 16852 9766 21742 9818
rect 21794 9766 21806 9818
rect 21858 9766 21870 9818
rect 21922 9766 21934 9818
rect 21986 9766 21998 9818
rect 22050 9766 22056 9818
rect 1104 9744 22056 9766
rect 1486 9664 1492 9716
rect 1544 9704 1550 9716
rect 2317 9707 2375 9713
rect 2317 9704 2329 9707
rect 1544 9676 2329 9704
rect 1544 9664 1550 9676
rect 2317 9673 2329 9676
rect 2363 9673 2375 9707
rect 2317 9667 2375 9673
rect 3237 9707 3295 9713
rect 3237 9673 3249 9707
rect 3283 9704 3295 9707
rect 3418 9704 3424 9716
rect 3283 9676 3424 9704
rect 3283 9673 3295 9676
rect 3237 9667 3295 9673
rect 3418 9664 3424 9676
rect 3476 9664 3482 9716
rect 4706 9704 4712 9716
rect 3988 9676 4712 9704
rect 2958 9596 2964 9648
rect 3016 9636 3022 9648
rect 3988 9636 4016 9676
rect 3016 9608 4016 9636
rect 4065 9639 4123 9645
rect 3016 9596 3022 9608
rect 4065 9605 4077 9639
rect 4111 9636 4123 9639
rect 4246 9636 4252 9648
rect 4111 9608 4252 9636
rect 4111 9605 4123 9608
rect 4065 9599 4123 9605
rect 4246 9596 4252 9608
rect 4304 9596 4310 9648
rect 2777 9571 2835 9577
rect 2777 9537 2789 9571
rect 2823 9568 2835 9571
rect 3970 9568 3976 9580
rect 2823 9540 3976 9568
rect 2823 9537 2835 9540
rect 2777 9531 2835 9537
rect 3970 9528 3976 9540
rect 4028 9528 4034 9580
rect 1394 9500 1400 9512
rect 1355 9472 1400 9500
rect 1394 9460 1400 9472
rect 1452 9460 1458 9512
rect 1673 9503 1731 9509
rect 1673 9469 1685 9503
rect 1719 9469 1731 9503
rect 3326 9500 3332 9512
rect 3287 9472 3332 9500
rect 1673 9463 1731 9469
rect 1688 9432 1716 9463
rect 3326 9460 3332 9472
rect 3384 9460 3390 9512
rect 3418 9460 3424 9512
rect 3476 9500 3482 9512
rect 3476 9472 3521 9500
rect 3476 9460 3482 9472
rect 4062 9460 4068 9512
rect 4120 9500 4126 9512
rect 4356 9509 4384 9676
rect 4706 9664 4712 9676
rect 4764 9664 4770 9716
rect 4801 9707 4859 9713
rect 4801 9673 4813 9707
rect 4847 9704 4859 9707
rect 5074 9704 5080 9716
rect 4847 9676 5080 9704
rect 4847 9673 4859 9676
rect 4801 9667 4859 9673
rect 5074 9664 5080 9676
rect 5132 9664 5138 9716
rect 8018 9664 8024 9716
rect 8076 9704 8082 9716
rect 13630 9704 13636 9716
rect 8076 9676 13636 9704
rect 8076 9664 8082 9676
rect 13630 9664 13636 9676
rect 13688 9664 13694 9716
rect 14476 9676 14688 9704
rect 10134 9645 10140 9648
rect 10128 9636 10140 9645
rect 5184 9608 8616 9636
rect 10095 9608 10140 9636
rect 4157 9503 4215 9509
rect 4157 9500 4169 9503
rect 4120 9472 4169 9500
rect 4120 9460 4126 9472
rect 4157 9469 4169 9472
rect 4203 9469 4215 9503
rect 4157 9463 4215 9469
rect 4341 9503 4399 9509
rect 4341 9469 4353 9503
rect 4387 9469 4399 9503
rect 4341 9463 4399 9469
rect 5184 9432 5212 9608
rect 5902 9528 5908 9580
rect 5960 9577 5966 9580
rect 5960 9568 5972 9577
rect 5960 9540 6005 9568
rect 5960 9531 5972 9540
rect 5960 9528 5966 9531
rect 6730 9528 6736 9580
rect 6788 9568 6794 9580
rect 7478 9571 7536 9577
rect 7478 9568 7490 9571
rect 6788 9540 7490 9568
rect 6788 9528 6794 9540
rect 7478 9537 7490 9540
rect 7524 9537 7536 9571
rect 7478 9531 7536 9537
rect 7745 9571 7803 9577
rect 7745 9537 7757 9571
rect 7791 9568 7803 9571
rect 7926 9568 7932 9580
rect 7791 9540 7932 9568
rect 7791 9537 7803 9540
rect 7745 9531 7803 9537
rect 7926 9528 7932 9540
rect 7984 9568 7990 9580
rect 8205 9571 8263 9577
rect 8205 9568 8217 9571
rect 7984 9540 8217 9568
rect 7984 9528 7990 9540
rect 8205 9537 8217 9540
rect 8251 9537 8263 9571
rect 8461 9571 8519 9577
rect 8461 9568 8473 9571
rect 8205 9531 8263 9537
rect 8312 9540 8473 9568
rect 6181 9503 6239 9509
rect 6181 9469 6193 9503
rect 6227 9500 6239 9503
rect 6362 9500 6368 9512
rect 6227 9472 6368 9500
rect 6227 9469 6239 9472
rect 6181 9463 6239 9469
rect 6362 9460 6368 9472
rect 6420 9460 6426 9512
rect 8312 9500 8340 9540
rect 8461 9537 8473 9540
rect 8507 9537 8519 9571
rect 8588 9568 8616 9608
rect 10128 9599 10140 9608
rect 10134 9596 10140 9599
rect 10192 9596 10198 9648
rect 12158 9596 12164 9648
rect 12216 9636 12222 9648
rect 14476 9636 14504 9676
rect 12216 9608 14504 9636
rect 12216 9596 12222 9608
rect 8588 9540 10916 9568
rect 8461 9531 8519 9537
rect 9766 9500 9772 9512
rect 7760 9472 8340 9500
rect 9324 9472 9772 9500
rect 7760 9444 7788 9472
rect 1688 9404 5212 9432
rect 7742 9392 7748 9444
rect 7800 9392 7806 9444
rect 2590 9364 2596 9376
rect 2551 9336 2596 9364
rect 2590 9324 2596 9336
rect 2648 9324 2654 9376
rect 2866 9364 2872 9376
rect 2827 9336 2872 9364
rect 2866 9324 2872 9336
rect 2924 9324 2930 9376
rect 3234 9324 3240 9376
rect 3292 9364 3298 9376
rect 3697 9367 3755 9373
rect 3697 9364 3709 9367
rect 3292 9336 3709 9364
rect 3292 9324 3298 9336
rect 3697 9333 3709 9336
rect 3743 9333 3755 9367
rect 3697 9327 3755 9333
rect 5994 9324 6000 9376
rect 6052 9364 6058 9376
rect 6365 9367 6423 9373
rect 6365 9364 6377 9367
rect 6052 9336 6377 9364
rect 6052 9324 6058 9336
rect 6365 9333 6377 9336
rect 6411 9333 6423 9367
rect 7926 9364 7932 9376
rect 7887 9336 7932 9364
rect 6365 9327 6423 9333
rect 7926 9324 7932 9336
rect 7984 9364 7990 9376
rect 8021 9367 8079 9373
rect 8021 9364 8033 9367
rect 7984 9336 8033 9364
rect 7984 9324 7990 9336
rect 8021 9333 8033 9336
rect 8067 9333 8079 9367
rect 8021 9327 8079 9333
rect 8110 9324 8116 9376
rect 8168 9364 8174 9376
rect 9324 9364 9352 9472
rect 9766 9460 9772 9472
rect 9824 9460 9830 9512
rect 9861 9503 9919 9509
rect 9861 9469 9873 9503
rect 9907 9469 9919 9503
rect 9861 9463 9919 9469
rect 9490 9392 9496 9444
rect 9548 9432 9554 9444
rect 9876 9432 9904 9463
rect 9548 9404 9904 9432
rect 10888 9432 10916 9540
rect 14550 9528 14556 9580
rect 14608 9568 14614 9580
rect 14660 9568 14688 9676
rect 17126 9674 17132 9716
rect 17052 9664 17132 9674
rect 17184 9664 17190 9716
rect 17405 9707 17463 9713
rect 17405 9673 17417 9707
rect 17451 9704 17463 9707
rect 17494 9704 17500 9716
rect 17451 9676 17500 9704
rect 17451 9673 17463 9676
rect 17405 9667 17463 9673
rect 17494 9664 17500 9676
rect 17552 9664 17558 9716
rect 19429 9707 19487 9713
rect 19429 9673 19441 9707
rect 19475 9704 19487 9707
rect 19518 9704 19524 9716
rect 19475 9676 19524 9704
rect 19475 9673 19487 9676
rect 19429 9667 19487 9673
rect 19518 9664 19524 9676
rect 19576 9664 19582 9716
rect 19889 9707 19947 9713
rect 19889 9673 19901 9707
rect 19935 9704 19947 9707
rect 20162 9704 20168 9716
rect 19935 9676 20168 9704
rect 19935 9673 19947 9676
rect 19889 9667 19947 9673
rect 20162 9664 20168 9676
rect 20220 9664 20226 9716
rect 20530 9664 20536 9716
rect 20588 9704 20594 9716
rect 20625 9707 20683 9713
rect 20625 9704 20637 9707
rect 20588 9676 20637 9704
rect 20588 9664 20594 9676
rect 20625 9673 20637 9676
rect 20671 9673 20683 9707
rect 20625 9667 20683 9673
rect 17052 9646 17172 9664
rect 14608 9540 14688 9568
rect 14717 9571 14775 9577
rect 14608 9528 14614 9540
rect 14717 9537 14729 9571
rect 14763 9568 14775 9571
rect 15010 9568 15016 9580
rect 14763 9540 15016 9568
rect 14763 9537 14775 9540
rect 14717 9531 14775 9537
rect 15010 9528 15016 9540
rect 15068 9528 15074 9580
rect 14461 9503 14519 9509
rect 14461 9500 14473 9503
rect 14292 9472 14473 9500
rect 10888 9404 12434 9432
rect 9548 9392 9554 9404
rect 9582 9364 9588 9376
rect 8168 9336 9352 9364
rect 9543 9336 9588 9364
rect 8168 9324 8174 9336
rect 9582 9324 9588 9336
rect 9640 9324 9646 9376
rect 9769 9367 9827 9373
rect 9769 9333 9781 9367
rect 9815 9364 9827 9367
rect 9876 9364 9904 9404
rect 10502 9364 10508 9376
rect 9815 9336 10508 9364
rect 9815 9333 9827 9336
rect 9769 9327 9827 9333
rect 10502 9324 10508 9336
rect 10560 9324 10566 9376
rect 11241 9367 11299 9373
rect 11241 9333 11253 9367
rect 11287 9364 11299 9367
rect 11698 9364 11704 9376
rect 11287 9336 11704 9364
rect 11287 9333 11299 9336
rect 11241 9327 11299 9333
rect 11698 9324 11704 9336
rect 11756 9324 11762 9376
rect 12406 9364 12434 9404
rect 13538 9364 13544 9376
rect 12406 9336 13544 9364
rect 13538 9324 13544 9336
rect 13596 9324 13602 9376
rect 13814 9324 13820 9376
rect 13872 9364 13878 9376
rect 14292 9373 14320 9472
rect 14461 9469 14473 9472
rect 14507 9469 14519 9503
rect 14461 9463 14519 9469
rect 15746 9460 15752 9512
rect 15804 9500 15810 9512
rect 17052 9500 17080 9646
rect 18138 9636 18144 9648
rect 18099 9608 18144 9636
rect 18138 9596 18144 9608
rect 18196 9596 18202 9648
rect 18892 9608 20116 9636
rect 18233 9571 18291 9577
rect 18233 9537 18245 9571
rect 18279 9537 18291 9571
rect 18233 9531 18291 9537
rect 17129 9503 17187 9509
rect 17129 9500 17141 9503
rect 15804 9472 16988 9500
rect 17052 9472 17141 9500
rect 15804 9460 15810 9472
rect 15933 9435 15991 9441
rect 15933 9432 15945 9435
rect 15396 9404 15945 9432
rect 14277 9367 14335 9373
rect 14277 9364 14289 9367
rect 13872 9336 14289 9364
rect 13872 9324 13878 9336
rect 14277 9333 14289 9336
rect 14323 9364 14335 9367
rect 15396 9364 15424 9404
rect 15933 9401 15945 9404
rect 15979 9432 15991 9435
rect 16390 9432 16396 9444
rect 15979 9404 16396 9432
rect 15979 9401 15991 9404
rect 15933 9395 15991 9401
rect 16390 9392 16396 9404
rect 16448 9392 16454 9444
rect 16960 9441 16988 9472
rect 17129 9469 17141 9472
rect 17175 9469 17187 9503
rect 17129 9463 17187 9469
rect 17313 9503 17371 9509
rect 17313 9469 17325 9503
rect 17359 9469 17371 9503
rect 17313 9463 17371 9469
rect 18049 9503 18107 9509
rect 18049 9469 18061 9503
rect 18095 9500 18107 9503
rect 18138 9500 18144 9512
rect 18095 9472 18144 9500
rect 18095 9469 18107 9472
rect 18049 9463 18107 9469
rect 16945 9435 17003 9441
rect 16945 9401 16957 9435
rect 16991 9432 17003 9435
rect 17328 9432 17356 9463
rect 18138 9460 18144 9472
rect 18196 9460 18202 9512
rect 16991 9404 17356 9432
rect 17773 9435 17831 9441
rect 16991 9401 17003 9404
rect 16945 9395 17003 9401
rect 17773 9401 17785 9435
rect 17819 9432 17831 9435
rect 18248 9432 18276 9531
rect 18892 9509 18920 9608
rect 19061 9571 19119 9577
rect 19061 9537 19073 9571
rect 19107 9537 19119 9571
rect 19061 9531 19119 9537
rect 18877 9503 18935 9509
rect 18877 9500 18889 9503
rect 17819 9404 18276 9432
rect 18340 9472 18889 9500
rect 17819 9401 17831 9404
rect 17773 9395 17831 9401
rect 14323 9336 15424 9364
rect 14323 9333 14335 9336
rect 14277 9327 14335 9333
rect 15470 9324 15476 9376
rect 15528 9364 15534 9376
rect 15841 9367 15899 9373
rect 15841 9364 15853 9367
rect 15528 9336 15853 9364
rect 15528 9324 15534 9336
rect 15841 9333 15853 9336
rect 15887 9364 15899 9367
rect 18340 9364 18368 9472
rect 18877 9469 18889 9472
rect 18923 9469 18935 9503
rect 18877 9463 18935 9469
rect 18969 9503 19027 9509
rect 18969 9469 18981 9503
rect 19015 9469 19027 9503
rect 18969 9463 19027 9469
rect 18601 9435 18659 9441
rect 18601 9401 18613 9435
rect 18647 9432 18659 9435
rect 18984 9432 19012 9463
rect 18647 9404 19012 9432
rect 18647 9401 18659 9404
rect 18601 9395 18659 9401
rect 15887 9336 18368 9364
rect 15887 9333 15899 9336
rect 15841 9327 15899 9333
rect 18506 9324 18512 9376
rect 18564 9364 18570 9376
rect 19076 9364 19104 9531
rect 20088 9509 20116 9608
rect 21269 9571 21327 9577
rect 21269 9537 21281 9571
rect 21315 9568 21327 9571
rect 21634 9568 21640 9580
rect 21315 9540 21640 9568
rect 21315 9537 21327 9540
rect 21269 9531 21327 9537
rect 21634 9528 21640 9540
rect 21692 9528 21698 9580
rect 19981 9503 20039 9509
rect 19981 9469 19993 9503
rect 20027 9469 20039 9503
rect 19981 9463 20039 9469
rect 20073 9503 20131 9509
rect 20073 9469 20085 9503
rect 20119 9469 20131 9503
rect 21542 9500 21548 9512
rect 21503 9472 21548 9500
rect 20073 9463 20131 9469
rect 19521 9435 19579 9441
rect 19521 9401 19533 9435
rect 19567 9432 19579 9435
rect 19610 9432 19616 9444
rect 19567 9404 19616 9432
rect 19567 9401 19579 9404
rect 19521 9395 19579 9401
rect 19610 9392 19616 9404
rect 19668 9392 19674 9444
rect 19996 9432 20024 9463
rect 21542 9460 21548 9472
rect 21600 9460 21606 9512
rect 20806 9432 20812 9444
rect 19996 9404 20812 9432
rect 20806 9392 20812 9404
rect 20864 9392 20870 9444
rect 18564 9336 19104 9364
rect 18564 9324 18570 9336
rect 1104 9274 21896 9296
rect 1104 9222 3549 9274
rect 3601 9222 3613 9274
rect 3665 9222 3677 9274
rect 3729 9222 3741 9274
rect 3793 9222 3805 9274
rect 3857 9222 8747 9274
rect 8799 9222 8811 9274
rect 8863 9222 8875 9274
rect 8927 9222 8939 9274
rect 8991 9222 9003 9274
rect 9055 9222 13945 9274
rect 13997 9222 14009 9274
rect 14061 9222 14073 9274
rect 14125 9222 14137 9274
rect 14189 9222 14201 9274
rect 14253 9222 19143 9274
rect 19195 9222 19207 9274
rect 19259 9222 19271 9274
rect 19323 9222 19335 9274
rect 19387 9222 19399 9274
rect 19451 9222 21896 9274
rect 1104 9200 21896 9222
rect 2409 9163 2467 9169
rect 2409 9129 2421 9163
rect 2455 9160 2467 9163
rect 2498 9160 2504 9172
rect 2455 9132 2504 9160
rect 2455 9129 2467 9132
rect 2409 9123 2467 9129
rect 2498 9120 2504 9132
rect 2556 9120 2562 9172
rect 6273 9163 6331 9169
rect 2746 9132 5856 9160
rect 2746 9092 2774 9132
rect 1964 9064 2774 9092
rect 5828 9092 5856 9132
rect 6273 9129 6285 9163
rect 6319 9160 6331 9163
rect 7374 9160 7380 9172
rect 6319 9132 7380 9160
rect 6319 9129 6331 9132
rect 6273 9123 6331 9129
rect 7374 9120 7380 9132
rect 7432 9120 7438 9172
rect 12158 9160 12164 9172
rect 7576 9132 12164 9160
rect 5828 9064 6408 9092
rect 1964 9033 1992 9064
rect 1949 9027 2007 9033
rect 1949 8993 1961 9027
rect 1995 8993 2007 9027
rect 2866 9024 2872 9036
rect 2827 8996 2872 9024
rect 1949 8987 2007 8993
rect 2866 8984 2872 8996
rect 2924 8984 2930 9036
rect 3053 9027 3111 9033
rect 3053 8993 3065 9027
rect 3099 9024 3111 9027
rect 6380 9024 6408 9064
rect 3099 8996 4844 9024
rect 6380 8996 6500 9024
rect 3099 8993 3111 8996
rect 3053 8987 3111 8993
rect 2222 8956 2228 8968
rect 2183 8928 2228 8956
rect 2222 8916 2228 8928
rect 2280 8956 2286 8968
rect 3237 8959 3295 8965
rect 3237 8956 3249 8959
rect 2280 8928 3249 8956
rect 2280 8916 2286 8928
rect 3237 8925 3249 8928
rect 3283 8925 3295 8959
rect 3237 8919 3295 8925
rect 2774 8780 2780 8832
rect 2832 8820 2838 8832
rect 4816 8820 4844 8996
rect 4893 8959 4951 8965
rect 4893 8925 4905 8959
rect 4939 8956 4951 8959
rect 6362 8956 6368 8968
rect 4939 8928 6368 8956
rect 4939 8925 4951 8928
rect 4893 8919 4951 8925
rect 6362 8916 6368 8928
rect 6420 8916 6426 8968
rect 6472 8956 6500 8996
rect 7576 8956 7604 9132
rect 12158 9120 12164 9132
rect 12216 9120 12222 9172
rect 13906 9160 13912 9172
rect 12544 9132 13912 9160
rect 7834 9092 7840 9104
rect 7795 9064 7840 9092
rect 7834 9052 7840 9064
rect 7892 9052 7898 9104
rect 7926 9052 7932 9104
rect 7984 9092 7990 9104
rect 8754 9092 8760 9104
rect 7984 9064 8760 9092
rect 7984 9052 7990 9064
rect 8754 9052 8760 9064
rect 8812 9092 8818 9104
rect 9033 9095 9091 9101
rect 9033 9092 9045 9095
rect 8812 9064 9045 9092
rect 8812 9052 8818 9064
rect 9033 9061 9045 9064
rect 9079 9092 9091 9095
rect 9490 9092 9496 9104
rect 9079 9064 9496 9092
rect 9079 9061 9091 9064
rect 9033 9055 9091 9061
rect 9490 9052 9496 9064
rect 9548 9052 9554 9104
rect 11974 9052 11980 9104
rect 12032 9092 12038 9104
rect 12544 9092 12572 9132
rect 13906 9120 13912 9132
rect 13964 9120 13970 9172
rect 15010 9120 15016 9172
rect 15068 9160 15074 9172
rect 15473 9163 15531 9169
rect 15473 9160 15485 9163
rect 15068 9132 15485 9160
rect 15068 9120 15074 9132
rect 15473 9129 15485 9132
rect 15519 9160 15531 9163
rect 18138 9160 18144 9172
rect 15519 9132 18144 9160
rect 15519 9129 15531 9132
rect 15473 9123 15531 9129
rect 18138 9120 18144 9132
rect 18196 9120 18202 9172
rect 18524 9132 19104 9160
rect 12032 9064 12572 9092
rect 16945 9095 17003 9101
rect 12032 9052 12038 9064
rect 16945 9061 16957 9095
rect 16991 9092 17003 9095
rect 17678 9092 17684 9104
rect 16991 9064 17684 9092
rect 16991 9061 17003 9064
rect 16945 9055 17003 9061
rect 17678 9052 17684 9064
rect 17736 9052 17742 9104
rect 17954 9092 17960 9104
rect 17915 9064 17960 9092
rect 17954 9052 17960 9064
rect 18012 9052 18018 9104
rect 8018 8984 8024 9036
rect 8076 9024 8082 9036
rect 18524 9033 18552 9132
rect 19076 9092 19104 9132
rect 19150 9120 19156 9172
rect 19208 9160 19214 9172
rect 19245 9163 19303 9169
rect 19245 9160 19257 9163
rect 19208 9132 19257 9160
rect 19208 9120 19214 9132
rect 19245 9129 19257 9132
rect 19291 9129 19303 9163
rect 19245 9123 19303 9129
rect 19334 9120 19340 9172
rect 19392 9160 19398 9172
rect 19978 9160 19984 9172
rect 19392 9132 19984 9160
rect 19392 9120 19398 9132
rect 19978 9120 19984 9132
rect 20036 9120 20042 9172
rect 20622 9160 20628 9172
rect 20583 9132 20628 9160
rect 20622 9120 20628 9132
rect 20680 9120 20686 9172
rect 20162 9092 20168 9104
rect 19076 9064 20168 9092
rect 20162 9052 20168 9064
rect 20220 9092 20226 9104
rect 20349 9095 20407 9101
rect 20349 9092 20361 9095
rect 20220 9064 20361 9092
rect 20220 9052 20226 9064
rect 20349 9061 20361 9064
rect 20395 9092 20407 9095
rect 20714 9092 20720 9104
rect 20395 9064 20720 9092
rect 20395 9061 20407 9064
rect 20349 9055 20407 9061
rect 20714 9052 20720 9064
rect 20772 9052 20778 9104
rect 8389 9027 8447 9033
rect 8389 9024 8401 9027
rect 8076 8996 8401 9024
rect 8076 8984 8082 8996
rect 8389 8993 8401 8996
rect 8435 8993 8447 9027
rect 17589 9027 17647 9033
rect 17589 9024 17601 9027
rect 8389 8987 8447 8993
rect 16592 8996 17601 9024
rect 8202 8956 8208 8968
rect 6472 8928 7604 8956
rect 8163 8928 8208 8956
rect 8202 8916 8208 8928
rect 8260 8916 8266 8968
rect 10238 8959 10296 8965
rect 10238 8925 10250 8959
rect 10284 8925 10296 8959
rect 10502 8956 10508 8968
rect 10463 8928 10508 8956
rect 10238 8919 10296 8925
rect 5166 8897 5172 8900
rect 5160 8888 5172 8897
rect 5127 8860 5172 8888
rect 5160 8851 5172 8860
rect 5166 8848 5172 8851
rect 5224 8848 5230 8900
rect 5718 8848 5724 8900
rect 5776 8888 5782 8900
rect 6610 8891 6668 8897
rect 6610 8888 6622 8891
rect 5776 8860 6622 8888
rect 5776 8848 5782 8860
rect 6610 8857 6622 8860
rect 6656 8857 6668 8891
rect 8846 8888 8852 8900
rect 6610 8851 6668 8857
rect 7668 8860 8852 8888
rect 7668 8820 7696 8860
rect 8846 8848 8852 8860
rect 8904 8888 8910 8900
rect 9582 8888 9588 8900
rect 8904 8860 9588 8888
rect 8904 8848 8910 8860
rect 9582 8848 9588 8860
rect 9640 8848 9646 8900
rect 10134 8848 10140 8900
rect 10192 8888 10198 8900
rect 10244 8888 10272 8919
rect 10502 8916 10508 8928
rect 10560 8956 10566 8968
rect 10597 8959 10655 8965
rect 10597 8956 10609 8959
rect 10560 8928 10609 8956
rect 10560 8916 10566 8928
rect 10597 8925 10609 8928
rect 10643 8925 10655 8959
rect 10597 8919 10655 8925
rect 10686 8916 10692 8968
rect 10744 8956 10750 8968
rect 10853 8959 10911 8965
rect 10853 8956 10865 8959
rect 10744 8928 10865 8956
rect 10744 8916 10750 8928
rect 10853 8925 10865 8928
rect 10899 8925 10911 8959
rect 13193 8959 13251 8965
rect 13193 8956 13205 8959
rect 10853 8919 10911 8925
rect 12995 8928 13205 8956
rect 12995 8888 13023 8928
rect 13193 8925 13205 8928
rect 13239 8956 13251 8959
rect 13354 8956 13360 8968
rect 13239 8928 13360 8956
rect 13239 8925 13251 8928
rect 13193 8919 13251 8925
rect 13354 8916 13360 8928
rect 13412 8916 13418 8968
rect 13449 8959 13507 8965
rect 13449 8925 13461 8959
rect 13495 8956 13507 8959
rect 14093 8959 14151 8965
rect 14093 8956 14105 8959
rect 13495 8928 14105 8956
rect 13495 8925 13507 8928
rect 13449 8919 13507 8925
rect 10192 8860 10272 8888
rect 11992 8860 13023 8888
rect 10192 8848 10198 8860
rect 2832 8792 2877 8820
rect 4816 8792 7696 8820
rect 2832 8780 2838 8792
rect 7742 8780 7748 8832
rect 7800 8820 7806 8832
rect 7800 8792 7845 8820
rect 7800 8780 7806 8792
rect 8110 8780 8116 8832
rect 8168 8820 8174 8832
rect 8297 8823 8355 8829
rect 8297 8820 8309 8823
rect 8168 8792 8309 8820
rect 8168 8780 8174 8792
rect 8297 8789 8309 8792
rect 8343 8789 8355 8823
rect 9122 8820 9128 8832
rect 9083 8792 9128 8820
rect 8297 8783 8355 8789
rect 9122 8780 9128 8792
rect 9180 8780 9186 8832
rect 11992 8829 12020 8860
rect 13832 8832 13860 8928
rect 14093 8925 14105 8928
rect 14139 8956 14151 8959
rect 15565 8959 15623 8965
rect 15565 8956 15577 8959
rect 14139 8928 15577 8956
rect 14139 8925 14151 8928
rect 14093 8919 14151 8925
rect 15565 8925 15577 8928
rect 15611 8925 15623 8959
rect 15565 8919 15623 8925
rect 15654 8916 15660 8968
rect 15712 8956 15718 8968
rect 15832 8959 15890 8965
rect 15832 8956 15844 8959
rect 15712 8928 15844 8956
rect 15712 8916 15718 8928
rect 15832 8925 15844 8928
rect 15878 8956 15890 8959
rect 16592 8956 16620 8996
rect 17589 8993 17601 8996
rect 17635 8993 17647 9027
rect 17589 8987 17647 8993
rect 18509 9027 18567 9033
rect 18509 8993 18521 9027
rect 18555 8993 18567 9027
rect 18509 8987 18567 8993
rect 19242 8984 19248 9036
rect 19300 9024 19306 9036
rect 19886 9024 19892 9036
rect 19300 8996 19748 9024
rect 19847 8996 19892 9024
rect 19300 8984 19306 8996
rect 15878 8928 16620 8956
rect 15878 8925 15890 8928
rect 15832 8919 15890 8925
rect 17402 8916 17408 8968
rect 17460 8956 17466 8968
rect 19334 8956 19340 8968
rect 17460 8928 19340 8956
rect 17460 8916 17466 8928
rect 19334 8916 19340 8928
rect 19392 8916 19398 8968
rect 14360 8891 14418 8897
rect 14360 8857 14372 8891
rect 14406 8888 14418 8891
rect 14458 8888 14464 8900
rect 14406 8860 14464 8888
rect 14406 8857 14418 8860
rect 14360 8851 14418 8857
rect 14458 8848 14464 8860
rect 14516 8848 14522 8900
rect 16942 8888 16948 8900
rect 14568 8860 16948 8888
rect 11977 8823 12035 8829
rect 11977 8789 11989 8823
rect 12023 8789 12035 8823
rect 11977 8783 12035 8789
rect 12069 8823 12127 8829
rect 12069 8789 12081 8823
rect 12115 8820 12127 8823
rect 12526 8820 12532 8832
rect 12115 8792 12532 8820
rect 12115 8789 12127 8792
rect 12069 8783 12127 8789
rect 12526 8780 12532 8792
rect 12584 8780 12590 8832
rect 13814 8820 13820 8832
rect 13775 8792 13820 8820
rect 13814 8780 13820 8792
rect 13872 8780 13878 8832
rect 13906 8780 13912 8832
rect 13964 8820 13970 8832
rect 14568 8820 14596 8860
rect 16942 8848 16948 8860
rect 17000 8848 17006 8900
rect 17494 8888 17500 8900
rect 17455 8860 17500 8888
rect 17494 8848 17500 8860
rect 17552 8848 17558 8900
rect 18138 8848 18144 8900
rect 18196 8888 18202 8900
rect 19426 8888 19432 8900
rect 18196 8860 19432 8888
rect 18196 8848 18202 8860
rect 19426 8848 19432 8860
rect 19484 8848 19490 8900
rect 19720 8888 19748 8996
rect 19886 8984 19892 8996
rect 19944 8984 19950 9036
rect 20990 9024 20996 9036
rect 20951 8996 20996 9024
rect 20990 8984 20996 8996
rect 21048 8984 21054 9036
rect 19978 8916 19984 8968
rect 20036 8956 20042 8968
rect 20441 8959 20499 8965
rect 20441 8956 20453 8959
rect 20036 8928 20453 8956
rect 20036 8916 20042 8928
rect 20441 8925 20453 8928
rect 20487 8925 20499 8959
rect 20441 8919 20499 8925
rect 20622 8916 20628 8968
rect 20680 8956 20686 8968
rect 20717 8959 20775 8965
rect 20717 8956 20729 8959
rect 20680 8928 20729 8956
rect 20680 8916 20686 8928
rect 20717 8925 20729 8928
rect 20763 8925 20775 8959
rect 20717 8919 20775 8925
rect 20165 8891 20223 8897
rect 20165 8888 20177 8891
rect 19720 8860 20177 8888
rect 20165 8857 20177 8860
rect 20211 8888 20223 8891
rect 20530 8888 20536 8900
rect 20211 8860 20536 8888
rect 20211 8857 20223 8860
rect 20165 8851 20223 8857
rect 20530 8848 20536 8860
rect 20588 8848 20594 8900
rect 17034 8820 17040 8832
rect 13964 8792 14596 8820
rect 16995 8792 17040 8820
rect 13964 8780 13970 8792
rect 17034 8780 17040 8792
rect 17092 8780 17098 8832
rect 17405 8823 17463 8829
rect 17405 8789 17417 8823
rect 17451 8820 17463 8823
rect 17586 8820 17592 8832
rect 17451 8792 17592 8820
rect 17451 8789 17463 8792
rect 17405 8783 17463 8789
rect 17586 8780 17592 8792
rect 17644 8780 17650 8832
rect 18322 8780 18328 8832
rect 18380 8820 18386 8832
rect 18598 8820 18604 8832
rect 18380 8792 18604 8820
rect 18380 8780 18386 8792
rect 18598 8780 18604 8792
rect 18656 8780 18662 8832
rect 18690 8780 18696 8832
rect 18748 8820 18754 8832
rect 18748 8792 18793 8820
rect 18748 8780 18754 8792
rect 18966 8780 18972 8832
rect 19024 8820 19030 8832
rect 19061 8823 19119 8829
rect 19061 8820 19073 8823
rect 19024 8792 19073 8820
rect 19024 8780 19030 8792
rect 19061 8789 19073 8792
rect 19107 8789 19119 8823
rect 19061 8783 19119 8789
rect 19518 8780 19524 8832
rect 19576 8820 19582 8832
rect 19613 8823 19671 8829
rect 19613 8820 19625 8823
rect 19576 8792 19625 8820
rect 19576 8780 19582 8792
rect 19613 8789 19625 8792
rect 19659 8789 19671 8823
rect 19613 8783 19671 8789
rect 19705 8823 19763 8829
rect 19705 8789 19717 8823
rect 19751 8820 19763 8823
rect 20070 8820 20076 8832
rect 19751 8792 20076 8820
rect 19751 8789 19763 8792
rect 19705 8783 19763 8789
rect 20070 8780 20076 8792
rect 20128 8780 20134 8832
rect 1104 8730 22056 8752
rect 1104 8678 6148 8730
rect 6200 8678 6212 8730
rect 6264 8678 6276 8730
rect 6328 8678 6340 8730
rect 6392 8678 6404 8730
rect 6456 8678 11346 8730
rect 11398 8678 11410 8730
rect 11462 8678 11474 8730
rect 11526 8678 11538 8730
rect 11590 8678 11602 8730
rect 11654 8678 16544 8730
rect 16596 8678 16608 8730
rect 16660 8678 16672 8730
rect 16724 8678 16736 8730
rect 16788 8678 16800 8730
rect 16852 8678 21742 8730
rect 21794 8678 21806 8730
rect 21858 8678 21870 8730
rect 21922 8678 21934 8730
rect 21986 8678 21998 8730
rect 22050 8678 22056 8730
rect 1104 8656 22056 8678
rect 1578 8616 1584 8628
rect 1539 8588 1584 8616
rect 1578 8576 1584 8588
rect 1636 8576 1642 8628
rect 2409 8619 2467 8625
rect 2409 8585 2421 8619
rect 2455 8616 2467 8619
rect 2774 8616 2780 8628
rect 2455 8588 2780 8616
rect 2455 8585 2467 8588
rect 2409 8579 2467 8585
rect 2774 8576 2780 8588
rect 2832 8576 2838 8628
rect 2866 8576 2872 8628
rect 2924 8616 2930 8628
rect 2924 8588 2969 8616
rect 2924 8576 2930 8588
rect 3142 8576 3148 8628
rect 3200 8616 3206 8628
rect 3237 8619 3295 8625
rect 3237 8616 3249 8619
rect 3200 8588 3249 8616
rect 3200 8576 3206 8588
rect 3237 8585 3249 8588
rect 3283 8585 3295 8619
rect 3237 8579 3295 8585
rect 3326 8576 3332 8628
rect 3384 8616 3390 8628
rect 3789 8619 3847 8625
rect 3789 8616 3801 8619
rect 3384 8588 3801 8616
rect 3384 8576 3390 8588
rect 3789 8585 3801 8588
rect 3835 8585 3847 8619
rect 3789 8579 3847 8585
rect 4249 8619 4307 8625
rect 4249 8585 4261 8619
rect 4295 8616 4307 8619
rect 7834 8616 7840 8628
rect 4295 8588 7840 8616
rect 4295 8585 4307 8588
rect 4249 8579 4307 8585
rect 7834 8576 7840 8588
rect 7892 8576 7898 8628
rect 11054 8576 11060 8628
rect 11112 8616 11118 8628
rect 11333 8619 11391 8625
rect 11333 8616 11345 8619
rect 11112 8588 11345 8616
rect 11112 8576 11118 8588
rect 11333 8585 11345 8588
rect 11379 8585 11391 8619
rect 11333 8579 11391 8585
rect 11422 8576 11428 8628
rect 11480 8616 11486 8628
rect 13449 8619 13507 8625
rect 13449 8616 13461 8619
rect 11480 8588 13461 8616
rect 11480 8576 11486 8588
rect 13449 8585 13461 8588
rect 13495 8616 13507 8619
rect 15654 8616 15660 8628
rect 13495 8588 15660 8616
rect 13495 8585 13507 8588
rect 13449 8579 13507 8585
rect 15654 8576 15660 8588
rect 15712 8576 15718 8628
rect 16574 8616 16580 8628
rect 16316 8588 16580 8616
rect 3605 8551 3663 8557
rect 3605 8548 3617 8551
rect 1412 8520 3617 8548
rect 1302 8440 1308 8492
rect 1360 8480 1366 8492
rect 1412 8489 1440 8520
rect 3605 8517 3617 8520
rect 3651 8517 3663 8551
rect 5626 8548 5632 8560
rect 3605 8511 3663 8517
rect 3988 8520 5632 8548
rect 1397 8483 1455 8489
rect 1397 8480 1409 8483
rect 1360 8452 1409 8480
rect 1360 8440 1366 8452
rect 1397 8449 1409 8452
rect 1443 8449 1455 8483
rect 2038 8480 2044 8492
rect 1999 8452 2044 8480
rect 1397 8443 1455 8449
rect 2038 8440 2044 8452
rect 2096 8440 2102 8492
rect 3988 8480 4016 8520
rect 5626 8508 5632 8520
rect 5684 8508 5690 8560
rect 6457 8551 6515 8557
rect 6457 8517 6469 8551
rect 6503 8548 6515 8551
rect 6546 8548 6552 8560
rect 6503 8520 6552 8548
rect 6503 8517 6515 8520
rect 6457 8511 6515 8517
rect 6546 8508 6552 8520
rect 6604 8548 6610 8560
rect 6641 8551 6699 8557
rect 6641 8548 6653 8551
rect 6604 8520 6653 8548
rect 6604 8508 6610 8520
rect 6641 8517 6653 8520
rect 6687 8548 6699 8551
rect 7193 8551 7251 8557
rect 7193 8548 7205 8551
rect 6687 8520 7205 8548
rect 6687 8517 6699 8520
rect 6641 8511 6699 8517
rect 7193 8517 7205 8520
rect 7239 8548 7251 8551
rect 10321 8551 10379 8557
rect 7239 8520 8708 8548
rect 7239 8517 7251 8520
rect 7193 8511 7251 8517
rect 4154 8480 4160 8492
rect 2608 8452 4016 8480
rect 4115 8452 4160 8480
rect 1765 8415 1823 8421
rect 1765 8381 1777 8415
rect 1811 8381 1823 8415
rect 1946 8412 1952 8424
rect 1907 8384 1952 8412
rect 1765 8375 1823 8381
rect 1780 8344 1808 8375
rect 1946 8372 1952 8384
rect 2004 8372 2010 8424
rect 2608 8421 2636 8452
rect 4154 8440 4160 8452
rect 4212 8440 4218 8492
rect 7374 8440 7380 8492
rect 7432 8480 7438 8492
rect 8680 8489 8708 8520
rect 10321 8517 10333 8551
rect 10367 8548 10379 8551
rect 10873 8551 10931 8557
rect 10873 8548 10885 8551
rect 10367 8520 10885 8548
rect 10367 8517 10379 8520
rect 10321 8511 10379 8517
rect 10873 8517 10885 8520
rect 10919 8548 10931 8551
rect 11146 8548 11152 8560
rect 10919 8520 11152 8548
rect 10919 8517 10931 8520
rect 10873 8511 10931 8517
rect 11146 8508 11152 8520
rect 11204 8508 11210 8560
rect 12336 8551 12394 8557
rect 12336 8517 12348 8551
rect 12382 8548 12394 8551
rect 12526 8548 12532 8560
rect 12382 8520 12532 8548
rect 12382 8517 12394 8520
rect 12336 8511 12394 8517
rect 12526 8508 12532 8520
rect 12584 8508 12590 8560
rect 13814 8508 13820 8560
rect 13872 8548 13878 8560
rect 16218 8551 16276 8557
rect 13872 8520 15056 8548
rect 13872 8508 13878 8520
rect 8398 8483 8456 8489
rect 8398 8480 8410 8483
rect 7432 8452 8410 8480
rect 7432 8440 7438 8452
rect 8398 8449 8410 8452
rect 8444 8449 8456 8483
rect 8398 8443 8456 8449
rect 8665 8483 8723 8489
rect 8665 8449 8677 8483
rect 8711 8480 8723 8483
rect 8754 8480 8760 8492
rect 8711 8452 8760 8480
rect 8711 8449 8723 8452
rect 8665 8443 8723 8449
rect 8754 8440 8760 8452
rect 8812 8440 8818 8492
rect 8846 8440 8852 8492
rect 8904 8480 8910 8492
rect 9013 8483 9071 8489
rect 9013 8480 9025 8483
rect 8904 8452 9025 8480
rect 8904 8440 8910 8452
rect 9013 8449 9025 8452
rect 9059 8449 9071 8483
rect 10962 8480 10968 8492
rect 10923 8452 10968 8480
rect 9013 8443 9071 8449
rect 10962 8440 10968 8452
rect 11020 8440 11026 8492
rect 14274 8440 14280 8492
rect 14332 8480 14338 8492
rect 15028 8489 15056 8520
rect 16218 8517 16230 8551
rect 16264 8548 16276 8551
rect 16316 8548 16344 8588
rect 16574 8576 16580 8588
rect 16632 8576 16638 8628
rect 17402 8616 17408 8628
rect 17363 8588 17408 8616
rect 17402 8576 17408 8588
rect 17460 8576 17466 8628
rect 17954 8616 17960 8628
rect 17915 8588 17960 8616
rect 17954 8576 17960 8588
rect 18012 8576 18018 8628
rect 18877 8619 18935 8625
rect 18877 8585 18889 8619
rect 18923 8585 18935 8619
rect 18877 8579 18935 8585
rect 19521 8619 19579 8625
rect 19521 8585 19533 8619
rect 19567 8616 19579 8619
rect 19981 8619 20039 8625
rect 19981 8616 19993 8619
rect 19567 8588 19993 8616
rect 19567 8585 19579 8588
rect 19521 8579 19579 8585
rect 19981 8585 19993 8588
rect 20027 8585 20039 8619
rect 20806 8616 20812 8628
rect 20767 8588 20812 8616
rect 19981 8579 20039 8585
rect 16264 8520 16344 8548
rect 16264 8517 16276 8520
rect 16218 8511 16276 8517
rect 16390 8508 16396 8560
rect 16448 8548 16454 8560
rect 16448 8520 16528 8548
rect 16448 8508 16454 8520
rect 16500 8489 16528 8520
rect 17310 8508 17316 8560
rect 17368 8548 17374 8560
rect 18892 8548 18920 8579
rect 20806 8576 20812 8588
rect 20864 8576 20870 8628
rect 17368 8520 18920 8548
rect 17368 8508 17374 8520
rect 18966 8508 18972 8560
rect 19024 8548 19030 8560
rect 21177 8551 21235 8557
rect 21177 8548 21189 8551
rect 19024 8520 21189 8548
rect 19024 8508 19030 8520
rect 21177 8517 21189 8520
rect 21223 8517 21235 8551
rect 21177 8511 21235 8517
rect 14757 8483 14815 8489
rect 14757 8480 14769 8483
rect 14332 8452 14769 8480
rect 14332 8440 14338 8452
rect 14757 8449 14769 8452
rect 14803 8480 14815 8483
rect 15013 8483 15071 8489
rect 14803 8452 14964 8480
rect 14803 8449 14815 8452
rect 14757 8443 14815 8449
rect 2593 8415 2651 8421
rect 2593 8381 2605 8415
rect 2639 8381 2651 8415
rect 2593 8375 2651 8381
rect 2774 8372 2780 8424
rect 2832 8412 2838 8424
rect 3326 8412 3332 8424
rect 2832 8384 2877 8412
rect 3287 8384 3332 8412
rect 2832 8372 2838 8384
rect 3326 8372 3332 8384
rect 3384 8372 3390 8424
rect 4062 8372 4068 8424
rect 4120 8412 4126 8424
rect 4341 8415 4399 8421
rect 4341 8412 4353 8415
rect 4120 8384 4353 8412
rect 4120 8372 4126 8384
rect 4341 8381 4353 8384
rect 4387 8381 4399 8415
rect 7650 8412 7656 8424
rect 4341 8375 4399 8381
rect 5092 8384 7656 8412
rect 3418 8344 3424 8356
rect 1780 8316 3424 8344
rect 3418 8304 3424 8316
rect 3476 8344 3482 8356
rect 5092 8344 5120 8384
rect 7650 8372 7656 8384
rect 7708 8372 7714 8424
rect 10689 8415 10747 8421
rect 10689 8412 10701 8415
rect 9784 8384 10701 8412
rect 3476 8316 5120 8344
rect 3476 8304 3482 8316
rect 5166 8304 5172 8356
rect 5224 8344 5230 8356
rect 7285 8347 7343 8353
rect 7285 8344 7297 8347
rect 5224 8316 7297 8344
rect 5224 8304 5230 8316
rect 7285 8313 7297 8316
rect 7331 8313 7343 8347
rect 9784 8344 9812 8384
rect 10689 8381 10701 8384
rect 10735 8381 10747 8415
rect 10689 8375 10747 8381
rect 11793 8415 11851 8421
rect 11793 8381 11805 8415
rect 11839 8412 11851 8415
rect 12069 8415 12127 8421
rect 12069 8412 12081 8415
rect 11839 8384 12081 8412
rect 11839 8381 11851 8384
rect 11793 8375 11851 8381
rect 10134 8344 10140 8356
rect 7285 8307 7343 8313
rect 9692 8316 9812 8344
rect 10047 8316 10140 8344
rect 2130 8236 2136 8288
rect 2188 8276 2194 8288
rect 4062 8276 4068 8288
rect 2188 8248 4068 8276
rect 2188 8236 2194 8248
rect 4062 8236 4068 8248
rect 4120 8236 4126 8288
rect 8478 8236 8484 8288
rect 8536 8276 8542 8288
rect 9692 8276 9720 8316
rect 10134 8304 10140 8316
rect 10192 8344 10198 8356
rect 10192 8316 10364 8344
rect 10192 8304 10198 8316
rect 8536 8248 9720 8276
rect 10336 8276 10364 8316
rect 10502 8304 10508 8356
rect 10560 8344 10566 8356
rect 11992 8344 12020 8384
rect 12069 8381 12081 8384
rect 12115 8381 12127 8415
rect 14936 8412 14964 8452
rect 15013 8449 15025 8483
rect 15059 8449 15071 8483
rect 16485 8483 16543 8489
rect 15013 8443 15071 8449
rect 15120 8452 16436 8480
rect 15120 8412 15148 8452
rect 14936 8384 15148 8412
rect 16408 8412 16436 8452
rect 16485 8449 16497 8483
rect 16531 8449 16543 8483
rect 17034 8480 17040 8492
rect 16995 8452 17040 8480
rect 16485 8443 16543 8449
rect 17034 8440 17040 8452
rect 17092 8440 17098 8492
rect 17865 8483 17923 8489
rect 17865 8449 17877 8483
rect 17911 8480 17923 8483
rect 18325 8483 18383 8489
rect 18325 8480 18337 8483
rect 17911 8452 18337 8480
rect 17911 8449 17923 8452
rect 17865 8443 17923 8449
rect 18325 8449 18337 8452
rect 18371 8449 18383 8483
rect 18325 8443 18383 8449
rect 18785 8483 18843 8489
rect 18785 8449 18797 8483
rect 18831 8480 18843 8483
rect 19061 8483 19119 8489
rect 19061 8480 19073 8483
rect 18831 8452 19073 8480
rect 18831 8449 18843 8452
rect 18785 8443 18843 8449
rect 19061 8449 19073 8452
rect 19107 8480 19119 8483
rect 19242 8480 19248 8492
rect 19107 8452 19248 8480
rect 19107 8449 19119 8452
rect 19061 8443 19119 8449
rect 19242 8440 19248 8452
rect 19300 8440 19306 8492
rect 19518 8440 19524 8492
rect 19576 8480 19582 8492
rect 20346 8480 20352 8492
rect 19576 8452 20352 8480
rect 19576 8440 19582 8452
rect 20346 8440 20352 8452
rect 20404 8440 20410 8492
rect 16761 8415 16819 8421
rect 16761 8412 16773 8415
rect 16408 8384 16773 8412
rect 12069 8375 12127 8381
rect 16761 8381 16773 8384
rect 16807 8381 16819 8415
rect 16942 8412 16948 8424
rect 16903 8384 16948 8412
rect 16761 8375 16819 8381
rect 16942 8372 16948 8384
rect 17000 8372 17006 8424
rect 18141 8415 18199 8421
rect 18141 8381 18153 8415
rect 18187 8381 18199 8415
rect 19610 8412 19616 8424
rect 19571 8384 19616 8412
rect 18141 8375 18199 8381
rect 10560 8316 12020 8344
rect 10560 8304 10566 8316
rect 11992 8288 12020 8316
rect 13633 8347 13691 8353
rect 13633 8313 13645 8347
rect 13679 8344 13691 8347
rect 13906 8344 13912 8356
rect 13679 8316 13912 8344
rect 13679 8313 13691 8316
rect 13633 8307 13691 8313
rect 13906 8304 13912 8316
rect 13964 8304 13970 8356
rect 15105 8347 15163 8353
rect 15105 8313 15117 8347
rect 15151 8344 15163 8347
rect 15194 8344 15200 8356
rect 15151 8316 15200 8344
rect 15151 8313 15163 8316
rect 15105 8307 15163 8313
rect 15194 8304 15200 8316
rect 15252 8304 15258 8356
rect 16574 8304 16580 8356
rect 16632 8344 16638 8356
rect 16632 8316 17724 8344
rect 16632 8304 16638 8316
rect 17696 8288 17724 8316
rect 10870 8276 10876 8288
rect 10336 8248 10876 8276
rect 8536 8236 8542 8248
rect 10870 8236 10876 8248
rect 10928 8236 10934 8288
rect 11974 8276 11980 8288
rect 11935 8248 11980 8276
rect 11974 8236 11980 8248
rect 12032 8236 12038 8288
rect 17494 8236 17500 8288
rect 17552 8276 17558 8288
rect 17552 8248 17597 8276
rect 17552 8236 17558 8248
rect 17678 8236 17684 8288
rect 17736 8276 17742 8288
rect 18156 8276 18184 8375
rect 19610 8372 19616 8384
rect 19668 8372 19674 8424
rect 19705 8415 19763 8421
rect 19705 8381 19717 8415
rect 19751 8381 19763 8415
rect 20438 8412 20444 8424
rect 20399 8384 20444 8412
rect 19705 8375 19763 8381
rect 18506 8304 18512 8356
rect 18564 8344 18570 8356
rect 19153 8347 19211 8353
rect 19153 8344 19165 8347
rect 18564 8316 19165 8344
rect 18564 8304 18570 8316
rect 19153 8313 19165 8316
rect 19199 8313 19211 8347
rect 19153 8307 19211 8313
rect 19426 8304 19432 8356
rect 19484 8344 19490 8356
rect 19720 8344 19748 8375
rect 20438 8372 20444 8384
rect 20496 8372 20502 8424
rect 20530 8372 20536 8424
rect 20588 8412 20594 8424
rect 21266 8412 21272 8424
rect 20588 8384 20633 8412
rect 21227 8384 21272 8412
rect 20588 8372 20594 8384
rect 21266 8372 21272 8384
rect 21324 8372 21330 8424
rect 21361 8415 21419 8421
rect 21361 8381 21373 8415
rect 21407 8381 21419 8415
rect 21361 8375 21419 8381
rect 21376 8344 21404 8375
rect 19484 8316 21404 8344
rect 19484 8304 19490 8316
rect 18690 8276 18696 8288
rect 17736 8248 18696 8276
rect 17736 8236 17742 8248
rect 18690 8236 18696 8248
rect 18748 8236 18754 8288
rect 1104 8186 21896 8208
rect 1104 8134 3549 8186
rect 3601 8134 3613 8186
rect 3665 8134 3677 8186
rect 3729 8134 3741 8186
rect 3793 8134 3805 8186
rect 3857 8134 8747 8186
rect 8799 8134 8811 8186
rect 8863 8134 8875 8186
rect 8927 8134 8939 8186
rect 8991 8134 9003 8186
rect 9055 8134 13945 8186
rect 13997 8134 14009 8186
rect 14061 8134 14073 8186
rect 14125 8134 14137 8186
rect 14189 8134 14201 8186
rect 14253 8134 19143 8186
rect 19195 8134 19207 8186
rect 19259 8134 19271 8186
rect 19323 8134 19335 8186
rect 19387 8134 19399 8186
rect 19451 8134 21896 8186
rect 1104 8112 21896 8134
rect 1394 8072 1400 8084
rect 1355 8044 1400 8072
rect 1394 8032 1400 8044
rect 1452 8032 1458 8084
rect 1946 8032 1952 8084
rect 2004 8072 2010 8084
rect 2409 8075 2467 8081
rect 2409 8072 2421 8075
rect 2004 8044 2421 8072
rect 2004 8032 2010 8044
rect 2409 8041 2421 8044
rect 2455 8041 2467 8075
rect 2409 8035 2467 8041
rect 2501 8075 2559 8081
rect 2501 8041 2513 8075
rect 2547 8072 2559 8075
rect 2774 8072 2780 8084
rect 2547 8044 2780 8072
rect 2547 8041 2559 8044
rect 2501 8035 2559 8041
rect 2774 8032 2780 8044
rect 2832 8032 2838 8084
rect 3513 8075 3571 8081
rect 3513 8041 3525 8075
rect 3559 8072 3571 8075
rect 3559 8044 10456 8072
rect 3559 8041 3571 8044
rect 3513 8035 3571 8041
rect 3970 7964 3976 8016
rect 4028 8004 4034 8016
rect 4341 8007 4399 8013
rect 4341 8004 4353 8007
rect 4028 7976 4353 8004
rect 4028 7964 4034 7976
rect 4341 7973 4353 7976
rect 4387 7973 4399 8007
rect 4341 7967 4399 7973
rect 4522 7964 4528 8016
rect 4580 8004 4586 8016
rect 5261 8007 5319 8013
rect 5261 8004 5273 8007
rect 4580 7976 5273 8004
rect 4580 7964 4586 7976
rect 5261 7973 5273 7976
rect 5307 7973 5319 8007
rect 5626 8004 5632 8016
rect 5587 7976 5632 8004
rect 5261 7967 5319 7973
rect 5626 7964 5632 7976
rect 5684 7964 5690 8016
rect 7374 8004 7380 8016
rect 7335 7976 7380 8004
rect 7374 7964 7380 7976
rect 7432 7964 7438 8016
rect 9674 8004 9680 8016
rect 9635 7976 9680 8004
rect 9674 7964 9680 7976
rect 9732 7964 9738 8016
rect 1857 7939 1915 7945
rect 1857 7905 1869 7939
rect 1903 7936 1915 7939
rect 2130 7936 2136 7948
rect 1903 7908 2136 7936
rect 1903 7905 1915 7908
rect 1857 7899 1915 7905
rect 2130 7896 2136 7908
rect 2188 7896 2194 7948
rect 2498 7896 2504 7948
rect 2556 7936 2562 7948
rect 3145 7939 3203 7945
rect 3145 7936 3157 7939
rect 2556 7908 3157 7936
rect 2556 7896 2562 7908
rect 3145 7905 3157 7908
rect 3191 7936 3203 7939
rect 4985 7939 5043 7945
rect 3191 7908 4844 7936
rect 3191 7905 3203 7908
rect 3145 7899 3203 7905
rect 2041 7871 2099 7877
rect 2041 7837 2053 7871
rect 2087 7868 2099 7871
rect 2682 7868 2688 7880
rect 2087 7840 2688 7868
rect 2087 7837 2099 7840
rect 2041 7831 2099 7837
rect 2682 7828 2688 7840
rect 2740 7828 2746 7880
rect 1949 7803 2007 7809
rect 1949 7769 1961 7803
rect 1995 7800 2007 7803
rect 2869 7803 2927 7809
rect 2869 7800 2881 7803
rect 1995 7772 2881 7800
rect 1995 7769 2007 7772
rect 1949 7763 2007 7769
rect 2869 7769 2881 7772
rect 2915 7800 2927 7803
rect 3050 7800 3056 7812
rect 2915 7772 3056 7800
rect 2915 7769 2927 7772
rect 2869 7763 2927 7769
rect 3050 7760 3056 7772
rect 3108 7760 3114 7812
rect 3418 7800 3424 7812
rect 3379 7772 3424 7800
rect 3418 7760 3424 7772
rect 3476 7800 3482 7812
rect 3789 7803 3847 7809
rect 3789 7800 3801 7803
rect 3476 7772 3801 7800
rect 3476 7760 3482 7772
rect 3789 7769 3801 7772
rect 3835 7769 3847 7803
rect 4816 7800 4844 7908
rect 4985 7905 4997 7939
rect 5031 7936 5043 7939
rect 5166 7936 5172 7948
rect 5031 7908 5172 7936
rect 5031 7905 5043 7908
rect 4985 7899 5043 7905
rect 5166 7896 5172 7908
rect 5224 7896 5230 7948
rect 9125 7939 9183 7945
rect 9125 7905 9137 7939
rect 9171 7936 9183 7939
rect 9398 7936 9404 7948
rect 9171 7908 9404 7936
rect 9171 7905 9183 7908
rect 9125 7899 9183 7905
rect 9398 7896 9404 7908
rect 9456 7896 9462 7948
rect 5537 7871 5595 7877
rect 5537 7837 5549 7871
rect 5583 7868 5595 7871
rect 6454 7868 6460 7880
rect 5583 7840 6460 7868
rect 5583 7837 5595 7840
rect 5537 7831 5595 7837
rect 6454 7828 6460 7840
rect 6512 7828 6518 7880
rect 7009 7871 7067 7877
rect 7009 7837 7021 7871
rect 7055 7868 7067 7871
rect 7285 7871 7343 7877
rect 7285 7868 7297 7871
rect 7055 7840 7297 7868
rect 7055 7837 7067 7840
rect 7009 7831 7067 7837
rect 7285 7837 7297 7840
rect 7331 7868 7343 7871
rect 8662 7868 8668 7880
rect 7331 7840 8668 7868
rect 7331 7837 7343 7840
rect 7285 7831 7343 7837
rect 8662 7828 8668 7840
rect 8720 7868 8726 7880
rect 8757 7871 8815 7877
rect 8757 7868 8769 7871
rect 8720 7840 8769 7868
rect 8720 7828 8726 7840
rect 8757 7837 8769 7840
rect 8803 7837 8815 7871
rect 8757 7831 8815 7837
rect 9217 7871 9275 7877
rect 9217 7837 9229 7871
rect 9263 7868 9275 7871
rect 9674 7868 9680 7880
rect 9263 7840 9680 7868
rect 9263 7837 9275 7840
rect 9217 7831 9275 7837
rect 9674 7828 9680 7840
rect 9732 7828 9738 7880
rect 6822 7809 6828 7812
rect 6764 7803 6828 7809
rect 6764 7800 6776 7803
rect 4816 7772 6776 7800
rect 3789 7763 3847 7769
rect 6764 7769 6776 7772
rect 6810 7769 6828 7803
rect 6764 7763 6828 7769
rect 6822 7760 6828 7763
rect 6880 7760 6886 7812
rect 8386 7760 8392 7812
rect 8444 7800 8450 7812
rect 8490 7803 8548 7809
rect 8490 7800 8502 7803
rect 8444 7772 8502 7800
rect 8444 7760 8450 7772
rect 8490 7769 8502 7772
rect 8536 7769 8548 7803
rect 10428 7800 10456 8044
rect 10502 8032 10508 8084
rect 10560 8032 10566 8084
rect 11057 8075 11115 8081
rect 11057 8041 11069 8075
rect 11103 8072 11115 8075
rect 11103 8044 16620 8072
rect 11103 8041 11115 8044
rect 11057 8035 11115 8041
rect 10520 8004 10548 8032
rect 11149 8007 11207 8013
rect 11149 8004 11161 8007
rect 10520 7976 11161 8004
rect 11149 7973 11161 7976
rect 11195 7973 11207 8007
rect 11149 7967 11207 7973
rect 14093 8007 14151 8013
rect 14093 7973 14105 8007
rect 14139 8004 14151 8007
rect 14274 8004 14280 8016
rect 14139 7976 14280 8004
rect 14139 7973 14151 7976
rect 14093 7967 14151 7973
rect 14274 7964 14280 7976
rect 14332 7964 14338 8016
rect 10505 7939 10563 7945
rect 10505 7905 10517 7939
rect 10551 7936 10563 7939
rect 11422 7936 11428 7948
rect 10551 7908 11428 7936
rect 10551 7905 10563 7908
rect 10505 7899 10563 7905
rect 11422 7896 11428 7908
rect 11480 7896 11486 7948
rect 16482 7936 16488 7948
rect 16443 7908 16488 7936
rect 16482 7896 16488 7908
rect 16540 7896 16546 7948
rect 16592 7945 16620 8044
rect 16942 8032 16948 8084
rect 17000 8072 17006 8084
rect 17129 8075 17187 8081
rect 17129 8072 17141 8075
rect 17000 8044 17141 8072
rect 17000 8032 17006 8044
rect 17129 8041 17141 8044
rect 17175 8041 17187 8075
rect 19610 8072 19616 8084
rect 19571 8044 19616 8072
rect 17129 8035 17187 8041
rect 19610 8032 19616 8044
rect 19668 8032 19674 8084
rect 20533 8075 20591 8081
rect 20533 8041 20545 8075
rect 20579 8072 20591 8075
rect 20622 8072 20628 8084
rect 20579 8044 20628 8072
rect 20579 8041 20591 8044
rect 20533 8035 20591 8041
rect 20622 8032 20628 8044
rect 20680 8032 20686 8084
rect 21266 8032 21272 8084
rect 21324 8072 21330 8084
rect 21361 8075 21419 8081
rect 21361 8072 21373 8075
rect 21324 8044 21373 8072
rect 21324 8032 21330 8044
rect 21361 8041 21373 8044
rect 21407 8041 21419 8075
rect 21542 8072 21548 8084
rect 21503 8044 21548 8072
rect 21361 8035 21419 8041
rect 21542 8032 21548 8044
rect 21600 8032 21606 8084
rect 16577 7939 16635 7945
rect 16577 7905 16589 7939
rect 16623 7905 16635 7939
rect 17681 7939 17739 7945
rect 17681 7936 17693 7939
rect 16577 7899 16635 7905
rect 16776 7908 17693 7936
rect 10594 7868 10600 7880
rect 10555 7840 10600 7868
rect 10594 7828 10600 7840
rect 10652 7828 10658 7880
rect 10689 7871 10747 7877
rect 10689 7837 10701 7871
rect 10735 7868 10747 7871
rect 11054 7868 11060 7880
rect 10735 7840 11060 7868
rect 10735 7837 10747 7840
rect 10689 7831 10747 7837
rect 11054 7828 11060 7840
rect 11112 7868 11118 7880
rect 11790 7868 11796 7880
rect 11112 7840 11796 7868
rect 11112 7828 11118 7840
rect 11790 7828 11796 7840
rect 11848 7828 11854 7880
rect 11974 7828 11980 7880
rect 12032 7868 12038 7880
rect 12529 7871 12587 7877
rect 12529 7868 12541 7871
rect 12032 7840 12541 7868
rect 12032 7828 12038 7840
rect 12529 7837 12541 7840
rect 12575 7868 12587 7871
rect 13449 7871 13507 7877
rect 13449 7868 13461 7871
rect 12575 7840 13461 7868
rect 12575 7837 12587 7840
rect 12529 7831 12587 7837
rect 13449 7837 13461 7840
rect 13495 7868 13507 7871
rect 13814 7868 13820 7880
rect 13495 7840 13820 7868
rect 13495 7837 13507 7840
rect 13449 7831 13507 7837
rect 13814 7828 13820 7840
rect 13872 7868 13878 7880
rect 15473 7871 15531 7877
rect 15473 7868 15485 7871
rect 13872 7840 15485 7868
rect 13872 7828 13878 7840
rect 15473 7837 15485 7840
rect 15519 7868 15531 7871
rect 15565 7871 15623 7877
rect 15565 7868 15577 7871
rect 15519 7840 15577 7868
rect 15519 7837 15531 7840
rect 15473 7831 15531 7837
rect 15565 7837 15577 7840
rect 15611 7837 15623 7871
rect 16666 7868 16672 7880
rect 16627 7840 16672 7868
rect 15565 7831 15623 7837
rect 16666 7828 16672 7840
rect 16724 7828 16730 7880
rect 12284 7803 12342 7809
rect 10428 7772 11284 7800
rect 8490 7763 8548 7769
rect 2961 7735 3019 7741
rect 2961 7701 2973 7735
rect 3007 7732 3019 7735
rect 3510 7732 3516 7744
rect 3007 7704 3516 7732
rect 3007 7701 3019 7704
rect 2961 7695 3019 7701
rect 3510 7692 3516 7704
rect 3568 7732 3574 7744
rect 4338 7732 4344 7744
rect 3568 7704 4344 7732
rect 3568 7692 3574 7704
rect 4338 7692 4344 7704
rect 4396 7692 4402 7744
rect 4706 7732 4712 7744
rect 4667 7704 4712 7732
rect 4706 7692 4712 7704
rect 4764 7692 4770 7744
rect 4801 7735 4859 7741
rect 4801 7701 4813 7735
rect 4847 7732 4859 7735
rect 5074 7732 5080 7744
rect 4847 7704 5080 7732
rect 4847 7701 4859 7704
rect 4801 7695 4859 7701
rect 5074 7692 5080 7704
rect 5132 7692 5138 7744
rect 5258 7692 5264 7744
rect 5316 7732 5322 7744
rect 6546 7732 6552 7744
rect 5316 7704 6552 7732
rect 5316 7692 5322 7704
rect 6546 7692 6552 7704
rect 6604 7692 6610 7744
rect 9309 7735 9367 7741
rect 9309 7701 9321 7735
rect 9355 7732 9367 7735
rect 9398 7732 9404 7744
rect 9355 7704 9404 7732
rect 9355 7701 9367 7704
rect 9309 7695 9367 7701
rect 9398 7692 9404 7704
rect 9456 7692 9462 7744
rect 11256 7732 11284 7772
rect 12284 7769 12296 7803
rect 12330 7800 12342 7803
rect 12986 7800 12992 7812
rect 12330 7772 12992 7800
rect 12330 7769 12342 7772
rect 12284 7763 12342 7769
rect 12986 7760 12992 7772
rect 13044 7800 13050 7812
rect 13722 7800 13728 7812
rect 13044 7772 13728 7800
rect 13044 7760 13050 7772
rect 13722 7760 13728 7772
rect 13780 7760 13786 7812
rect 15194 7760 15200 7812
rect 15252 7809 15258 7812
rect 15252 7800 15264 7809
rect 16390 7800 16396 7812
rect 15252 7772 16396 7800
rect 15252 7763 15264 7772
rect 15252 7760 15258 7763
rect 16390 7760 16396 7772
rect 16448 7800 16454 7812
rect 16776 7800 16804 7908
rect 17681 7905 17693 7908
rect 17727 7905 17739 7939
rect 17681 7899 17739 7905
rect 18601 7939 18659 7945
rect 18601 7905 18613 7939
rect 18647 7936 18659 7939
rect 18690 7936 18696 7948
rect 18647 7908 18696 7936
rect 18647 7905 18659 7908
rect 18601 7899 18659 7905
rect 18690 7896 18696 7908
rect 18748 7896 18754 7948
rect 20162 7936 20168 7948
rect 20123 7908 20168 7936
rect 20162 7896 20168 7908
rect 20220 7936 20226 7948
rect 20717 7939 20775 7945
rect 20717 7936 20729 7939
rect 20220 7908 20729 7936
rect 20220 7896 20226 7908
rect 20717 7905 20729 7908
rect 20763 7905 20775 7939
rect 20717 7899 20775 7905
rect 17770 7868 17776 7880
rect 16448 7772 16804 7800
rect 16960 7840 17776 7868
rect 16448 7760 16454 7772
rect 16960 7732 16988 7840
rect 17770 7828 17776 7840
rect 17828 7828 17834 7880
rect 18046 7828 18052 7880
rect 18104 7868 18110 7880
rect 20990 7868 20996 7880
rect 18104 7840 20996 7868
rect 18104 7828 18110 7840
rect 20990 7828 20996 7840
rect 21048 7828 21054 7880
rect 17589 7803 17647 7809
rect 17589 7800 17601 7803
rect 17052 7772 17601 7800
rect 17052 7741 17080 7772
rect 17589 7769 17601 7772
rect 17635 7769 17647 7803
rect 17589 7763 17647 7769
rect 17862 7760 17868 7812
rect 17920 7800 17926 7812
rect 18325 7803 18383 7809
rect 18325 7800 18337 7803
rect 17920 7772 18337 7800
rect 17920 7760 17926 7772
rect 18325 7769 18337 7772
rect 18371 7769 18383 7803
rect 18325 7763 18383 7769
rect 18782 7760 18788 7812
rect 18840 7800 18846 7812
rect 20901 7803 20959 7809
rect 20901 7800 20913 7803
rect 18840 7772 20913 7800
rect 18840 7760 18846 7772
rect 20901 7769 20913 7772
rect 20947 7800 20959 7803
rect 21082 7800 21088 7812
rect 20947 7772 21088 7800
rect 20947 7769 20959 7772
rect 20901 7763 20959 7769
rect 21082 7760 21088 7772
rect 21140 7760 21146 7812
rect 11256 7704 16988 7732
rect 17037 7735 17095 7741
rect 17037 7701 17049 7735
rect 17083 7701 17095 7735
rect 17037 7695 17095 7701
rect 17497 7735 17555 7741
rect 17497 7701 17509 7735
rect 17543 7732 17555 7735
rect 17770 7732 17776 7744
rect 17543 7704 17776 7732
rect 17543 7701 17555 7704
rect 17497 7695 17555 7701
rect 17770 7692 17776 7704
rect 17828 7692 17834 7744
rect 17954 7732 17960 7744
rect 17915 7704 17960 7732
rect 17954 7692 17960 7704
rect 18012 7692 18018 7744
rect 18414 7732 18420 7744
rect 18375 7704 18420 7732
rect 18414 7692 18420 7704
rect 18472 7732 18478 7744
rect 18598 7732 18604 7744
rect 18472 7704 18604 7732
rect 18472 7692 18478 7704
rect 18598 7692 18604 7704
rect 18656 7692 18662 7744
rect 19978 7732 19984 7744
rect 19939 7704 19984 7732
rect 19978 7692 19984 7704
rect 20036 7692 20042 7744
rect 20073 7735 20131 7741
rect 20073 7701 20085 7735
rect 20119 7732 20131 7735
rect 20254 7732 20260 7744
rect 20119 7704 20260 7732
rect 20119 7701 20131 7704
rect 20073 7695 20131 7701
rect 20254 7692 20260 7704
rect 20312 7692 20318 7744
rect 1104 7642 22056 7664
rect 1104 7590 6148 7642
rect 6200 7590 6212 7642
rect 6264 7590 6276 7642
rect 6328 7590 6340 7642
rect 6392 7590 6404 7642
rect 6456 7590 11346 7642
rect 11398 7590 11410 7642
rect 11462 7590 11474 7642
rect 11526 7590 11538 7642
rect 11590 7590 11602 7642
rect 11654 7590 16544 7642
rect 16596 7590 16608 7642
rect 16660 7590 16672 7642
rect 16724 7590 16736 7642
rect 16788 7590 16800 7642
rect 16852 7590 21742 7642
rect 21794 7590 21806 7642
rect 21858 7590 21870 7642
rect 21922 7590 21934 7642
rect 21986 7590 21998 7642
rect 22050 7590 22056 7642
rect 1104 7568 22056 7590
rect 2866 7488 2872 7540
rect 2924 7528 2930 7540
rect 3145 7531 3203 7537
rect 3145 7528 3157 7531
rect 2924 7500 3157 7528
rect 2924 7488 2930 7500
rect 3145 7497 3157 7500
rect 3191 7497 3203 7531
rect 3145 7491 3203 7497
rect 3513 7531 3571 7537
rect 3513 7497 3525 7531
rect 3559 7497 3571 7531
rect 3513 7491 3571 7497
rect 2406 7420 2412 7472
rect 2464 7460 2470 7472
rect 3528 7460 3556 7491
rect 4154 7488 4160 7540
rect 4212 7528 4218 7540
rect 4249 7531 4307 7537
rect 4249 7528 4261 7531
rect 4212 7500 4261 7528
rect 4212 7488 4218 7500
rect 4249 7497 4261 7500
rect 4295 7497 4307 7531
rect 4249 7491 4307 7497
rect 4522 7488 4528 7540
rect 4580 7528 4586 7540
rect 4617 7531 4675 7537
rect 4617 7528 4629 7531
rect 4580 7500 4629 7528
rect 4580 7488 4586 7500
rect 4617 7497 4629 7500
rect 4663 7497 4675 7531
rect 5074 7528 5080 7540
rect 5035 7500 5080 7528
rect 4617 7491 4675 7497
rect 5074 7488 5080 7500
rect 5132 7488 5138 7540
rect 5442 7528 5448 7540
rect 5403 7500 5448 7528
rect 5442 7488 5448 7500
rect 5500 7488 5506 7540
rect 5534 7488 5540 7540
rect 5592 7528 5598 7540
rect 6730 7528 6736 7540
rect 5592 7500 6736 7528
rect 5592 7488 5598 7500
rect 6730 7488 6736 7500
rect 6788 7488 6794 7540
rect 8202 7488 8208 7540
rect 8260 7528 8266 7540
rect 8941 7531 8999 7537
rect 8941 7528 8953 7531
rect 8260 7500 8953 7528
rect 8260 7488 8266 7500
rect 8941 7497 8953 7500
rect 8987 7497 8999 7531
rect 9398 7528 9404 7540
rect 9359 7500 9404 7528
rect 8941 7491 8999 7497
rect 9398 7488 9404 7500
rect 9456 7488 9462 7540
rect 9953 7531 10011 7537
rect 9953 7497 9965 7531
rect 9999 7528 10011 7531
rect 10321 7531 10379 7537
rect 10321 7528 10333 7531
rect 9999 7500 10333 7528
rect 9999 7497 10011 7500
rect 9953 7491 10011 7497
rect 10321 7497 10333 7500
rect 10367 7497 10379 7531
rect 10321 7491 10379 7497
rect 10689 7531 10747 7537
rect 10689 7497 10701 7531
rect 10735 7528 10747 7531
rect 11054 7528 11060 7540
rect 10735 7500 11060 7528
rect 10735 7497 10747 7500
rect 10689 7491 10747 7497
rect 11054 7488 11060 7500
rect 11112 7488 11118 7540
rect 11241 7531 11299 7537
rect 11241 7497 11253 7531
rect 11287 7528 11299 7531
rect 11974 7528 11980 7540
rect 11287 7500 11980 7528
rect 11287 7497 11299 7500
rect 11241 7491 11299 7497
rect 11974 7488 11980 7500
rect 12032 7488 12038 7540
rect 16853 7531 16911 7537
rect 16853 7497 16865 7531
rect 16899 7528 16911 7531
rect 17034 7528 17040 7540
rect 16899 7500 17040 7528
rect 16899 7497 16911 7500
rect 16853 7491 16911 7497
rect 17034 7488 17040 7500
rect 17092 7488 17098 7540
rect 17221 7531 17279 7537
rect 17221 7497 17233 7531
rect 17267 7528 17279 7531
rect 17494 7528 17500 7540
rect 17267 7500 17500 7528
rect 17267 7497 17279 7500
rect 17221 7491 17279 7497
rect 17494 7488 17500 7500
rect 17552 7488 17558 7540
rect 17770 7488 17776 7540
rect 17828 7528 17834 7540
rect 18141 7531 18199 7537
rect 18141 7528 18153 7531
rect 17828 7500 18153 7528
rect 17828 7488 17834 7500
rect 18141 7497 18153 7500
rect 18187 7497 18199 7531
rect 18141 7491 18199 7497
rect 20625 7531 20683 7537
rect 20625 7497 20637 7531
rect 20671 7528 20683 7531
rect 20898 7528 20904 7540
rect 20671 7500 20904 7528
rect 20671 7497 20683 7500
rect 20625 7491 20683 7497
rect 20898 7488 20904 7500
rect 20956 7488 20962 7540
rect 2464 7432 3556 7460
rect 2464 7420 2470 7432
rect 3878 7420 3884 7472
rect 3936 7460 3942 7472
rect 4062 7460 4068 7472
rect 3936 7432 4068 7460
rect 3936 7420 3942 7432
rect 4062 7420 4068 7432
rect 4120 7420 4126 7472
rect 4709 7463 4767 7469
rect 4709 7429 4721 7463
rect 4755 7460 4767 7463
rect 5258 7460 5264 7472
rect 4755 7432 5264 7460
rect 4755 7429 4767 7432
rect 4709 7423 4767 7429
rect 5258 7420 5264 7432
rect 5316 7420 5322 7472
rect 5350 7420 5356 7472
rect 5408 7460 5414 7472
rect 5997 7463 6055 7469
rect 5408 7432 5672 7460
rect 5408 7420 5414 7432
rect 2777 7395 2835 7401
rect 2777 7361 2789 7395
rect 2823 7392 2835 7395
rect 3237 7395 3295 7401
rect 3237 7392 3249 7395
rect 2823 7364 3249 7392
rect 2823 7361 2835 7364
rect 2777 7355 2835 7361
rect 3237 7361 3249 7364
rect 3283 7361 3295 7395
rect 3237 7355 3295 7361
rect 3697 7395 3755 7401
rect 3697 7361 3709 7395
rect 3743 7392 3755 7395
rect 3743 7364 3924 7392
rect 3743 7361 3755 7364
rect 3697 7355 3755 7361
rect 1946 7324 1952 7336
rect 1907 7296 1952 7324
rect 1946 7284 1952 7296
rect 2004 7284 2010 7336
rect 2222 7324 2228 7336
rect 2183 7296 2228 7324
rect 2222 7284 2228 7296
rect 2280 7284 2286 7336
rect 2498 7324 2504 7336
rect 2459 7296 2504 7324
rect 2498 7284 2504 7296
rect 2556 7284 2562 7336
rect 2590 7284 2596 7336
rect 2648 7324 2654 7336
rect 2685 7327 2743 7333
rect 2685 7324 2697 7327
rect 2648 7296 2697 7324
rect 2648 7284 2654 7296
rect 2685 7293 2697 7296
rect 2731 7293 2743 7327
rect 2685 7287 2743 7293
rect 3896 7197 3924 7364
rect 4798 7284 4804 7336
rect 4856 7324 4862 7336
rect 5537 7327 5595 7333
rect 4856 7296 4901 7324
rect 4856 7284 4862 7296
rect 5537 7293 5549 7327
rect 5583 7293 5595 7327
rect 5644 7324 5672 7432
rect 5997 7429 6009 7463
rect 6043 7460 6055 7463
rect 6546 7460 6552 7472
rect 6043 7432 6552 7460
rect 6043 7429 6055 7432
rect 5997 7423 6055 7429
rect 6546 7420 6552 7432
rect 6604 7420 6610 7472
rect 8386 7420 8392 7472
rect 8444 7460 8450 7472
rect 9122 7460 9128 7472
rect 8444 7432 9128 7460
rect 8444 7420 8450 7432
rect 9122 7420 9128 7432
rect 9180 7460 9186 7472
rect 9180 7432 10088 7460
rect 9180 7420 9186 7432
rect 8573 7395 8631 7401
rect 8573 7361 8585 7395
rect 8619 7392 8631 7395
rect 9033 7395 9091 7401
rect 9033 7392 9045 7395
rect 8619 7364 9045 7392
rect 8619 7361 8631 7364
rect 8573 7355 8631 7361
rect 9033 7361 9045 7364
rect 9079 7361 9091 7395
rect 9858 7392 9864 7404
rect 9819 7364 9864 7392
rect 9033 7355 9091 7361
rect 9858 7352 9864 7364
rect 9916 7352 9922 7404
rect 5721 7327 5779 7333
rect 5721 7324 5733 7327
rect 5644 7296 5733 7324
rect 5537 7287 5595 7293
rect 5721 7293 5733 7296
rect 5767 7324 5779 7327
rect 7374 7324 7380 7336
rect 5767 7296 7380 7324
rect 5767 7293 5779 7296
rect 5721 7287 5779 7293
rect 5552 7256 5580 7287
rect 7374 7284 7380 7296
rect 7432 7284 7438 7336
rect 8478 7284 8484 7336
rect 8536 7324 8542 7336
rect 10060 7333 10088 7432
rect 10594 7420 10600 7472
rect 10652 7460 10658 7472
rect 10781 7463 10839 7469
rect 10781 7460 10793 7463
rect 10652 7432 10793 7460
rect 10652 7420 10658 7432
rect 10781 7429 10793 7432
rect 10827 7429 10839 7463
rect 10781 7423 10839 7429
rect 17313 7463 17371 7469
rect 17313 7429 17325 7463
rect 17359 7460 17371 7463
rect 17954 7460 17960 7472
rect 17359 7432 17960 7460
rect 17359 7429 17371 7432
rect 17313 7423 17371 7429
rect 17954 7420 17960 7432
rect 18012 7420 18018 7472
rect 18046 7420 18052 7472
rect 18104 7460 18110 7472
rect 18509 7463 18567 7469
rect 18509 7460 18521 7463
rect 18104 7432 18521 7460
rect 18104 7420 18110 7432
rect 18509 7429 18521 7432
rect 18555 7429 18567 7463
rect 18509 7423 18567 7429
rect 18601 7463 18659 7469
rect 18601 7429 18613 7463
rect 18647 7460 18659 7463
rect 20346 7460 20352 7472
rect 18647 7432 20352 7460
rect 18647 7429 18659 7432
rect 18601 7423 18659 7429
rect 20346 7420 20352 7432
rect 20404 7420 20410 7472
rect 20441 7395 20499 7401
rect 20441 7392 20453 7395
rect 20088 7364 20453 7392
rect 8757 7327 8815 7333
rect 8757 7324 8769 7327
rect 8536 7296 8769 7324
rect 8536 7284 8542 7296
rect 8757 7293 8769 7296
rect 8803 7293 8815 7327
rect 8757 7287 8815 7293
rect 10045 7327 10103 7333
rect 10045 7293 10057 7327
rect 10091 7293 10103 7327
rect 10045 7287 10103 7293
rect 10870 7284 10876 7336
rect 10928 7324 10934 7336
rect 10928 7296 10973 7324
rect 10928 7284 10934 7296
rect 16390 7284 16396 7336
rect 16448 7324 16454 7336
rect 17405 7327 17463 7333
rect 17405 7324 17417 7327
rect 16448 7296 17417 7324
rect 16448 7284 16454 7296
rect 17405 7293 17417 7296
rect 17451 7293 17463 7327
rect 18690 7324 18696 7336
rect 18651 7296 18696 7324
rect 17405 7287 17463 7293
rect 18690 7284 18696 7296
rect 18748 7284 18754 7336
rect 8846 7256 8852 7268
rect 5552 7228 8852 7256
rect 8846 7216 8852 7228
rect 8904 7216 8910 7268
rect 9030 7216 9036 7268
rect 9088 7256 9094 7268
rect 9493 7259 9551 7265
rect 9493 7256 9505 7259
rect 9088 7228 9505 7256
rect 9088 7216 9094 7228
rect 9493 7225 9505 7228
rect 9539 7225 9551 7259
rect 9493 7219 9551 7225
rect 3881 7191 3939 7197
rect 3881 7157 3893 7191
rect 3927 7188 3939 7191
rect 4154 7188 4160 7200
rect 3927 7160 4160 7188
rect 3927 7157 3939 7160
rect 3881 7151 3939 7157
rect 4154 7148 4160 7160
rect 4212 7148 4218 7200
rect 8202 7188 8208 7200
rect 8163 7160 8208 7188
rect 8202 7148 8208 7160
rect 8260 7188 8266 7200
rect 9766 7188 9772 7200
rect 8260 7160 9772 7188
rect 8260 7148 8266 7160
rect 9766 7148 9772 7160
rect 9824 7148 9830 7200
rect 17770 7188 17776 7200
rect 17731 7160 17776 7188
rect 17770 7148 17776 7160
rect 17828 7188 17834 7200
rect 20088 7188 20116 7364
rect 20441 7361 20453 7364
rect 20487 7361 20499 7395
rect 20441 7355 20499 7361
rect 20530 7352 20536 7404
rect 20588 7392 20594 7404
rect 20993 7395 21051 7401
rect 20993 7392 21005 7395
rect 20588 7364 21005 7392
rect 20588 7352 20594 7364
rect 20993 7361 21005 7364
rect 21039 7361 21051 7395
rect 20993 7355 21051 7361
rect 20165 7327 20223 7333
rect 20165 7293 20177 7327
rect 20211 7324 20223 7327
rect 20714 7324 20720 7336
rect 20211 7296 20720 7324
rect 20211 7293 20223 7296
rect 20165 7287 20223 7293
rect 20714 7284 20720 7296
rect 20772 7284 20778 7336
rect 20257 7191 20315 7197
rect 20257 7188 20269 7191
rect 17828 7160 20269 7188
rect 17828 7148 17834 7160
rect 20257 7157 20269 7160
rect 20303 7157 20315 7191
rect 20257 7151 20315 7157
rect 1104 7098 21896 7120
rect 1104 7046 3549 7098
rect 3601 7046 3613 7098
rect 3665 7046 3677 7098
rect 3729 7046 3741 7098
rect 3793 7046 3805 7098
rect 3857 7046 8747 7098
rect 8799 7046 8811 7098
rect 8863 7046 8875 7098
rect 8927 7046 8939 7098
rect 8991 7046 9003 7098
rect 9055 7046 13945 7098
rect 13997 7046 14009 7098
rect 14061 7046 14073 7098
rect 14125 7046 14137 7098
rect 14189 7046 14201 7098
rect 14253 7046 19143 7098
rect 19195 7046 19207 7098
rect 19259 7046 19271 7098
rect 19323 7046 19335 7098
rect 19387 7046 19399 7098
rect 19451 7046 21896 7098
rect 1104 7024 21896 7046
rect 4985 6987 5043 6993
rect 4985 6953 4997 6987
rect 5031 6984 5043 6987
rect 5442 6984 5448 6996
rect 5031 6956 5448 6984
rect 5031 6953 5043 6956
rect 4985 6947 5043 6953
rect 5442 6944 5448 6956
rect 5500 6944 5506 6996
rect 9674 6984 9680 6996
rect 9635 6956 9680 6984
rect 9674 6944 9680 6956
rect 9732 6944 9738 6996
rect 9766 6944 9772 6996
rect 9824 6984 9830 6996
rect 17770 6984 17776 6996
rect 9824 6956 17776 6984
rect 9824 6944 9830 6956
rect 17770 6944 17776 6956
rect 17828 6944 17834 6996
rect 1949 6919 2007 6925
rect 1949 6885 1961 6919
rect 1995 6914 2007 6919
rect 1995 6886 2029 6914
rect 1995 6885 2007 6886
rect 1949 6879 2007 6885
rect 1578 6808 1584 6860
rect 1636 6848 1642 6860
rect 1964 6848 1992 6879
rect 2774 6876 2780 6928
rect 2832 6916 2838 6928
rect 3602 6916 3608 6928
rect 2832 6888 3608 6916
rect 2832 6876 2838 6888
rect 3602 6876 3608 6888
rect 3660 6876 3666 6928
rect 5902 6876 5908 6928
rect 5960 6916 5966 6928
rect 20901 6919 20959 6925
rect 20901 6916 20913 6919
rect 5960 6888 9904 6916
rect 5960 6876 5966 6888
rect 9876 6860 9904 6888
rect 12406 6888 12664 6916
rect 1636 6820 1992 6848
rect 1636 6808 1642 6820
rect 2130 6808 2136 6860
rect 2188 6848 2194 6860
rect 2593 6851 2651 6857
rect 2593 6848 2605 6851
rect 2188 6820 2605 6848
rect 2188 6808 2194 6820
rect 2593 6817 2605 6820
rect 2639 6817 2651 6851
rect 2593 6811 2651 6817
rect 2958 6808 2964 6860
rect 3016 6848 3022 6860
rect 3513 6851 3571 6857
rect 3513 6848 3525 6851
rect 3016 6820 3525 6848
rect 3016 6808 3022 6820
rect 3513 6817 3525 6820
rect 3559 6817 3571 6851
rect 3970 6848 3976 6860
rect 3931 6820 3976 6848
rect 3513 6811 3571 6817
rect 1394 6740 1400 6792
rect 1452 6780 1458 6792
rect 1489 6783 1547 6789
rect 1489 6780 1501 6783
rect 1452 6752 1501 6780
rect 1452 6740 1458 6752
rect 1489 6749 1501 6752
rect 1535 6749 1547 6783
rect 1489 6743 1547 6749
rect 1670 6740 1676 6792
rect 1728 6780 1734 6792
rect 1765 6783 1823 6789
rect 1765 6780 1777 6783
rect 1728 6752 1777 6780
rect 1728 6740 1734 6752
rect 1765 6749 1777 6752
rect 1811 6749 1823 6783
rect 1765 6743 1823 6749
rect 2409 6783 2467 6789
rect 2409 6749 2421 6783
rect 2455 6780 2467 6783
rect 3326 6780 3332 6792
rect 2455 6752 3332 6780
rect 2455 6749 2467 6752
rect 2409 6743 2467 6749
rect 1780 6712 1808 6743
rect 3326 6740 3332 6752
rect 3384 6740 3390 6792
rect 3528 6780 3556 6811
rect 3970 6808 3976 6820
rect 4028 6808 4034 6860
rect 4062 6808 4068 6860
rect 4120 6808 4126 6860
rect 4430 6848 4436 6860
rect 4391 6820 4436 6848
rect 4430 6808 4436 6820
rect 4488 6848 4494 6860
rect 5534 6848 5540 6860
rect 4488 6820 5540 6848
rect 4488 6808 4494 6820
rect 5534 6808 5540 6820
rect 5592 6808 5598 6860
rect 5629 6851 5687 6857
rect 5629 6817 5641 6851
rect 5675 6817 5687 6851
rect 5629 6811 5687 6817
rect 3878 6780 3884 6792
rect 3528 6752 3884 6780
rect 3878 6740 3884 6752
rect 3936 6740 3942 6792
rect 4080 6780 4108 6808
rect 3988 6752 4108 6780
rect 4525 6783 4583 6789
rect 3988 6724 4016 6752
rect 4525 6749 4537 6783
rect 4571 6780 4583 6783
rect 4798 6780 4804 6792
rect 4571 6752 4804 6780
rect 4571 6749 4583 6752
rect 4525 6743 4583 6749
rect 4798 6740 4804 6752
rect 4856 6780 4862 6792
rect 4982 6780 4988 6792
rect 4856 6752 4988 6780
rect 4856 6740 4862 6752
rect 4982 6740 4988 6752
rect 5040 6740 5046 6792
rect 5258 6740 5264 6792
rect 5316 6780 5322 6792
rect 5644 6780 5672 6811
rect 5718 6808 5724 6860
rect 5776 6848 5782 6860
rect 6457 6851 6515 6857
rect 6457 6848 6469 6851
rect 5776 6820 6469 6848
rect 5776 6808 5782 6820
rect 6457 6817 6469 6820
rect 6503 6848 6515 6851
rect 8386 6848 8392 6860
rect 6503 6820 8392 6848
rect 6503 6817 6515 6820
rect 6457 6811 6515 6817
rect 8386 6808 8392 6820
rect 8444 6808 8450 6860
rect 8478 6808 8484 6860
rect 8536 6848 8542 6860
rect 9033 6851 9091 6857
rect 9033 6848 9045 6851
rect 8536 6820 9045 6848
rect 8536 6808 8542 6820
rect 9033 6817 9045 6820
rect 9079 6817 9091 6851
rect 9033 6811 9091 6817
rect 9858 6808 9864 6860
rect 9916 6848 9922 6860
rect 10413 6851 10471 6857
rect 10413 6848 10425 6851
rect 9916 6820 10425 6848
rect 9916 6808 9922 6820
rect 10413 6817 10425 6820
rect 10459 6848 10471 6851
rect 12406 6848 12434 6888
rect 12526 6848 12532 6860
rect 10459 6820 12434 6848
rect 12487 6820 12532 6848
rect 10459 6817 10471 6820
rect 10413 6811 10471 6817
rect 12526 6808 12532 6820
rect 12584 6808 12590 6860
rect 12636 6848 12664 6888
rect 20272 6888 20913 6916
rect 15378 6848 15384 6860
rect 12636 6820 15384 6848
rect 15378 6808 15384 6820
rect 15436 6808 15442 6860
rect 18230 6808 18236 6860
rect 18288 6848 18294 6860
rect 20272 6848 20300 6888
rect 20901 6885 20913 6888
rect 20947 6885 20959 6919
rect 20901 6879 20959 6885
rect 18288 6820 20300 6848
rect 20349 6851 20407 6857
rect 18288 6808 18294 6820
rect 20349 6817 20361 6851
rect 20395 6848 20407 6851
rect 20622 6848 20628 6860
rect 20395 6820 20628 6848
rect 20395 6817 20407 6820
rect 20349 6811 20407 6817
rect 20622 6808 20628 6820
rect 20680 6848 20686 6860
rect 21269 6851 21327 6857
rect 20680 6820 21128 6848
rect 20680 6808 20686 6820
rect 6365 6783 6423 6789
rect 6365 6780 6377 6783
rect 5316 6752 5672 6780
rect 5736 6752 6377 6780
rect 5316 6740 5322 6752
rect 3789 6715 3847 6721
rect 3789 6712 3801 6715
rect 1780 6684 3801 6712
rect 3789 6681 3801 6684
rect 3835 6681 3847 6715
rect 3789 6675 3847 6681
rect 3970 6672 3976 6724
rect 4028 6672 4034 6724
rect 4062 6672 4068 6724
rect 4120 6712 4126 6724
rect 5445 6715 5503 6721
rect 5445 6712 5457 6715
rect 4120 6684 5457 6712
rect 4120 6672 4126 6684
rect 5445 6681 5457 6684
rect 5491 6712 5503 6715
rect 5736 6712 5764 6752
rect 6365 6749 6377 6752
rect 6411 6749 6423 6783
rect 16942 6780 16948 6792
rect 6365 6743 6423 6749
rect 12406 6752 16948 6780
rect 5491 6684 5764 6712
rect 6273 6715 6331 6721
rect 5491 6681 5503 6684
rect 5445 6675 5503 6681
rect 6273 6681 6285 6715
rect 6319 6712 6331 6715
rect 6733 6715 6791 6721
rect 6733 6712 6745 6715
rect 6319 6684 6745 6712
rect 6319 6681 6331 6684
rect 6273 6675 6331 6681
rect 6733 6681 6745 6684
rect 6779 6681 6791 6715
rect 9769 6715 9827 6721
rect 9769 6712 9781 6715
rect 6733 6675 6791 6681
rect 9232 6684 9781 6712
rect 9232 6656 9260 6684
rect 9769 6681 9781 6684
rect 9815 6712 9827 6715
rect 12406 6712 12434 6752
rect 16942 6740 16948 6752
rect 17000 6740 17006 6792
rect 20533 6783 20591 6789
rect 20533 6749 20545 6783
rect 20579 6780 20591 6783
rect 20806 6780 20812 6792
rect 20579 6752 20812 6780
rect 20579 6749 20591 6752
rect 20533 6743 20591 6749
rect 20806 6740 20812 6752
rect 20864 6740 20870 6792
rect 21100 6789 21128 6820
rect 21269 6817 21281 6851
rect 21315 6848 21327 6851
rect 22370 6848 22376 6860
rect 21315 6820 22376 6848
rect 21315 6817 21327 6820
rect 21269 6811 21327 6817
rect 22370 6808 22376 6820
rect 22428 6808 22434 6860
rect 21085 6783 21143 6789
rect 21085 6749 21097 6783
rect 21131 6749 21143 6783
rect 21450 6780 21456 6792
rect 21411 6752 21456 6780
rect 21085 6743 21143 6749
rect 21450 6740 21456 6752
rect 21508 6740 21514 6792
rect 9815 6684 12434 6712
rect 12805 6715 12863 6721
rect 9815 6681 9827 6684
rect 9769 6675 9827 6681
rect 12805 6681 12817 6715
rect 12851 6712 12863 6715
rect 13265 6715 13323 6721
rect 13265 6712 13277 6715
rect 12851 6684 13277 6712
rect 12851 6681 12863 6684
rect 12805 6675 12863 6681
rect 13265 6681 13277 6684
rect 13311 6681 13323 6715
rect 13265 6675 13323 6681
rect 14642 6672 14648 6724
rect 14700 6712 14706 6724
rect 18506 6712 18512 6724
rect 14700 6684 18512 6712
rect 14700 6672 14706 6684
rect 18506 6672 18512 6684
rect 18564 6672 18570 6724
rect 20165 6715 20223 6721
rect 20165 6681 20177 6715
rect 20211 6712 20223 6715
rect 21468 6712 21496 6740
rect 20211 6684 21496 6712
rect 20211 6681 20223 6684
rect 20165 6675 20223 6681
rect 1578 6644 1584 6656
rect 1539 6616 1584 6644
rect 1578 6604 1584 6616
rect 1636 6604 1642 6656
rect 2038 6644 2044 6656
rect 1999 6616 2044 6644
rect 2038 6604 2044 6616
rect 2096 6604 2102 6656
rect 2130 6604 2136 6656
rect 2188 6644 2194 6656
rect 2501 6647 2559 6653
rect 2501 6644 2513 6647
rect 2188 6616 2513 6644
rect 2188 6604 2194 6616
rect 2501 6613 2513 6616
rect 2547 6644 2559 6647
rect 2590 6644 2596 6656
rect 2547 6616 2596 6644
rect 2547 6613 2559 6616
rect 2501 6607 2559 6613
rect 2590 6604 2596 6616
rect 2648 6604 2654 6656
rect 2866 6644 2872 6656
rect 2827 6616 2872 6644
rect 2866 6604 2872 6616
rect 2924 6604 2930 6656
rect 3234 6644 3240 6656
rect 3195 6616 3240 6644
rect 3234 6604 3240 6616
rect 3292 6604 3298 6656
rect 3329 6647 3387 6653
rect 3329 6613 3341 6647
rect 3375 6644 3387 6647
rect 3510 6644 3516 6656
rect 3375 6616 3516 6644
rect 3375 6613 3387 6616
rect 3329 6607 3387 6613
rect 3510 6604 3516 6616
rect 3568 6604 3574 6656
rect 4614 6604 4620 6656
rect 4672 6644 4678 6656
rect 4672 6616 4717 6644
rect 4672 6604 4678 6616
rect 4890 6604 4896 6656
rect 4948 6644 4954 6656
rect 5077 6647 5135 6653
rect 5077 6644 5089 6647
rect 4948 6616 5089 6644
rect 4948 6604 4954 6616
rect 5077 6613 5089 6616
rect 5123 6613 5135 6647
rect 5077 6607 5135 6613
rect 5258 6604 5264 6656
rect 5316 6644 5322 6656
rect 5537 6647 5595 6653
rect 5537 6644 5549 6647
rect 5316 6616 5549 6644
rect 5316 6604 5322 6616
rect 5537 6613 5549 6616
rect 5583 6613 5595 6647
rect 5902 6644 5908 6656
rect 5863 6616 5908 6644
rect 5537 6607 5595 6613
rect 5902 6604 5908 6616
rect 5960 6604 5966 6656
rect 9214 6644 9220 6656
rect 9175 6616 9220 6644
rect 9214 6604 9220 6616
rect 9272 6604 9278 6656
rect 9306 6604 9312 6656
rect 9364 6644 9370 6656
rect 12710 6644 12716 6656
rect 9364 6616 9409 6644
rect 12671 6616 12716 6644
rect 9364 6604 9370 6616
rect 12710 6604 12716 6616
rect 12768 6604 12774 6656
rect 13173 6647 13231 6653
rect 13173 6613 13185 6647
rect 13219 6644 13231 6647
rect 19794 6644 19800 6656
rect 13219 6616 19800 6644
rect 13219 6613 13231 6616
rect 13173 6607 13231 6613
rect 19794 6604 19800 6616
rect 19852 6604 19858 6656
rect 20622 6644 20628 6656
rect 20583 6616 20628 6644
rect 20622 6604 20628 6616
rect 20680 6604 20686 6656
rect 1104 6554 22056 6576
rect 1104 6502 6148 6554
rect 6200 6502 6212 6554
rect 6264 6502 6276 6554
rect 6328 6502 6340 6554
rect 6392 6502 6404 6554
rect 6456 6502 11346 6554
rect 11398 6502 11410 6554
rect 11462 6502 11474 6554
rect 11526 6502 11538 6554
rect 11590 6502 11602 6554
rect 11654 6502 16544 6554
rect 16596 6502 16608 6554
rect 16660 6502 16672 6554
rect 16724 6502 16736 6554
rect 16788 6502 16800 6554
rect 16852 6502 21742 6554
rect 21794 6502 21806 6554
rect 21858 6502 21870 6554
rect 21922 6502 21934 6554
rect 21986 6502 21998 6554
rect 22050 6502 22056 6554
rect 1104 6480 22056 6502
rect 2222 6400 2228 6452
rect 2280 6440 2286 6452
rect 2593 6443 2651 6449
rect 2593 6440 2605 6443
rect 2280 6412 2605 6440
rect 2280 6400 2286 6412
rect 2593 6409 2605 6412
rect 2639 6409 2651 6443
rect 2593 6403 2651 6409
rect 3145 6443 3203 6449
rect 3145 6409 3157 6443
rect 3191 6440 3203 6443
rect 3326 6440 3332 6452
rect 3191 6412 3332 6440
rect 3191 6409 3203 6412
rect 3145 6403 3203 6409
rect 3326 6400 3332 6412
rect 3384 6400 3390 6452
rect 3510 6440 3516 6452
rect 3471 6412 3516 6440
rect 3510 6400 3516 6412
rect 3568 6400 3574 6452
rect 4706 6400 4712 6452
rect 4764 6440 4770 6452
rect 4893 6443 4951 6449
rect 4893 6440 4905 6443
rect 4764 6412 4905 6440
rect 4764 6400 4770 6412
rect 4893 6409 4905 6412
rect 4939 6409 4951 6443
rect 4893 6403 4951 6409
rect 5261 6443 5319 6449
rect 5261 6409 5273 6443
rect 5307 6440 5319 6443
rect 5902 6440 5908 6452
rect 5307 6412 5908 6440
rect 5307 6409 5319 6412
rect 5261 6403 5319 6409
rect 5902 6400 5908 6412
rect 5960 6400 5966 6452
rect 11701 6443 11759 6449
rect 11701 6409 11713 6443
rect 11747 6440 11759 6443
rect 11974 6440 11980 6452
rect 11747 6412 11980 6440
rect 11747 6409 11759 6412
rect 11701 6403 11759 6409
rect 11974 6400 11980 6412
rect 12032 6400 12038 6452
rect 12710 6440 12716 6452
rect 12671 6412 12716 6440
rect 12710 6400 12716 6412
rect 12768 6400 12774 6452
rect 14185 6443 14243 6449
rect 14185 6409 14197 6443
rect 14231 6409 14243 6443
rect 14642 6440 14648 6452
rect 14603 6412 14648 6440
rect 14185 6403 14243 6409
rect 2958 6332 2964 6384
rect 3016 6372 3022 6384
rect 3053 6375 3111 6381
rect 3053 6372 3065 6375
rect 3016 6344 3065 6372
rect 3016 6332 3022 6344
rect 3053 6341 3065 6344
rect 3099 6341 3111 6375
rect 3053 6335 3111 6341
rect 3602 6332 3608 6384
rect 3660 6372 3666 6384
rect 3973 6375 4031 6381
rect 3973 6372 3985 6375
rect 3660 6344 3985 6372
rect 3660 6332 3666 6344
rect 3973 6341 3985 6344
rect 4019 6341 4031 6375
rect 3973 6335 4031 6341
rect 4522 6332 4528 6384
rect 4580 6372 4586 6384
rect 9214 6372 9220 6384
rect 4580 6344 9220 6372
rect 4580 6332 4586 6344
rect 9214 6332 9220 6344
rect 9272 6332 9278 6384
rect 12069 6375 12127 6381
rect 12069 6341 12081 6375
rect 12115 6372 12127 6375
rect 14200 6372 14228 6403
rect 14642 6400 14648 6412
rect 14700 6400 14706 6452
rect 15473 6443 15531 6449
rect 15473 6409 15485 6443
rect 15519 6440 15531 6443
rect 20622 6440 20628 6452
rect 15519 6412 20628 6440
rect 15519 6409 15531 6412
rect 15473 6403 15531 6409
rect 20622 6400 20628 6412
rect 20680 6400 20686 6452
rect 15378 6372 15384 6384
rect 12115 6344 14228 6372
rect 14384 6344 14780 6372
rect 15291 6344 15384 6372
rect 12115 6341 12127 6344
rect 12069 6335 12127 6341
rect 2590 6264 2596 6316
rect 2648 6304 2654 6316
rect 2774 6304 2780 6316
rect 2648 6276 2780 6304
rect 2648 6264 2654 6276
rect 2774 6264 2780 6276
rect 2832 6264 2838 6316
rect 3326 6304 3332 6316
rect 3160 6276 3332 6304
rect 3160 6248 3188 6276
rect 3326 6264 3332 6276
rect 3384 6304 3390 6316
rect 3384 6276 4200 6304
rect 3384 6264 3390 6276
rect 1949 6239 2007 6245
rect 1949 6205 1961 6239
rect 1995 6205 2007 6239
rect 2222 6236 2228 6248
rect 2183 6208 2228 6236
rect 1949 6199 2007 6205
rect 1964 6168 1992 6199
rect 2222 6196 2228 6208
rect 2280 6196 2286 6248
rect 2314 6196 2320 6248
rect 2372 6236 2378 6248
rect 2961 6239 3019 6245
rect 2372 6208 2417 6236
rect 2372 6196 2378 6208
rect 2961 6205 2973 6239
rect 3007 6236 3019 6239
rect 3142 6236 3148 6248
rect 3007 6208 3148 6236
rect 3007 6205 3019 6208
rect 2961 6199 3019 6205
rect 3142 6196 3148 6208
rect 3200 6196 3206 6248
rect 4062 6236 4068 6248
rect 4023 6208 4068 6236
rect 4062 6196 4068 6208
rect 4120 6196 4126 6248
rect 4172 6245 4200 6276
rect 4798 6264 4804 6316
rect 4856 6304 4862 6316
rect 4856 6276 5856 6304
rect 4856 6264 4862 6276
rect 4157 6239 4215 6245
rect 4157 6205 4169 6239
rect 4203 6205 4215 6239
rect 5350 6236 5356 6248
rect 5311 6208 5356 6236
rect 4157 6199 4215 6205
rect 5350 6196 5356 6208
rect 5408 6196 5414 6248
rect 5442 6196 5448 6248
rect 5500 6236 5506 6248
rect 5828 6245 5856 6276
rect 10502 6264 10508 6316
rect 10560 6304 10566 6316
rect 13078 6304 13084 6316
rect 10560 6276 12296 6304
rect 13039 6276 13084 6304
rect 10560 6264 10566 6276
rect 5813 6239 5871 6245
rect 5500 6208 5545 6236
rect 5500 6196 5506 6208
rect 5813 6205 5825 6239
rect 5859 6236 5871 6239
rect 5902 6236 5908 6248
rect 5859 6208 5908 6236
rect 5859 6205 5871 6208
rect 5813 6199 5871 6205
rect 5902 6196 5908 6208
rect 5960 6196 5966 6248
rect 12268 6245 12296 6276
rect 13078 6264 13084 6276
rect 13136 6264 13142 6316
rect 13722 6264 13728 6316
rect 13780 6304 13786 6316
rect 14384 6304 14412 6344
rect 14550 6304 14556 6316
rect 13780 6276 14412 6304
rect 14511 6276 14556 6304
rect 13780 6264 13786 6276
rect 14550 6264 14556 6276
rect 14608 6264 14614 6316
rect 12161 6239 12219 6245
rect 12161 6205 12173 6239
rect 12207 6205 12219 6239
rect 12161 6199 12219 6205
rect 12253 6239 12311 6245
rect 12253 6205 12265 6239
rect 12299 6205 12311 6239
rect 13170 6236 13176 6248
rect 13131 6208 13176 6236
rect 12253 6199 12311 6205
rect 8202 6168 8208 6180
rect 1964 6140 8208 6168
rect 8202 6128 8208 6140
rect 8260 6128 8266 6180
rect 12176 6168 12204 6199
rect 13170 6196 13176 6208
rect 13228 6196 13234 6248
rect 13354 6236 13360 6248
rect 13315 6208 13360 6236
rect 13354 6196 13360 6208
rect 13412 6196 13418 6248
rect 14090 6236 14096 6248
rect 14003 6208 14096 6236
rect 14090 6196 14096 6208
rect 14148 6236 14154 6248
rect 14642 6236 14648 6248
rect 14148 6208 14648 6236
rect 14148 6196 14154 6208
rect 14642 6196 14648 6208
rect 14700 6196 14706 6248
rect 14752 6245 14780 6344
rect 15378 6332 15384 6344
rect 15436 6372 15442 6384
rect 15933 6375 15991 6381
rect 15933 6372 15945 6375
rect 15436 6344 15945 6372
rect 15436 6332 15442 6344
rect 15933 6341 15945 6344
rect 15979 6372 15991 6375
rect 20530 6372 20536 6384
rect 15979 6344 20536 6372
rect 15979 6341 15991 6344
rect 15933 6335 15991 6341
rect 20530 6332 20536 6344
rect 20588 6332 20594 6384
rect 16942 6264 16948 6316
rect 17000 6304 17006 6316
rect 20993 6307 21051 6313
rect 20993 6304 21005 6307
rect 17000 6276 21005 6304
rect 17000 6264 17006 6276
rect 20993 6273 21005 6276
rect 21039 6273 21051 6307
rect 20993 6267 21051 6273
rect 14737 6239 14795 6245
rect 14737 6205 14749 6239
rect 14783 6236 14795 6239
rect 15565 6239 15623 6245
rect 15565 6236 15577 6239
rect 14783 6208 15577 6236
rect 14783 6205 14795 6208
rect 14737 6199 14795 6205
rect 15565 6205 15577 6208
rect 15611 6205 15623 6239
rect 15565 6199 15623 6205
rect 20625 6239 20683 6245
rect 20625 6205 20637 6239
rect 20671 6236 20683 6239
rect 20714 6236 20720 6248
rect 20671 6208 20720 6236
rect 20671 6205 20683 6208
rect 20625 6199 20683 6205
rect 20714 6196 20720 6208
rect 20772 6196 20778 6248
rect 15013 6171 15071 6177
rect 15013 6168 15025 6171
rect 12176 6140 15025 6168
rect 15013 6137 15025 6140
rect 15059 6137 15071 6171
rect 15013 6131 15071 6137
rect 3142 6060 3148 6112
rect 3200 6100 3206 6112
rect 3605 6103 3663 6109
rect 3605 6100 3617 6103
rect 3200 6072 3617 6100
rect 3200 6060 3206 6072
rect 3605 6069 3617 6072
rect 3651 6069 3663 6103
rect 3605 6063 3663 6069
rect 1104 6010 21896 6032
rect 1104 5958 3549 6010
rect 3601 5958 3613 6010
rect 3665 5958 3677 6010
rect 3729 5958 3741 6010
rect 3793 5958 3805 6010
rect 3857 5958 8747 6010
rect 8799 5958 8811 6010
rect 8863 5958 8875 6010
rect 8927 5958 8939 6010
rect 8991 5958 9003 6010
rect 9055 5958 13945 6010
rect 13997 5958 14009 6010
rect 14061 5958 14073 6010
rect 14125 5958 14137 6010
rect 14189 5958 14201 6010
rect 14253 5958 19143 6010
rect 19195 5958 19207 6010
rect 19259 5958 19271 6010
rect 19323 5958 19335 6010
rect 19387 5958 19399 6010
rect 19451 5958 21896 6010
rect 1104 5936 21896 5958
rect 1762 5896 1768 5908
rect 1723 5868 1768 5896
rect 1762 5856 1768 5868
rect 1820 5856 1826 5908
rect 3234 5856 3240 5908
rect 3292 5896 3298 5908
rect 3329 5899 3387 5905
rect 3329 5896 3341 5899
rect 3292 5868 3341 5896
rect 3292 5856 3298 5868
rect 3329 5865 3341 5868
rect 3375 5865 3387 5899
rect 5350 5896 5356 5908
rect 5311 5868 5356 5896
rect 3329 5859 3387 5865
rect 5350 5856 5356 5868
rect 5408 5856 5414 5908
rect 13170 5856 13176 5908
rect 13228 5896 13234 5908
rect 21085 5899 21143 5905
rect 21085 5896 21097 5899
rect 13228 5868 21097 5896
rect 13228 5856 13234 5868
rect 21085 5865 21097 5868
rect 21131 5865 21143 5899
rect 21085 5859 21143 5865
rect 2866 5828 2872 5840
rect 2608 5800 2872 5828
rect 2406 5760 2412 5772
rect 2367 5732 2412 5760
rect 2406 5720 2412 5732
rect 2464 5720 2470 5772
rect 1394 5692 1400 5704
rect 1355 5664 1400 5692
rect 1394 5652 1400 5664
rect 1452 5652 1458 5704
rect 2225 5627 2283 5633
rect 2225 5593 2237 5627
rect 2271 5624 2283 5627
rect 2608 5624 2636 5800
rect 2866 5788 2872 5800
rect 2924 5788 2930 5840
rect 2777 5763 2835 5769
rect 2777 5729 2789 5763
rect 2823 5760 2835 5763
rect 2823 5732 3096 5760
rect 2823 5729 2835 5732
rect 2777 5723 2835 5729
rect 2271 5596 2636 5624
rect 2271 5593 2283 5596
rect 2225 5587 2283 5593
rect 2682 5584 2688 5636
rect 2740 5624 2746 5636
rect 2961 5627 3019 5633
rect 2961 5624 2973 5627
rect 2740 5596 2973 5624
rect 2740 5584 2746 5596
rect 2961 5593 2973 5596
rect 3007 5593 3019 5627
rect 3068 5624 3096 5732
rect 4430 5720 4436 5772
rect 4488 5760 4494 5772
rect 4709 5763 4767 5769
rect 4709 5760 4721 5763
rect 4488 5732 4721 5760
rect 4488 5720 4494 5732
rect 4709 5729 4721 5732
rect 4755 5729 4767 5763
rect 14550 5760 14556 5772
rect 14511 5732 14556 5760
rect 4709 5723 4767 5729
rect 14550 5720 14556 5732
rect 14608 5720 14614 5772
rect 20809 5763 20867 5769
rect 20809 5729 20821 5763
rect 20855 5760 20867 5763
rect 20855 5732 21588 5760
rect 20855 5729 20867 5732
rect 20809 5723 20867 5729
rect 21560 5704 21588 5732
rect 20993 5695 21051 5701
rect 20993 5661 21005 5695
rect 21039 5692 21051 5695
rect 21266 5692 21272 5704
rect 21039 5664 21272 5692
rect 21039 5661 21051 5664
rect 20993 5655 21051 5661
rect 21266 5652 21272 5664
rect 21324 5652 21330 5704
rect 21542 5692 21548 5704
rect 21503 5664 21548 5692
rect 21542 5652 21548 5664
rect 21600 5652 21606 5704
rect 3326 5624 3332 5636
rect 3068 5596 3332 5624
rect 2961 5587 3019 5593
rect 3326 5584 3332 5596
rect 3384 5584 3390 5636
rect 3510 5584 3516 5636
rect 3568 5624 3574 5636
rect 4893 5627 4951 5633
rect 4893 5624 4905 5627
rect 3568 5596 4905 5624
rect 3568 5584 3574 5596
rect 4893 5593 4905 5596
rect 4939 5624 4951 5627
rect 5258 5624 5264 5636
rect 4939 5596 5264 5624
rect 4939 5593 4951 5596
rect 4893 5587 4951 5593
rect 5258 5584 5264 5596
rect 5316 5584 5322 5636
rect 10962 5584 10968 5636
rect 11020 5624 11026 5636
rect 11020 5596 21404 5624
rect 11020 5584 11026 5596
rect 1578 5556 1584 5568
rect 1539 5528 1584 5556
rect 1578 5516 1584 5528
rect 1636 5516 1642 5568
rect 2130 5556 2136 5568
rect 2091 5528 2136 5556
rect 2130 5516 2136 5528
rect 2188 5516 2194 5568
rect 2866 5556 2872 5568
rect 2779 5528 2872 5556
rect 2866 5516 2872 5528
rect 2924 5556 2930 5568
rect 3970 5556 3976 5568
rect 2924 5528 3976 5556
rect 2924 5516 2930 5528
rect 3970 5516 3976 5528
rect 4028 5556 4034 5568
rect 21376 5565 21404 5596
rect 4985 5559 5043 5565
rect 4985 5556 4997 5559
rect 4028 5528 4997 5556
rect 4028 5516 4034 5528
rect 4985 5525 4997 5528
rect 5031 5525 5043 5559
rect 4985 5519 5043 5525
rect 21361 5559 21419 5565
rect 21361 5525 21373 5559
rect 21407 5525 21419 5559
rect 21361 5519 21419 5525
rect 1104 5466 22056 5488
rect 1104 5414 6148 5466
rect 6200 5414 6212 5466
rect 6264 5414 6276 5466
rect 6328 5414 6340 5466
rect 6392 5414 6404 5466
rect 6456 5414 11346 5466
rect 11398 5414 11410 5466
rect 11462 5414 11474 5466
rect 11526 5414 11538 5466
rect 11590 5414 11602 5466
rect 11654 5414 16544 5466
rect 16596 5414 16608 5466
rect 16660 5414 16672 5466
rect 16724 5414 16736 5466
rect 16788 5414 16800 5466
rect 16852 5414 21742 5466
rect 21794 5414 21806 5466
rect 21858 5414 21870 5466
rect 21922 5414 21934 5466
rect 21986 5414 21998 5466
rect 22050 5414 22056 5466
rect 1104 5392 22056 5414
rect 1581 5355 1639 5361
rect 1581 5321 1593 5355
rect 1627 5352 1639 5355
rect 1670 5352 1676 5364
rect 1627 5324 1676 5352
rect 1627 5321 1639 5324
rect 1581 5315 1639 5321
rect 1670 5312 1676 5324
rect 1728 5312 1734 5364
rect 2130 5312 2136 5364
rect 2188 5352 2194 5364
rect 2409 5355 2467 5361
rect 2409 5352 2421 5355
rect 2188 5324 2421 5352
rect 2188 5312 2194 5324
rect 2409 5321 2421 5324
rect 2455 5321 2467 5355
rect 2409 5315 2467 5321
rect 2774 5312 2780 5364
rect 2832 5352 2838 5364
rect 2832 5324 2877 5352
rect 2832 5312 2838 5324
rect 2958 5312 2964 5364
rect 3016 5352 3022 5364
rect 3510 5352 3516 5364
rect 3016 5324 3516 5352
rect 3016 5312 3022 5324
rect 3510 5312 3516 5324
rect 3568 5312 3574 5364
rect 18414 5312 18420 5364
rect 18472 5352 18478 5364
rect 21361 5355 21419 5361
rect 21361 5352 21373 5355
rect 18472 5324 21373 5352
rect 18472 5312 18478 5324
rect 21361 5321 21373 5324
rect 21407 5321 21419 5355
rect 21361 5315 21419 5321
rect 2041 5287 2099 5293
rect 2041 5253 2053 5287
rect 2087 5284 2099 5287
rect 2314 5284 2320 5296
rect 2087 5256 2320 5284
rect 2087 5253 2099 5256
rect 2041 5247 2099 5253
rect 2314 5244 2320 5256
rect 2372 5244 2378 5296
rect 1394 5216 1400 5228
rect 1355 5188 1400 5216
rect 1394 5176 1400 5188
rect 1452 5216 1458 5228
rect 2869 5219 2927 5225
rect 2869 5216 2881 5219
rect 1452 5188 2881 5216
rect 1452 5176 1458 5188
rect 2869 5185 2881 5188
rect 2915 5185 2927 5219
rect 2869 5179 2927 5185
rect 21269 5219 21327 5225
rect 21269 5185 21281 5219
rect 21315 5216 21327 5219
rect 21542 5216 21548 5228
rect 21315 5188 21548 5216
rect 21315 5185 21327 5188
rect 21269 5179 21327 5185
rect 21542 5176 21548 5188
rect 21600 5176 21606 5228
rect 1857 5151 1915 5157
rect 1857 5117 1869 5151
rect 1903 5117 1915 5151
rect 1857 5111 1915 5117
rect 1949 5151 2007 5157
rect 1949 5117 1961 5151
rect 1995 5148 2007 5151
rect 3142 5148 3148 5160
rect 1995 5120 3148 5148
rect 1995 5117 2007 5120
rect 1949 5111 2007 5117
rect 1872 5012 1900 5111
rect 3142 5108 3148 5120
rect 3200 5108 3206 5160
rect 2222 5040 2228 5092
rect 2280 5080 2286 5092
rect 2501 5083 2559 5089
rect 2501 5080 2513 5083
rect 2280 5052 2513 5080
rect 2280 5040 2286 5052
rect 2501 5049 2513 5052
rect 2547 5049 2559 5083
rect 2501 5043 2559 5049
rect 3878 5012 3884 5024
rect 1872 4984 3884 5012
rect 3878 4972 3884 4984
rect 3936 4972 3942 5024
rect 1104 4922 21896 4944
rect 1104 4870 3549 4922
rect 3601 4870 3613 4922
rect 3665 4870 3677 4922
rect 3729 4870 3741 4922
rect 3793 4870 3805 4922
rect 3857 4870 8747 4922
rect 8799 4870 8811 4922
rect 8863 4870 8875 4922
rect 8927 4870 8939 4922
rect 8991 4870 9003 4922
rect 9055 4870 13945 4922
rect 13997 4870 14009 4922
rect 14061 4870 14073 4922
rect 14125 4870 14137 4922
rect 14189 4870 14201 4922
rect 14253 4870 19143 4922
rect 19195 4870 19207 4922
rect 19259 4870 19271 4922
rect 19323 4870 19335 4922
rect 19387 4870 19399 4922
rect 19451 4870 21896 4922
rect 1104 4848 21896 4870
rect 1581 4811 1639 4817
rect 1581 4777 1593 4811
rect 1627 4808 1639 4811
rect 2038 4808 2044 4820
rect 1627 4780 2044 4808
rect 1627 4777 1639 4780
rect 1581 4771 1639 4777
rect 2038 4768 2044 4780
rect 2096 4768 2102 4820
rect 2133 4811 2191 4817
rect 2133 4777 2145 4811
rect 2179 4808 2191 4811
rect 2682 4808 2688 4820
rect 2179 4780 2688 4808
rect 2179 4777 2191 4780
rect 2133 4771 2191 4777
rect 2682 4768 2688 4780
rect 2740 4768 2746 4820
rect 1857 4743 1915 4749
rect 1857 4709 1869 4743
rect 1903 4740 1915 4743
rect 4062 4740 4068 4752
rect 1903 4712 4068 4740
rect 1903 4709 1915 4712
rect 1857 4703 1915 4709
rect 4062 4700 4068 4712
rect 4120 4700 4126 4752
rect 20990 4672 20996 4684
rect 20951 4644 20996 4672
rect 20990 4632 20996 4644
rect 21048 4632 21054 4684
rect 1394 4604 1400 4616
rect 1355 4576 1400 4604
rect 1394 4564 1400 4576
rect 1452 4564 1458 4616
rect 1670 4604 1676 4616
rect 1631 4576 1676 4604
rect 1670 4564 1676 4576
rect 1728 4564 1734 4616
rect 1946 4604 1952 4616
rect 1907 4576 1952 4604
rect 1946 4564 1952 4576
rect 2004 4604 2010 4616
rect 2225 4607 2283 4613
rect 2225 4604 2237 4607
rect 2004 4576 2237 4604
rect 2004 4564 2010 4576
rect 2225 4573 2237 4576
rect 2271 4573 2283 4607
rect 2225 4567 2283 4573
rect 20625 4607 20683 4613
rect 20625 4573 20637 4607
rect 20671 4604 20683 4607
rect 20714 4604 20720 4616
rect 20671 4576 20720 4604
rect 20671 4573 20683 4576
rect 20625 4567 20683 4573
rect 20714 4564 20720 4576
rect 20772 4564 20778 4616
rect 1104 4378 22056 4400
rect 1104 4326 6148 4378
rect 6200 4326 6212 4378
rect 6264 4326 6276 4378
rect 6328 4326 6340 4378
rect 6392 4326 6404 4378
rect 6456 4326 11346 4378
rect 11398 4326 11410 4378
rect 11462 4326 11474 4378
rect 11526 4326 11538 4378
rect 11590 4326 11602 4378
rect 11654 4326 16544 4378
rect 16596 4326 16608 4378
rect 16660 4326 16672 4378
rect 16724 4326 16736 4378
rect 16788 4326 16800 4378
rect 16852 4326 21742 4378
rect 21794 4326 21806 4378
rect 21858 4326 21870 4378
rect 21922 4326 21934 4378
rect 21986 4326 21998 4378
rect 22050 4326 22056 4378
rect 1104 4304 22056 4326
rect 1394 4224 1400 4276
rect 1452 4224 1458 4276
rect 1670 4264 1676 4276
rect 1631 4236 1676 4264
rect 1670 4224 1676 4236
rect 1728 4224 1734 4276
rect 21082 4264 21088 4276
rect 21043 4236 21088 4264
rect 21082 4224 21088 4236
rect 21140 4224 21146 4276
rect 1412 4196 1440 4224
rect 1857 4199 1915 4205
rect 1857 4196 1869 4199
rect 1412 4168 1869 4196
rect 1857 4165 1869 4168
rect 1903 4165 1915 4199
rect 1857 4159 1915 4165
rect 1394 4128 1400 4140
rect 1355 4100 1400 4128
rect 1394 4088 1400 4100
rect 1452 4128 1458 4140
rect 2041 4131 2099 4137
rect 2041 4128 2053 4131
rect 1452 4100 2053 4128
rect 1452 4088 1458 4100
rect 2041 4097 2053 4100
rect 2087 4097 2099 4131
rect 2041 4091 2099 4097
rect 20993 4131 21051 4137
rect 20993 4097 21005 4131
rect 21039 4128 21051 4131
rect 21266 4128 21272 4140
rect 21039 4100 21272 4128
rect 21039 4097 21051 4100
rect 20993 4091 21051 4097
rect 21266 4088 21272 4100
rect 21324 4088 21330 4140
rect 21542 4128 21548 4140
rect 21503 4100 21548 4128
rect 21542 4088 21548 4100
rect 21600 4088 21606 4140
rect 20809 4063 20867 4069
rect 20809 4029 20821 4063
rect 20855 4060 20867 4063
rect 21560 4060 21588 4088
rect 20855 4032 21588 4060
rect 20855 4029 20867 4032
rect 20809 4023 20867 4029
rect 1581 3995 1639 4001
rect 1581 3961 1593 3995
rect 1627 3992 1639 3995
rect 2866 3992 2872 4004
rect 1627 3964 2872 3992
rect 1627 3961 1639 3964
rect 1581 3955 1639 3961
rect 2866 3952 2872 3964
rect 2924 3952 2930 4004
rect 18322 3952 18328 4004
rect 18380 3992 18386 4004
rect 21361 3995 21419 4001
rect 21361 3992 21373 3995
rect 18380 3964 21373 3992
rect 18380 3952 18386 3964
rect 21361 3961 21373 3964
rect 21407 3961 21419 3995
rect 21361 3955 21419 3961
rect 1104 3834 21896 3856
rect 1104 3782 3549 3834
rect 3601 3782 3613 3834
rect 3665 3782 3677 3834
rect 3729 3782 3741 3834
rect 3793 3782 3805 3834
rect 3857 3782 8747 3834
rect 8799 3782 8811 3834
rect 8863 3782 8875 3834
rect 8927 3782 8939 3834
rect 8991 3782 9003 3834
rect 9055 3782 13945 3834
rect 13997 3782 14009 3834
rect 14061 3782 14073 3834
rect 14125 3782 14137 3834
rect 14189 3782 14201 3834
rect 14253 3782 19143 3834
rect 19195 3782 19207 3834
rect 19259 3782 19271 3834
rect 19323 3782 19335 3834
rect 19387 3782 19399 3834
rect 19451 3782 21896 3834
rect 1104 3760 21896 3782
rect 1581 3723 1639 3729
rect 1581 3689 1593 3723
rect 1627 3720 1639 3723
rect 3050 3720 3056 3732
rect 1627 3692 3056 3720
rect 1627 3689 1639 3692
rect 1581 3683 1639 3689
rect 3050 3680 3056 3692
rect 3108 3680 3114 3732
rect 20346 3680 20352 3732
rect 20404 3720 20410 3732
rect 21361 3723 21419 3729
rect 21361 3720 21373 3723
rect 20404 3692 21373 3720
rect 20404 3680 20410 3692
rect 21361 3689 21373 3692
rect 21407 3689 21419 3723
rect 21361 3683 21419 3689
rect 1394 3516 1400 3528
rect 1355 3488 1400 3516
rect 1394 3476 1400 3488
rect 1452 3516 1458 3528
rect 1673 3519 1731 3525
rect 1673 3516 1685 3519
rect 1452 3488 1685 3516
rect 1452 3476 1458 3488
rect 1673 3485 1685 3488
rect 1719 3485 1731 3519
rect 1673 3479 1731 3485
rect 21269 3519 21327 3525
rect 21269 3485 21281 3519
rect 21315 3516 21327 3519
rect 21542 3516 21548 3528
rect 21315 3488 21548 3516
rect 21315 3485 21327 3488
rect 21269 3479 21327 3485
rect 21542 3476 21548 3488
rect 21600 3476 21606 3528
rect 1670 3340 1676 3392
rect 1728 3380 1734 3392
rect 1857 3383 1915 3389
rect 1857 3380 1869 3383
rect 1728 3352 1869 3380
rect 1728 3340 1734 3352
rect 1857 3349 1869 3352
rect 1903 3349 1915 3383
rect 1857 3343 1915 3349
rect 1104 3290 22056 3312
rect 1104 3238 6148 3290
rect 6200 3238 6212 3290
rect 6264 3238 6276 3290
rect 6328 3238 6340 3290
rect 6392 3238 6404 3290
rect 6456 3238 11346 3290
rect 11398 3238 11410 3290
rect 11462 3238 11474 3290
rect 11526 3238 11538 3290
rect 11590 3238 11602 3290
rect 11654 3238 16544 3290
rect 16596 3238 16608 3290
rect 16660 3238 16672 3290
rect 16724 3238 16736 3290
rect 16788 3238 16800 3290
rect 16852 3238 21742 3290
rect 21794 3238 21806 3290
rect 21858 3238 21870 3290
rect 21922 3238 21934 3290
rect 21986 3238 21998 3290
rect 22050 3238 22056 3290
rect 1104 3216 22056 3238
rect 1581 3179 1639 3185
rect 1581 3145 1593 3179
rect 1627 3145 1639 3179
rect 1854 3176 1860 3188
rect 1815 3148 1860 3176
rect 1581 3139 1639 3145
rect 1596 3108 1624 3139
rect 1854 3136 1860 3148
rect 1912 3136 1918 3188
rect 2133 3179 2191 3185
rect 2133 3145 2145 3179
rect 2179 3176 2191 3179
rect 3418 3176 3424 3188
rect 2179 3148 3424 3176
rect 2179 3145 2191 3148
rect 2133 3139 2191 3145
rect 3418 3136 3424 3148
rect 3476 3136 3482 3188
rect 5994 3136 6000 3188
rect 6052 3176 6058 3188
rect 6181 3179 6239 3185
rect 6181 3176 6193 3179
rect 6052 3148 6193 3176
rect 6052 3136 6058 3148
rect 6181 3145 6193 3148
rect 6227 3145 6239 3179
rect 6181 3139 6239 3145
rect 20438 3136 20444 3188
rect 20496 3176 20502 3188
rect 21361 3179 21419 3185
rect 21361 3176 21373 3179
rect 20496 3148 21373 3176
rect 20496 3136 20502 3148
rect 21361 3145 21373 3148
rect 21407 3145 21419 3179
rect 21361 3139 21419 3145
rect 2958 3108 2964 3120
rect 1596 3080 2964 3108
rect 2958 3068 2964 3080
rect 3016 3068 3022 3120
rect 1394 3040 1400 3052
rect 1355 3012 1400 3040
rect 1394 3000 1400 3012
rect 1452 3000 1458 3052
rect 1670 3040 1676 3052
rect 1631 3012 1676 3040
rect 1670 3000 1676 3012
rect 1728 3000 1734 3052
rect 1949 3043 2007 3049
rect 1949 3009 1961 3043
rect 1995 3040 2007 3043
rect 5997 3043 6055 3049
rect 1995 3012 2544 3040
rect 1995 3009 2007 3012
rect 1949 3003 2007 3009
rect 1412 2972 1440 3000
rect 2409 2975 2467 2981
rect 2409 2972 2421 2975
rect 1412 2944 2421 2972
rect 2409 2941 2421 2944
rect 2455 2941 2467 2975
rect 2409 2935 2467 2941
rect 2225 2839 2283 2845
rect 2225 2805 2237 2839
rect 2271 2836 2283 2839
rect 2516 2836 2544 3012
rect 5997 3009 6009 3043
rect 6043 3040 6055 3043
rect 8662 3040 8668 3052
rect 6043 3012 8668 3040
rect 6043 3009 6055 3012
rect 5997 3003 6055 3009
rect 8662 3000 8668 3012
rect 8720 3000 8726 3052
rect 9125 3043 9183 3049
rect 9125 3009 9137 3043
rect 9171 3040 9183 3043
rect 16114 3040 16120 3052
rect 9171 3012 16120 3040
rect 9171 3009 9183 3012
rect 9125 3003 9183 3009
rect 16114 3000 16120 3012
rect 16172 3000 16178 3052
rect 17037 3043 17095 3049
rect 17037 3009 17049 3043
rect 17083 3040 17095 3043
rect 20622 3040 20628 3052
rect 17083 3012 20628 3040
rect 17083 3009 17095 3012
rect 17037 3003 17095 3009
rect 20622 3000 20628 3012
rect 20680 3000 20686 3052
rect 20993 3043 21051 3049
rect 20993 3009 21005 3043
rect 21039 3040 21051 3043
rect 21266 3040 21272 3052
rect 21039 3012 21272 3040
rect 21039 3009 21051 3012
rect 20993 3003 21051 3009
rect 21266 3000 21272 3012
rect 21324 3000 21330 3052
rect 21542 3040 21548 3052
rect 21503 3012 21548 3040
rect 21542 3000 21548 3012
rect 21600 3000 21606 3052
rect 20809 2975 20867 2981
rect 20809 2941 20821 2975
rect 20855 2972 20867 2975
rect 21560 2972 21588 3000
rect 20855 2944 21588 2972
rect 20855 2941 20867 2944
rect 20809 2935 20867 2941
rect 5810 2864 5816 2916
rect 5868 2904 5874 2916
rect 8941 2907 8999 2913
rect 8941 2904 8953 2907
rect 5868 2876 8953 2904
rect 5868 2864 5874 2876
rect 8941 2873 8953 2876
rect 8987 2873 8999 2907
rect 16850 2904 16856 2916
rect 16811 2876 16856 2904
rect 8941 2867 8999 2873
rect 16850 2864 16856 2876
rect 16908 2864 16914 2916
rect 19978 2864 19984 2916
rect 20036 2904 20042 2916
rect 21085 2907 21143 2913
rect 21085 2904 21097 2907
rect 20036 2876 21097 2904
rect 20036 2864 20042 2876
rect 21085 2873 21097 2876
rect 21131 2873 21143 2907
rect 21085 2867 21143 2873
rect 2774 2836 2780 2848
rect 2271 2808 2780 2836
rect 2271 2805 2283 2808
rect 2225 2799 2283 2805
rect 2774 2796 2780 2808
rect 2832 2796 2838 2848
rect 20254 2796 20260 2848
rect 20312 2836 20318 2848
rect 20714 2836 20720 2848
rect 20312 2808 20720 2836
rect 20312 2796 20318 2808
rect 20714 2796 20720 2808
rect 20772 2796 20778 2848
rect 1104 2746 21896 2768
rect 1104 2694 3549 2746
rect 3601 2694 3613 2746
rect 3665 2694 3677 2746
rect 3729 2694 3741 2746
rect 3793 2694 3805 2746
rect 3857 2694 8747 2746
rect 8799 2694 8811 2746
rect 8863 2694 8875 2746
rect 8927 2694 8939 2746
rect 8991 2694 9003 2746
rect 9055 2694 13945 2746
rect 13997 2694 14009 2746
rect 14061 2694 14073 2746
rect 14125 2694 14137 2746
rect 14189 2694 14201 2746
rect 14253 2694 19143 2746
rect 19195 2694 19207 2746
rect 19259 2694 19271 2746
rect 19323 2694 19335 2746
rect 19387 2694 19399 2746
rect 19451 2694 21896 2746
rect 1104 2672 21896 2694
rect 2501 2635 2559 2641
rect 2501 2601 2513 2635
rect 2547 2632 2559 2635
rect 6546 2632 6552 2644
rect 2547 2604 6552 2632
rect 2547 2601 2559 2604
rect 2501 2595 2559 2601
rect 6546 2592 6552 2604
rect 6604 2592 6610 2644
rect 8662 2592 8668 2644
rect 8720 2632 8726 2644
rect 11517 2635 11575 2641
rect 11517 2632 11529 2635
rect 8720 2604 11529 2632
rect 8720 2592 8726 2604
rect 11517 2601 11529 2604
rect 11563 2601 11575 2635
rect 16114 2632 16120 2644
rect 16075 2604 16120 2632
rect 11517 2595 11575 2601
rect 16114 2592 16120 2604
rect 16172 2592 16178 2644
rect 20622 2592 20628 2644
rect 20680 2632 20686 2644
rect 20717 2635 20775 2641
rect 20717 2632 20729 2635
rect 20680 2604 20729 2632
rect 20680 2592 20686 2604
rect 20717 2601 20729 2604
rect 20763 2601 20775 2635
rect 20717 2595 20775 2601
rect 20806 2592 20812 2644
rect 20864 2632 20870 2644
rect 21085 2635 21143 2641
rect 21085 2632 21097 2635
rect 20864 2604 21097 2632
rect 20864 2592 20870 2604
rect 21085 2601 21097 2604
rect 21131 2601 21143 2635
rect 21085 2595 21143 2601
rect 20257 2567 20315 2573
rect 20257 2533 20269 2567
rect 20303 2564 20315 2567
rect 20303 2536 21588 2564
rect 20303 2533 20315 2536
rect 20257 2527 20315 2533
rect 1949 2499 2007 2505
rect 1949 2465 1961 2499
rect 1995 2496 2007 2499
rect 4614 2496 4620 2508
rect 1995 2468 4620 2496
rect 1995 2465 2007 2468
rect 1949 2459 2007 2465
rect 4614 2456 4620 2468
rect 4672 2456 4678 2508
rect 20441 2499 20499 2505
rect 20441 2465 20453 2499
rect 20487 2496 20499 2499
rect 20487 2468 21312 2496
rect 20487 2465 20499 2468
rect 20441 2459 20499 2465
rect 21284 2440 21312 2468
rect 21560 2440 21588 2536
rect 2222 2428 2228 2440
rect 2183 2400 2228 2428
rect 2222 2388 2228 2400
rect 2280 2388 2286 2440
rect 2314 2388 2320 2440
rect 2372 2428 2378 2440
rect 2593 2431 2651 2437
rect 2593 2428 2605 2431
rect 2372 2400 2605 2428
rect 2372 2388 2378 2400
rect 2593 2397 2605 2400
rect 2639 2397 2651 2431
rect 2593 2391 2651 2397
rect 6730 2388 6736 2440
rect 6788 2428 6794 2440
rect 7193 2431 7251 2437
rect 7193 2428 7205 2431
rect 6788 2400 7205 2428
rect 6788 2388 6794 2400
rect 7193 2397 7205 2400
rect 7239 2397 7251 2431
rect 7193 2391 7251 2397
rect 11701 2431 11759 2437
rect 11701 2397 11713 2431
rect 11747 2397 11759 2431
rect 16301 2431 16359 2437
rect 16301 2428 16313 2431
rect 11701 2391 11759 2397
rect 16040 2400 16313 2428
rect 2240 2360 2268 2388
rect 2777 2363 2835 2369
rect 2777 2360 2789 2363
rect 2240 2332 2789 2360
rect 2777 2329 2789 2332
rect 2823 2329 2835 2363
rect 2777 2323 2835 2329
rect 11716 2304 11744 2391
rect 16040 2304 16068 2400
rect 16301 2397 16313 2400
rect 16347 2397 16359 2431
rect 16301 2391 16359 2397
rect 20622 2388 20628 2440
rect 20680 2428 20686 2440
rect 20901 2431 20959 2437
rect 20901 2428 20913 2431
rect 20680 2400 20913 2428
rect 20680 2388 20686 2400
rect 20901 2397 20913 2400
rect 20947 2397 20959 2431
rect 21266 2428 21272 2440
rect 21227 2400 21272 2428
rect 20901 2391 20959 2397
rect 21266 2388 21272 2400
rect 21324 2388 21330 2440
rect 21542 2428 21548 2440
rect 21503 2400 21548 2428
rect 21542 2388 21548 2400
rect 21600 2388 21606 2440
rect 20162 2320 20168 2372
rect 20220 2360 20226 2372
rect 20220 2332 21404 2360
rect 20220 2320 20226 2332
rect 6822 2252 6828 2304
rect 6880 2292 6886 2304
rect 7009 2295 7067 2301
rect 7009 2292 7021 2295
rect 6880 2264 7021 2292
rect 6880 2252 6886 2264
rect 7009 2261 7021 2264
rect 7055 2261 7067 2295
rect 7009 2255 7067 2261
rect 11698 2252 11704 2304
rect 11756 2292 11762 2304
rect 11793 2295 11851 2301
rect 11793 2292 11805 2295
rect 11756 2264 11805 2292
rect 11756 2252 11762 2264
rect 11793 2261 11805 2264
rect 11839 2261 11851 2295
rect 16022 2292 16028 2304
rect 15983 2264 16028 2292
rect 11793 2255 11851 2261
rect 16022 2252 16028 2264
rect 16080 2252 16086 2304
rect 20622 2292 20628 2304
rect 20583 2264 20628 2292
rect 20622 2252 20628 2264
rect 20680 2252 20686 2304
rect 21376 2301 21404 2332
rect 21361 2295 21419 2301
rect 21361 2261 21373 2295
rect 21407 2261 21419 2295
rect 21361 2255 21419 2261
rect 1104 2202 22056 2224
rect 1104 2150 6148 2202
rect 6200 2150 6212 2202
rect 6264 2150 6276 2202
rect 6328 2150 6340 2202
rect 6392 2150 6404 2202
rect 6456 2150 11346 2202
rect 11398 2150 11410 2202
rect 11462 2150 11474 2202
rect 11526 2150 11538 2202
rect 11590 2150 11602 2202
rect 11654 2150 16544 2202
rect 16596 2150 16608 2202
rect 16660 2150 16672 2202
rect 16724 2150 16736 2202
rect 16788 2150 16800 2202
rect 16852 2150 21742 2202
rect 21794 2150 21806 2202
rect 21858 2150 21870 2202
rect 21922 2150 21934 2202
rect 21986 2150 21998 2202
rect 22050 2150 22056 2202
rect 1104 2128 22056 2150
<< via1 >>
rect 8944 20816 8996 20868
rect 15568 20816 15620 20868
rect 6148 20646 6200 20698
rect 6212 20646 6264 20698
rect 6276 20646 6328 20698
rect 6340 20646 6392 20698
rect 6404 20646 6456 20698
rect 11346 20646 11398 20698
rect 11410 20646 11462 20698
rect 11474 20646 11526 20698
rect 11538 20646 11590 20698
rect 11602 20646 11654 20698
rect 16544 20646 16596 20698
rect 16608 20646 16660 20698
rect 16672 20646 16724 20698
rect 16736 20646 16788 20698
rect 16800 20646 16852 20698
rect 21742 20646 21794 20698
rect 21806 20646 21858 20698
rect 21870 20646 21922 20698
rect 21934 20646 21986 20698
rect 21998 20646 22050 20698
rect 5540 20587 5592 20596
rect 5540 20553 5549 20587
rect 5549 20553 5583 20587
rect 5583 20553 5592 20587
rect 5540 20544 5592 20553
rect 5724 20544 5776 20596
rect 6000 20544 6052 20596
rect 7380 20544 7432 20596
rect 8944 20544 8996 20596
rect 9036 20544 9088 20596
rect 9220 20544 9272 20596
rect 4252 20476 4304 20528
rect 4528 20476 4580 20528
rect 1676 20451 1728 20460
rect 1676 20417 1685 20451
rect 1685 20417 1719 20451
rect 1719 20417 1728 20451
rect 1676 20408 1728 20417
rect 2044 20408 2096 20460
rect 2872 20408 2924 20460
rect 3240 20340 3292 20392
rect 3516 20408 3568 20460
rect 5448 20476 5500 20528
rect 6828 20476 6880 20528
rect 7012 20476 7064 20528
rect 5540 20408 5592 20460
rect 5816 20408 5868 20460
rect 6368 20451 6420 20460
rect 6368 20417 6377 20451
rect 6377 20417 6411 20451
rect 6411 20417 6420 20451
rect 6368 20408 6420 20417
rect 7104 20408 7156 20460
rect 7564 20476 7616 20528
rect 7840 20408 7892 20460
rect 8300 20476 8352 20528
rect 8024 20451 8076 20460
rect 8024 20417 8033 20451
rect 8033 20417 8067 20451
rect 8067 20417 8076 20451
rect 8024 20408 8076 20417
rect 8392 20408 8444 20460
rect 9772 20544 9824 20596
rect 10508 20544 10560 20596
rect 3976 20340 4028 20392
rect 4344 20340 4396 20392
rect 4712 20340 4764 20392
rect 8116 20340 8168 20392
rect 9588 20408 9640 20460
rect 13084 20476 13136 20528
rect 9864 20451 9916 20460
rect 9864 20417 9873 20451
rect 9873 20417 9907 20451
rect 9907 20417 9916 20451
rect 9864 20408 9916 20417
rect 8668 20340 8720 20392
rect 11060 20451 11112 20460
rect 11060 20417 11069 20451
rect 11069 20417 11103 20451
rect 11103 20417 11112 20451
rect 11060 20408 11112 20417
rect 11244 20408 11296 20460
rect 11980 20408 12032 20460
rect 12256 20408 12308 20460
rect 12808 20451 12860 20460
rect 12808 20417 12817 20451
rect 12817 20417 12851 20451
rect 12851 20417 12860 20451
rect 12808 20408 12860 20417
rect 13636 20408 13688 20460
rect 10232 20383 10284 20392
rect 10232 20349 10241 20383
rect 10241 20349 10275 20383
rect 10275 20349 10284 20383
rect 10232 20340 10284 20349
rect 10416 20383 10468 20392
rect 10416 20349 10425 20383
rect 10425 20349 10459 20383
rect 10459 20349 10468 20383
rect 10416 20340 10468 20349
rect 12532 20340 12584 20392
rect 12992 20340 13044 20392
rect 15108 20476 15160 20528
rect 14280 20408 14332 20460
rect 15200 20408 15252 20460
rect 2688 20272 2740 20324
rect 5724 20272 5776 20324
rect 8576 20272 8628 20324
rect 9404 20272 9456 20324
rect 9680 20272 9732 20324
rect 9864 20272 9916 20324
rect 10784 20272 10836 20324
rect 13912 20340 13964 20392
rect 14464 20340 14516 20392
rect 14740 20340 14792 20392
rect 14832 20340 14884 20392
rect 16028 20544 16080 20596
rect 16948 20544 17000 20596
rect 17960 20544 18012 20596
rect 18696 20544 18748 20596
rect 20076 20544 20128 20596
rect 15568 20476 15620 20528
rect 19064 20476 19116 20528
rect 15660 20408 15712 20460
rect 16120 20451 16172 20460
rect 16120 20417 16129 20451
rect 16129 20417 16163 20451
rect 16163 20417 16172 20451
rect 16120 20408 16172 20417
rect 16212 20408 16264 20460
rect 16856 20408 16908 20460
rect 17408 20451 17460 20460
rect 17408 20417 17417 20451
rect 17417 20417 17451 20451
rect 17451 20417 17460 20451
rect 17408 20408 17460 20417
rect 17776 20451 17828 20460
rect 17776 20417 17785 20451
rect 17785 20417 17819 20451
rect 17819 20417 17828 20451
rect 17776 20408 17828 20417
rect 18144 20451 18196 20460
rect 18144 20417 18153 20451
rect 18153 20417 18187 20451
rect 18187 20417 18196 20451
rect 18144 20408 18196 20417
rect 18880 20408 18932 20460
rect 18972 20408 19024 20460
rect 19616 20451 19668 20460
rect 19616 20417 19625 20451
rect 19625 20417 19659 20451
rect 19659 20417 19668 20451
rect 19616 20408 19668 20417
rect 19984 20451 20036 20460
rect 19984 20417 19993 20451
rect 19993 20417 20027 20451
rect 20027 20417 20036 20451
rect 19984 20408 20036 20417
rect 20352 20451 20404 20460
rect 20352 20417 20361 20451
rect 20361 20417 20395 20451
rect 20395 20417 20404 20451
rect 20352 20408 20404 20417
rect 13820 20272 13872 20324
rect 15292 20272 15344 20324
rect 16580 20272 16632 20324
rect 17500 20272 17552 20324
rect 1492 20247 1544 20256
rect 1492 20213 1501 20247
rect 1501 20213 1535 20247
rect 1535 20213 1544 20247
rect 1492 20204 1544 20213
rect 4896 20247 4948 20256
rect 4896 20213 4905 20247
rect 4905 20213 4939 20247
rect 4939 20213 4948 20247
rect 4896 20204 4948 20213
rect 5264 20204 5316 20256
rect 6828 20247 6880 20256
rect 6828 20213 6837 20247
rect 6837 20213 6871 20247
rect 6871 20213 6880 20247
rect 6828 20204 6880 20213
rect 7196 20204 7248 20256
rect 7472 20204 7524 20256
rect 7656 20247 7708 20256
rect 7656 20213 7665 20247
rect 7665 20213 7699 20247
rect 7699 20213 7708 20247
rect 7656 20204 7708 20213
rect 8208 20247 8260 20256
rect 8208 20213 8217 20247
rect 8217 20213 8251 20247
rect 8251 20213 8260 20247
rect 8208 20204 8260 20213
rect 8300 20247 8352 20256
rect 8300 20213 8309 20247
rect 8309 20213 8343 20247
rect 8343 20213 8352 20247
rect 8300 20204 8352 20213
rect 8484 20204 8536 20256
rect 9312 20204 9364 20256
rect 9496 20204 9548 20256
rect 9956 20204 10008 20256
rect 12164 20204 12216 20256
rect 13912 20247 13964 20256
rect 13912 20213 13921 20247
rect 13921 20213 13955 20247
rect 13955 20213 13964 20247
rect 13912 20204 13964 20213
rect 14188 20204 14240 20256
rect 17132 20204 17184 20256
rect 18696 20204 18748 20256
rect 19708 20340 19760 20392
rect 21364 20408 21416 20460
rect 19340 20272 19392 20324
rect 19432 20204 19484 20256
rect 20444 20204 20496 20256
rect 3549 20102 3601 20154
rect 3613 20102 3665 20154
rect 3677 20102 3729 20154
rect 3741 20102 3793 20154
rect 3805 20102 3857 20154
rect 8747 20102 8799 20154
rect 8811 20102 8863 20154
rect 8875 20102 8927 20154
rect 8939 20102 8991 20154
rect 9003 20102 9055 20154
rect 13945 20102 13997 20154
rect 14009 20102 14061 20154
rect 14073 20102 14125 20154
rect 14137 20102 14189 20154
rect 14201 20102 14253 20154
rect 19143 20102 19195 20154
rect 19207 20102 19259 20154
rect 19271 20102 19323 20154
rect 19335 20102 19387 20154
rect 19399 20102 19451 20154
rect 1860 20043 1912 20052
rect 1860 20009 1869 20043
rect 1869 20009 1903 20043
rect 1903 20009 1912 20043
rect 1860 20000 1912 20009
rect 2780 20000 2832 20052
rect 3056 20043 3108 20052
rect 3056 20009 3065 20043
rect 3065 20009 3099 20043
rect 3099 20009 3108 20043
rect 3056 20000 3108 20009
rect 3240 20000 3292 20052
rect 3516 20000 3568 20052
rect 7104 20000 7156 20052
rect 8668 20000 8720 20052
rect 10416 20000 10468 20052
rect 10600 20043 10652 20052
rect 10600 20009 10609 20043
rect 10609 20009 10643 20043
rect 10643 20009 10652 20043
rect 10600 20000 10652 20009
rect 14280 20000 14332 20052
rect 14556 20000 14608 20052
rect 15752 20000 15804 20052
rect 16856 20043 16908 20052
rect 4712 19932 4764 19984
rect 7564 19932 7616 19984
rect 8484 19932 8536 19984
rect 9404 19932 9456 19984
rect 9588 19932 9640 19984
rect 10140 19932 10192 19984
rect 10876 19932 10928 19984
rect 2228 19796 2280 19848
rect 2320 19728 2372 19780
rect 2504 19796 2556 19848
rect 2872 19839 2924 19848
rect 2872 19805 2881 19839
rect 2881 19805 2915 19839
rect 2915 19805 2924 19839
rect 2872 19796 2924 19805
rect 3148 19796 3200 19848
rect 1492 19703 1544 19712
rect 1492 19669 1501 19703
rect 1501 19669 1535 19703
rect 1535 19669 1544 19703
rect 1492 19660 1544 19669
rect 3240 19660 3292 19712
rect 3884 19796 3936 19848
rect 4252 19839 4304 19848
rect 4252 19805 4261 19839
rect 4261 19805 4295 19839
rect 4295 19805 4304 19839
rect 4252 19796 4304 19805
rect 4620 19839 4672 19848
rect 4620 19805 4629 19839
rect 4629 19805 4663 19839
rect 4663 19805 4672 19839
rect 4620 19796 4672 19805
rect 4988 19839 5040 19848
rect 4712 19728 4764 19780
rect 4160 19660 4212 19712
rect 4436 19703 4488 19712
rect 4436 19669 4445 19703
rect 4445 19669 4479 19703
rect 4479 19669 4488 19703
rect 4436 19660 4488 19669
rect 4988 19805 4997 19839
rect 4997 19805 5031 19839
rect 5031 19805 5040 19839
rect 4988 19796 5040 19805
rect 6000 19839 6052 19848
rect 6000 19805 6009 19839
rect 6009 19805 6043 19839
rect 6043 19805 6052 19839
rect 6000 19796 6052 19805
rect 7288 19864 7340 19916
rect 9772 19864 9824 19916
rect 10048 19864 10100 19916
rect 10232 19864 10284 19916
rect 10784 19864 10836 19916
rect 12072 19864 12124 19916
rect 13360 19864 13412 19916
rect 4896 19728 4948 19780
rect 5172 19660 5224 19712
rect 5632 19728 5684 19780
rect 6828 19796 6880 19848
rect 9680 19796 9732 19848
rect 7748 19728 7800 19780
rect 8944 19728 8996 19780
rect 9404 19728 9456 19780
rect 10324 19796 10376 19848
rect 11888 19796 11940 19848
rect 12440 19839 12492 19848
rect 12440 19805 12449 19839
rect 12449 19805 12483 19839
rect 12483 19805 12492 19839
rect 12440 19796 12492 19805
rect 12624 19796 12676 19848
rect 12716 19839 12768 19848
rect 12716 19805 12725 19839
rect 12725 19805 12759 19839
rect 12759 19805 12768 19839
rect 13452 19839 13504 19848
rect 12716 19796 12768 19805
rect 13452 19805 13461 19839
rect 13461 19805 13495 19839
rect 13495 19805 13504 19839
rect 13452 19796 13504 19805
rect 13544 19796 13596 19848
rect 13820 19796 13872 19848
rect 14832 19796 14884 19848
rect 15200 19932 15252 19984
rect 16856 20009 16865 20043
rect 16865 20009 16899 20043
rect 16899 20009 16908 20043
rect 16856 20000 16908 20009
rect 17408 20043 17460 20052
rect 17408 20009 17417 20043
rect 17417 20009 17451 20043
rect 17451 20009 17460 20043
rect 17408 20000 17460 20009
rect 17776 20043 17828 20052
rect 17776 20009 17785 20043
rect 17785 20009 17819 20043
rect 17819 20009 17828 20043
rect 17776 20000 17828 20009
rect 18236 20000 18288 20052
rect 18880 20043 18932 20052
rect 18880 20009 18889 20043
rect 18889 20009 18923 20043
rect 18923 20009 18932 20043
rect 18880 20000 18932 20009
rect 19892 20043 19944 20052
rect 19892 20009 19901 20043
rect 19901 20009 19935 20043
rect 19935 20009 19944 20043
rect 19892 20000 19944 20009
rect 20260 20043 20312 20052
rect 20260 20009 20269 20043
rect 20269 20009 20303 20043
rect 20303 20009 20312 20043
rect 20260 20000 20312 20009
rect 20812 20000 20864 20052
rect 15016 19864 15068 19916
rect 16120 19864 16172 19916
rect 15292 19796 15344 19848
rect 16304 19839 16356 19848
rect 7012 19660 7064 19712
rect 7380 19660 7432 19712
rect 8116 19660 8168 19712
rect 9036 19660 9088 19712
rect 9680 19660 9732 19712
rect 11796 19728 11848 19780
rect 12348 19728 12400 19780
rect 13176 19660 13228 19712
rect 14556 19703 14608 19712
rect 14556 19669 14565 19703
rect 14565 19669 14599 19703
rect 14599 19669 14608 19703
rect 16304 19805 16313 19839
rect 16313 19805 16347 19839
rect 16347 19805 16356 19839
rect 16304 19796 16356 19805
rect 16396 19839 16448 19848
rect 16396 19805 16405 19839
rect 16405 19805 16439 19839
rect 16439 19805 16448 19839
rect 16396 19796 16448 19805
rect 16948 19796 17000 19848
rect 17224 19839 17276 19848
rect 17224 19805 17233 19839
rect 17233 19805 17267 19839
rect 17267 19805 17276 19839
rect 21180 19932 21232 19984
rect 17224 19796 17276 19805
rect 14556 19660 14608 19669
rect 14832 19660 14884 19712
rect 14924 19660 14976 19712
rect 15752 19660 15804 19712
rect 18052 19839 18104 19848
rect 18052 19805 18061 19839
rect 18061 19805 18095 19839
rect 18095 19805 18104 19839
rect 18604 19839 18656 19848
rect 18052 19796 18104 19805
rect 18604 19805 18613 19839
rect 18613 19805 18647 19839
rect 18647 19805 18656 19839
rect 18604 19796 18656 19805
rect 18788 19796 18840 19848
rect 19708 19796 19760 19848
rect 20260 19796 20312 19848
rect 20996 19796 21048 19848
rect 20720 19728 20772 19780
rect 19800 19660 19852 19712
rect 20168 19660 20220 19712
rect 21456 19703 21508 19712
rect 21456 19669 21465 19703
rect 21465 19669 21499 19703
rect 21499 19669 21508 19703
rect 21456 19660 21508 19669
rect 6148 19558 6200 19610
rect 6212 19558 6264 19610
rect 6276 19558 6328 19610
rect 6340 19558 6392 19610
rect 6404 19558 6456 19610
rect 11346 19558 11398 19610
rect 11410 19558 11462 19610
rect 11474 19558 11526 19610
rect 11538 19558 11590 19610
rect 11602 19558 11654 19610
rect 16544 19558 16596 19610
rect 16608 19558 16660 19610
rect 16672 19558 16724 19610
rect 16736 19558 16788 19610
rect 16800 19558 16852 19610
rect 21742 19558 21794 19610
rect 21806 19558 21858 19610
rect 21870 19558 21922 19610
rect 21934 19558 21986 19610
rect 21998 19558 22050 19610
rect 2320 19456 2372 19508
rect 2872 19499 2924 19508
rect 2872 19465 2881 19499
rect 2881 19465 2915 19499
rect 2915 19465 2924 19499
rect 2872 19456 2924 19465
rect 3240 19499 3292 19508
rect 2228 19388 2280 19440
rect 3240 19465 3249 19499
rect 3249 19465 3283 19499
rect 3283 19465 3292 19499
rect 3240 19456 3292 19465
rect 3332 19456 3384 19508
rect 3976 19499 4028 19508
rect 3976 19465 3985 19499
rect 3985 19465 4019 19499
rect 4019 19465 4028 19499
rect 3976 19456 4028 19465
rect 4988 19456 5040 19508
rect 5080 19456 5132 19508
rect 7932 19456 7984 19508
rect 8484 19456 8536 19508
rect 9220 19456 9272 19508
rect 9680 19456 9732 19508
rect 12348 19456 12400 19508
rect 12624 19499 12676 19508
rect 12624 19465 12633 19499
rect 12633 19465 12667 19499
rect 12667 19465 12676 19499
rect 12624 19456 12676 19465
rect 12808 19499 12860 19508
rect 12808 19465 12817 19499
rect 12817 19465 12851 19499
rect 12851 19465 12860 19499
rect 12808 19456 12860 19465
rect 13360 19499 13412 19508
rect 13360 19465 13369 19499
rect 13369 19465 13403 19499
rect 13403 19465 13412 19499
rect 13360 19456 13412 19465
rect 15016 19499 15068 19508
rect 15016 19465 15025 19499
rect 15025 19465 15059 19499
rect 15059 19465 15068 19499
rect 15016 19456 15068 19465
rect 15660 19499 15712 19508
rect 3056 19388 3108 19440
rect 2044 19363 2096 19372
rect 2044 19329 2053 19363
rect 2053 19329 2087 19363
rect 2087 19329 2096 19363
rect 2044 19320 2096 19329
rect 2320 19363 2372 19372
rect 2320 19329 2329 19363
rect 2329 19329 2363 19363
rect 2363 19329 2372 19363
rect 2320 19320 2372 19329
rect 1860 19227 1912 19236
rect 1860 19193 1869 19227
rect 1869 19193 1903 19227
rect 1903 19193 1912 19227
rect 1860 19184 1912 19193
rect 1492 19159 1544 19168
rect 1492 19125 1501 19159
rect 1501 19125 1535 19159
rect 1535 19125 1544 19159
rect 1492 19116 1544 19125
rect 2964 19320 3016 19372
rect 3240 19320 3292 19372
rect 3332 19320 3384 19372
rect 2872 19252 2924 19304
rect 5908 19388 5960 19440
rect 7104 19388 7156 19440
rect 3792 19363 3844 19372
rect 3792 19329 3801 19363
rect 3801 19329 3835 19363
rect 3835 19329 3844 19363
rect 3792 19320 3844 19329
rect 3976 19320 4028 19372
rect 5172 19320 5224 19372
rect 6736 19320 6788 19372
rect 7564 19363 7616 19372
rect 7564 19329 7582 19363
rect 7582 19329 7616 19363
rect 8300 19431 8352 19440
rect 8300 19397 8309 19431
rect 8309 19397 8343 19431
rect 8343 19397 8352 19431
rect 8300 19388 8352 19397
rect 7564 19320 7616 19329
rect 4160 19252 4212 19304
rect 4344 19252 4396 19304
rect 4712 19295 4764 19304
rect 4712 19261 4721 19295
rect 4721 19261 4755 19295
rect 4755 19261 4764 19295
rect 4712 19252 4764 19261
rect 4896 19295 4948 19304
rect 4896 19261 4905 19295
rect 4905 19261 4939 19295
rect 4939 19261 4948 19295
rect 4896 19252 4948 19261
rect 5632 19295 5684 19304
rect 5632 19261 5641 19295
rect 5641 19261 5675 19295
rect 5675 19261 5684 19295
rect 5632 19252 5684 19261
rect 8116 19320 8168 19372
rect 8668 19363 8720 19372
rect 8668 19329 8702 19363
rect 8702 19329 8720 19363
rect 8668 19320 8720 19329
rect 9036 19320 9088 19372
rect 11888 19388 11940 19440
rect 15660 19465 15669 19499
rect 15669 19465 15703 19499
rect 15703 19465 15712 19499
rect 15660 19456 15712 19465
rect 16212 19456 16264 19508
rect 17224 19456 17276 19508
rect 18144 19499 18196 19508
rect 3608 19184 3660 19236
rect 4160 19159 4212 19168
rect 4160 19125 4169 19159
rect 4169 19125 4203 19159
rect 4203 19125 4212 19159
rect 4160 19116 4212 19125
rect 6000 19184 6052 19236
rect 6644 19184 6696 19236
rect 4804 19116 4856 19168
rect 5356 19159 5408 19168
rect 5356 19125 5365 19159
rect 5365 19125 5399 19159
rect 5399 19125 5408 19159
rect 5356 19116 5408 19125
rect 6184 19159 6236 19168
rect 6184 19125 6193 19159
rect 6193 19125 6227 19159
rect 6227 19125 6236 19159
rect 6184 19116 6236 19125
rect 6552 19116 6604 19168
rect 7932 19116 7984 19168
rect 8116 19159 8168 19168
rect 8116 19125 8125 19159
rect 8125 19125 8159 19159
rect 8159 19125 8168 19159
rect 8116 19116 8168 19125
rect 10048 19320 10100 19372
rect 11980 19363 12032 19372
rect 9772 19227 9824 19236
rect 9772 19193 9781 19227
rect 9781 19193 9815 19227
rect 9815 19193 9824 19227
rect 9772 19184 9824 19193
rect 9680 19116 9732 19168
rect 11704 19295 11756 19304
rect 11704 19261 11713 19295
rect 11713 19261 11747 19295
rect 11747 19261 11756 19295
rect 11704 19252 11756 19261
rect 11980 19329 11989 19363
rect 11989 19329 12023 19363
rect 12023 19329 12032 19363
rect 11980 19320 12032 19329
rect 12072 19320 12124 19372
rect 12256 19252 12308 19304
rect 10968 19184 11020 19236
rect 14464 19363 14516 19372
rect 14464 19329 14482 19363
rect 14482 19329 14516 19363
rect 14464 19320 14516 19329
rect 14924 19320 14976 19372
rect 15200 19363 15252 19372
rect 15200 19329 15209 19363
rect 15209 19329 15243 19363
rect 15243 19329 15252 19363
rect 15200 19320 15252 19329
rect 15660 19320 15712 19372
rect 15844 19320 15896 19372
rect 17132 19363 17184 19372
rect 17132 19329 17141 19363
rect 17141 19329 17175 19363
rect 17175 19329 17184 19363
rect 17132 19320 17184 19329
rect 18144 19465 18153 19499
rect 18153 19465 18187 19499
rect 18187 19465 18196 19499
rect 18144 19456 18196 19465
rect 18604 19499 18656 19508
rect 18604 19465 18613 19499
rect 18613 19465 18647 19499
rect 18647 19465 18656 19499
rect 18604 19456 18656 19465
rect 18972 19456 19024 19508
rect 19064 19456 19116 19508
rect 19984 19456 20036 19508
rect 20260 19499 20312 19508
rect 20260 19465 20269 19499
rect 20269 19465 20303 19499
rect 20303 19465 20312 19499
rect 20260 19456 20312 19465
rect 20904 19456 20956 19508
rect 21088 19499 21140 19508
rect 21088 19465 21097 19499
rect 21097 19465 21131 19499
rect 21131 19465 21140 19499
rect 21088 19456 21140 19465
rect 17960 19388 18012 19440
rect 19800 19388 19852 19440
rect 11152 19116 11204 19168
rect 11796 19116 11848 19168
rect 14372 19116 14424 19168
rect 16396 19252 16448 19304
rect 16856 19295 16908 19304
rect 16856 19261 16865 19295
rect 16865 19261 16899 19295
rect 16899 19261 16908 19295
rect 16856 19252 16908 19261
rect 17040 19295 17092 19304
rect 17040 19261 17049 19295
rect 17049 19261 17083 19295
rect 17083 19261 17092 19295
rect 17040 19252 17092 19261
rect 14832 19184 14884 19236
rect 16028 19227 16080 19236
rect 16028 19193 16037 19227
rect 16037 19193 16071 19227
rect 16071 19193 16080 19227
rect 16028 19184 16080 19193
rect 18420 19363 18472 19372
rect 18420 19329 18429 19363
rect 18429 19329 18463 19363
rect 18463 19329 18472 19363
rect 18420 19320 18472 19329
rect 18880 19320 18932 19372
rect 19524 19320 19576 19372
rect 19984 19363 20036 19372
rect 19984 19329 19993 19363
rect 19993 19329 20027 19363
rect 20027 19329 20036 19363
rect 19984 19320 20036 19329
rect 20904 19363 20956 19372
rect 18236 19252 18288 19304
rect 20904 19329 20913 19363
rect 20913 19329 20947 19363
rect 20947 19329 20956 19363
rect 20904 19320 20956 19329
rect 21272 19363 21324 19372
rect 21272 19329 21281 19363
rect 21281 19329 21315 19363
rect 21315 19329 21324 19363
rect 21272 19320 21324 19329
rect 18144 19184 18196 19236
rect 19524 19227 19576 19236
rect 19524 19193 19533 19227
rect 19533 19193 19567 19227
rect 19567 19193 19576 19227
rect 19524 19184 19576 19193
rect 20812 19184 20864 19236
rect 20168 19159 20220 19168
rect 20168 19125 20177 19159
rect 20177 19125 20211 19159
rect 20211 19125 20220 19159
rect 20168 19116 20220 19125
rect 21456 19159 21508 19168
rect 21456 19125 21465 19159
rect 21465 19125 21499 19159
rect 21499 19125 21508 19159
rect 21456 19116 21508 19125
rect 3549 19014 3601 19066
rect 3613 19014 3665 19066
rect 3677 19014 3729 19066
rect 3741 19014 3793 19066
rect 3805 19014 3857 19066
rect 8747 19014 8799 19066
rect 8811 19014 8863 19066
rect 8875 19014 8927 19066
rect 8939 19014 8991 19066
rect 9003 19014 9055 19066
rect 13945 19014 13997 19066
rect 14009 19014 14061 19066
rect 14073 19014 14125 19066
rect 14137 19014 14189 19066
rect 14201 19014 14253 19066
rect 19143 19014 19195 19066
rect 19207 19014 19259 19066
rect 19271 19014 19323 19066
rect 19335 19014 19387 19066
rect 19399 19014 19451 19066
rect 2044 18912 2096 18964
rect 2412 18912 2464 18964
rect 1860 18844 1912 18896
rect 1768 18776 1820 18828
rect 2412 18819 2464 18828
rect 2044 18708 2096 18760
rect 2412 18785 2421 18819
rect 2421 18785 2455 18819
rect 2455 18785 2464 18819
rect 2412 18776 2464 18785
rect 3976 18912 4028 18964
rect 4896 18955 4948 18964
rect 4896 18921 4905 18955
rect 4905 18921 4939 18955
rect 4939 18921 4948 18955
rect 4896 18912 4948 18921
rect 2688 18844 2740 18896
rect 3240 18844 3292 18896
rect 3332 18844 3384 18896
rect 4988 18844 5040 18896
rect 6644 18912 6696 18964
rect 10968 18912 11020 18964
rect 11428 18912 11480 18964
rect 13452 18912 13504 18964
rect 13636 18955 13688 18964
rect 13636 18921 13645 18955
rect 13645 18921 13679 18955
rect 13679 18921 13688 18955
rect 13636 18912 13688 18921
rect 14096 18912 14148 18964
rect 14372 18912 14424 18964
rect 14464 18912 14516 18964
rect 16856 18912 16908 18964
rect 17040 18912 17092 18964
rect 20904 18912 20956 18964
rect 21548 18912 21600 18964
rect 5632 18844 5684 18896
rect 6276 18844 6328 18896
rect 6460 18844 6512 18896
rect 6552 18776 6604 18828
rect 7564 18776 7616 18828
rect 3976 18708 4028 18760
rect 1492 18615 1544 18624
rect 1492 18581 1501 18615
rect 1501 18581 1535 18615
rect 1535 18581 1544 18615
rect 1492 18572 1544 18581
rect 4436 18683 4488 18692
rect 3516 18615 3568 18624
rect 3516 18581 3525 18615
rect 3525 18581 3559 18615
rect 3559 18581 3568 18615
rect 3516 18572 3568 18581
rect 4436 18649 4445 18683
rect 4445 18649 4479 18683
rect 4479 18649 4488 18683
rect 4436 18640 4488 18649
rect 6184 18708 6236 18760
rect 4804 18572 4856 18624
rect 5172 18615 5224 18624
rect 5172 18581 5181 18615
rect 5181 18581 5215 18615
rect 5215 18581 5224 18615
rect 5172 18572 5224 18581
rect 6552 18640 6604 18692
rect 8760 18751 8812 18760
rect 8760 18717 8769 18751
rect 8769 18717 8803 18751
rect 8803 18717 8812 18751
rect 8760 18708 8812 18717
rect 9496 18708 9548 18760
rect 9220 18640 9272 18692
rect 9036 18572 9088 18624
rect 9680 18844 9732 18896
rect 11336 18844 11388 18896
rect 16580 18887 16632 18896
rect 16580 18853 16589 18887
rect 16589 18853 16623 18887
rect 16623 18853 16632 18887
rect 16580 18844 16632 18853
rect 17132 18844 17184 18896
rect 11888 18751 11940 18760
rect 11888 18717 11897 18751
rect 11897 18717 11931 18751
rect 11931 18717 11940 18751
rect 11888 18708 11940 18717
rect 12440 18708 12492 18760
rect 13268 18708 13320 18760
rect 14096 18751 14148 18760
rect 14096 18717 14105 18751
rect 14105 18717 14139 18751
rect 14139 18717 14148 18751
rect 14096 18708 14148 18717
rect 17960 18751 18012 18760
rect 17960 18717 17969 18751
rect 17969 18717 18003 18751
rect 18003 18717 18012 18751
rect 17960 18708 18012 18717
rect 9772 18640 9824 18692
rect 11336 18640 11388 18692
rect 16580 18640 16632 18692
rect 17224 18640 17276 18692
rect 21272 18844 21324 18896
rect 22284 18776 22336 18828
rect 20628 18751 20680 18760
rect 20628 18717 20637 18751
rect 20637 18717 20671 18751
rect 20671 18717 20680 18751
rect 20628 18708 20680 18717
rect 20812 18708 20864 18760
rect 21272 18751 21324 18760
rect 21272 18717 21281 18751
rect 21281 18717 21315 18751
rect 21315 18717 21324 18751
rect 21272 18708 21324 18717
rect 13452 18572 13504 18624
rect 18328 18572 18380 18624
rect 20352 18572 20404 18624
rect 21456 18615 21508 18624
rect 21456 18581 21465 18615
rect 21465 18581 21499 18615
rect 21499 18581 21508 18615
rect 21456 18572 21508 18581
rect 6148 18470 6200 18522
rect 6212 18470 6264 18522
rect 6276 18470 6328 18522
rect 6340 18470 6392 18522
rect 6404 18470 6456 18522
rect 11346 18470 11398 18522
rect 11410 18470 11462 18522
rect 11474 18470 11526 18522
rect 11538 18470 11590 18522
rect 11602 18470 11654 18522
rect 16544 18470 16596 18522
rect 16608 18470 16660 18522
rect 16672 18470 16724 18522
rect 16736 18470 16788 18522
rect 16800 18470 16852 18522
rect 21742 18470 21794 18522
rect 21806 18470 21858 18522
rect 21870 18470 21922 18522
rect 21934 18470 21986 18522
rect 21998 18470 22050 18522
rect 1676 18368 1728 18420
rect 2688 18368 2740 18420
rect 3148 18368 3200 18420
rect 3884 18411 3936 18420
rect 3884 18377 3893 18411
rect 3893 18377 3927 18411
rect 3927 18377 3936 18411
rect 3884 18368 3936 18377
rect 4068 18411 4120 18420
rect 4068 18377 4077 18411
rect 4077 18377 4111 18411
rect 4111 18377 4120 18411
rect 4068 18368 4120 18377
rect 4528 18411 4580 18420
rect 4528 18377 4537 18411
rect 4537 18377 4571 18411
rect 4571 18377 4580 18411
rect 4528 18368 4580 18377
rect 4620 18368 4672 18420
rect 5448 18368 5500 18420
rect 5908 18368 5960 18420
rect 1400 18300 1452 18352
rect 1952 18232 2004 18284
rect 2964 18300 3016 18352
rect 3976 18300 4028 18352
rect 5816 18300 5868 18352
rect 1308 18096 1360 18148
rect 1860 18096 1912 18148
rect 2412 18232 2464 18284
rect 3424 18232 3476 18284
rect 4712 18164 4764 18216
rect 6644 18300 6696 18352
rect 7932 18368 7984 18420
rect 8668 18368 8720 18420
rect 9588 18368 9640 18420
rect 8576 18343 8628 18352
rect 8576 18309 8585 18343
rect 8585 18309 8619 18343
rect 8619 18309 8628 18343
rect 8576 18300 8628 18309
rect 9496 18343 9548 18352
rect 9496 18309 9530 18343
rect 9530 18309 9548 18343
rect 9496 18300 9548 18309
rect 10232 18300 10284 18352
rect 10600 18300 10652 18352
rect 8760 18232 8812 18284
rect 11888 18300 11940 18352
rect 10876 18232 10928 18284
rect 13176 18232 13228 18284
rect 10692 18207 10744 18216
rect 10692 18173 10701 18207
rect 10701 18173 10735 18207
rect 10735 18173 10744 18207
rect 10692 18164 10744 18173
rect 11796 18207 11848 18216
rect 11796 18173 11805 18207
rect 11805 18173 11839 18207
rect 11839 18173 11848 18207
rect 11796 18164 11848 18173
rect 12440 18164 12492 18216
rect 14372 18300 14424 18352
rect 16304 18368 16356 18420
rect 18420 18368 18472 18420
rect 21272 18368 21324 18420
rect 14832 18232 14884 18284
rect 18052 18300 18104 18352
rect 15752 18275 15804 18284
rect 15752 18241 15761 18275
rect 15761 18241 15795 18275
rect 15795 18241 15804 18275
rect 15752 18232 15804 18241
rect 17408 18275 17460 18284
rect 17408 18241 17417 18275
rect 17417 18241 17451 18275
rect 17451 18241 17460 18275
rect 17408 18232 17460 18241
rect 20536 18275 20588 18284
rect 20536 18241 20545 18275
rect 20545 18241 20579 18275
rect 20579 18241 20588 18275
rect 20536 18232 20588 18241
rect 2504 18096 2556 18148
rect 2872 18139 2924 18148
rect 2872 18105 2881 18139
rect 2881 18105 2915 18139
rect 2915 18105 2924 18139
rect 2872 18096 2924 18105
rect 3148 18096 3200 18148
rect 3240 18096 3292 18148
rect 1492 18071 1544 18080
rect 1492 18037 1501 18071
rect 1501 18037 1535 18071
rect 1535 18037 1544 18071
rect 1492 18028 1544 18037
rect 2688 18071 2740 18080
rect 2688 18037 2697 18071
rect 2697 18037 2731 18071
rect 2731 18037 2740 18071
rect 2688 18028 2740 18037
rect 3332 18071 3384 18080
rect 3332 18037 3341 18071
rect 3341 18037 3375 18071
rect 3375 18037 3384 18071
rect 3332 18028 3384 18037
rect 4068 18028 4120 18080
rect 6000 18096 6052 18148
rect 6644 18096 6696 18148
rect 8300 18096 8352 18148
rect 9036 18028 9088 18080
rect 9496 18028 9548 18080
rect 10508 18028 10560 18080
rect 12808 18028 12860 18080
rect 15568 18164 15620 18216
rect 18420 18207 18472 18216
rect 18420 18173 18429 18207
rect 18429 18173 18463 18207
rect 18463 18173 18472 18207
rect 18420 18164 18472 18173
rect 19892 18164 19944 18216
rect 21180 18232 21232 18284
rect 18328 18096 18380 18148
rect 20720 18096 20772 18148
rect 18052 18071 18104 18080
rect 18052 18037 18061 18071
rect 18061 18037 18095 18071
rect 18095 18037 18104 18071
rect 18052 18028 18104 18037
rect 21456 18071 21508 18080
rect 21456 18037 21465 18071
rect 21465 18037 21499 18071
rect 21499 18037 21508 18071
rect 21456 18028 21508 18037
rect 3549 17926 3601 17978
rect 3613 17926 3665 17978
rect 3677 17926 3729 17978
rect 3741 17926 3793 17978
rect 3805 17926 3857 17978
rect 8747 17926 8799 17978
rect 8811 17926 8863 17978
rect 8875 17926 8927 17978
rect 8939 17926 8991 17978
rect 9003 17926 9055 17978
rect 13945 17926 13997 17978
rect 14009 17926 14061 17978
rect 14073 17926 14125 17978
rect 14137 17926 14189 17978
rect 14201 17926 14253 17978
rect 19143 17926 19195 17978
rect 19207 17926 19259 17978
rect 19271 17926 19323 17978
rect 19335 17926 19387 17978
rect 19399 17926 19451 17978
rect 2044 17824 2096 17876
rect 2320 17824 2372 17876
rect 2596 17867 2648 17876
rect 2596 17833 2605 17867
rect 2605 17833 2639 17867
rect 2639 17833 2648 17867
rect 2596 17824 2648 17833
rect 6000 17824 6052 17876
rect 6920 17824 6972 17876
rect 7380 17824 7432 17876
rect 7840 17824 7892 17876
rect 8392 17824 8444 17876
rect 8760 17867 8812 17876
rect 8760 17833 8769 17867
rect 8769 17833 8803 17867
rect 8803 17833 8812 17867
rect 8760 17824 8812 17833
rect 9128 17824 9180 17876
rect 9864 17824 9916 17876
rect 10416 17867 10468 17876
rect 10416 17833 10425 17867
rect 10425 17833 10459 17867
rect 10459 17833 10468 17867
rect 10416 17824 10468 17833
rect 11152 17824 11204 17876
rect 12072 17824 12124 17876
rect 12624 17824 12676 17876
rect 8024 17756 8076 17808
rect 2596 17688 2648 17740
rect 8208 17731 8260 17740
rect 8208 17697 8217 17731
rect 8217 17697 8251 17731
rect 8251 17697 8260 17731
rect 8208 17688 8260 17697
rect 10508 17756 10560 17808
rect 11520 17756 11572 17808
rect 15568 17824 15620 17876
rect 15752 17824 15804 17876
rect 20536 17824 20588 17876
rect 14556 17756 14608 17808
rect 16948 17756 17000 17808
rect 17500 17756 17552 17808
rect 9772 17688 9824 17740
rect 10048 17688 10100 17740
rect 11244 17688 11296 17740
rect 11704 17688 11756 17740
rect 12164 17731 12216 17740
rect 12164 17697 12173 17731
rect 12173 17697 12207 17731
rect 12207 17697 12216 17731
rect 12164 17688 12216 17697
rect 14004 17688 14056 17740
rect 15844 17688 15896 17740
rect 17592 17688 17644 17740
rect 18788 17731 18840 17740
rect 18788 17697 18797 17731
rect 18797 17697 18831 17731
rect 18831 17697 18840 17731
rect 18788 17688 18840 17697
rect 1584 17620 1636 17672
rect 2044 17663 2096 17672
rect 2044 17629 2053 17663
rect 2053 17629 2087 17663
rect 2087 17629 2096 17663
rect 2044 17620 2096 17629
rect 2320 17663 2372 17672
rect 2320 17629 2329 17663
rect 2329 17629 2363 17663
rect 2363 17629 2372 17663
rect 2320 17620 2372 17629
rect 2228 17552 2280 17604
rect 6828 17595 6880 17604
rect 6828 17561 6846 17595
rect 6846 17561 6880 17595
rect 7656 17620 7708 17672
rect 8024 17620 8076 17672
rect 8760 17620 8812 17672
rect 6828 17552 6880 17561
rect 1492 17527 1544 17536
rect 1492 17493 1501 17527
rect 1501 17493 1535 17527
rect 1535 17493 1544 17527
rect 1492 17484 1544 17493
rect 1860 17527 1912 17536
rect 1860 17493 1869 17527
rect 1869 17493 1903 17527
rect 1903 17493 1912 17527
rect 1860 17484 1912 17493
rect 5080 17484 5132 17536
rect 6644 17484 6696 17536
rect 8208 17552 8260 17604
rect 8576 17552 8628 17604
rect 9404 17552 9456 17604
rect 7748 17484 7800 17536
rect 11980 17552 12032 17604
rect 12624 17552 12676 17604
rect 9680 17484 9732 17536
rect 10140 17484 10192 17536
rect 10600 17484 10652 17536
rect 10968 17484 11020 17536
rect 11520 17527 11572 17536
rect 11520 17493 11529 17527
rect 11529 17493 11563 17527
rect 11563 17493 11572 17527
rect 11520 17484 11572 17493
rect 11796 17484 11848 17536
rect 12072 17484 12124 17536
rect 13728 17620 13780 17672
rect 15752 17663 15804 17672
rect 15752 17629 15761 17663
rect 15761 17629 15795 17663
rect 15795 17629 15804 17663
rect 15752 17620 15804 17629
rect 16304 17663 16356 17672
rect 16304 17629 16313 17663
rect 16313 17629 16347 17663
rect 16347 17629 16356 17663
rect 16304 17620 16356 17629
rect 18052 17620 18104 17672
rect 13176 17527 13228 17536
rect 13176 17493 13185 17527
rect 13185 17493 13219 17527
rect 13219 17493 13228 17527
rect 13176 17484 13228 17493
rect 14372 17527 14424 17536
rect 14372 17493 14381 17527
rect 14381 17493 14415 17527
rect 14415 17493 14424 17527
rect 14372 17484 14424 17493
rect 15476 17595 15528 17604
rect 15476 17561 15494 17595
rect 15494 17561 15528 17595
rect 15476 17552 15528 17561
rect 17684 17552 17736 17604
rect 18420 17620 18472 17672
rect 19800 17663 19852 17672
rect 19800 17629 19809 17663
rect 19809 17629 19843 17663
rect 19843 17629 19852 17663
rect 19800 17620 19852 17629
rect 20628 17620 20680 17672
rect 21272 17663 21324 17672
rect 21272 17629 21281 17663
rect 21281 17629 21315 17663
rect 21315 17629 21324 17663
rect 21272 17620 21324 17629
rect 16948 17527 17000 17536
rect 16948 17493 16957 17527
rect 16957 17493 16991 17527
rect 16991 17493 17000 17527
rect 16948 17484 17000 17493
rect 17224 17484 17276 17536
rect 17408 17527 17460 17536
rect 17408 17493 17417 17527
rect 17417 17493 17451 17527
rect 17451 17493 17460 17527
rect 17408 17484 17460 17493
rect 18144 17484 18196 17536
rect 21088 17527 21140 17536
rect 21088 17493 21097 17527
rect 21097 17493 21131 17527
rect 21131 17493 21140 17527
rect 21088 17484 21140 17493
rect 21456 17527 21508 17536
rect 21456 17493 21465 17527
rect 21465 17493 21499 17527
rect 21499 17493 21508 17527
rect 21456 17484 21508 17493
rect 6148 17382 6200 17434
rect 6212 17382 6264 17434
rect 6276 17382 6328 17434
rect 6340 17382 6392 17434
rect 6404 17382 6456 17434
rect 11346 17382 11398 17434
rect 11410 17382 11462 17434
rect 11474 17382 11526 17434
rect 11538 17382 11590 17434
rect 11602 17382 11654 17434
rect 16544 17382 16596 17434
rect 16608 17382 16660 17434
rect 16672 17382 16724 17434
rect 16736 17382 16788 17434
rect 16800 17382 16852 17434
rect 21742 17382 21794 17434
rect 21806 17382 21858 17434
rect 21870 17382 21922 17434
rect 21934 17382 21986 17434
rect 21998 17382 22050 17434
rect 4344 17280 4396 17332
rect 9404 17280 9456 17332
rect 9680 17323 9732 17332
rect 9680 17289 9689 17323
rect 9689 17289 9723 17323
rect 9723 17289 9732 17323
rect 9680 17280 9732 17289
rect 10692 17280 10744 17332
rect 11888 17280 11940 17332
rect 14556 17280 14608 17332
rect 14832 17280 14884 17332
rect 15844 17280 15896 17332
rect 16304 17280 16356 17332
rect 17684 17280 17736 17332
rect 19892 17323 19944 17332
rect 19892 17289 19901 17323
rect 19901 17289 19935 17323
rect 19935 17289 19944 17323
rect 19892 17280 19944 17289
rect 2228 17144 2280 17196
rect 4160 17187 4212 17196
rect 4160 17153 4169 17187
rect 4169 17153 4203 17187
rect 4203 17153 4212 17187
rect 4160 17144 4212 17153
rect 4712 17144 4764 17196
rect 5080 17187 5132 17196
rect 5080 17153 5114 17187
rect 5114 17153 5132 17187
rect 5080 17144 5132 17153
rect 5356 17144 5408 17196
rect 7564 17212 7616 17264
rect 11612 17212 11664 17264
rect 12072 17255 12124 17264
rect 12072 17221 12081 17255
rect 12081 17221 12115 17255
rect 12115 17221 12124 17255
rect 12072 17212 12124 17221
rect 17408 17212 17460 17264
rect 17776 17212 17828 17264
rect 6644 17187 6696 17196
rect 6644 17153 6653 17187
rect 6653 17153 6687 17187
rect 6687 17153 6696 17187
rect 6644 17144 6696 17153
rect 6736 17144 6788 17196
rect 1492 16983 1544 16992
rect 1492 16949 1501 16983
rect 1501 16949 1535 16983
rect 1535 16949 1544 16983
rect 1492 16940 1544 16949
rect 3240 16940 3292 16992
rect 8300 17144 8352 17196
rect 11796 17144 11848 17196
rect 11980 17187 12032 17196
rect 11980 17153 11989 17187
rect 11989 17153 12023 17187
rect 12023 17153 12032 17187
rect 11980 17144 12032 17153
rect 12440 17187 12492 17196
rect 12440 17153 12449 17187
rect 12449 17153 12483 17187
rect 12483 17153 12492 17187
rect 12440 17144 12492 17153
rect 13084 17144 13136 17196
rect 15200 17144 15252 17196
rect 15752 17144 15804 17196
rect 17040 17187 17092 17196
rect 17040 17153 17049 17187
rect 17049 17153 17083 17187
rect 17083 17153 17092 17187
rect 17040 17144 17092 17153
rect 17868 17187 17920 17196
rect 17868 17153 17877 17187
rect 17877 17153 17911 17187
rect 17911 17153 17920 17187
rect 17868 17144 17920 17153
rect 18236 17144 18288 17196
rect 20536 17144 20588 17196
rect 8208 17119 8260 17128
rect 8208 17085 8217 17119
rect 8217 17085 8251 17119
rect 8251 17085 8260 17119
rect 8208 17076 8260 17085
rect 9772 17076 9824 17128
rect 10232 17076 10284 17128
rect 10600 17119 10652 17128
rect 10600 17085 10609 17119
rect 10609 17085 10643 17119
rect 10643 17085 10652 17119
rect 10600 17076 10652 17085
rect 12164 17119 12216 17128
rect 12164 17085 12173 17119
rect 12173 17085 12207 17119
rect 12207 17085 12216 17119
rect 12164 17076 12216 17085
rect 15384 17076 15436 17128
rect 17132 17119 17184 17128
rect 6184 16983 6236 16992
rect 6184 16949 6193 16983
rect 6193 16949 6227 16983
rect 6227 16949 6236 16983
rect 6184 16940 6236 16949
rect 6552 16940 6604 16992
rect 6828 16940 6880 16992
rect 7932 16940 7984 16992
rect 10048 17008 10100 17060
rect 14004 17008 14056 17060
rect 17132 17085 17141 17119
rect 17141 17085 17175 17119
rect 17175 17085 17184 17119
rect 17132 17076 17184 17085
rect 17316 17119 17368 17128
rect 17316 17085 17325 17119
rect 17325 17085 17359 17119
rect 17359 17085 17368 17119
rect 17316 17076 17368 17085
rect 17684 17076 17736 17128
rect 10140 16940 10192 16992
rect 11152 16940 11204 16992
rect 13636 16940 13688 16992
rect 14556 16940 14608 16992
rect 19800 16940 19852 16992
rect 21456 16983 21508 16992
rect 21456 16949 21465 16983
rect 21465 16949 21499 16983
rect 21499 16949 21508 16983
rect 21456 16940 21508 16949
rect 3549 16838 3601 16890
rect 3613 16838 3665 16890
rect 3677 16838 3729 16890
rect 3741 16838 3793 16890
rect 3805 16838 3857 16890
rect 8747 16838 8799 16890
rect 8811 16838 8863 16890
rect 8875 16838 8927 16890
rect 8939 16838 8991 16890
rect 9003 16838 9055 16890
rect 13945 16838 13997 16890
rect 14009 16838 14061 16890
rect 14073 16838 14125 16890
rect 14137 16838 14189 16890
rect 14201 16838 14253 16890
rect 19143 16838 19195 16890
rect 19207 16838 19259 16890
rect 19271 16838 19323 16890
rect 19335 16838 19387 16890
rect 19399 16838 19451 16890
rect 2320 16736 2372 16788
rect 4160 16736 4212 16788
rect 6644 16736 6696 16788
rect 8208 16779 8260 16788
rect 8208 16745 8217 16779
rect 8217 16745 8251 16779
rect 8251 16745 8260 16779
rect 8208 16736 8260 16745
rect 2964 16668 3016 16720
rect 2872 16643 2924 16652
rect 2872 16609 2881 16643
rect 2881 16609 2915 16643
rect 2915 16609 2924 16643
rect 2872 16600 2924 16609
rect 5356 16600 5408 16652
rect 6552 16600 6604 16652
rect 11888 16736 11940 16788
rect 3240 16532 3292 16584
rect 4160 16532 4212 16584
rect 6184 16532 6236 16584
rect 10140 16532 10192 16584
rect 10876 16575 10928 16584
rect 10876 16541 10885 16575
rect 10885 16541 10919 16575
rect 10919 16541 10928 16575
rect 10876 16532 10928 16541
rect 11244 16532 11296 16584
rect 11796 16532 11848 16584
rect 13636 16736 13688 16788
rect 13728 16736 13780 16788
rect 13544 16711 13596 16720
rect 13544 16677 13553 16711
rect 13553 16677 13587 16711
rect 13587 16677 13596 16711
rect 13544 16668 13596 16677
rect 17868 16736 17920 16788
rect 18144 16736 18196 16788
rect 20628 16779 20680 16788
rect 20628 16745 20637 16779
rect 20637 16745 20671 16779
rect 20671 16745 20680 16779
rect 20628 16736 20680 16745
rect 13360 16575 13412 16584
rect 13360 16541 13369 16575
rect 13369 16541 13403 16575
rect 13403 16541 13412 16575
rect 13360 16532 13412 16541
rect 2320 16464 2372 16516
rect 4896 16464 4948 16516
rect 8392 16464 8444 16516
rect 10784 16464 10836 16516
rect 12348 16464 12400 16516
rect 16948 16668 17000 16720
rect 18788 16668 18840 16720
rect 13636 16532 13688 16584
rect 17500 16532 17552 16584
rect 18052 16600 18104 16652
rect 17684 16464 17736 16516
rect 18144 16532 18196 16584
rect 19616 16600 19668 16652
rect 1492 16439 1544 16448
rect 1492 16405 1501 16439
rect 1501 16405 1535 16439
rect 1535 16405 1544 16439
rect 1492 16396 1544 16405
rect 2412 16439 2464 16448
rect 2412 16405 2421 16439
rect 2421 16405 2455 16439
rect 2455 16405 2464 16439
rect 2412 16396 2464 16405
rect 8024 16439 8076 16448
rect 8024 16405 8033 16439
rect 8033 16405 8067 16439
rect 8067 16405 8076 16439
rect 8024 16396 8076 16405
rect 9220 16396 9272 16448
rect 11060 16439 11112 16448
rect 11060 16405 11069 16439
rect 11069 16405 11103 16439
rect 11103 16405 11112 16439
rect 11060 16396 11112 16405
rect 11244 16396 11296 16448
rect 15108 16396 15160 16448
rect 15384 16396 15436 16448
rect 16396 16439 16448 16448
rect 16396 16405 16405 16439
rect 16405 16405 16439 16439
rect 16439 16405 16448 16439
rect 16396 16396 16448 16405
rect 16488 16396 16540 16448
rect 17316 16396 17368 16448
rect 17776 16439 17828 16448
rect 17776 16405 17785 16439
rect 17785 16405 17819 16439
rect 17819 16405 17828 16439
rect 17776 16396 17828 16405
rect 18604 16439 18656 16448
rect 18604 16405 18613 16439
rect 18613 16405 18647 16439
rect 18647 16405 18656 16439
rect 20812 16532 20864 16584
rect 18604 16396 18656 16405
rect 20996 16439 21048 16448
rect 20996 16405 21005 16439
rect 21005 16405 21039 16439
rect 21039 16405 21048 16439
rect 21456 16439 21508 16448
rect 20996 16396 21048 16405
rect 21456 16405 21465 16439
rect 21465 16405 21499 16439
rect 21499 16405 21508 16439
rect 21456 16396 21508 16405
rect 6148 16294 6200 16346
rect 6212 16294 6264 16346
rect 6276 16294 6328 16346
rect 6340 16294 6392 16346
rect 6404 16294 6456 16346
rect 11346 16294 11398 16346
rect 11410 16294 11462 16346
rect 11474 16294 11526 16346
rect 11538 16294 11590 16346
rect 11602 16294 11654 16346
rect 16544 16294 16596 16346
rect 16608 16294 16660 16346
rect 16672 16294 16724 16346
rect 16736 16294 16788 16346
rect 16800 16294 16852 16346
rect 21742 16294 21794 16346
rect 21806 16294 21858 16346
rect 21870 16294 21922 16346
rect 21934 16294 21986 16346
rect 21998 16294 22050 16346
rect 2136 16235 2188 16244
rect 2136 16201 2145 16235
rect 2145 16201 2179 16235
rect 2179 16201 2188 16235
rect 2136 16192 2188 16201
rect 2320 16192 2372 16244
rect 4160 16192 4212 16244
rect 4712 16192 4764 16244
rect 3976 16124 4028 16176
rect 1492 15895 1544 15904
rect 1492 15861 1501 15895
rect 1501 15861 1535 15895
rect 1535 15861 1544 15895
rect 1492 15852 1544 15861
rect 1952 16056 2004 16108
rect 2320 16099 2372 16108
rect 2320 16065 2329 16099
rect 2329 16065 2363 16099
rect 2363 16065 2372 16099
rect 2320 16056 2372 16065
rect 2780 16099 2832 16108
rect 2780 16065 2789 16099
rect 2789 16065 2823 16099
rect 2823 16065 2832 16099
rect 2780 16056 2832 16065
rect 4068 16056 4120 16108
rect 5448 16056 5500 16108
rect 6644 16192 6696 16244
rect 11152 16192 11204 16244
rect 11336 16235 11388 16244
rect 11336 16201 11345 16235
rect 11345 16201 11379 16235
rect 11379 16201 11388 16235
rect 11336 16192 11388 16201
rect 11520 16192 11572 16244
rect 12716 16192 12768 16244
rect 13728 16235 13780 16244
rect 13728 16201 13737 16235
rect 13737 16201 13771 16235
rect 13771 16201 13780 16235
rect 13728 16192 13780 16201
rect 14648 16192 14700 16244
rect 15108 16192 15160 16244
rect 16304 16192 16356 16244
rect 16396 16192 16448 16244
rect 17224 16192 17276 16244
rect 17960 16192 18012 16244
rect 20536 16235 20588 16244
rect 11244 16124 11296 16176
rect 2964 16031 3016 16040
rect 2964 15997 2973 16031
rect 2973 15997 3007 16031
rect 3007 15997 3016 16031
rect 2964 15988 3016 15997
rect 1860 15963 1912 15972
rect 1860 15929 1869 15963
rect 1869 15929 1903 15963
rect 1903 15929 1912 15963
rect 1860 15920 1912 15929
rect 5356 16031 5408 16040
rect 5356 15997 5365 16031
rect 5365 15997 5399 16031
rect 5399 15997 5408 16031
rect 5356 15988 5408 15997
rect 6276 15988 6328 16040
rect 7196 16056 7248 16108
rect 8208 16056 8260 16108
rect 10048 16056 10100 16108
rect 10140 16056 10192 16108
rect 12072 16099 12124 16108
rect 12072 16065 12081 16099
rect 12081 16065 12115 16099
rect 12115 16065 12124 16099
rect 12072 16056 12124 16065
rect 9220 16031 9272 16040
rect 9220 15997 9229 16031
rect 9229 15997 9263 16031
rect 9263 15997 9272 16031
rect 9220 15988 9272 15997
rect 10692 16031 10744 16040
rect 6368 15920 6420 15972
rect 10692 15997 10701 16031
rect 10701 15997 10735 16031
rect 10735 15997 10744 16031
rect 10692 15988 10744 15997
rect 11980 15988 12032 16040
rect 16212 16124 16264 16176
rect 20536 16201 20545 16235
rect 20545 16201 20579 16235
rect 20579 16201 20588 16235
rect 20536 16192 20588 16201
rect 21180 16192 21232 16244
rect 22376 16124 22428 16176
rect 13728 16056 13780 16108
rect 13912 16056 13964 16108
rect 15476 16056 15528 16108
rect 18788 16056 18840 16108
rect 20260 16056 20312 16108
rect 20904 16099 20956 16108
rect 2320 15852 2372 15904
rect 2964 15852 3016 15904
rect 3332 15852 3384 15904
rect 7564 15852 7616 15904
rect 9864 15852 9916 15904
rect 10784 15852 10836 15904
rect 11612 15852 11664 15904
rect 12072 15852 12124 15904
rect 12900 15852 12952 15904
rect 13544 15852 13596 15904
rect 17040 15920 17092 15972
rect 17592 15988 17644 16040
rect 18144 16031 18196 16040
rect 18144 15997 18153 16031
rect 18153 15997 18187 16031
rect 18187 15997 18196 16031
rect 18144 15988 18196 15997
rect 20904 16065 20913 16099
rect 20913 16065 20947 16099
rect 20947 16065 20956 16099
rect 20904 16056 20956 16065
rect 21364 16056 21416 16108
rect 18604 15963 18656 15972
rect 18604 15929 18613 15963
rect 18613 15929 18647 15963
rect 18647 15929 18656 15963
rect 18604 15920 18656 15929
rect 21088 15963 21140 15972
rect 21088 15929 21097 15963
rect 21097 15929 21131 15963
rect 21131 15929 21140 15963
rect 21088 15920 21140 15929
rect 15200 15895 15252 15904
rect 15200 15861 15209 15895
rect 15209 15861 15243 15895
rect 15243 15861 15252 15895
rect 15200 15852 15252 15861
rect 15752 15852 15804 15904
rect 20168 15895 20220 15904
rect 20168 15861 20177 15895
rect 20177 15861 20211 15895
rect 20211 15861 20220 15895
rect 20168 15852 20220 15861
rect 21456 15895 21508 15904
rect 21456 15861 21465 15895
rect 21465 15861 21499 15895
rect 21499 15861 21508 15895
rect 21456 15852 21508 15861
rect 3549 15750 3601 15802
rect 3613 15750 3665 15802
rect 3677 15750 3729 15802
rect 3741 15750 3793 15802
rect 3805 15750 3857 15802
rect 8747 15750 8799 15802
rect 8811 15750 8863 15802
rect 8875 15750 8927 15802
rect 8939 15750 8991 15802
rect 9003 15750 9055 15802
rect 13945 15750 13997 15802
rect 14009 15750 14061 15802
rect 14073 15750 14125 15802
rect 14137 15750 14189 15802
rect 14201 15750 14253 15802
rect 19143 15750 19195 15802
rect 19207 15750 19259 15802
rect 19271 15750 19323 15802
rect 19335 15750 19387 15802
rect 19399 15750 19451 15802
rect 1952 15691 2004 15700
rect 1952 15657 1961 15691
rect 1961 15657 1995 15691
rect 1995 15657 2004 15691
rect 1952 15648 2004 15657
rect 2228 15691 2280 15700
rect 2228 15657 2237 15691
rect 2237 15657 2271 15691
rect 2271 15657 2280 15691
rect 2228 15648 2280 15657
rect 5448 15691 5500 15700
rect 5448 15657 5457 15691
rect 5457 15657 5491 15691
rect 5491 15657 5500 15691
rect 5448 15648 5500 15657
rect 6276 15691 6328 15700
rect 6276 15657 6285 15691
rect 6285 15657 6319 15691
rect 6319 15657 6328 15691
rect 6276 15648 6328 15657
rect 6368 15648 6420 15700
rect 10048 15691 10100 15700
rect 10048 15657 10057 15691
rect 10057 15657 10091 15691
rect 10091 15657 10100 15691
rect 10048 15648 10100 15657
rect 10876 15691 10928 15700
rect 10876 15657 10885 15691
rect 10885 15657 10919 15691
rect 10919 15657 10928 15691
rect 10876 15648 10928 15657
rect 11060 15648 11112 15700
rect 11980 15691 12032 15700
rect 2044 15580 2096 15632
rect 5448 15512 5500 15564
rect 6552 15512 6604 15564
rect 1676 15487 1728 15496
rect 1676 15453 1685 15487
rect 1685 15453 1719 15487
rect 1719 15453 1728 15487
rect 1676 15444 1728 15453
rect 2412 15487 2464 15496
rect 2412 15453 2421 15487
rect 2421 15453 2455 15487
rect 2455 15453 2464 15487
rect 2412 15444 2464 15453
rect 4620 15376 4672 15428
rect 6644 15444 6696 15496
rect 6552 15376 6604 15428
rect 7748 15376 7800 15428
rect 1492 15351 1544 15360
rect 1492 15317 1501 15351
rect 1501 15317 1535 15351
rect 1535 15317 1544 15351
rect 1492 15308 1544 15317
rect 4528 15351 4580 15360
rect 4528 15317 4537 15351
rect 4537 15317 4571 15351
rect 4571 15317 4580 15351
rect 4528 15308 4580 15317
rect 11520 15580 11572 15632
rect 7932 15512 7984 15564
rect 10232 15512 10284 15564
rect 11336 15555 11388 15564
rect 11336 15521 11345 15555
rect 11345 15521 11379 15555
rect 11379 15521 11388 15555
rect 11336 15512 11388 15521
rect 9312 15487 9364 15496
rect 9312 15453 9321 15487
rect 9321 15453 9355 15487
rect 9355 15453 9364 15487
rect 9312 15444 9364 15453
rect 8208 15376 8260 15428
rect 10140 15444 10192 15496
rect 11060 15444 11112 15496
rect 11980 15657 11989 15691
rect 11989 15657 12023 15691
rect 12023 15657 12032 15691
rect 11980 15648 12032 15657
rect 13728 15648 13780 15700
rect 12164 15512 12216 15564
rect 13084 15512 13136 15564
rect 15476 15648 15528 15700
rect 12348 15487 12400 15496
rect 12072 15376 12124 15428
rect 9864 15308 9916 15360
rect 10600 15308 10652 15360
rect 11612 15308 11664 15360
rect 11888 15308 11940 15360
rect 12348 15453 12357 15487
rect 12357 15453 12391 15487
rect 12391 15453 12400 15487
rect 12348 15444 12400 15453
rect 17132 15648 17184 15700
rect 18144 15648 18196 15700
rect 20260 15691 20312 15700
rect 20260 15657 20269 15691
rect 20269 15657 20303 15691
rect 20303 15657 20312 15691
rect 20260 15648 20312 15657
rect 21272 15648 21324 15700
rect 21548 15648 21600 15700
rect 16948 15487 17000 15496
rect 16948 15453 16957 15487
rect 16957 15453 16991 15487
rect 16991 15453 17000 15487
rect 16948 15444 17000 15453
rect 21640 15580 21692 15632
rect 17592 15555 17644 15564
rect 17592 15521 17601 15555
rect 17601 15521 17635 15555
rect 17635 15521 17644 15555
rect 17592 15512 17644 15521
rect 14372 15419 14424 15428
rect 14372 15385 14406 15419
rect 14406 15385 14424 15419
rect 14372 15376 14424 15385
rect 17960 15444 18012 15496
rect 20996 15444 21048 15496
rect 18144 15376 18196 15428
rect 18880 15376 18932 15428
rect 20720 15376 20772 15428
rect 18420 15308 18472 15360
rect 22100 15376 22152 15428
rect 6148 15206 6200 15258
rect 6212 15206 6264 15258
rect 6276 15206 6328 15258
rect 6340 15206 6392 15258
rect 6404 15206 6456 15258
rect 11346 15206 11398 15258
rect 11410 15206 11462 15258
rect 11474 15206 11526 15258
rect 11538 15206 11590 15258
rect 11602 15206 11654 15258
rect 16544 15206 16596 15258
rect 16608 15206 16660 15258
rect 16672 15206 16724 15258
rect 16736 15206 16788 15258
rect 16800 15206 16852 15258
rect 21742 15206 21794 15258
rect 21806 15206 21858 15258
rect 21870 15206 21922 15258
rect 21934 15206 21986 15258
rect 21998 15206 22050 15258
rect 1676 15104 1728 15156
rect 2412 15104 2464 15156
rect 4436 15104 4488 15156
rect 4528 15104 4580 15156
rect 6644 15147 6696 15156
rect 6644 15113 6653 15147
rect 6653 15113 6687 15147
rect 6687 15113 6696 15147
rect 6644 15104 6696 15113
rect 1952 15011 2004 15020
rect 1952 14977 1961 15011
rect 1961 14977 1995 15011
rect 1995 14977 2004 15011
rect 1952 14968 2004 14977
rect 5080 15036 5132 15088
rect 6552 15036 6604 15088
rect 2780 14968 2832 15020
rect 4344 15011 4396 15020
rect 2504 14832 2556 14884
rect 4344 14977 4353 15011
rect 4353 14977 4387 15011
rect 4387 14977 4396 15011
rect 4344 14968 4396 14977
rect 7564 14968 7616 15020
rect 8024 14968 8076 15020
rect 9128 15104 9180 15156
rect 8576 15079 8628 15088
rect 8576 15045 8585 15079
rect 8585 15045 8619 15079
rect 8619 15045 8628 15079
rect 8576 15036 8628 15045
rect 8208 14968 8260 15020
rect 11336 15104 11388 15156
rect 13728 15147 13780 15156
rect 13728 15113 13737 15147
rect 13737 15113 13771 15147
rect 13771 15113 13780 15147
rect 13728 15104 13780 15113
rect 10324 14968 10376 15020
rect 12808 14968 12860 15020
rect 13728 14968 13780 15020
rect 15476 15104 15528 15156
rect 16948 15104 17000 15156
rect 20720 15147 20772 15156
rect 20720 15113 20729 15147
rect 20729 15113 20763 15147
rect 20763 15113 20772 15147
rect 20720 15104 20772 15113
rect 20904 15104 20956 15156
rect 18144 15036 18196 15088
rect 5356 14943 5408 14952
rect 5356 14909 5365 14943
rect 5365 14909 5399 14943
rect 5399 14909 5408 14943
rect 5356 14900 5408 14909
rect 18972 15011 19024 15020
rect 18972 14977 18981 15011
rect 18981 14977 19015 15011
rect 19015 14977 19024 15011
rect 18972 14968 19024 14977
rect 19524 14968 19576 15020
rect 4896 14832 4948 14884
rect 5540 14832 5592 14884
rect 1492 14807 1544 14816
rect 1492 14773 1501 14807
rect 1501 14773 1535 14807
rect 1535 14773 1544 14807
rect 1492 14764 1544 14773
rect 4160 14764 4212 14816
rect 6736 14807 6788 14816
rect 6736 14773 6745 14807
rect 6745 14773 6779 14807
rect 6779 14773 6788 14807
rect 6736 14764 6788 14773
rect 8116 14832 8168 14884
rect 15384 14900 15436 14952
rect 15752 14900 15804 14952
rect 17224 14943 17276 14952
rect 17224 14909 17233 14943
rect 17233 14909 17267 14943
rect 17267 14909 17276 14943
rect 17224 14900 17276 14909
rect 19064 14943 19116 14952
rect 19064 14909 19073 14943
rect 19073 14909 19107 14943
rect 19107 14909 19116 14943
rect 19064 14900 19116 14909
rect 20904 14968 20956 15020
rect 11704 14832 11756 14884
rect 17960 14832 18012 14884
rect 18696 14832 18748 14884
rect 8300 14764 8352 14816
rect 8668 14764 8720 14816
rect 11520 14807 11572 14816
rect 11520 14773 11529 14807
rect 11529 14773 11563 14807
rect 11563 14773 11572 14807
rect 11520 14764 11572 14773
rect 12992 14764 13044 14816
rect 21180 14807 21232 14816
rect 21180 14773 21189 14807
rect 21189 14773 21223 14807
rect 21223 14773 21232 14807
rect 21180 14764 21232 14773
rect 21456 14807 21508 14816
rect 21456 14773 21465 14807
rect 21465 14773 21499 14807
rect 21499 14773 21508 14807
rect 21456 14764 21508 14773
rect 3549 14662 3601 14714
rect 3613 14662 3665 14714
rect 3677 14662 3729 14714
rect 3741 14662 3793 14714
rect 3805 14662 3857 14714
rect 8747 14662 8799 14714
rect 8811 14662 8863 14714
rect 8875 14662 8927 14714
rect 8939 14662 8991 14714
rect 9003 14662 9055 14714
rect 13945 14662 13997 14714
rect 14009 14662 14061 14714
rect 14073 14662 14125 14714
rect 14137 14662 14189 14714
rect 14201 14662 14253 14714
rect 19143 14662 19195 14714
rect 19207 14662 19259 14714
rect 19271 14662 19323 14714
rect 19335 14662 19387 14714
rect 19399 14662 19451 14714
rect 1952 14560 2004 14612
rect 4344 14560 4396 14612
rect 4712 14492 4764 14544
rect 5356 14492 5408 14544
rect 5448 14424 5500 14476
rect 7748 14560 7800 14612
rect 9128 14603 9180 14612
rect 9128 14569 9137 14603
rect 9137 14569 9171 14603
rect 9171 14569 9180 14603
rect 9128 14560 9180 14569
rect 11060 14560 11112 14612
rect 11336 14603 11388 14612
rect 11336 14569 11345 14603
rect 11345 14569 11379 14603
rect 11379 14569 11388 14603
rect 11336 14560 11388 14569
rect 13728 14560 13780 14612
rect 14372 14560 14424 14612
rect 8576 14424 8628 14476
rect 13912 14492 13964 14544
rect 15476 14467 15528 14476
rect 1768 14356 1820 14408
rect 2044 14399 2096 14408
rect 2044 14365 2053 14399
rect 2053 14365 2087 14399
rect 2087 14365 2096 14399
rect 2044 14356 2096 14365
rect 3424 14356 3476 14408
rect 4160 14399 4212 14408
rect 4160 14365 4169 14399
rect 4169 14365 4203 14399
rect 4203 14365 4212 14399
rect 4160 14356 4212 14365
rect 5540 14399 5592 14408
rect 5540 14365 5549 14399
rect 5549 14365 5583 14399
rect 5583 14365 5592 14399
rect 5540 14356 5592 14365
rect 6644 14356 6696 14408
rect 7472 14356 7524 14408
rect 8300 14356 8352 14408
rect 15476 14433 15485 14467
rect 15485 14433 15519 14467
rect 15519 14433 15528 14467
rect 15476 14424 15528 14433
rect 17224 14560 17276 14612
rect 19064 14560 19116 14612
rect 18696 14424 18748 14476
rect 20996 14560 21048 14612
rect 19800 14467 19852 14476
rect 1492 14263 1544 14272
rect 1492 14229 1501 14263
rect 1501 14229 1535 14263
rect 1535 14229 1544 14263
rect 1492 14220 1544 14229
rect 1860 14263 1912 14272
rect 1860 14229 1869 14263
rect 1869 14229 1903 14263
rect 1903 14229 1912 14263
rect 1860 14220 1912 14229
rect 4528 14220 4580 14272
rect 5356 14220 5408 14272
rect 6000 14263 6052 14272
rect 6000 14229 6009 14263
rect 6009 14229 6043 14263
rect 6043 14229 6052 14263
rect 6000 14220 6052 14229
rect 6736 14288 6788 14340
rect 10048 14288 10100 14340
rect 10692 14288 10744 14340
rect 9404 14220 9456 14272
rect 11520 14288 11572 14340
rect 15568 14356 15620 14408
rect 16396 14356 16448 14408
rect 16028 14288 16080 14340
rect 19064 14356 19116 14408
rect 19800 14433 19809 14467
rect 19809 14433 19843 14467
rect 19843 14433 19852 14467
rect 19800 14424 19852 14433
rect 20628 14399 20680 14408
rect 20628 14365 20637 14399
rect 20637 14365 20671 14399
rect 20671 14365 20680 14399
rect 20628 14356 20680 14365
rect 20996 14356 21048 14408
rect 17868 14220 17920 14272
rect 18512 14288 18564 14340
rect 19524 14220 19576 14272
rect 20076 14263 20128 14272
rect 20076 14229 20085 14263
rect 20085 14229 20119 14263
rect 20119 14229 20128 14263
rect 20076 14220 20128 14229
rect 21088 14263 21140 14272
rect 21088 14229 21097 14263
rect 21097 14229 21131 14263
rect 21131 14229 21140 14263
rect 21088 14220 21140 14229
rect 21456 14263 21508 14272
rect 21456 14229 21465 14263
rect 21465 14229 21499 14263
rect 21499 14229 21508 14263
rect 21456 14220 21508 14229
rect 6148 14118 6200 14170
rect 6212 14118 6264 14170
rect 6276 14118 6328 14170
rect 6340 14118 6392 14170
rect 6404 14118 6456 14170
rect 11346 14118 11398 14170
rect 11410 14118 11462 14170
rect 11474 14118 11526 14170
rect 11538 14118 11590 14170
rect 11602 14118 11654 14170
rect 16544 14118 16596 14170
rect 16608 14118 16660 14170
rect 16672 14118 16724 14170
rect 16736 14118 16788 14170
rect 16800 14118 16852 14170
rect 21742 14118 21794 14170
rect 21806 14118 21858 14170
rect 21870 14118 21922 14170
rect 21934 14118 21986 14170
rect 21998 14118 22050 14170
rect 1584 14016 1636 14068
rect 4528 14059 4580 14068
rect 4528 14025 4537 14059
rect 4537 14025 4571 14059
rect 4571 14025 4580 14059
rect 4528 14016 4580 14025
rect 4896 14059 4948 14068
rect 4896 14025 4905 14059
rect 4905 14025 4939 14059
rect 4939 14025 4948 14059
rect 4896 14016 4948 14025
rect 5356 14059 5408 14068
rect 5356 14025 5365 14059
rect 5365 14025 5399 14059
rect 5399 14025 5408 14059
rect 5356 14016 5408 14025
rect 6184 14059 6236 14068
rect 6184 14025 6193 14059
rect 6193 14025 6227 14059
rect 6227 14025 6236 14059
rect 6184 14016 6236 14025
rect 4988 13948 5040 14000
rect 1676 13923 1728 13932
rect 1676 13889 1685 13923
rect 1685 13889 1719 13923
rect 1719 13889 1728 13923
rect 1676 13880 1728 13889
rect 4160 13923 4212 13932
rect 1492 13719 1544 13728
rect 1492 13685 1501 13719
rect 1501 13685 1535 13719
rect 1535 13685 1544 13719
rect 1492 13676 1544 13685
rect 4160 13889 4169 13923
rect 4169 13889 4203 13923
rect 4203 13889 4212 13923
rect 4160 13880 4212 13889
rect 6092 13880 6144 13932
rect 6644 14016 6696 14068
rect 6644 13923 6696 13932
rect 6644 13889 6678 13923
rect 6678 13889 6696 13923
rect 6644 13880 6696 13889
rect 8484 13923 8536 13932
rect 8484 13889 8493 13923
rect 8493 13889 8527 13923
rect 8527 13889 8536 13923
rect 8484 13880 8536 13889
rect 8576 13880 8628 13932
rect 11060 13948 11112 14000
rect 13360 14016 13412 14068
rect 13728 14016 13780 14068
rect 5448 13855 5500 13864
rect 5448 13821 5457 13855
rect 5457 13821 5491 13855
rect 5491 13821 5500 13855
rect 5448 13812 5500 13821
rect 13820 13948 13872 14000
rect 13912 13880 13964 13932
rect 14280 14016 14332 14068
rect 15016 14016 15068 14068
rect 16396 14016 16448 14068
rect 18236 14059 18288 14068
rect 18236 14025 18245 14059
rect 18245 14025 18279 14059
rect 18279 14025 18288 14059
rect 18236 14016 18288 14025
rect 18880 14016 18932 14068
rect 19064 14059 19116 14068
rect 19064 14025 19073 14059
rect 19073 14025 19107 14059
rect 19107 14025 19116 14059
rect 19064 14016 19116 14025
rect 16580 13948 16632 14000
rect 14464 13923 14516 13932
rect 14464 13889 14498 13923
rect 14498 13889 14516 13923
rect 14464 13880 14516 13889
rect 15016 13880 15068 13932
rect 16948 13880 17000 13932
rect 15844 13855 15896 13864
rect 4712 13744 4764 13796
rect 15844 13821 15853 13855
rect 15853 13821 15887 13855
rect 15887 13821 15896 13855
rect 15844 13812 15896 13821
rect 17132 13855 17184 13864
rect 17132 13821 17141 13855
rect 17141 13821 17175 13855
rect 17175 13821 17184 13855
rect 17132 13812 17184 13821
rect 18236 13880 18288 13932
rect 18972 13948 19024 14000
rect 20076 14016 20128 14068
rect 7564 13676 7616 13728
rect 7748 13719 7800 13728
rect 7748 13685 7757 13719
rect 7757 13685 7791 13719
rect 7791 13685 7800 13719
rect 7748 13676 7800 13685
rect 7932 13676 7984 13728
rect 10324 13676 10376 13728
rect 13176 13744 13228 13796
rect 15752 13744 15804 13796
rect 18144 13812 18196 13864
rect 18604 13855 18656 13864
rect 17684 13744 17736 13796
rect 18604 13821 18613 13855
rect 18613 13821 18647 13855
rect 18647 13821 18656 13855
rect 18604 13812 18656 13821
rect 19800 13880 19852 13932
rect 21272 13923 21324 13932
rect 21272 13889 21281 13923
rect 21281 13889 21315 13923
rect 21315 13889 21324 13923
rect 21272 13880 21324 13889
rect 18972 13744 19024 13796
rect 11704 13676 11756 13728
rect 12440 13676 12492 13728
rect 15476 13676 15528 13728
rect 16028 13719 16080 13728
rect 16028 13685 16037 13719
rect 16037 13685 16071 13719
rect 16071 13685 16080 13719
rect 16028 13676 16080 13685
rect 21548 13744 21600 13796
rect 19708 13676 19760 13728
rect 21456 13719 21508 13728
rect 21456 13685 21465 13719
rect 21465 13685 21499 13719
rect 21499 13685 21508 13719
rect 21456 13676 21508 13685
rect 3549 13574 3601 13626
rect 3613 13574 3665 13626
rect 3677 13574 3729 13626
rect 3741 13574 3793 13626
rect 3805 13574 3857 13626
rect 8747 13574 8799 13626
rect 8811 13574 8863 13626
rect 8875 13574 8927 13626
rect 8939 13574 8991 13626
rect 9003 13574 9055 13626
rect 13945 13574 13997 13626
rect 14009 13574 14061 13626
rect 14073 13574 14125 13626
rect 14137 13574 14189 13626
rect 14201 13574 14253 13626
rect 19143 13574 19195 13626
rect 19207 13574 19259 13626
rect 19271 13574 19323 13626
rect 19335 13574 19387 13626
rect 19399 13574 19451 13626
rect 1676 13472 1728 13524
rect 2780 13472 2832 13524
rect 5540 13472 5592 13524
rect 6184 13515 6236 13524
rect 6184 13481 6193 13515
rect 6193 13481 6227 13515
rect 6227 13481 6236 13515
rect 6184 13472 6236 13481
rect 3056 13404 3108 13456
rect 6092 13404 6144 13456
rect 8484 13472 8536 13524
rect 5632 13336 5684 13388
rect 6000 13336 6052 13388
rect 7748 13379 7800 13388
rect 7748 13345 7757 13379
rect 7757 13345 7791 13379
rect 7791 13345 7800 13379
rect 7748 13336 7800 13345
rect 7932 13336 7984 13388
rect 10324 13447 10376 13456
rect 10324 13413 10333 13447
rect 10333 13413 10367 13447
rect 10367 13413 10376 13447
rect 10324 13404 10376 13413
rect 1400 13311 1452 13320
rect 1400 13277 1409 13311
rect 1409 13277 1443 13311
rect 1443 13277 1452 13311
rect 1400 13268 1452 13277
rect 2320 13268 2372 13320
rect 3976 13268 4028 13320
rect 5356 13200 5408 13252
rect 7104 13200 7156 13252
rect 2228 13175 2280 13184
rect 2228 13141 2237 13175
rect 2237 13141 2271 13175
rect 2271 13141 2280 13175
rect 2228 13132 2280 13141
rect 4436 13175 4488 13184
rect 4436 13141 4445 13175
rect 4445 13141 4479 13175
rect 4479 13141 4488 13175
rect 4436 13132 4488 13141
rect 5448 13132 5500 13184
rect 6828 13132 6880 13184
rect 8116 13268 8168 13320
rect 8208 13268 8260 13320
rect 7288 13200 7340 13252
rect 9772 13268 9824 13320
rect 13176 13472 13228 13524
rect 18236 13515 18288 13524
rect 14372 13379 14424 13388
rect 14372 13345 14381 13379
rect 14381 13345 14415 13379
rect 14415 13345 14424 13379
rect 14372 13336 14424 13345
rect 12716 13311 12768 13320
rect 12716 13277 12725 13311
rect 12725 13277 12759 13311
rect 12759 13277 12768 13311
rect 12716 13268 12768 13277
rect 16580 13404 16632 13456
rect 15476 13379 15528 13388
rect 15476 13345 15485 13379
rect 15485 13345 15519 13379
rect 15519 13345 15528 13379
rect 15476 13336 15528 13345
rect 15568 13379 15620 13388
rect 15568 13345 15577 13379
rect 15577 13345 15611 13379
rect 15611 13345 15620 13379
rect 18236 13481 18245 13515
rect 18245 13481 18279 13515
rect 18279 13481 18288 13515
rect 18236 13472 18288 13481
rect 20996 13515 21048 13524
rect 20996 13481 21005 13515
rect 21005 13481 21039 13515
rect 21039 13481 21048 13515
rect 20996 13472 21048 13481
rect 21364 13472 21416 13524
rect 15568 13336 15620 13345
rect 17592 13379 17644 13388
rect 17592 13345 17601 13379
rect 17601 13345 17635 13379
rect 17635 13345 17644 13379
rect 17592 13336 17644 13345
rect 18972 13379 19024 13388
rect 18972 13345 18981 13379
rect 18981 13345 19015 13379
rect 19015 13345 19024 13379
rect 18972 13336 19024 13345
rect 15844 13268 15896 13320
rect 17868 13311 17920 13320
rect 17868 13277 17877 13311
rect 17877 13277 17911 13311
rect 17911 13277 17920 13311
rect 17868 13268 17920 13277
rect 18696 13268 18748 13320
rect 7564 13132 7616 13184
rect 8300 13132 8352 13184
rect 9680 13132 9732 13184
rect 9772 13132 9824 13184
rect 11244 13132 11296 13184
rect 11704 13200 11756 13252
rect 12348 13200 12400 13252
rect 12256 13132 12308 13184
rect 13176 13175 13228 13184
rect 13176 13141 13185 13175
rect 13185 13141 13219 13175
rect 13219 13141 13228 13175
rect 13176 13132 13228 13141
rect 14924 13175 14976 13184
rect 14924 13141 14933 13175
rect 14933 13141 14967 13175
rect 14967 13141 14976 13175
rect 14924 13132 14976 13141
rect 21364 13336 21416 13388
rect 15568 13132 15620 13184
rect 16028 13132 16080 13184
rect 17040 13175 17092 13184
rect 17040 13141 17049 13175
rect 17049 13141 17083 13175
rect 17083 13141 17092 13175
rect 17040 13132 17092 13141
rect 17132 13175 17184 13184
rect 17132 13141 17141 13175
rect 17141 13141 17175 13175
rect 17175 13141 17184 13175
rect 17776 13175 17828 13184
rect 17132 13132 17184 13141
rect 17776 13141 17785 13175
rect 17785 13141 17819 13175
rect 17819 13141 17828 13175
rect 17776 13132 17828 13141
rect 21548 13311 21600 13320
rect 21548 13277 21557 13311
rect 21557 13277 21591 13311
rect 21591 13277 21600 13311
rect 21548 13268 21600 13277
rect 20812 13132 20864 13184
rect 21640 13132 21692 13184
rect 6148 13030 6200 13082
rect 6212 13030 6264 13082
rect 6276 13030 6328 13082
rect 6340 13030 6392 13082
rect 6404 13030 6456 13082
rect 11346 13030 11398 13082
rect 11410 13030 11462 13082
rect 11474 13030 11526 13082
rect 11538 13030 11590 13082
rect 11602 13030 11654 13082
rect 16544 13030 16596 13082
rect 16608 13030 16660 13082
rect 16672 13030 16724 13082
rect 16736 13030 16788 13082
rect 16800 13030 16852 13082
rect 21742 13030 21794 13082
rect 21806 13030 21858 13082
rect 21870 13030 21922 13082
rect 21934 13030 21986 13082
rect 21998 13030 22050 13082
rect 2320 12971 2372 12980
rect 2320 12937 2329 12971
rect 2329 12937 2363 12971
rect 2363 12937 2372 12971
rect 2320 12928 2372 12937
rect 5540 12928 5592 12980
rect 6000 12928 6052 12980
rect 6828 12928 6880 12980
rect 8300 12971 8352 12980
rect 2504 12835 2556 12844
rect 2504 12801 2513 12835
rect 2513 12801 2547 12835
rect 2547 12801 2556 12835
rect 2504 12792 2556 12801
rect 3056 12835 3108 12844
rect 3056 12801 3065 12835
rect 3065 12801 3099 12835
rect 3099 12801 3108 12835
rect 3056 12792 3108 12801
rect 3148 12792 3200 12844
rect 2228 12767 2280 12776
rect 2228 12733 2237 12767
rect 2237 12733 2271 12767
rect 2271 12733 2280 12767
rect 2228 12724 2280 12733
rect 5356 12792 5408 12844
rect 4896 12767 4948 12776
rect 3424 12656 3476 12708
rect 3976 12588 4028 12640
rect 4896 12733 4905 12767
rect 4905 12733 4939 12767
rect 4939 12733 4948 12767
rect 4896 12724 4948 12733
rect 5448 12699 5500 12708
rect 5448 12665 5457 12699
rect 5457 12665 5491 12699
rect 5491 12665 5500 12699
rect 5448 12656 5500 12665
rect 7012 12860 7064 12912
rect 7196 12860 7248 12912
rect 6368 12792 6420 12844
rect 7748 12835 7800 12844
rect 7748 12801 7757 12835
rect 7757 12801 7791 12835
rect 7791 12801 7800 12835
rect 7748 12792 7800 12801
rect 8300 12937 8309 12971
rect 8309 12937 8343 12971
rect 8343 12937 8352 12971
rect 8300 12928 8352 12937
rect 8668 12928 8720 12980
rect 9496 12971 9548 12980
rect 9496 12937 9505 12971
rect 9505 12937 9539 12971
rect 9539 12937 9548 12971
rect 9496 12928 9548 12937
rect 9680 12928 9732 12980
rect 9772 12928 9824 12980
rect 8760 12903 8812 12912
rect 8760 12869 8769 12903
rect 8769 12869 8803 12903
rect 8803 12869 8812 12903
rect 8760 12860 8812 12869
rect 10140 12928 10192 12980
rect 11244 12928 11296 12980
rect 11888 12971 11940 12980
rect 11888 12937 11897 12971
rect 11897 12937 11931 12971
rect 11931 12937 11940 12971
rect 12256 12971 12308 12980
rect 11888 12928 11940 12937
rect 12256 12937 12265 12971
rect 12265 12937 12299 12971
rect 12299 12937 12308 12971
rect 12256 12928 12308 12937
rect 12624 12928 12676 12980
rect 17040 12928 17092 12980
rect 18604 12928 18656 12980
rect 20720 12928 20772 12980
rect 20996 12971 21048 12980
rect 20996 12937 21005 12971
rect 21005 12937 21039 12971
rect 21039 12937 21048 12971
rect 20996 12928 21048 12937
rect 12440 12860 12492 12912
rect 6092 12767 6144 12776
rect 6092 12733 6101 12767
rect 6101 12733 6135 12767
rect 6135 12733 6144 12767
rect 6092 12724 6144 12733
rect 7840 12724 7892 12776
rect 9312 12792 9364 12844
rect 6276 12588 6328 12640
rect 9404 12767 9456 12776
rect 9404 12733 9413 12767
rect 9413 12733 9447 12767
rect 9447 12733 9456 12767
rect 9404 12724 9456 12733
rect 10140 12767 10192 12776
rect 10140 12733 10149 12767
rect 10149 12733 10183 12767
rect 10183 12733 10192 12767
rect 10140 12724 10192 12733
rect 12164 12792 12216 12844
rect 11704 12767 11756 12776
rect 11704 12733 11713 12767
rect 11713 12733 11747 12767
rect 11747 12733 11756 12767
rect 11704 12724 11756 12733
rect 11888 12724 11940 12776
rect 12716 12835 12768 12844
rect 12716 12801 12725 12835
rect 12725 12801 12759 12835
rect 12759 12801 12768 12835
rect 16212 12903 16264 12912
rect 12716 12792 12768 12801
rect 12992 12835 13044 12844
rect 12992 12801 13026 12835
rect 13026 12801 13044 12835
rect 12992 12792 13044 12801
rect 13360 12792 13412 12844
rect 15752 12835 15804 12844
rect 16212 12869 16221 12903
rect 16221 12869 16255 12903
rect 16255 12869 16264 12903
rect 16212 12860 16264 12869
rect 15752 12801 15770 12835
rect 15770 12801 15804 12835
rect 15752 12792 15804 12801
rect 17500 12792 17552 12844
rect 16764 12767 16816 12776
rect 16764 12733 16773 12767
rect 16773 12733 16807 12767
rect 16807 12733 16816 12767
rect 16764 12724 16816 12733
rect 18972 12792 19024 12844
rect 19524 12792 19576 12844
rect 21088 12835 21140 12844
rect 21088 12801 21097 12835
rect 21097 12801 21131 12835
rect 21131 12801 21140 12835
rect 21088 12792 21140 12801
rect 21456 12835 21508 12844
rect 21456 12801 21465 12835
rect 21465 12801 21499 12835
rect 21499 12801 21508 12835
rect 21456 12792 21508 12801
rect 18420 12767 18472 12776
rect 18420 12733 18429 12767
rect 18429 12733 18463 12767
rect 18463 12733 18472 12767
rect 18420 12724 18472 12733
rect 20260 12767 20312 12776
rect 8300 12588 8352 12640
rect 9496 12588 9548 12640
rect 9680 12588 9732 12640
rect 10968 12588 11020 12640
rect 12624 12656 12676 12708
rect 12164 12588 12216 12640
rect 12900 12588 12952 12640
rect 13636 12588 13688 12640
rect 14464 12588 14516 12640
rect 17040 12656 17092 12708
rect 20260 12733 20269 12767
rect 20269 12733 20303 12767
rect 20303 12733 20312 12767
rect 20260 12724 20312 12733
rect 20720 12656 20772 12708
rect 17592 12588 17644 12640
rect 3549 12486 3601 12538
rect 3613 12486 3665 12538
rect 3677 12486 3729 12538
rect 3741 12486 3793 12538
rect 3805 12486 3857 12538
rect 8747 12486 8799 12538
rect 8811 12486 8863 12538
rect 8875 12486 8927 12538
rect 8939 12486 8991 12538
rect 9003 12486 9055 12538
rect 13945 12486 13997 12538
rect 14009 12486 14061 12538
rect 14073 12486 14125 12538
rect 14137 12486 14189 12538
rect 14201 12486 14253 12538
rect 19143 12486 19195 12538
rect 19207 12486 19259 12538
rect 19271 12486 19323 12538
rect 19335 12486 19387 12538
rect 19399 12486 19451 12538
rect 2044 12384 2096 12436
rect 3056 12384 3108 12436
rect 3884 12427 3936 12436
rect 1676 12359 1728 12368
rect 1676 12325 1685 12359
rect 1685 12325 1719 12359
rect 1719 12325 1728 12359
rect 1676 12316 1728 12325
rect 3884 12393 3893 12427
rect 3893 12393 3927 12427
rect 3927 12393 3936 12427
rect 3884 12384 3936 12393
rect 4436 12427 4488 12436
rect 4436 12393 4445 12427
rect 4445 12393 4479 12427
rect 4479 12393 4488 12427
rect 4436 12384 4488 12393
rect 6368 12384 6420 12436
rect 5724 12316 5776 12368
rect 9496 12384 9548 12436
rect 9772 12427 9824 12436
rect 9772 12393 9781 12427
rect 9781 12393 9815 12427
rect 9815 12393 9824 12427
rect 9772 12384 9824 12393
rect 1492 12223 1544 12232
rect 1492 12189 1501 12223
rect 1501 12189 1535 12223
rect 1535 12189 1544 12223
rect 1492 12180 1544 12189
rect 1952 12180 2004 12232
rect 2964 12180 3016 12232
rect 4896 12180 4948 12232
rect 6092 12248 6144 12300
rect 6736 12248 6788 12300
rect 7104 12248 7156 12300
rect 8024 12316 8076 12368
rect 8116 12291 8168 12300
rect 8116 12257 8125 12291
rect 8125 12257 8159 12291
rect 8159 12257 8168 12291
rect 8116 12248 8168 12257
rect 8300 12291 8352 12300
rect 8300 12257 8309 12291
rect 8309 12257 8343 12291
rect 8343 12257 8352 12291
rect 8300 12248 8352 12257
rect 9220 12291 9272 12300
rect 9220 12257 9229 12291
rect 9229 12257 9263 12291
rect 9263 12257 9272 12291
rect 9220 12248 9272 12257
rect 10324 12384 10376 12436
rect 12992 12384 13044 12436
rect 13176 12427 13228 12436
rect 13176 12393 13185 12427
rect 13185 12393 13219 12427
rect 13219 12393 13228 12427
rect 13176 12384 13228 12393
rect 1860 12155 1912 12164
rect 1860 12121 1869 12155
rect 1869 12121 1903 12155
rect 1903 12121 1912 12155
rect 1860 12112 1912 12121
rect 2688 12044 2740 12096
rect 4896 12087 4948 12096
rect 4896 12053 4905 12087
rect 4905 12053 4939 12087
rect 4939 12053 4948 12087
rect 4896 12044 4948 12053
rect 5080 12044 5132 12096
rect 5356 12044 5408 12096
rect 6000 12087 6052 12096
rect 6000 12053 6009 12087
rect 6009 12053 6043 12087
rect 6043 12053 6052 12087
rect 6000 12044 6052 12053
rect 6644 12180 6696 12232
rect 7840 12180 7892 12232
rect 8392 12223 8444 12232
rect 8392 12189 8401 12223
rect 8401 12189 8435 12223
rect 8435 12189 8444 12223
rect 8392 12180 8444 12189
rect 7380 12112 7432 12164
rect 7656 12112 7708 12164
rect 6736 12044 6788 12096
rect 8668 12044 8720 12096
rect 9312 12112 9364 12164
rect 10324 12248 10376 12300
rect 10508 12248 10560 12300
rect 12348 12248 12400 12300
rect 12808 12316 12860 12368
rect 16764 12384 16816 12436
rect 15384 12316 15436 12368
rect 18696 12384 18748 12436
rect 18880 12384 18932 12436
rect 22100 12384 22152 12436
rect 9496 12180 9548 12232
rect 9956 12180 10008 12232
rect 10784 12180 10836 12232
rect 9772 12112 9824 12164
rect 11704 12112 11756 12164
rect 12532 12112 12584 12164
rect 10600 12087 10652 12096
rect 10600 12053 10609 12087
rect 10609 12053 10643 12087
rect 10643 12053 10652 12087
rect 10600 12044 10652 12053
rect 10876 12044 10928 12096
rect 11060 12087 11112 12096
rect 11060 12053 11069 12087
rect 11069 12053 11103 12087
rect 11103 12053 11112 12087
rect 11060 12044 11112 12053
rect 12164 12087 12216 12096
rect 12164 12053 12173 12087
rect 12173 12053 12207 12087
rect 12207 12053 12216 12087
rect 12164 12044 12216 12053
rect 12256 12087 12308 12096
rect 12256 12053 12265 12087
rect 12265 12053 12299 12087
rect 12299 12053 12308 12087
rect 17040 12248 17092 12300
rect 17500 12291 17552 12300
rect 17500 12257 17509 12291
rect 17509 12257 17543 12291
rect 17543 12257 17552 12291
rect 17500 12248 17552 12257
rect 19616 12316 19668 12368
rect 18420 12248 18472 12300
rect 21456 12316 21508 12368
rect 17868 12180 17920 12232
rect 20260 12180 20312 12232
rect 14004 12112 14056 12164
rect 18880 12112 18932 12164
rect 20536 12155 20588 12164
rect 12256 12044 12308 12053
rect 14188 12044 14240 12096
rect 17132 12044 17184 12096
rect 17224 12044 17276 12096
rect 17868 12044 17920 12096
rect 18144 12087 18196 12096
rect 18144 12053 18153 12087
rect 18153 12053 18187 12087
rect 18187 12053 18196 12087
rect 18144 12044 18196 12053
rect 18328 12044 18380 12096
rect 19708 12087 19760 12096
rect 19708 12053 19717 12087
rect 19717 12053 19751 12087
rect 19751 12053 19760 12087
rect 19708 12044 19760 12053
rect 20536 12121 20545 12155
rect 20545 12121 20579 12155
rect 20579 12121 20588 12155
rect 20536 12112 20588 12121
rect 21456 12155 21508 12164
rect 21456 12121 21465 12155
rect 21465 12121 21499 12155
rect 21499 12121 21508 12155
rect 21456 12112 21508 12121
rect 6148 11942 6200 11994
rect 6212 11942 6264 11994
rect 6276 11942 6328 11994
rect 6340 11942 6392 11994
rect 6404 11942 6456 11994
rect 11346 11942 11398 11994
rect 11410 11942 11462 11994
rect 11474 11942 11526 11994
rect 11538 11942 11590 11994
rect 11602 11942 11654 11994
rect 16544 11942 16596 11994
rect 16608 11942 16660 11994
rect 16672 11942 16724 11994
rect 16736 11942 16788 11994
rect 16800 11942 16852 11994
rect 21742 11942 21794 11994
rect 21806 11942 21858 11994
rect 21870 11942 21922 11994
rect 21934 11942 21986 11994
rect 21998 11942 22050 11994
rect 1768 11840 1820 11892
rect 4252 11840 4304 11892
rect 5724 11883 5776 11892
rect 5724 11849 5733 11883
rect 5733 11849 5767 11883
rect 5767 11849 5776 11883
rect 5724 11840 5776 11849
rect 1400 11704 1452 11756
rect 4804 11772 4856 11824
rect 6644 11840 6696 11892
rect 7748 11840 7800 11892
rect 10876 11883 10928 11892
rect 1308 11636 1360 11688
rect 1676 11679 1728 11688
rect 1676 11645 1685 11679
rect 1685 11645 1719 11679
rect 1719 11645 1728 11679
rect 1676 11636 1728 11645
rect 2136 11747 2188 11756
rect 2136 11713 2145 11747
rect 2145 11713 2179 11747
rect 2179 11713 2188 11747
rect 2136 11704 2188 11713
rect 5264 11704 5316 11756
rect 2596 11636 2648 11688
rect 5632 11636 5684 11688
rect 6092 11704 6144 11756
rect 6276 11704 6328 11756
rect 6644 11747 6696 11756
rect 6644 11713 6678 11747
rect 6678 11713 6696 11747
rect 6644 11704 6696 11713
rect 10876 11849 10885 11883
rect 10885 11849 10919 11883
rect 10919 11849 10928 11883
rect 10876 11840 10928 11849
rect 14280 11883 14332 11892
rect 10508 11772 10560 11824
rect 10600 11772 10652 11824
rect 12164 11815 12216 11824
rect 12164 11781 12198 11815
rect 12198 11781 12216 11815
rect 12164 11772 12216 11781
rect 9128 11747 9180 11756
rect 8300 11679 8352 11688
rect 8300 11645 8309 11679
rect 8309 11645 8343 11679
rect 8343 11645 8352 11679
rect 8300 11636 8352 11645
rect 8116 11568 8168 11620
rect 4068 11500 4120 11552
rect 5448 11500 5500 11552
rect 5632 11500 5684 11552
rect 7012 11500 7064 11552
rect 8024 11500 8076 11552
rect 8668 11543 8720 11552
rect 8668 11509 8677 11543
rect 8677 11509 8711 11543
rect 8711 11509 8720 11543
rect 8668 11500 8720 11509
rect 9128 11713 9137 11747
rect 9137 11713 9171 11747
rect 9171 11713 9180 11747
rect 9128 11704 9180 11713
rect 9404 11747 9456 11756
rect 9404 11713 9438 11747
rect 9438 11713 9456 11747
rect 9404 11704 9456 11713
rect 9680 11704 9732 11756
rect 10784 11679 10836 11688
rect 10784 11645 10793 11679
rect 10793 11645 10827 11679
rect 10827 11645 10836 11679
rect 10784 11636 10836 11645
rect 13268 11704 13320 11756
rect 14280 11849 14289 11883
rect 14289 11849 14323 11883
rect 14323 11849 14332 11883
rect 14280 11840 14332 11849
rect 17776 11840 17828 11892
rect 18328 11883 18380 11892
rect 18328 11849 18337 11883
rect 18337 11849 18371 11883
rect 18371 11849 18380 11883
rect 18328 11840 18380 11849
rect 20536 11840 20588 11892
rect 21364 11883 21416 11892
rect 21364 11849 21373 11883
rect 21373 11849 21407 11883
rect 21407 11849 21416 11883
rect 21364 11840 21416 11849
rect 16120 11772 16172 11824
rect 17316 11772 17368 11824
rect 15568 11704 15620 11756
rect 17132 11704 17184 11756
rect 18696 11747 18748 11756
rect 18696 11713 18705 11747
rect 18705 11713 18739 11747
rect 18739 11713 18748 11747
rect 18696 11704 18748 11713
rect 19248 11772 19300 11824
rect 20812 11772 20864 11824
rect 21548 11747 21600 11756
rect 21548 11713 21557 11747
rect 21557 11713 21591 11747
rect 21591 11713 21600 11747
rect 21548 11704 21600 11713
rect 11888 11679 11940 11688
rect 10416 11500 10468 11552
rect 11612 11500 11664 11552
rect 11888 11645 11897 11679
rect 11897 11645 11931 11679
rect 11931 11645 11940 11679
rect 11888 11636 11940 11645
rect 15660 11679 15712 11688
rect 15660 11645 15669 11679
rect 15669 11645 15703 11679
rect 15703 11645 15712 11679
rect 15660 11636 15712 11645
rect 17592 11636 17644 11688
rect 17960 11636 18012 11688
rect 18880 11679 18932 11688
rect 18880 11645 18889 11679
rect 18889 11645 18923 11679
rect 18923 11645 18932 11679
rect 18880 11636 18932 11645
rect 19064 11636 19116 11688
rect 19800 11679 19852 11688
rect 19800 11645 19809 11679
rect 19809 11645 19843 11679
rect 19843 11645 19852 11679
rect 19800 11636 19852 11645
rect 19984 11679 20036 11688
rect 19984 11645 19993 11679
rect 19993 11645 20027 11679
rect 20027 11645 20036 11679
rect 19984 11636 20036 11645
rect 21364 11636 21416 11688
rect 14280 11568 14332 11620
rect 18236 11568 18288 11620
rect 18328 11568 18380 11620
rect 19248 11568 19300 11620
rect 21456 11568 21508 11620
rect 12992 11500 13044 11552
rect 13360 11500 13412 11552
rect 16580 11500 16632 11552
rect 17776 11500 17828 11552
rect 20168 11500 20220 11552
rect 21088 11543 21140 11552
rect 21088 11509 21097 11543
rect 21097 11509 21131 11543
rect 21131 11509 21140 11543
rect 21088 11500 21140 11509
rect 3549 11398 3601 11450
rect 3613 11398 3665 11450
rect 3677 11398 3729 11450
rect 3741 11398 3793 11450
rect 3805 11398 3857 11450
rect 8747 11398 8799 11450
rect 8811 11398 8863 11450
rect 8875 11398 8927 11450
rect 8939 11398 8991 11450
rect 9003 11398 9055 11450
rect 13945 11398 13997 11450
rect 14009 11398 14061 11450
rect 14073 11398 14125 11450
rect 14137 11398 14189 11450
rect 14201 11398 14253 11450
rect 19143 11398 19195 11450
rect 19207 11398 19259 11450
rect 19271 11398 19323 11450
rect 19335 11398 19387 11450
rect 19399 11398 19451 11450
rect 1952 11339 2004 11348
rect 1952 11305 1961 11339
rect 1961 11305 1995 11339
rect 1995 11305 2004 11339
rect 1952 11296 2004 11305
rect 6920 11296 6972 11348
rect 7288 11339 7340 11348
rect 7288 11305 7297 11339
rect 7297 11305 7331 11339
rect 7331 11305 7340 11339
rect 7288 11296 7340 11305
rect 9128 11296 9180 11348
rect 5908 11228 5960 11280
rect 2228 11092 2280 11144
rect 3240 11092 3292 11144
rect 4344 11092 4396 11144
rect 5172 11160 5224 11212
rect 8484 11160 8536 11212
rect 11612 11296 11664 11348
rect 4804 11135 4856 11144
rect 4804 11101 4813 11135
rect 4813 11101 4847 11135
rect 4847 11101 4856 11135
rect 4804 11092 4856 11101
rect 6552 11092 6604 11144
rect 12256 11160 12308 11212
rect 13820 11228 13872 11280
rect 9220 11135 9272 11144
rect 9220 11101 9254 11135
rect 9254 11101 9272 11135
rect 9220 11092 9272 11101
rect 1492 11067 1544 11076
rect 1492 11033 1501 11067
rect 1501 11033 1535 11067
rect 1535 11033 1544 11067
rect 1492 11024 1544 11033
rect 3332 11024 3384 11076
rect 5080 11024 5132 11076
rect 6276 11024 6328 11076
rect 8116 11024 8168 11076
rect 8300 11024 8352 11076
rect 10784 11092 10836 11144
rect 11704 11092 11756 11144
rect 14740 11296 14792 11348
rect 16948 11296 17000 11348
rect 17132 11339 17184 11348
rect 17132 11305 17141 11339
rect 17141 11305 17175 11339
rect 17175 11305 17184 11339
rect 17132 11296 17184 11305
rect 17316 11339 17368 11348
rect 17316 11305 17325 11339
rect 17325 11305 17359 11339
rect 17359 11305 17368 11339
rect 17316 11296 17368 11305
rect 18696 11296 18748 11348
rect 20168 11339 20220 11348
rect 20168 11305 20177 11339
rect 20177 11305 20211 11339
rect 20211 11305 20220 11339
rect 20168 11296 20220 11305
rect 20812 11296 20864 11348
rect 21180 11296 21232 11348
rect 15568 11228 15620 11280
rect 17684 11228 17736 11280
rect 18788 11228 18840 11280
rect 16212 11203 16264 11212
rect 16212 11169 16221 11203
rect 16221 11169 16255 11203
rect 16255 11169 16264 11203
rect 16212 11160 16264 11169
rect 16580 11203 16632 11212
rect 16580 11169 16589 11203
rect 16589 11169 16623 11203
rect 16623 11169 16632 11203
rect 16580 11160 16632 11169
rect 17960 11160 18012 11212
rect 18696 11160 18748 11212
rect 19064 11160 19116 11212
rect 19800 11203 19852 11212
rect 19800 11169 19809 11203
rect 19809 11169 19843 11203
rect 19843 11169 19852 11203
rect 19800 11160 19852 11169
rect 21180 11160 21232 11212
rect 9404 11024 9456 11076
rect 2044 10999 2096 11008
rect 2044 10965 2053 10999
rect 2053 10965 2087 10999
rect 2087 10965 2096 10999
rect 2412 10999 2464 11008
rect 2044 10956 2096 10965
rect 2412 10965 2421 10999
rect 2421 10965 2455 10999
rect 2455 10965 2464 10999
rect 2412 10956 2464 10965
rect 2780 10956 2832 11008
rect 4252 10999 4304 11008
rect 4252 10965 4261 10999
rect 4261 10965 4295 10999
rect 4295 10965 4304 10999
rect 4252 10956 4304 10965
rect 13084 11024 13136 11076
rect 14096 11135 14148 11144
rect 14096 11101 14105 11135
rect 14105 11101 14139 11135
rect 14139 11101 14148 11135
rect 14096 11092 14148 11101
rect 18420 11092 18472 11144
rect 18604 11092 18656 11144
rect 14464 11024 14516 11076
rect 16212 11024 16264 11076
rect 17960 11024 18012 11076
rect 18328 11024 18380 11076
rect 19984 11092 20036 11144
rect 19248 11024 19300 11076
rect 20352 11024 20404 11076
rect 20536 11067 20588 11076
rect 20536 11033 20545 11067
rect 20545 11033 20579 11067
rect 20579 11033 20588 11067
rect 20996 11092 21048 11144
rect 21456 11135 21508 11144
rect 21456 11101 21465 11135
rect 21465 11101 21499 11135
rect 21499 11101 21508 11135
rect 21456 11092 21508 11101
rect 21088 11067 21140 11076
rect 20536 11024 20588 11033
rect 21088 11033 21097 11067
rect 21097 11033 21131 11067
rect 21131 11033 21140 11067
rect 21088 11024 21140 11033
rect 16396 10956 16448 11008
rect 19432 10956 19484 11008
rect 19892 10956 19944 11008
rect 6148 10854 6200 10906
rect 6212 10854 6264 10906
rect 6276 10854 6328 10906
rect 6340 10854 6392 10906
rect 6404 10854 6456 10906
rect 11346 10854 11398 10906
rect 11410 10854 11462 10906
rect 11474 10854 11526 10906
rect 11538 10854 11590 10906
rect 11602 10854 11654 10906
rect 16544 10854 16596 10906
rect 16608 10854 16660 10906
rect 16672 10854 16724 10906
rect 16736 10854 16788 10906
rect 16800 10854 16852 10906
rect 21742 10854 21794 10906
rect 21806 10854 21858 10906
rect 21870 10854 21922 10906
rect 21934 10854 21986 10906
rect 21998 10854 22050 10906
rect 2044 10752 2096 10804
rect 2228 10795 2280 10804
rect 2228 10761 2237 10795
rect 2237 10761 2271 10795
rect 2271 10761 2280 10795
rect 2228 10752 2280 10761
rect 2412 10752 2464 10804
rect 2780 10795 2832 10804
rect 2780 10761 2789 10795
rect 2789 10761 2823 10795
rect 2823 10761 2832 10795
rect 2780 10752 2832 10761
rect 3976 10752 4028 10804
rect 4160 10752 4212 10804
rect 4620 10752 4672 10804
rect 4712 10752 4764 10804
rect 10140 10752 10192 10804
rect 10416 10752 10468 10804
rect 12256 10795 12308 10804
rect 12256 10761 12265 10795
rect 12265 10761 12299 10795
rect 12299 10761 12308 10795
rect 12256 10752 12308 10761
rect 14096 10752 14148 10804
rect 15660 10752 15712 10804
rect 16764 10752 16816 10804
rect 17040 10752 17092 10804
rect 18144 10752 18196 10804
rect 19708 10752 19760 10804
rect 19892 10752 19944 10804
rect 20628 10752 20680 10804
rect 20812 10795 20864 10804
rect 20812 10761 20821 10795
rect 20821 10761 20855 10795
rect 20855 10761 20864 10795
rect 20812 10752 20864 10761
rect 1768 10616 1820 10668
rect 2688 10659 2740 10668
rect 2688 10625 2697 10659
rect 2697 10625 2731 10659
rect 2731 10625 2740 10659
rect 2688 10616 2740 10625
rect 5172 10684 5224 10736
rect 7380 10684 7432 10736
rect 12164 10684 12216 10736
rect 15384 10727 15436 10736
rect 15384 10693 15402 10727
rect 15402 10693 15436 10727
rect 15384 10684 15436 10693
rect 2964 10591 3016 10600
rect 2964 10557 2973 10591
rect 2973 10557 3007 10591
rect 3007 10557 3016 10591
rect 2964 10548 3016 10557
rect 3884 10591 3936 10600
rect 3884 10557 3893 10591
rect 3893 10557 3927 10591
rect 3927 10557 3936 10591
rect 3884 10548 3936 10557
rect 4160 10548 4212 10600
rect 4804 10591 4856 10600
rect 4804 10557 4813 10591
rect 4813 10557 4847 10591
rect 4847 10557 4856 10591
rect 4804 10548 4856 10557
rect 5080 10548 5132 10600
rect 6552 10480 6604 10532
rect 3424 10455 3476 10464
rect 3424 10421 3433 10455
rect 3433 10421 3467 10455
rect 3467 10421 3476 10455
rect 3424 10412 3476 10421
rect 4252 10455 4304 10464
rect 4252 10421 4261 10455
rect 4261 10421 4295 10455
rect 4295 10421 4304 10455
rect 4252 10412 4304 10421
rect 5172 10455 5224 10464
rect 5172 10421 5181 10455
rect 5181 10421 5215 10455
rect 5215 10421 5224 10455
rect 5172 10412 5224 10421
rect 6368 10455 6420 10464
rect 6368 10421 6377 10455
rect 6377 10421 6411 10455
rect 6411 10421 6420 10455
rect 6368 10412 6420 10421
rect 10784 10616 10836 10668
rect 17408 10616 17460 10668
rect 18328 10616 18380 10668
rect 19616 10684 19668 10736
rect 14648 10548 14700 10600
rect 15660 10591 15712 10600
rect 15660 10557 15669 10591
rect 15669 10557 15703 10591
rect 15703 10557 15712 10591
rect 15660 10548 15712 10557
rect 16396 10548 16448 10600
rect 17040 10591 17092 10600
rect 17040 10557 17049 10591
rect 17049 10557 17083 10591
rect 17083 10557 17092 10591
rect 17040 10548 17092 10557
rect 17224 10591 17276 10600
rect 17224 10557 17233 10591
rect 17233 10557 17267 10591
rect 17267 10557 17276 10591
rect 17224 10548 17276 10557
rect 18880 10548 18932 10600
rect 19432 10659 19484 10668
rect 19432 10625 19441 10659
rect 19441 10625 19475 10659
rect 19475 10625 19484 10659
rect 19432 10616 19484 10625
rect 19984 10616 20036 10668
rect 20076 10616 20128 10668
rect 21456 10659 21508 10668
rect 21456 10625 21465 10659
rect 21465 10625 21499 10659
rect 21499 10625 21508 10659
rect 21456 10616 21508 10625
rect 14464 10412 14516 10464
rect 18696 10480 18748 10532
rect 16396 10412 16448 10464
rect 18880 10412 18932 10464
rect 20812 10548 20864 10600
rect 20720 10480 20772 10532
rect 20628 10412 20680 10464
rect 3549 10310 3601 10362
rect 3613 10310 3665 10362
rect 3677 10310 3729 10362
rect 3741 10310 3793 10362
rect 3805 10310 3857 10362
rect 8747 10310 8799 10362
rect 8811 10310 8863 10362
rect 8875 10310 8927 10362
rect 8939 10310 8991 10362
rect 9003 10310 9055 10362
rect 13945 10310 13997 10362
rect 14009 10310 14061 10362
rect 14073 10310 14125 10362
rect 14137 10310 14189 10362
rect 14201 10310 14253 10362
rect 19143 10310 19195 10362
rect 19207 10310 19259 10362
rect 19271 10310 19323 10362
rect 19335 10310 19387 10362
rect 19399 10310 19451 10362
rect 2320 10251 2372 10260
rect 2320 10217 2329 10251
rect 2329 10217 2363 10251
rect 2363 10217 2372 10251
rect 2320 10208 2372 10217
rect 2688 10208 2740 10260
rect 3884 10208 3936 10260
rect 5172 10208 5224 10260
rect 10232 10208 10284 10260
rect 17224 10208 17276 10260
rect 17408 10251 17460 10260
rect 17408 10217 17417 10251
rect 17417 10217 17451 10251
rect 17451 10217 17460 10251
rect 17408 10208 17460 10217
rect 18328 10251 18380 10260
rect 18328 10217 18337 10251
rect 18337 10217 18371 10251
rect 18371 10217 18380 10251
rect 18328 10208 18380 10217
rect 2228 10140 2280 10192
rect 4160 10140 4212 10192
rect 5724 10183 5776 10192
rect 5724 10149 5733 10183
rect 5733 10149 5767 10183
rect 5767 10149 5776 10183
rect 5724 10140 5776 10149
rect 13084 10183 13136 10192
rect 13084 10149 13093 10183
rect 13093 10149 13127 10183
rect 13127 10149 13136 10183
rect 13084 10140 13136 10149
rect 19156 10208 19208 10260
rect 2044 10115 2096 10124
rect 2044 10081 2053 10115
rect 2053 10081 2087 10115
rect 2087 10081 2096 10115
rect 2044 10072 2096 10081
rect 3056 10072 3108 10124
rect 3332 10115 3384 10124
rect 3332 10081 3341 10115
rect 3341 10081 3375 10115
rect 3375 10081 3384 10115
rect 3332 10072 3384 10081
rect 4804 10072 4856 10124
rect 1492 10047 1544 10056
rect 1492 10013 1501 10047
rect 1501 10013 1535 10047
rect 1535 10013 1544 10047
rect 1492 10004 1544 10013
rect 2136 10047 2188 10056
rect 2136 10013 2145 10047
rect 2145 10013 2179 10047
rect 2179 10013 2188 10047
rect 2136 10004 2188 10013
rect 1860 9979 1912 9988
rect 1860 9945 1869 9979
rect 1869 9945 1903 9979
rect 1903 9945 1912 9979
rect 1860 9936 1912 9945
rect 1952 9868 2004 9920
rect 3976 10004 4028 10056
rect 4436 10047 4488 10056
rect 4436 10013 4445 10047
rect 4445 10013 4479 10047
rect 4479 10013 4488 10047
rect 4436 10004 4488 10013
rect 5172 10004 5224 10056
rect 4620 9936 4672 9988
rect 15660 10115 15712 10124
rect 6552 10004 6604 10056
rect 8024 9936 8076 9988
rect 15660 10081 15669 10115
rect 15669 10081 15703 10115
rect 15703 10081 15712 10115
rect 15660 10072 15712 10081
rect 16580 10115 16632 10124
rect 16580 10081 16589 10115
rect 16589 10081 16623 10115
rect 16623 10081 16632 10115
rect 16580 10072 16632 10081
rect 16856 10115 16908 10124
rect 16856 10081 16865 10115
rect 16865 10081 16899 10115
rect 16899 10081 16908 10115
rect 16856 10072 16908 10081
rect 17040 10072 17092 10124
rect 19800 10208 19852 10260
rect 19984 10251 20036 10260
rect 19984 10217 19993 10251
rect 19993 10217 20027 10251
rect 20027 10217 20036 10251
rect 19984 10208 20036 10217
rect 21272 10208 21324 10260
rect 21364 10251 21416 10260
rect 21364 10217 21373 10251
rect 21373 10217 21407 10251
rect 21407 10217 21416 10251
rect 21364 10208 21416 10217
rect 19432 10140 19484 10192
rect 20628 10115 20680 10124
rect 12256 10004 12308 10056
rect 18512 10004 18564 10056
rect 18788 10004 18840 10056
rect 11980 9979 12032 9988
rect 11980 9945 11992 9979
rect 11992 9945 12032 9979
rect 11980 9936 12032 9945
rect 12164 9936 12216 9988
rect 15384 9979 15436 9988
rect 4344 9911 4396 9920
rect 4344 9877 4353 9911
rect 4353 9877 4387 9911
rect 4387 9877 4396 9911
rect 4344 9868 4396 9877
rect 4712 9868 4764 9920
rect 6368 9868 6420 9920
rect 6736 9868 6788 9920
rect 9772 9868 9824 9920
rect 9956 9911 10008 9920
rect 9956 9877 9965 9911
rect 9965 9877 9999 9911
rect 9999 9877 10008 9911
rect 15384 9945 15402 9979
rect 15402 9945 15436 9979
rect 15384 9936 15436 9945
rect 20628 10081 20637 10115
rect 20637 10081 20671 10115
rect 20671 10081 20680 10115
rect 20628 10072 20680 10081
rect 19524 10047 19576 10056
rect 19524 10013 19533 10047
rect 19533 10013 19567 10047
rect 19567 10013 19576 10047
rect 19524 10004 19576 10013
rect 19708 10004 19760 10056
rect 21456 10047 21508 10056
rect 9956 9868 10008 9877
rect 16764 9868 16816 9920
rect 17224 9868 17276 9920
rect 17960 9868 18012 9920
rect 20444 9936 20496 9988
rect 20628 9936 20680 9988
rect 21456 10013 21465 10047
rect 21465 10013 21499 10047
rect 21499 10013 21508 10047
rect 21456 10004 21508 10013
rect 19616 9911 19668 9920
rect 19616 9877 19625 9911
rect 19625 9877 19659 9911
rect 19659 9877 19668 9911
rect 20168 9911 20220 9920
rect 19616 9868 19668 9877
rect 20168 9877 20177 9911
rect 20177 9877 20211 9911
rect 20211 9877 20220 9911
rect 20168 9868 20220 9877
rect 20536 9911 20588 9920
rect 20536 9877 20545 9911
rect 20545 9877 20579 9911
rect 20579 9877 20588 9911
rect 20536 9868 20588 9877
rect 6148 9766 6200 9818
rect 6212 9766 6264 9818
rect 6276 9766 6328 9818
rect 6340 9766 6392 9818
rect 6404 9766 6456 9818
rect 11346 9766 11398 9818
rect 11410 9766 11462 9818
rect 11474 9766 11526 9818
rect 11538 9766 11590 9818
rect 11602 9766 11654 9818
rect 16544 9766 16596 9818
rect 16608 9766 16660 9818
rect 16672 9766 16724 9818
rect 16736 9766 16788 9818
rect 16800 9766 16852 9818
rect 21742 9766 21794 9818
rect 21806 9766 21858 9818
rect 21870 9766 21922 9818
rect 21934 9766 21986 9818
rect 21998 9766 22050 9818
rect 1492 9664 1544 9716
rect 3424 9664 3476 9716
rect 2964 9596 3016 9648
rect 4252 9596 4304 9648
rect 3976 9528 4028 9580
rect 1400 9503 1452 9512
rect 1400 9469 1409 9503
rect 1409 9469 1443 9503
rect 1443 9469 1452 9503
rect 1400 9460 1452 9469
rect 3332 9503 3384 9512
rect 3332 9469 3341 9503
rect 3341 9469 3375 9503
rect 3375 9469 3384 9503
rect 3332 9460 3384 9469
rect 3424 9503 3476 9512
rect 3424 9469 3433 9503
rect 3433 9469 3467 9503
rect 3467 9469 3476 9503
rect 3424 9460 3476 9469
rect 4068 9460 4120 9512
rect 4712 9664 4764 9716
rect 5080 9664 5132 9716
rect 8024 9664 8076 9716
rect 13636 9664 13688 9716
rect 10140 9639 10192 9648
rect 5908 9571 5960 9580
rect 5908 9537 5926 9571
rect 5926 9537 5960 9571
rect 5908 9528 5960 9537
rect 6736 9528 6788 9580
rect 7932 9528 7984 9580
rect 6368 9460 6420 9512
rect 10140 9605 10174 9639
rect 10174 9605 10192 9639
rect 10140 9596 10192 9605
rect 12164 9596 12216 9648
rect 7748 9392 7800 9444
rect 2596 9367 2648 9376
rect 2596 9333 2605 9367
rect 2605 9333 2639 9367
rect 2639 9333 2648 9367
rect 2596 9324 2648 9333
rect 2872 9367 2924 9376
rect 2872 9333 2881 9367
rect 2881 9333 2915 9367
rect 2915 9333 2924 9367
rect 2872 9324 2924 9333
rect 3240 9324 3292 9376
rect 6000 9324 6052 9376
rect 7932 9367 7984 9376
rect 7932 9333 7941 9367
rect 7941 9333 7975 9367
rect 7975 9333 7984 9367
rect 7932 9324 7984 9333
rect 8116 9324 8168 9376
rect 9772 9460 9824 9512
rect 9496 9392 9548 9444
rect 14556 9528 14608 9580
rect 17132 9664 17184 9716
rect 17500 9664 17552 9716
rect 19524 9664 19576 9716
rect 20168 9664 20220 9716
rect 20536 9664 20588 9716
rect 15016 9528 15068 9580
rect 9588 9367 9640 9376
rect 9588 9333 9597 9367
rect 9597 9333 9631 9367
rect 9631 9333 9640 9367
rect 9588 9324 9640 9333
rect 10508 9324 10560 9376
rect 11704 9324 11756 9376
rect 13544 9324 13596 9376
rect 13820 9324 13872 9376
rect 15752 9460 15804 9512
rect 18144 9639 18196 9648
rect 18144 9605 18153 9639
rect 18153 9605 18187 9639
rect 18187 9605 18196 9639
rect 18144 9596 18196 9605
rect 16396 9392 16448 9444
rect 18144 9460 18196 9512
rect 15476 9324 15528 9376
rect 18512 9324 18564 9376
rect 21640 9528 21692 9580
rect 21548 9503 21600 9512
rect 19616 9392 19668 9444
rect 21548 9469 21557 9503
rect 21557 9469 21591 9503
rect 21591 9469 21600 9503
rect 21548 9460 21600 9469
rect 20812 9392 20864 9444
rect 3549 9222 3601 9274
rect 3613 9222 3665 9274
rect 3677 9222 3729 9274
rect 3741 9222 3793 9274
rect 3805 9222 3857 9274
rect 8747 9222 8799 9274
rect 8811 9222 8863 9274
rect 8875 9222 8927 9274
rect 8939 9222 8991 9274
rect 9003 9222 9055 9274
rect 13945 9222 13997 9274
rect 14009 9222 14061 9274
rect 14073 9222 14125 9274
rect 14137 9222 14189 9274
rect 14201 9222 14253 9274
rect 19143 9222 19195 9274
rect 19207 9222 19259 9274
rect 19271 9222 19323 9274
rect 19335 9222 19387 9274
rect 19399 9222 19451 9274
rect 2504 9120 2556 9172
rect 7380 9120 7432 9172
rect 2872 9027 2924 9036
rect 2872 8993 2881 9027
rect 2881 8993 2915 9027
rect 2915 8993 2924 9027
rect 2872 8984 2924 8993
rect 2228 8959 2280 8968
rect 2228 8925 2237 8959
rect 2237 8925 2271 8959
rect 2271 8925 2280 8959
rect 2228 8916 2280 8925
rect 2780 8823 2832 8832
rect 2780 8789 2789 8823
rect 2789 8789 2823 8823
rect 2823 8789 2832 8823
rect 6368 8959 6420 8968
rect 6368 8925 6377 8959
rect 6377 8925 6411 8959
rect 6411 8925 6420 8959
rect 6368 8916 6420 8925
rect 12164 9120 12216 9172
rect 7840 9095 7892 9104
rect 7840 9061 7849 9095
rect 7849 9061 7883 9095
rect 7883 9061 7892 9095
rect 7840 9052 7892 9061
rect 7932 9052 7984 9104
rect 8760 9095 8812 9104
rect 8760 9061 8769 9095
rect 8769 9061 8803 9095
rect 8803 9061 8812 9095
rect 8760 9052 8812 9061
rect 9496 9052 9548 9104
rect 11980 9052 12032 9104
rect 13912 9120 13964 9172
rect 15016 9120 15068 9172
rect 18144 9120 18196 9172
rect 17684 9052 17736 9104
rect 17960 9095 18012 9104
rect 17960 9061 17969 9095
rect 17969 9061 18003 9095
rect 18003 9061 18012 9095
rect 17960 9052 18012 9061
rect 8024 8984 8076 9036
rect 19156 9120 19208 9172
rect 19340 9120 19392 9172
rect 19984 9120 20036 9172
rect 20628 9163 20680 9172
rect 20628 9129 20637 9163
rect 20637 9129 20671 9163
rect 20671 9129 20680 9163
rect 20628 9120 20680 9129
rect 20168 9052 20220 9104
rect 20720 9052 20772 9104
rect 8208 8959 8260 8968
rect 8208 8925 8217 8959
rect 8217 8925 8251 8959
rect 8251 8925 8260 8959
rect 8208 8916 8260 8925
rect 10508 8959 10560 8968
rect 5172 8891 5224 8900
rect 5172 8857 5206 8891
rect 5206 8857 5224 8891
rect 5172 8848 5224 8857
rect 5724 8848 5776 8900
rect 8852 8848 8904 8900
rect 9588 8848 9640 8900
rect 10140 8848 10192 8900
rect 10508 8925 10517 8959
rect 10517 8925 10551 8959
rect 10551 8925 10560 8959
rect 10508 8916 10560 8925
rect 10692 8916 10744 8968
rect 13360 8916 13412 8968
rect 2780 8780 2832 8789
rect 7748 8823 7800 8832
rect 7748 8789 7757 8823
rect 7757 8789 7791 8823
rect 7791 8789 7800 8823
rect 7748 8780 7800 8789
rect 8116 8780 8168 8832
rect 9128 8823 9180 8832
rect 9128 8789 9137 8823
rect 9137 8789 9171 8823
rect 9171 8789 9180 8823
rect 9128 8780 9180 8789
rect 15660 8916 15712 8968
rect 19248 8984 19300 9036
rect 19892 9027 19944 9036
rect 17408 8916 17460 8968
rect 19340 8916 19392 8968
rect 14464 8848 14516 8900
rect 12532 8780 12584 8832
rect 13820 8823 13872 8832
rect 13820 8789 13829 8823
rect 13829 8789 13863 8823
rect 13863 8789 13872 8823
rect 13820 8780 13872 8789
rect 13912 8780 13964 8832
rect 16948 8848 17000 8900
rect 17500 8891 17552 8900
rect 17500 8857 17509 8891
rect 17509 8857 17543 8891
rect 17543 8857 17552 8891
rect 17500 8848 17552 8857
rect 18144 8848 18196 8900
rect 19432 8848 19484 8900
rect 19892 8993 19901 9027
rect 19901 8993 19935 9027
rect 19935 8993 19944 9027
rect 19892 8984 19944 8993
rect 20996 9027 21048 9036
rect 20996 8993 21005 9027
rect 21005 8993 21039 9027
rect 21039 8993 21048 9027
rect 20996 8984 21048 8993
rect 19984 8916 20036 8968
rect 20628 8916 20680 8968
rect 20536 8848 20588 8900
rect 17040 8823 17092 8832
rect 17040 8789 17049 8823
rect 17049 8789 17083 8823
rect 17083 8789 17092 8823
rect 17040 8780 17092 8789
rect 17592 8780 17644 8832
rect 18328 8780 18380 8832
rect 18604 8823 18656 8832
rect 18604 8789 18613 8823
rect 18613 8789 18647 8823
rect 18647 8789 18656 8823
rect 18604 8780 18656 8789
rect 18696 8823 18748 8832
rect 18696 8789 18705 8823
rect 18705 8789 18739 8823
rect 18739 8789 18748 8823
rect 18696 8780 18748 8789
rect 18972 8780 19024 8832
rect 19524 8780 19576 8832
rect 20076 8780 20128 8832
rect 6148 8678 6200 8730
rect 6212 8678 6264 8730
rect 6276 8678 6328 8730
rect 6340 8678 6392 8730
rect 6404 8678 6456 8730
rect 11346 8678 11398 8730
rect 11410 8678 11462 8730
rect 11474 8678 11526 8730
rect 11538 8678 11590 8730
rect 11602 8678 11654 8730
rect 16544 8678 16596 8730
rect 16608 8678 16660 8730
rect 16672 8678 16724 8730
rect 16736 8678 16788 8730
rect 16800 8678 16852 8730
rect 21742 8678 21794 8730
rect 21806 8678 21858 8730
rect 21870 8678 21922 8730
rect 21934 8678 21986 8730
rect 21998 8678 22050 8730
rect 1584 8619 1636 8628
rect 1584 8585 1593 8619
rect 1593 8585 1627 8619
rect 1627 8585 1636 8619
rect 1584 8576 1636 8585
rect 2780 8576 2832 8628
rect 2872 8619 2924 8628
rect 2872 8585 2881 8619
rect 2881 8585 2915 8619
rect 2915 8585 2924 8619
rect 2872 8576 2924 8585
rect 3148 8576 3200 8628
rect 3332 8576 3384 8628
rect 7840 8576 7892 8628
rect 11060 8576 11112 8628
rect 11428 8576 11480 8628
rect 15660 8576 15712 8628
rect 1308 8440 1360 8492
rect 2044 8483 2096 8492
rect 2044 8449 2053 8483
rect 2053 8449 2087 8483
rect 2087 8449 2096 8483
rect 2044 8440 2096 8449
rect 5632 8508 5684 8560
rect 6552 8508 6604 8560
rect 4160 8483 4212 8492
rect 1952 8415 2004 8424
rect 1952 8381 1961 8415
rect 1961 8381 1995 8415
rect 1995 8381 2004 8415
rect 1952 8372 2004 8381
rect 4160 8449 4169 8483
rect 4169 8449 4203 8483
rect 4203 8449 4212 8483
rect 4160 8440 4212 8449
rect 7380 8440 7432 8492
rect 11152 8508 11204 8560
rect 12532 8508 12584 8560
rect 13820 8508 13872 8560
rect 8760 8483 8812 8492
rect 8760 8449 8769 8483
rect 8769 8449 8803 8483
rect 8803 8449 8812 8483
rect 8760 8440 8812 8449
rect 8852 8440 8904 8492
rect 10968 8483 11020 8492
rect 10968 8449 10977 8483
rect 10977 8449 11011 8483
rect 11011 8449 11020 8483
rect 10968 8440 11020 8449
rect 14280 8440 14332 8492
rect 16580 8576 16632 8628
rect 17408 8619 17460 8628
rect 17408 8585 17417 8619
rect 17417 8585 17451 8619
rect 17451 8585 17460 8619
rect 17408 8576 17460 8585
rect 17960 8619 18012 8628
rect 17960 8585 17969 8619
rect 17969 8585 18003 8619
rect 18003 8585 18012 8619
rect 17960 8576 18012 8585
rect 20812 8619 20864 8628
rect 16396 8508 16448 8560
rect 17316 8508 17368 8560
rect 20812 8585 20821 8619
rect 20821 8585 20855 8619
rect 20855 8585 20864 8619
rect 20812 8576 20864 8585
rect 18972 8508 19024 8560
rect 2780 8415 2832 8424
rect 2780 8381 2789 8415
rect 2789 8381 2823 8415
rect 2823 8381 2832 8415
rect 3332 8415 3384 8424
rect 2780 8372 2832 8381
rect 3332 8381 3341 8415
rect 3341 8381 3375 8415
rect 3375 8381 3384 8415
rect 3332 8372 3384 8381
rect 4068 8372 4120 8424
rect 3424 8304 3476 8356
rect 7656 8372 7708 8424
rect 5172 8304 5224 8356
rect 10140 8347 10192 8356
rect 2136 8236 2188 8288
rect 4068 8236 4120 8288
rect 8484 8236 8536 8288
rect 10140 8313 10149 8347
rect 10149 8313 10183 8347
rect 10183 8313 10192 8347
rect 10140 8304 10192 8313
rect 10508 8347 10560 8356
rect 10508 8313 10517 8347
rect 10517 8313 10551 8347
rect 10551 8313 10560 8347
rect 17040 8483 17092 8492
rect 17040 8449 17049 8483
rect 17049 8449 17083 8483
rect 17083 8449 17092 8483
rect 17040 8440 17092 8449
rect 19248 8440 19300 8492
rect 19524 8440 19576 8492
rect 20352 8483 20404 8492
rect 20352 8449 20361 8483
rect 20361 8449 20395 8483
rect 20395 8449 20404 8483
rect 20352 8440 20404 8449
rect 16948 8415 17000 8424
rect 16948 8381 16957 8415
rect 16957 8381 16991 8415
rect 16991 8381 17000 8415
rect 16948 8372 17000 8381
rect 19616 8415 19668 8424
rect 10508 8304 10560 8313
rect 13912 8304 13964 8356
rect 15200 8304 15252 8356
rect 16580 8304 16632 8356
rect 10876 8236 10928 8288
rect 11980 8279 12032 8288
rect 11980 8245 11989 8279
rect 11989 8245 12023 8279
rect 12023 8245 12032 8279
rect 11980 8236 12032 8245
rect 17500 8279 17552 8288
rect 17500 8245 17509 8279
rect 17509 8245 17543 8279
rect 17543 8245 17552 8279
rect 17500 8236 17552 8245
rect 17684 8236 17736 8288
rect 19616 8381 19625 8415
rect 19625 8381 19659 8415
rect 19659 8381 19668 8415
rect 19616 8372 19668 8381
rect 20444 8415 20496 8424
rect 18512 8304 18564 8356
rect 19432 8304 19484 8356
rect 20444 8381 20453 8415
rect 20453 8381 20487 8415
rect 20487 8381 20496 8415
rect 20444 8372 20496 8381
rect 20536 8415 20588 8424
rect 20536 8381 20545 8415
rect 20545 8381 20579 8415
rect 20579 8381 20588 8415
rect 21272 8415 21324 8424
rect 20536 8372 20588 8381
rect 21272 8381 21281 8415
rect 21281 8381 21315 8415
rect 21315 8381 21324 8415
rect 21272 8372 21324 8381
rect 18696 8236 18748 8288
rect 3549 8134 3601 8186
rect 3613 8134 3665 8186
rect 3677 8134 3729 8186
rect 3741 8134 3793 8186
rect 3805 8134 3857 8186
rect 8747 8134 8799 8186
rect 8811 8134 8863 8186
rect 8875 8134 8927 8186
rect 8939 8134 8991 8186
rect 9003 8134 9055 8186
rect 13945 8134 13997 8186
rect 14009 8134 14061 8186
rect 14073 8134 14125 8186
rect 14137 8134 14189 8186
rect 14201 8134 14253 8186
rect 19143 8134 19195 8186
rect 19207 8134 19259 8186
rect 19271 8134 19323 8186
rect 19335 8134 19387 8186
rect 19399 8134 19451 8186
rect 1400 8075 1452 8084
rect 1400 8041 1409 8075
rect 1409 8041 1443 8075
rect 1443 8041 1452 8075
rect 1400 8032 1452 8041
rect 1952 8032 2004 8084
rect 2780 8032 2832 8084
rect 3976 7964 4028 8016
rect 4528 7964 4580 8016
rect 5632 8007 5684 8016
rect 5632 7973 5641 8007
rect 5641 7973 5675 8007
rect 5675 7973 5684 8007
rect 5632 7964 5684 7973
rect 7380 8007 7432 8016
rect 7380 7973 7389 8007
rect 7389 7973 7423 8007
rect 7423 7973 7432 8007
rect 7380 7964 7432 7973
rect 9680 8007 9732 8016
rect 9680 7973 9689 8007
rect 9689 7973 9723 8007
rect 9723 7973 9732 8007
rect 9680 7964 9732 7973
rect 2136 7896 2188 7948
rect 2504 7896 2556 7948
rect 2688 7828 2740 7880
rect 3056 7760 3108 7812
rect 3424 7803 3476 7812
rect 3424 7769 3433 7803
rect 3433 7769 3467 7803
rect 3467 7769 3476 7803
rect 3424 7760 3476 7769
rect 5172 7896 5224 7948
rect 9404 7896 9456 7948
rect 6460 7828 6512 7880
rect 8668 7828 8720 7880
rect 9680 7828 9732 7880
rect 6828 7760 6880 7812
rect 8392 7760 8444 7812
rect 10508 8032 10560 8084
rect 14280 7964 14332 8016
rect 11428 7896 11480 7948
rect 16488 7939 16540 7948
rect 16488 7905 16497 7939
rect 16497 7905 16531 7939
rect 16531 7905 16540 7939
rect 16488 7896 16540 7905
rect 16948 8032 17000 8084
rect 19616 8075 19668 8084
rect 19616 8041 19625 8075
rect 19625 8041 19659 8075
rect 19659 8041 19668 8075
rect 19616 8032 19668 8041
rect 20628 8032 20680 8084
rect 21272 8032 21324 8084
rect 21548 8075 21600 8084
rect 21548 8041 21557 8075
rect 21557 8041 21591 8075
rect 21591 8041 21600 8075
rect 21548 8032 21600 8041
rect 10600 7871 10652 7880
rect 10600 7837 10609 7871
rect 10609 7837 10643 7871
rect 10643 7837 10652 7871
rect 10600 7828 10652 7837
rect 11060 7828 11112 7880
rect 11796 7828 11848 7880
rect 11980 7828 12032 7880
rect 13820 7871 13872 7880
rect 13820 7837 13829 7871
rect 13829 7837 13863 7871
rect 13863 7837 13872 7871
rect 13820 7828 13872 7837
rect 16672 7871 16724 7880
rect 16672 7837 16681 7871
rect 16681 7837 16715 7871
rect 16715 7837 16724 7871
rect 16672 7828 16724 7837
rect 3516 7692 3568 7744
rect 4344 7692 4396 7744
rect 4712 7735 4764 7744
rect 4712 7701 4721 7735
rect 4721 7701 4755 7735
rect 4755 7701 4764 7735
rect 4712 7692 4764 7701
rect 5080 7692 5132 7744
rect 5264 7692 5316 7744
rect 6552 7692 6604 7744
rect 9404 7692 9456 7744
rect 12992 7760 13044 7812
rect 13728 7760 13780 7812
rect 15200 7803 15252 7812
rect 15200 7769 15218 7803
rect 15218 7769 15252 7803
rect 15200 7760 15252 7769
rect 16396 7760 16448 7812
rect 18696 7896 18748 7948
rect 20168 7939 20220 7948
rect 20168 7905 20177 7939
rect 20177 7905 20211 7939
rect 20211 7905 20220 7939
rect 20168 7896 20220 7905
rect 17776 7828 17828 7880
rect 18052 7828 18104 7880
rect 20996 7871 21048 7880
rect 20996 7837 21005 7871
rect 21005 7837 21039 7871
rect 21039 7837 21048 7871
rect 20996 7828 21048 7837
rect 17868 7760 17920 7812
rect 18788 7760 18840 7812
rect 21088 7760 21140 7812
rect 17776 7692 17828 7744
rect 17960 7735 18012 7744
rect 17960 7701 17969 7735
rect 17969 7701 18003 7735
rect 18003 7701 18012 7735
rect 17960 7692 18012 7701
rect 18420 7735 18472 7744
rect 18420 7701 18429 7735
rect 18429 7701 18463 7735
rect 18463 7701 18472 7735
rect 18420 7692 18472 7701
rect 18604 7692 18656 7744
rect 19984 7735 20036 7744
rect 19984 7701 19993 7735
rect 19993 7701 20027 7735
rect 20027 7701 20036 7735
rect 19984 7692 20036 7701
rect 20260 7692 20312 7744
rect 6148 7590 6200 7642
rect 6212 7590 6264 7642
rect 6276 7590 6328 7642
rect 6340 7590 6392 7642
rect 6404 7590 6456 7642
rect 11346 7590 11398 7642
rect 11410 7590 11462 7642
rect 11474 7590 11526 7642
rect 11538 7590 11590 7642
rect 11602 7590 11654 7642
rect 16544 7590 16596 7642
rect 16608 7590 16660 7642
rect 16672 7590 16724 7642
rect 16736 7590 16788 7642
rect 16800 7590 16852 7642
rect 21742 7590 21794 7642
rect 21806 7590 21858 7642
rect 21870 7590 21922 7642
rect 21934 7590 21986 7642
rect 21998 7590 22050 7642
rect 2872 7488 2924 7540
rect 2412 7420 2464 7472
rect 4160 7488 4212 7540
rect 4528 7488 4580 7540
rect 5080 7531 5132 7540
rect 5080 7497 5089 7531
rect 5089 7497 5123 7531
rect 5123 7497 5132 7531
rect 5080 7488 5132 7497
rect 5448 7531 5500 7540
rect 5448 7497 5457 7531
rect 5457 7497 5491 7531
rect 5491 7497 5500 7531
rect 5448 7488 5500 7497
rect 5540 7488 5592 7540
rect 6736 7488 6788 7540
rect 8208 7488 8260 7540
rect 9404 7531 9456 7540
rect 9404 7497 9413 7531
rect 9413 7497 9447 7531
rect 9447 7497 9456 7531
rect 9404 7488 9456 7497
rect 11060 7488 11112 7540
rect 11980 7488 12032 7540
rect 17040 7488 17092 7540
rect 17500 7488 17552 7540
rect 17776 7488 17828 7540
rect 20904 7488 20956 7540
rect 3884 7420 3936 7472
rect 4068 7420 4120 7472
rect 5264 7420 5316 7472
rect 5356 7420 5408 7472
rect 1952 7327 2004 7336
rect 1952 7293 1961 7327
rect 1961 7293 1995 7327
rect 1995 7293 2004 7327
rect 1952 7284 2004 7293
rect 2228 7327 2280 7336
rect 2228 7293 2237 7327
rect 2237 7293 2271 7327
rect 2271 7293 2280 7327
rect 2228 7284 2280 7293
rect 2504 7327 2556 7336
rect 2504 7293 2513 7327
rect 2513 7293 2547 7327
rect 2547 7293 2556 7327
rect 2504 7284 2556 7293
rect 2596 7284 2648 7336
rect 4804 7327 4856 7336
rect 4804 7293 4813 7327
rect 4813 7293 4847 7327
rect 4847 7293 4856 7327
rect 4804 7284 4856 7293
rect 6552 7420 6604 7472
rect 8392 7420 8444 7472
rect 9128 7420 9180 7472
rect 9864 7395 9916 7404
rect 9864 7361 9873 7395
rect 9873 7361 9907 7395
rect 9907 7361 9916 7395
rect 9864 7352 9916 7361
rect 7380 7284 7432 7336
rect 8484 7284 8536 7336
rect 10600 7420 10652 7472
rect 17960 7420 18012 7472
rect 18052 7420 18104 7472
rect 20352 7420 20404 7472
rect 10876 7327 10928 7336
rect 10876 7293 10885 7327
rect 10885 7293 10919 7327
rect 10919 7293 10928 7327
rect 10876 7284 10928 7293
rect 16396 7284 16448 7336
rect 18696 7327 18748 7336
rect 18696 7293 18705 7327
rect 18705 7293 18739 7327
rect 18739 7293 18748 7327
rect 18696 7284 18748 7293
rect 8852 7216 8904 7268
rect 9036 7216 9088 7268
rect 4160 7148 4212 7200
rect 8208 7191 8260 7200
rect 8208 7157 8217 7191
rect 8217 7157 8251 7191
rect 8251 7157 8260 7191
rect 8208 7148 8260 7157
rect 9772 7148 9824 7200
rect 17776 7191 17828 7200
rect 17776 7157 17785 7191
rect 17785 7157 17819 7191
rect 17819 7157 17828 7191
rect 20536 7352 20588 7404
rect 20720 7327 20772 7336
rect 20720 7293 20729 7327
rect 20729 7293 20763 7327
rect 20763 7293 20772 7327
rect 20720 7284 20772 7293
rect 17776 7148 17828 7157
rect 3549 7046 3601 7098
rect 3613 7046 3665 7098
rect 3677 7046 3729 7098
rect 3741 7046 3793 7098
rect 3805 7046 3857 7098
rect 8747 7046 8799 7098
rect 8811 7046 8863 7098
rect 8875 7046 8927 7098
rect 8939 7046 8991 7098
rect 9003 7046 9055 7098
rect 13945 7046 13997 7098
rect 14009 7046 14061 7098
rect 14073 7046 14125 7098
rect 14137 7046 14189 7098
rect 14201 7046 14253 7098
rect 19143 7046 19195 7098
rect 19207 7046 19259 7098
rect 19271 7046 19323 7098
rect 19335 7046 19387 7098
rect 19399 7046 19451 7098
rect 5448 6944 5500 6996
rect 9680 6987 9732 6996
rect 9680 6953 9689 6987
rect 9689 6953 9723 6987
rect 9723 6953 9732 6987
rect 9680 6944 9732 6953
rect 9772 6944 9824 6996
rect 17776 6944 17828 6996
rect 1584 6808 1636 6860
rect 2780 6876 2832 6928
rect 3608 6876 3660 6928
rect 5908 6876 5960 6928
rect 2136 6808 2188 6860
rect 2964 6808 3016 6860
rect 3976 6851 4028 6860
rect 1400 6740 1452 6792
rect 1676 6740 1728 6792
rect 3332 6740 3384 6792
rect 3976 6817 3985 6851
rect 3985 6817 4019 6851
rect 4019 6817 4028 6851
rect 3976 6808 4028 6817
rect 4068 6808 4120 6860
rect 4436 6851 4488 6860
rect 4436 6817 4445 6851
rect 4445 6817 4479 6851
rect 4479 6817 4488 6851
rect 4436 6808 4488 6817
rect 5540 6808 5592 6860
rect 3884 6740 3936 6792
rect 4804 6740 4856 6792
rect 4988 6740 5040 6792
rect 5264 6740 5316 6792
rect 5724 6808 5776 6860
rect 8392 6808 8444 6860
rect 8484 6808 8536 6860
rect 9864 6808 9916 6860
rect 12532 6851 12584 6860
rect 12532 6817 12541 6851
rect 12541 6817 12575 6851
rect 12575 6817 12584 6851
rect 12532 6808 12584 6817
rect 15384 6808 15436 6860
rect 18236 6808 18288 6860
rect 20628 6808 20680 6860
rect 3976 6672 4028 6724
rect 4068 6672 4120 6724
rect 16948 6740 17000 6792
rect 20812 6783 20864 6792
rect 20812 6749 20821 6783
rect 20821 6749 20855 6783
rect 20855 6749 20864 6783
rect 20812 6740 20864 6749
rect 22376 6808 22428 6860
rect 21456 6783 21508 6792
rect 21456 6749 21465 6783
rect 21465 6749 21499 6783
rect 21499 6749 21508 6783
rect 21456 6740 21508 6749
rect 14648 6672 14700 6724
rect 18512 6672 18564 6724
rect 1584 6647 1636 6656
rect 1584 6613 1593 6647
rect 1593 6613 1627 6647
rect 1627 6613 1636 6647
rect 1584 6604 1636 6613
rect 2044 6647 2096 6656
rect 2044 6613 2053 6647
rect 2053 6613 2087 6647
rect 2087 6613 2096 6647
rect 2044 6604 2096 6613
rect 2136 6604 2188 6656
rect 2596 6604 2648 6656
rect 2872 6647 2924 6656
rect 2872 6613 2881 6647
rect 2881 6613 2915 6647
rect 2915 6613 2924 6647
rect 2872 6604 2924 6613
rect 3240 6647 3292 6656
rect 3240 6613 3249 6647
rect 3249 6613 3283 6647
rect 3283 6613 3292 6647
rect 3240 6604 3292 6613
rect 3516 6604 3568 6656
rect 4620 6647 4672 6656
rect 4620 6613 4629 6647
rect 4629 6613 4663 6647
rect 4663 6613 4672 6647
rect 4620 6604 4672 6613
rect 4896 6604 4948 6656
rect 5264 6604 5316 6656
rect 5908 6647 5960 6656
rect 5908 6613 5917 6647
rect 5917 6613 5951 6647
rect 5951 6613 5960 6647
rect 5908 6604 5960 6613
rect 9220 6647 9272 6656
rect 9220 6613 9229 6647
rect 9229 6613 9263 6647
rect 9263 6613 9272 6647
rect 9220 6604 9272 6613
rect 9312 6647 9364 6656
rect 9312 6613 9321 6647
rect 9321 6613 9355 6647
rect 9355 6613 9364 6647
rect 12716 6647 12768 6656
rect 9312 6604 9364 6613
rect 12716 6613 12725 6647
rect 12725 6613 12759 6647
rect 12759 6613 12768 6647
rect 12716 6604 12768 6613
rect 19800 6604 19852 6656
rect 20628 6647 20680 6656
rect 20628 6613 20637 6647
rect 20637 6613 20671 6647
rect 20671 6613 20680 6647
rect 20628 6604 20680 6613
rect 6148 6502 6200 6554
rect 6212 6502 6264 6554
rect 6276 6502 6328 6554
rect 6340 6502 6392 6554
rect 6404 6502 6456 6554
rect 11346 6502 11398 6554
rect 11410 6502 11462 6554
rect 11474 6502 11526 6554
rect 11538 6502 11590 6554
rect 11602 6502 11654 6554
rect 16544 6502 16596 6554
rect 16608 6502 16660 6554
rect 16672 6502 16724 6554
rect 16736 6502 16788 6554
rect 16800 6502 16852 6554
rect 21742 6502 21794 6554
rect 21806 6502 21858 6554
rect 21870 6502 21922 6554
rect 21934 6502 21986 6554
rect 21998 6502 22050 6554
rect 2228 6400 2280 6452
rect 3332 6400 3384 6452
rect 3516 6443 3568 6452
rect 3516 6409 3525 6443
rect 3525 6409 3559 6443
rect 3559 6409 3568 6443
rect 3516 6400 3568 6409
rect 4712 6400 4764 6452
rect 5908 6400 5960 6452
rect 11980 6400 12032 6452
rect 12716 6443 12768 6452
rect 12716 6409 12725 6443
rect 12725 6409 12759 6443
rect 12759 6409 12768 6443
rect 12716 6400 12768 6409
rect 14648 6443 14700 6452
rect 2964 6332 3016 6384
rect 3608 6332 3660 6384
rect 4528 6332 4580 6384
rect 9220 6332 9272 6384
rect 14648 6409 14657 6443
rect 14657 6409 14691 6443
rect 14691 6409 14700 6443
rect 14648 6400 14700 6409
rect 20628 6400 20680 6452
rect 15384 6375 15436 6384
rect 2596 6264 2648 6316
rect 2780 6264 2832 6316
rect 3332 6264 3384 6316
rect 2228 6239 2280 6248
rect 2228 6205 2237 6239
rect 2237 6205 2271 6239
rect 2271 6205 2280 6239
rect 2228 6196 2280 6205
rect 2320 6239 2372 6248
rect 2320 6205 2329 6239
rect 2329 6205 2363 6239
rect 2363 6205 2372 6239
rect 2320 6196 2372 6205
rect 3148 6196 3200 6248
rect 4068 6239 4120 6248
rect 4068 6205 4077 6239
rect 4077 6205 4111 6239
rect 4111 6205 4120 6239
rect 4068 6196 4120 6205
rect 4804 6264 4856 6316
rect 5356 6239 5408 6248
rect 5356 6205 5365 6239
rect 5365 6205 5399 6239
rect 5399 6205 5408 6239
rect 5356 6196 5408 6205
rect 5448 6239 5500 6248
rect 5448 6205 5457 6239
rect 5457 6205 5491 6239
rect 5491 6205 5500 6239
rect 10508 6264 10560 6316
rect 13084 6307 13136 6316
rect 5448 6196 5500 6205
rect 5908 6196 5960 6248
rect 13084 6273 13093 6307
rect 13093 6273 13127 6307
rect 13127 6273 13136 6307
rect 13084 6264 13136 6273
rect 13728 6264 13780 6316
rect 14556 6307 14608 6316
rect 14556 6273 14565 6307
rect 14565 6273 14599 6307
rect 14599 6273 14608 6307
rect 14556 6264 14608 6273
rect 13176 6239 13228 6248
rect 8208 6128 8260 6180
rect 13176 6205 13185 6239
rect 13185 6205 13219 6239
rect 13219 6205 13228 6239
rect 13176 6196 13228 6205
rect 13360 6239 13412 6248
rect 13360 6205 13369 6239
rect 13369 6205 13403 6239
rect 13403 6205 13412 6239
rect 13360 6196 13412 6205
rect 14096 6239 14148 6248
rect 14096 6205 14105 6239
rect 14105 6205 14139 6239
rect 14139 6205 14148 6239
rect 14096 6196 14148 6205
rect 14648 6196 14700 6248
rect 15384 6341 15393 6375
rect 15393 6341 15427 6375
rect 15427 6341 15436 6375
rect 15384 6332 15436 6341
rect 20536 6332 20588 6384
rect 16948 6264 17000 6316
rect 20720 6239 20772 6248
rect 20720 6205 20729 6239
rect 20729 6205 20763 6239
rect 20763 6205 20772 6239
rect 20720 6196 20772 6205
rect 3148 6060 3200 6112
rect 3549 5958 3601 6010
rect 3613 5958 3665 6010
rect 3677 5958 3729 6010
rect 3741 5958 3793 6010
rect 3805 5958 3857 6010
rect 8747 5958 8799 6010
rect 8811 5958 8863 6010
rect 8875 5958 8927 6010
rect 8939 5958 8991 6010
rect 9003 5958 9055 6010
rect 13945 5958 13997 6010
rect 14009 5958 14061 6010
rect 14073 5958 14125 6010
rect 14137 5958 14189 6010
rect 14201 5958 14253 6010
rect 19143 5958 19195 6010
rect 19207 5958 19259 6010
rect 19271 5958 19323 6010
rect 19335 5958 19387 6010
rect 19399 5958 19451 6010
rect 1768 5899 1820 5908
rect 1768 5865 1777 5899
rect 1777 5865 1811 5899
rect 1811 5865 1820 5899
rect 1768 5856 1820 5865
rect 3240 5856 3292 5908
rect 5356 5899 5408 5908
rect 5356 5865 5365 5899
rect 5365 5865 5399 5899
rect 5399 5865 5408 5899
rect 5356 5856 5408 5865
rect 13176 5856 13228 5908
rect 2412 5763 2464 5772
rect 2412 5729 2421 5763
rect 2421 5729 2455 5763
rect 2455 5729 2464 5763
rect 2412 5720 2464 5729
rect 1400 5695 1452 5704
rect 1400 5661 1409 5695
rect 1409 5661 1443 5695
rect 1443 5661 1452 5695
rect 1400 5652 1452 5661
rect 2872 5788 2924 5840
rect 2688 5584 2740 5636
rect 4436 5720 4488 5772
rect 14556 5763 14608 5772
rect 14556 5729 14565 5763
rect 14565 5729 14599 5763
rect 14599 5729 14608 5763
rect 14556 5720 14608 5729
rect 21272 5695 21324 5704
rect 21272 5661 21281 5695
rect 21281 5661 21315 5695
rect 21315 5661 21324 5695
rect 21272 5652 21324 5661
rect 21548 5695 21600 5704
rect 21548 5661 21557 5695
rect 21557 5661 21591 5695
rect 21591 5661 21600 5695
rect 21548 5652 21600 5661
rect 3332 5584 3384 5636
rect 3516 5584 3568 5636
rect 5264 5584 5316 5636
rect 10968 5584 11020 5636
rect 1584 5559 1636 5568
rect 1584 5525 1593 5559
rect 1593 5525 1627 5559
rect 1627 5525 1636 5559
rect 1584 5516 1636 5525
rect 2136 5559 2188 5568
rect 2136 5525 2145 5559
rect 2145 5525 2179 5559
rect 2179 5525 2188 5559
rect 2136 5516 2188 5525
rect 2872 5559 2924 5568
rect 2872 5525 2881 5559
rect 2881 5525 2915 5559
rect 2915 5525 2924 5559
rect 2872 5516 2924 5525
rect 3976 5516 4028 5568
rect 6148 5414 6200 5466
rect 6212 5414 6264 5466
rect 6276 5414 6328 5466
rect 6340 5414 6392 5466
rect 6404 5414 6456 5466
rect 11346 5414 11398 5466
rect 11410 5414 11462 5466
rect 11474 5414 11526 5466
rect 11538 5414 11590 5466
rect 11602 5414 11654 5466
rect 16544 5414 16596 5466
rect 16608 5414 16660 5466
rect 16672 5414 16724 5466
rect 16736 5414 16788 5466
rect 16800 5414 16852 5466
rect 21742 5414 21794 5466
rect 21806 5414 21858 5466
rect 21870 5414 21922 5466
rect 21934 5414 21986 5466
rect 21998 5414 22050 5466
rect 1676 5312 1728 5364
rect 2136 5312 2188 5364
rect 2780 5355 2832 5364
rect 2780 5321 2789 5355
rect 2789 5321 2823 5355
rect 2823 5321 2832 5355
rect 2780 5312 2832 5321
rect 2964 5312 3016 5364
rect 3516 5312 3568 5364
rect 18420 5312 18472 5364
rect 2320 5244 2372 5296
rect 1400 5219 1452 5228
rect 1400 5185 1409 5219
rect 1409 5185 1443 5219
rect 1443 5185 1452 5219
rect 1400 5176 1452 5185
rect 21548 5219 21600 5228
rect 21548 5185 21557 5219
rect 21557 5185 21591 5219
rect 21591 5185 21600 5219
rect 21548 5176 21600 5185
rect 3148 5108 3200 5160
rect 2228 5040 2280 5092
rect 3884 4972 3936 5024
rect 3549 4870 3601 4922
rect 3613 4870 3665 4922
rect 3677 4870 3729 4922
rect 3741 4870 3793 4922
rect 3805 4870 3857 4922
rect 8747 4870 8799 4922
rect 8811 4870 8863 4922
rect 8875 4870 8927 4922
rect 8939 4870 8991 4922
rect 9003 4870 9055 4922
rect 13945 4870 13997 4922
rect 14009 4870 14061 4922
rect 14073 4870 14125 4922
rect 14137 4870 14189 4922
rect 14201 4870 14253 4922
rect 19143 4870 19195 4922
rect 19207 4870 19259 4922
rect 19271 4870 19323 4922
rect 19335 4870 19387 4922
rect 19399 4870 19451 4922
rect 2044 4768 2096 4820
rect 2688 4768 2740 4820
rect 4068 4700 4120 4752
rect 20996 4675 21048 4684
rect 20996 4641 21005 4675
rect 21005 4641 21039 4675
rect 21039 4641 21048 4675
rect 20996 4632 21048 4641
rect 1400 4607 1452 4616
rect 1400 4573 1409 4607
rect 1409 4573 1443 4607
rect 1443 4573 1452 4607
rect 1400 4564 1452 4573
rect 1676 4607 1728 4616
rect 1676 4573 1685 4607
rect 1685 4573 1719 4607
rect 1719 4573 1728 4607
rect 1676 4564 1728 4573
rect 1952 4607 2004 4616
rect 1952 4573 1961 4607
rect 1961 4573 1995 4607
rect 1995 4573 2004 4607
rect 1952 4564 2004 4573
rect 20720 4607 20772 4616
rect 20720 4573 20729 4607
rect 20729 4573 20763 4607
rect 20763 4573 20772 4607
rect 20720 4564 20772 4573
rect 6148 4326 6200 4378
rect 6212 4326 6264 4378
rect 6276 4326 6328 4378
rect 6340 4326 6392 4378
rect 6404 4326 6456 4378
rect 11346 4326 11398 4378
rect 11410 4326 11462 4378
rect 11474 4326 11526 4378
rect 11538 4326 11590 4378
rect 11602 4326 11654 4378
rect 16544 4326 16596 4378
rect 16608 4326 16660 4378
rect 16672 4326 16724 4378
rect 16736 4326 16788 4378
rect 16800 4326 16852 4378
rect 21742 4326 21794 4378
rect 21806 4326 21858 4378
rect 21870 4326 21922 4378
rect 21934 4326 21986 4378
rect 21998 4326 22050 4378
rect 1400 4224 1452 4276
rect 1676 4267 1728 4276
rect 1676 4233 1685 4267
rect 1685 4233 1719 4267
rect 1719 4233 1728 4267
rect 1676 4224 1728 4233
rect 21088 4267 21140 4276
rect 21088 4233 21097 4267
rect 21097 4233 21131 4267
rect 21131 4233 21140 4267
rect 21088 4224 21140 4233
rect 1400 4131 1452 4140
rect 1400 4097 1409 4131
rect 1409 4097 1443 4131
rect 1443 4097 1452 4131
rect 1400 4088 1452 4097
rect 21272 4131 21324 4140
rect 21272 4097 21281 4131
rect 21281 4097 21315 4131
rect 21315 4097 21324 4131
rect 21272 4088 21324 4097
rect 21548 4131 21600 4140
rect 21548 4097 21557 4131
rect 21557 4097 21591 4131
rect 21591 4097 21600 4131
rect 21548 4088 21600 4097
rect 2872 3952 2924 4004
rect 18328 3952 18380 4004
rect 3549 3782 3601 3834
rect 3613 3782 3665 3834
rect 3677 3782 3729 3834
rect 3741 3782 3793 3834
rect 3805 3782 3857 3834
rect 8747 3782 8799 3834
rect 8811 3782 8863 3834
rect 8875 3782 8927 3834
rect 8939 3782 8991 3834
rect 9003 3782 9055 3834
rect 13945 3782 13997 3834
rect 14009 3782 14061 3834
rect 14073 3782 14125 3834
rect 14137 3782 14189 3834
rect 14201 3782 14253 3834
rect 19143 3782 19195 3834
rect 19207 3782 19259 3834
rect 19271 3782 19323 3834
rect 19335 3782 19387 3834
rect 19399 3782 19451 3834
rect 3056 3680 3108 3732
rect 20352 3680 20404 3732
rect 1400 3519 1452 3528
rect 1400 3485 1409 3519
rect 1409 3485 1443 3519
rect 1443 3485 1452 3519
rect 1400 3476 1452 3485
rect 21548 3519 21600 3528
rect 21548 3485 21557 3519
rect 21557 3485 21591 3519
rect 21591 3485 21600 3519
rect 21548 3476 21600 3485
rect 1676 3340 1728 3392
rect 6148 3238 6200 3290
rect 6212 3238 6264 3290
rect 6276 3238 6328 3290
rect 6340 3238 6392 3290
rect 6404 3238 6456 3290
rect 11346 3238 11398 3290
rect 11410 3238 11462 3290
rect 11474 3238 11526 3290
rect 11538 3238 11590 3290
rect 11602 3238 11654 3290
rect 16544 3238 16596 3290
rect 16608 3238 16660 3290
rect 16672 3238 16724 3290
rect 16736 3238 16788 3290
rect 16800 3238 16852 3290
rect 21742 3238 21794 3290
rect 21806 3238 21858 3290
rect 21870 3238 21922 3290
rect 21934 3238 21986 3290
rect 21998 3238 22050 3290
rect 1860 3179 1912 3188
rect 1860 3145 1869 3179
rect 1869 3145 1903 3179
rect 1903 3145 1912 3179
rect 1860 3136 1912 3145
rect 3424 3136 3476 3188
rect 6000 3136 6052 3188
rect 20444 3136 20496 3188
rect 2964 3068 3016 3120
rect 1400 3043 1452 3052
rect 1400 3009 1409 3043
rect 1409 3009 1443 3043
rect 1443 3009 1452 3043
rect 1400 3000 1452 3009
rect 1676 3043 1728 3052
rect 1676 3009 1685 3043
rect 1685 3009 1719 3043
rect 1719 3009 1728 3043
rect 1676 3000 1728 3009
rect 8668 3000 8720 3052
rect 16120 3000 16172 3052
rect 20628 3000 20680 3052
rect 21272 3043 21324 3052
rect 21272 3009 21281 3043
rect 21281 3009 21315 3043
rect 21315 3009 21324 3043
rect 21272 3000 21324 3009
rect 21548 3043 21600 3052
rect 21548 3009 21557 3043
rect 21557 3009 21591 3043
rect 21591 3009 21600 3043
rect 21548 3000 21600 3009
rect 5816 2864 5868 2916
rect 16856 2907 16908 2916
rect 16856 2873 16865 2907
rect 16865 2873 16899 2907
rect 16899 2873 16908 2907
rect 16856 2864 16908 2873
rect 19984 2864 20036 2916
rect 2780 2796 2832 2848
rect 20260 2796 20312 2848
rect 20720 2796 20772 2848
rect 3549 2694 3601 2746
rect 3613 2694 3665 2746
rect 3677 2694 3729 2746
rect 3741 2694 3793 2746
rect 3805 2694 3857 2746
rect 8747 2694 8799 2746
rect 8811 2694 8863 2746
rect 8875 2694 8927 2746
rect 8939 2694 8991 2746
rect 9003 2694 9055 2746
rect 13945 2694 13997 2746
rect 14009 2694 14061 2746
rect 14073 2694 14125 2746
rect 14137 2694 14189 2746
rect 14201 2694 14253 2746
rect 19143 2694 19195 2746
rect 19207 2694 19259 2746
rect 19271 2694 19323 2746
rect 19335 2694 19387 2746
rect 19399 2694 19451 2746
rect 6552 2592 6604 2644
rect 8668 2592 8720 2644
rect 16120 2635 16172 2644
rect 16120 2601 16129 2635
rect 16129 2601 16163 2635
rect 16163 2601 16172 2635
rect 16120 2592 16172 2601
rect 20628 2592 20680 2644
rect 20812 2592 20864 2644
rect 4620 2456 4672 2508
rect 2228 2431 2280 2440
rect 2228 2397 2237 2431
rect 2237 2397 2271 2431
rect 2271 2397 2280 2431
rect 2228 2388 2280 2397
rect 2320 2431 2372 2440
rect 2320 2397 2329 2431
rect 2329 2397 2363 2431
rect 2363 2397 2372 2431
rect 2320 2388 2372 2397
rect 6736 2388 6788 2440
rect 20628 2388 20680 2440
rect 21272 2431 21324 2440
rect 21272 2397 21281 2431
rect 21281 2397 21315 2431
rect 21315 2397 21324 2431
rect 21272 2388 21324 2397
rect 21548 2431 21600 2440
rect 21548 2397 21557 2431
rect 21557 2397 21591 2431
rect 21591 2397 21600 2431
rect 21548 2388 21600 2397
rect 20168 2320 20220 2372
rect 6828 2252 6880 2304
rect 11704 2252 11756 2304
rect 16028 2295 16080 2304
rect 16028 2261 16037 2295
rect 16037 2261 16071 2295
rect 16071 2261 16080 2295
rect 16028 2252 16080 2261
rect 20628 2295 20680 2304
rect 20628 2261 20637 2295
rect 20637 2261 20671 2295
rect 20671 2261 20680 2295
rect 20628 2252 20680 2261
rect 6148 2150 6200 2202
rect 6212 2150 6264 2202
rect 6276 2150 6328 2202
rect 6340 2150 6392 2202
rect 6404 2150 6456 2202
rect 11346 2150 11398 2202
rect 11410 2150 11462 2202
rect 11474 2150 11526 2202
rect 11538 2150 11590 2202
rect 11602 2150 11654 2202
rect 16544 2150 16596 2202
rect 16608 2150 16660 2202
rect 16672 2150 16724 2202
rect 16736 2150 16788 2202
rect 16800 2150 16852 2202
rect 21742 2150 21794 2202
rect 21806 2150 21858 2202
rect 21870 2150 21922 2202
rect 21934 2150 21986 2202
rect 21998 2150 22050 2202
<< metal2 >>
rect 1674 22200 1730 23000
rect 2042 22200 2098 23000
rect 2410 22200 2466 23000
rect 2778 22200 2834 23000
rect 3146 22200 3202 23000
rect 3514 22200 3570 23000
rect 3882 22200 3938 23000
rect 4250 22200 4306 23000
rect 4618 22200 4674 23000
rect 4986 22200 5042 23000
rect 5354 22200 5410 23000
rect 5722 22200 5778 23000
rect 6090 22200 6146 23000
rect 6458 22200 6514 23000
rect 6826 22200 6882 23000
rect 7194 22200 7250 23000
rect 7562 22200 7618 23000
rect 7930 22200 7986 23000
rect 8298 22200 8354 23000
rect 8404 22222 8616 22250
rect 1688 20618 1716 22200
rect 1688 20590 1808 20618
rect 1676 20460 1728 20466
rect 1676 20402 1728 20408
rect 1492 20256 1544 20262
rect 1492 20198 1544 20204
rect 1504 20097 1532 20198
rect 1490 20088 1546 20097
rect 1490 20023 1546 20032
rect 1492 19712 1544 19718
rect 1490 19680 1492 19689
rect 1544 19680 1546 19689
rect 1490 19615 1546 19624
rect 1492 19168 1544 19174
rect 1492 19110 1544 19116
rect 1504 18873 1532 19110
rect 1490 18864 1546 18873
rect 1490 18799 1546 18808
rect 1492 18624 1544 18630
rect 1492 18566 1544 18572
rect 1504 18465 1532 18566
rect 1490 18456 1546 18465
rect 1688 18426 1716 20402
rect 1780 18834 1808 20590
rect 1858 20496 1914 20505
rect 2056 20466 2084 22200
rect 1858 20431 1914 20440
rect 2044 20460 2096 20466
rect 1872 20058 1900 20431
rect 2096 20420 2176 20448
rect 2044 20402 2096 20408
rect 1860 20052 1912 20058
rect 1860 19994 1912 20000
rect 2044 19372 2096 19378
rect 2044 19314 2096 19320
rect 1858 19272 1914 19281
rect 1858 19207 1860 19216
rect 1912 19207 1914 19216
rect 1860 19178 1912 19184
rect 2056 18970 2084 19314
rect 2044 18964 2096 18970
rect 2044 18906 2096 18912
rect 1860 18896 1912 18902
rect 1860 18838 1912 18844
rect 1768 18828 1820 18834
rect 1768 18770 1820 18776
rect 1490 18391 1546 18400
rect 1676 18420 1728 18426
rect 1676 18362 1728 18368
rect 1400 18352 1452 18358
rect 1400 18294 1452 18300
rect 1308 18148 1360 18154
rect 1308 18090 1360 18096
rect 1320 11694 1348 18090
rect 1412 13410 1440 18294
rect 1872 18154 1900 18838
rect 2044 18760 2096 18766
rect 2044 18702 2096 18708
rect 1952 18284 2004 18290
rect 1952 18226 2004 18232
rect 1860 18148 1912 18154
rect 1860 18090 1912 18096
rect 1492 18080 1544 18086
rect 1490 18048 1492 18057
rect 1544 18048 1546 18057
rect 1490 17983 1546 17992
rect 1964 17762 1992 18226
rect 2056 17882 2084 18702
rect 2148 17898 2176 20420
rect 2424 19938 2452 22200
rect 2792 21026 2820 22200
rect 3054 21312 3110 21321
rect 3054 21247 3110 21256
rect 2792 20998 2912 21026
rect 2778 20904 2834 20913
rect 2778 20839 2834 20848
rect 2688 20324 2740 20330
rect 2688 20266 2740 20272
rect 2424 19910 2544 19938
rect 2516 19854 2544 19910
rect 2228 19848 2280 19854
rect 2228 19790 2280 19796
rect 2504 19848 2556 19854
rect 2556 19796 2636 19802
rect 2504 19790 2636 19796
rect 2240 19446 2268 19790
rect 2320 19780 2372 19786
rect 2516 19774 2636 19790
rect 2320 19722 2372 19728
rect 2332 19514 2360 19722
rect 2320 19508 2372 19514
rect 2320 19450 2372 19456
rect 2228 19440 2280 19446
rect 2228 19382 2280 19388
rect 2320 19372 2372 19378
rect 2320 19314 2372 19320
rect 2044 17876 2096 17882
rect 2148 17870 2268 17898
rect 2332 17882 2360 19314
rect 2412 18964 2464 18970
rect 2412 18906 2464 18912
rect 2424 18834 2452 18906
rect 2412 18828 2464 18834
rect 2412 18770 2464 18776
rect 2412 18284 2464 18290
rect 2412 18226 2464 18232
rect 2044 17818 2096 17824
rect 1964 17734 2176 17762
rect 1584 17672 1636 17678
rect 2044 17672 2096 17678
rect 1584 17614 1636 17620
rect 1858 17640 1914 17649
rect 1492 17536 1544 17542
rect 1492 17478 1544 17484
rect 1504 17241 1532 17478
rect 1490 17232 1546 17241
rect 1490 17167 1546 17176
rect 1492 16992 1544 16998
rect 1492 16934 1544 16940
rect 1504 16833 1532 16934
rect 1490 16824 1546 16833
rect 1490 16759 1546 16768
rect 1492 16448 1544 16454
rect 1490 16416 1492 16425
rect 1544 16416 1546 16425
rect 1490 16351 1546 16360
rect 1492 15904 1544 15910
rect 1492 15846 1544 15852
rect 1504 15609 1532 15846
rect 1490 15600 1546 15609
rect 1490 15535 1546 15544
rect 1492 15360 1544 15366
rect 1492 15302 1544 15308
rect 1504 15201 1532 15302
rect 1490 15192 1546 15201
rect 1490 15127 1546 15136
rect 1492 14816 1544 14822
rect 1490 14784 1492 14793
rect 1544 14784 1546 14793
rect 1490 14719 1546 14728
rect 1492 14272 1544 14278
rect 1492 14214 1544 14220
rect 1504 13977 1532 14214
rect 1596 14074 1624 17614
rect 2044 17614 2096 17620
rect 1858 17575 1914 17584
rect 1872 17542 1900 17575
rect 1860 17536 1912 17542
rect 1860 17478 1912 17484
rect 1766 16552 1822 16561
rect 1766 16487 1822 16496
rect 1676 15496 1728 15502
rect 1676 15438 1728 15444
rect 1688 15162 1716 15438
rect 1676 15156 1728 15162
rect 1676 15098 1728 15104
rect 1780 14498 1808 16487
rect 1952 16108 2004 16114
rect 1952 16050 2004 16056
rect 1858 16008 1914 16017
rect 1858 15943 1860 15952
rect 1912 15943 1914 15952
rect 1860 15914 1912 15920
rect 1964 15706 1992 16050
rect 1952 15700 2004 15706
rect 1952 15642 2004 15648
rect 2056 15638 2084 17614
rect 2148 16250 2176 17734
rect 2240 17610 2268 17870
rect 2320 17876 2372 17882
rect 2320 17818 2372 17824
rect 2320 17672 2372 17678
rect 2320 17614 2372 17620
rect 2228 17604 2280 17610
rect 2228 17546 2280 17552
rect 2228 17196 2280 17202
rect 2228 17138 2280 17144
rect 2136 16244 2188 16250
rect 2136 16186 2188 16192
rect 2240 15706 2268 17138
rect 2332 16794 2360 17614
rect 2320 16788 2372 16794
rect 2320 16730 2372 16736
rect 2424 16561 2452 18226
rect 2504 18148 2556 18154
rect 2504 18090 2556 18096
rect 2410 16552 2466 16561
rect 2320 16516 2372 16522
rect 2410 16487 2466 16496
rect 2320 16458 2372 16464
rect 2332 16250 2360 16458
rect 2412 16448 2464 16454
rect 2412 16390 2464 16396
rect 2320 16244 2372 16250
rect 2320 16186 2372 16192
rect 2320 16108 2372 16114
rect 2424 16096 2452 16390
rect 2372 16068 2452 16096
rect 2320 16050 2372 16056
rect 2332 16017 2360 16050
rect 2318 16008 2374 16017
rect 2318 15943 2374 15952
rect 2320 15904 2372 15910
rect 2320 15846 2372 15852
rect 2228 15700 2280 15706
rect 2228 15642 2280 15648
rect 2044 15632 2096 15638
rect 2044 15574 2096 15580
rect 1952 15020 2004 15026
rect 1952 14962 2004 14968
rect 1964 14618 1992 14962
rect 1952 14612 2004 14618
rect 1952 14554 2004 14560
rect 1780 14470 1992 14498
rect 1768 14408 1820 14414
rect 1768 14350 1820 14356
rect 1858 14376 1914 14385
rect 1584 14068 1636 14074
rect 1584 14010 1636 14016
rect 1490 13968 1546 13977
rect 1490 13903 1546 13912
rect 1676 13932 1728 13938
rect 1676 13874 1728 13880
rect 1492 13728 1544 13734
rect 1492 13670 1544 13676
rect 1504 13569 1532 13670
rect 1490 13560 1546 13569
rect 1688 13530 1716 13874
rect 1490 13495 1546 13504
rect 1676 13524 1728 13530
rect 1676 13466 1728 13472
rect 1412 13382 1624 13410
rect 1400 13320 1452 13326
rect 1400 13262 1452 13268
rect 1412 13161 1440 13262
rect 1398 13152 1454 13161
rect 1398 13087 1454 13096
rect 1490 12336 1546 12345
rect 1490 12271 1546 12280
rect 1504 12238 1532 12271
rect 1492 12232 1544 12238
rect 1492 12174 1544 12180
rect 1400 11756 1452 11762
rect 1400 11698 1452 11704
rect 1308 11688 1360 11694
rect 1308 11630 1360 11636
rect 1412 10713 1440 11698
rect 1490 11112 1546 11121
rect 1490 11047 1492 11056
rect 1544 11047 1546 11056
rect 1492 11018 1544 11024
rect 1398 10704 1454 10713
rect 1398 10639 1454 10648
rect 1490 10296 1546 10305
rect 1490 10231 1546 10240
rect 1504 10062 1532 10231
rect 1492 10056 1544 10062
rect 1492 9998 1544 10004
rect 1504 9722 1532 9998
rect 1492 9716 1544 9722
rect 1492 9658 1544 9664
rect 1400 9512 1452 9518
rect 1400 9454 1452 9460
rect 1412 9081 1440 9454
rect 1398 9072 1454 9081
rect 1398 9007 1454 9016
rect 1308 8492 1360 8498
rect 1308 8434 1360 8440
rect 1320 8265 1348 8434
rect 1306 8256 1362 8265
rect 1306 8191 1362 8200
rect 1412 8090 1440 9007
rect 1596 8634 1624 13382
rect 1676 12368 1728 12374
rect 1674 12336 1676 12345
rect 1728 12336 1730 12345
rect 1674 12271 1730 12280
rect 1780 11898 1808 14350
rect 1858 14311 1914 14320
rect 1872 14278 1900 14311
rect 1860 14272 1912 14278
rect 1860 14214 1912 14220
rect 1964 12322 1992 14470
rect 2044 14408 2096 14414
rect 2044 14350 2096 14356
rect 2056 12442 2084 14350
rect 2332 13410 2360 15846
rect 2412 15496 2464 15502
rect 2412 15438 2464 15444
rect 2424 15162 2452 15438
rect 2412 15156 2464 15162
rect 2412 15098 2464 15104
rect 2516 14890 2544 18090
rect 2608 17882 2636 19774
rect 2700 18902 2728 20266
rect 2792 20058 2820 20839
rect 2884 20466 2912 20998
rect 2872 20460 2924 20466
rect 2872 20402 2924 20408
rect 3068 20058 3096 21247
rect 2780 20052 2832 20058
rect 2780 19994 2832 20000
rect 3056 20052 3108 20058
rect 3056 19994 3108 20000
rect 3160 19854 3188 22200
rect 3528 20466 3556 22200
rect 3516 20460 3568 20466
rect 3436 20420 3516 20448
rect 3240 20392 3292 20398
rect 3240 20334 3292 20340
rect 3330 20360 3386 20369
rect 3252 20058 3280 20334
rect 3330 20295 3386 20304
rect 3240 20052 3292 20058
rect 3240 19994 3292 20000
rect 2872 19848 2924 19854
rect 2872 19790 2924 19796
rect 3148 19848 3200 19854
rect 3148 19790 3200 19796
rect 2884 19514 2912 19790
rect 2872 19508 2924 19514
rect 2872 19450 2924 19456
rect 3056 19440 3108 19446
rect 3056 19382 3108 19388
rect 2964 19372 3016 19378
rect 2964 19314 3016 19320
rect 2872 19304 2924 19310
rect 2870 19272 2872 19281
rect 2924 19272 2926 19281
rect 2870 19207 2926 19216
rect 2688 18896 2740 18902
rect 2688 18838 2740 18844
rect 2688 18420 2740 18426
rect 2688 18362 2740 18368
rect 2700 18193 2728 18362
rect 2778 18320 2834 18329
rect 2778 18255 2834 18264
rect 2686 18184 2742 18193
rect 2686 18119 2742 18128
rect 2688 18080 2740 18086
rect 2792 18034 2820 18255
rect 2884 18154 2912 19207
rect 2976 18358 3004 19314
rect 2964 18352 3016 18358
rect 2964 18294 3016 18300
rect 2872 18148 2924 18154
rect 2872 18090 2924 18096
rect 2740 18028 2820 18034
rect 2688 18022 2820 18028
rect 2700 18006 2820 18022
rect 2596 17876 2648 17882
rect 2596 17818 2648 17824
rect 2596 17740 2648 17746
rect 2596 17682 2648 17688
rect 2504 14884 2556 14890
rect 2504 14826 2556 14832
rect 2332 13382 2452 13410
rect 2320 13320 2372 13326
rect 2320 13262 2372 13268
rect 2228 13184 2280 13190
rect 2228 13126 2280 13132
rect 2240 12782 2268 13126
rect 2332 12986 2360 13262
rect 2320 12980 2372 12986
rect 2320 12922 2372 12928
rect 2228 12776 2280 12782
rect 2226 12744 2228 12753
rect 2280 12744 2282 12753
rect 2226 12679 2282 12688
rect 2044 12436 2096 12442
rect 2044 12378 2096 12384
rect 1964 12294 2084 12322
rect 1952 12232 2004 12238
rect 1952 12174 2004 12180
rect 1860 12164 1912 12170
rect 1860 12106 1912 12112
rect 1872 11937 1900 12106
rect 1858 11928 1914 11937
rect 1768 11892 1820 11898
rect 1858 11863 1914 11872
rect 1768 11834 1820 11840
rect 1676 11688 1728 11694
rect 1674 11656 1676 11665
rect 1728 11656 1730 11665
rect 1674 11591 1730 11600
rect 1964 11354 1992 12174
rect 1952 11348 2004 11354
rect 1952 11290 2004 11296
rect 2056 11098 2084 12294
rect 2136 11756 2188 11762
rect 2136 11698 2188 11704
rect 2148 11529 2176 11698
rect 2134 11520 2190 11529
rect 2134 11455 2190 11464
rect 1688 11070 2084 11098
rect 2228 11144 2280 11150
rect 2424 11098 2452 13382
rect 2504 12844 2556 12850
rect 2504 12786 2556 12792
rect 2228 11086 2280 11092
rect 1584 8628 1636 8634
rect 1584 8570 1636 8576
rect 1688 8514 1716 11070
rect 2044 11008 2096 11014
rect 2044 10950 2096 10956
rect 2056 10810 2084 10950
rect 2240 10810 2268 11086
rect 2332 11070 2452 11098
rect 2044 10804 2096 10810
rect 2044 10746 2096 10752
rect 2228 10804 2280 10810
rect 2228 10746 2280 10752
rect 2332 10690 2360 11070
rect 2412 11008 2464 11014
rect 2412 10950 2464 10956
rect 2424 10810 2452 10950
rect 2412 10804 2464 10810
rect 2412 10746 2464 10752
rect 1768 10668 1820 10674
rect 2332 10662 2452 10690
rect 1768 10610 1820 10616
rect 1504 8486 1716 8514
rect 1400 8084 1452 8090
rect 1400 8026 1452 8032
rect 1398 7848 1454 7857
rect 1398 7783 1454 7792
rect 1412 6798 1440 7783
rect 1504 6882 1532 8486
rect 1504 6866 1624 6882
rect 1504 6860 1636 6866
rect 1504 6854 1584 6860
rect 1584 6802 1636 6808
rect 1400 6792 1452 6798
rect 1676 6792 1728 6798
rect 1400 6734 1452 6740
rect 1582 6760 1638 6769
rect 1676 6734 1728 6740
rect 1582 6695 1638 6704
rect 1596 6662 1624 6695
rect 1584 6656 1636 6662
rect 1688 6633 1716 6734
rect 1584 6598 1636 6604
rect 1674 6624 1730 6633
rect 1674 6559 1730 6568
rect 1780 5914 1808 10610
rect 2318 10568 2374 10577
rect 2318 10503 2374 10512
rect 2332 10266 2360 10503
rect 2320 10260 2372 10266
rect 2320 10202 2372 10208
rect 2228 10192 2280 10198
rect 2042 10160 2098 10169
rect 2228 10134 2280 10140
rect 2042 10095 2044 10104
rect 2096 10095 2098 10104
rect 2044 10066 2096 10072
rect 2136 10056 2188 10062
rect 2136 9998 2188 10004
rect 1860 9988 1912 9994
rect 1860 9930 1912 9936
rect 1872 9489 1900 9930
rect 1952 9920 2004 9926
rect 2148 9897 2176 9998
rect 1952 9862 2004 9868
rect 2134 9888 2190 9897
rect 1858 9480 1914 9489
rect 1858 9415 1914 9424
rect 1964 9330 1992 9862
rect 2134 9823 2190 9832
rect 2240 9625 2268 10134
rect 2226 9616 2282 9625
rect 2226 9551 2282 9560
rect 1872 9302 1992 9330
rect 1768 5908 1820 5914
rect 1768 5850 1820 5856
rect 1398 5808 1454 5817
rect 1398 5743 1454 5752
rect 1674 5808 1730 5817
rect 1674 5743 1730 5752
rect 1412 5710 1440 5743
rect 1400 5704 1452 5710
rect 1400 5646 1452 5652
rect 1582 5672 1638 5681
rect 1582 5607 1638 5616
rect 1596 5574 1624 5607
rect 1584 5568 1636 5574
rect 1584 5510 1636 5516
rect 1398 5400 1454 5409
rect 1688 5370 1716 5743
rect 1398 5335 1454 5344
rect 1676 5364 1728 5370
rect 1412 5234 1440 5335
rect 1676 5306 1728 5312
rect 1400 5228 1452 5234
rect 1400 5170 1452 5176
rect 1398 4992 1454 5001
rect 1398 4927 1454 4936
rect 1412 4622 1440 4927
rect 1400 4616 1452 4622
rect 1676 4616 1728 4622
rect 1400 4558 1452 4564
rect 1674 4584 1676 4593
rect 1728 4584 1730 4593
rect 1412 4282 1440 4558
rect 1674 4519 1730 4528
rect 1688 4282 1716 4519
rect 1400 4276 1452 4282
rect 1400 4218 1452 4224
rect 1676 4276 1728 4282
rect 1676 4218 1728 4224
rect 1400 4140 1452 4146
rect 1400 4082 1452 4088
rect 1412 3777 1440 4082
rect 1398 3768 1454 3777
rect 1398 3703 1454 3712
rect 1400 3528 1452 3534
rect 1400 3470 1452 3476
rect 1412 3369 1440 3470
rect 1676 3392 1728 3398
rect 1398 3360 1454 3369
rect 1676 3334 1728 3340
rect 1398 3295 1454 3304
rect 1688 3058 1716 3334
rect 1872 3194 1900 9302
rect 2228 8968 2280 8974
rect 2228 8910 2280 8916
rect 2240 8673 2268 8910
rect 2226 8664 2282 8673
rect 2226 8599 2282 8608
rect 2044 8492 2096 8498
rect 2044 8434 2096 8440
rect 1952 8424 2004 8430
rect 1952 8366 2004 8372
rect 1964 8090 1992 8366
rect 1952 8084 2004 8090
rect 1952 8026 2004 8032
rect 1952 7336 2004 7342
rect 1952 7278 2004 7284
rect 1964 6361 1992 7278
rect 2056 6662 2084 8434
rect 2136 8288 2188 8294
rect 2136 8230 2188 8236
rect 2148 7954 2176 8230
rect 2136 7948 2188 7954
rect 2136 7890 2188 7896
rect 2148 6866 2176 7890
rect 2424 7478 2452 10662
rect 2516 9178 2544 12786
rect 2608 11778 2636 17682
rect 2964 16720 3016 16726
rect 2964 16662 3016 16668
rect 2872 16652 2924 16658
rect 2872 16594 2924 16600
rect 2778 16144 2834 16153
rect 2778 16079 2780 16088
rect 2832 16079 2834 16088
rect 2780 16050 2832 16056
rect 2780 15020 2832 15026
rect 2780 14962 2832 14968
rect 2792 13530 2820 14962
rect 2780 13524 2832 13530
rect 2780 13466 2832 13472
rect 2686 12200 2742 12209
rect 2686 12135 2742 12144
rect 2700 12102 2728 12135
rect 2688 12096 2740 12102
rect 2688 12038 2740 12044
rect 2608 11750 2728 11778
rect 2596 11688 2648 11694
rect 2596 11630 2648 11636
rect 2608 9382 2636 11630
rect 2700 10849 2728 11750
rect 2780 11008 2832 11014
rect 2780 10950 2832 10956
rect 2686 10840 2742 10849
rect 2792 10810 2820 10950
rect 2686 10775 2742 10784
rect 2780 10804 2832 10810
rect 2780 10746 2832 10752
rect 2688 10668 2740 10674
rect 2688 10610 2740 10616
rect 2700 10266 2728 10610
rect 2688 10260 2740 10266
rect 2688 10202 2740 10208
rect 2884 9466 2912 16594
rect 2976 16046 3004 16662
rect 2964 16040 3016 16046
rect 2964 15982 3016 15988
rect 2964 15904 3016 15910
rect 2964 15846 3016 15852
rect 2976 12238 3004 15846
rect 3068 13462 3096 19382
rect 3160 18426 3188 19790
rect 3240 19712 3292 19718
rect 3240 19654 3292 19660
rect 3252 19514 3280 19654
rect 3344 19514 3372 20295
rect 3240 19508 3292 19514
rect 3240 19450 3292 19456
rect 3332 19508 3384 19514
rect 3332 19450 3384 19456
rect 3240 19372 3292 19378
rect 3240 19314 3292 19320
rect 3332 19372 3384 19378
rect 3332 19314 3384 19320
rect 3252 19009 3280 19314
rect 3238 19000 3294 19009
rect 3238 18935 3294 18944
rect 3344 18902 3372 19314
rect 3240 18896 3292 18902
rect 3240 18838 3292 18844
rect 3332 18896 3384 18902
rect 3332 18838 3384 18844
rect 3148 18420 3200 18426
rect 3148 18362 3200 18368
rect 3252 18154 3280 18838
rect 3330 18728 3386 18737
rect 3330 18663 3386 18672
rect 3148 18148 3200 18154
rect 3148 18090 3200 18096
rect 3240 18148 3292 18154
rect 3240 18090 3292 18096
rect 3160 16436 3188 18090
rect 3344 18086 3372 18663
rect 3436 18290 3464 20420
rect 3516 20402 3568 20408
rect 3549 20156 3857 20165
rect 3549 20154 3555 20156
rect 3611 20154 3635 20156
rect 3691 20154 3715 20156
rect 3771 20154 3795 20156
rect 3851 20154 3857 20156
rect 3611 20102 3613 20154
rect 3793 20102 3795 20154
rect 3549 20100 3555 20102
rect 3611 20100 3635 20102
rect 3691 20100 3715 20102
rect 3771 20100 3795 20102
rect 3851 20100 3857 20102
rect 3549 20091 3857 20100
rect 3516 20052 3568 20058
rect 3516 19994 3568 20000
rect 3528 19334 3556 19994
rect 3896 19854 3924 22200
rect 4264 20534 4292 22200
rect 4252 20528 4304 20534
rect 4252 20470 4304 20476
rect 4528 20528 4580 20534
rect 4528 20470 4580 20476
rect 3976 20392 4028 20398
rect 4344 20392 4396 20398
rect 4028 20352 4108 20380
rect 3976 20334 4028 20340
rect 3974 20088 4030 20097
rect 3974 20023 4030 20032
rect 3884 19848 3936 19854
rect 3884 19790 3936 19796
rect 3790 19408 3846 19417
rect 3790 19343 3792 19352
rect 3528 19306 3648 19334
rect 3844 19343 3846 19352
rect 3792 19314 3844 19320
rect 3620 19242 3648 19306
rect 3608 19236 3660 19242
rect 3608 19178 3660 19184
rect 3549 19068 3857 19077
rect 3549 19066 3555 19068
rect 3611 19066 3635 19068
rect 3691 19066 3715 19068
rect 3771 19066 3795 19068
rect 3851 19066 3857 19068
rect 3611 19014 3613 19066
rect 3793 19014 3795 19066
rect 3549 19012 3555 19014
rect 3611 19012 3635 19014
rect 3691 19012 3715 19014
rect 3771 19012 3795 19014
rect 3851 19012 3857 19014
rect 3549 19003 3857 19012
rect 3514 18728 3570 18737
rect 3514 18663 3570 18672
rect 3528 18630 3556 18663
rect 3516 18624 3568 18630
rect 3516 18566 3568 18572
rect 3896 18426 3924 19790
rect 3988 19514 4016 20023
rect 3976 19508 4028 19514
rect 3976 19450 4028 19456
rect 3976 19372 4028 19378
rect 3976 19314 4028 19320
rect 3988 18970 4016 19314
rect 3976 18964 4028 18970
rect 3976 18906 4028 18912
rect 3976 18760 4028 18766
rect 3976 18702 4028 18708
rect 3884 18420 3936 18426
rect 3884 18362 3936 18368
rect 3988 18358 4016 18702
rect 4080 18426 4108 20352
rect 4344 20334 4396 20340
rect 4252 19848 4304 19854
rect 4252 19790 4304 19796
rect 4160 19712 4212 19718
rect 4160 19654 4212 19660
rect 4172 19310 4200 19654
rect 4160 19304 4212 19310
rect 4160 19246 4212 19252
rect 4160 19168 4212 19174
rect 4158 19136 4160 19145
rect 4212 19136 4214 19145
rect 4158 19071 4214 19080
rect 4068 18420 4120 18426
rect 4068 18362 4120 18368
rect 3976 18352 4028 18358
rect 3976 18294 4028 18300
rect 3424 18284 3476 18290
rect 3424 18226 3476 18232
rect 3332 18080 3384 18086
rect 3332 18022 3384 18028
rect 3240 16992 3292 16998
rect 3240 16934 3292 16940
rect 3252 16590 3280 16934
rect 3240 16584 3292 16590
rect 3240 16526 3292 16532
rect 3160 16408 3280 16436
rect 3056 13456 3108 13462
rect 3056 13398 3108 13404
rect 3056 12844 3108 12850
rect 3056 12786 3108 12792
rect 3148 12844 3200 12850
rect 3148 12786 3200 12792
rect 3068 12442 3096 12786
rect 3056 12436 3108 12442
rect 3056 12378 3108 12384
rect 2964 12232 3016 12238
rect 2964 12174 3016 12180
rect 2964 10600 3016 10606
rect 2964 10542 3016 10548
rect 2976 9654 3004 10542
rect 3056 10124 3108 10130
rect 3056 10066 3108 10072
rect 2964 9648 3016 9654
rect 2964 9590 3016 9596
rect 2792 9438 2912 9466
rect 2596 9376 2648 9382
rect 2596 9318 2648 9324
rect 2504 9172 2556 9178
rect 2504 9114 2556 9120
rect 2792 8922 2820 9438
rect 2872 9376 2924 9382
rect 2872 9318 2924 9324
rect 2884 9042 2912 9318
rect 2872 9036 2924 9042
rect 2872 8978 2924 8984
rect 2700 8894 2820 8922
rect 2504 7948 2556 7954
rect 2504 7890 2556 7896
rect 2412 7472 2464 7478
rect 2412 7414 2464 7420
rect 2516 7342 2544 7890
rect 2700 7886 2728 8894
rect 2780 8832 2832 8838
rect 2780 8774 2832 8780
rect 2792 8634 2820 8774
rect 2780 8628 2832 8634
rect 2780 8570 2832 8576
rect 2872 8628 2924 8634
rect 2872 8570 2924 8576
rect 2780 8424 2832 8430
rect 2780 8366 2832 8372
rect 2792 8090 2820 8366
rect 2780 8084 2832 8090
rect 2780 8026 2832 8032
rect 2688 7880 2740 7886
rect 2688 7822 2740 7828
rect 2228 7336 2280 7342
rect 2504 7336 2556 7342
rect 2228 7278 2280 7284
rect 2410 7304 2466 7313
rect 2240 7041 2268 7278
rect 2504 7278 2556 7284
rect 2596 7336 2648 7342
rect 2596 7278 2648 7284
rect 2410 7239 2466 7248
rect 2226 7032 2282 7041
rect 2226 6967 2282 6976
rect 2136 6860 2188 6866
rect 2136 6802 2188 6808
rect 2044 6656 2096 6662
rect 2044 6598 2096 6604
rect 2136 6656 2188 6662
rect 2136 6598 2188 6604
rect 2148 6474 2176 6598
rect 2056 6446 2176 6474
rect 2240 6458 2268 6967
rect 2228 6452 2280 6458
rect 1950 6352 2006 6361
rect 1950 6287 2006 6296
rect 2056 4826 2084 6446
rect 2228 6394 2280 6400
rect 2228 6248 2280 6254
rect 2226 6216 2228 6225
rect 2320 6248 2372 6254
rect 2280 6216 2282 6225
rect 2320 6190 2372 6196
rect 2226 6151 2282 6160
rect 2136 5568 2188 5574
rect 2136 5510 2188 5516
rect 2148 5370 2176 5510
rect 2136 5364 2188 5370
rect 2136 5306 2188 5312
rect 2240 5098 2268 6151
rect 2332 5302 2360 6190
rect 2424 5778 2452 7239
rect 2608 6662 2636 7278
rect 2596 6656 2648 6662
rect 2596 6598 2648 6604
rect 2608 6322 2636 6598
rect 2596 6316 2648 6322
rect 2596 6258 2648 6264
rect 2412 5772 2464 5778
rect 2412 5714 2464 5720
rect 2700 5642 2728 7822
rect 2884 7546 2912 8570
rect 2872 7540 2924 7546
rect 2872 7482 2924 7488
rect 2780 6928 2832 6934
rect 2780 6870 2832 6876
rect 2792 6322 2820 6870
rect 2976 6866 3004 9590
rect 3068 7970 3096 10066
rect 3160 8634 3188 12786
rect 3252 11257 3280 16408
rect 3344 15910 3372 18022
rect 3549 17980 3857 17989
rect 3549 17978 3555 17980
rect 3611 17978 3635 17980
rect 3691 17978 3715 17980
rect 3771 17978 3795 17980
rect 3851 17978 3857 17980
rect 3611 17926 3613 17978
rect 3793 17926 3795 17978
rect 3549 17924 3555 17926
rect 3611 17924 3635 17926
rect 3691 17924 3715 17926
rect 3771 17924 3795 17926
rect 3851 17924 3857 17926
rect 3549 17915 3857 17924
rect 3549 16892 3857 16901
rect 3549 16890 3555 16892
rect 3611 16890 3635 16892
rect 3691 16890 3715 16892
rect 3771 16890 3795 16892
rect 3851 16890 3857 16892
rect 3611 16838 3613 16890
rect 3793 16838 3795 16890
rect 3549 16836 3555 16838
rect 3611 16836 3635 16838
rect 3691 16836 3715 16838
rect 3771 16836 3795 16838
rect 3851 16836 3857 16838
rect 3549 16827 3857 16836
rect 3988 16182 4016 18294
rect 4068 18080 4120 18086
rect 4066 18048 4068 18057
rect 4120 18048 4122 18057
rect 4066 17983 4122 17992
rect 4160 17196 4212 17202
rect 4160 17138 4212 17144
rect 4172 16794 4200 17138
rect 4160 16788 4212 16794
rect 4160 16730 4212 16736
rect 4160 16584 4212 16590
rect 4160 16526 4212 16532
rect 4172 16250 4200 16526
rect 4160 16244 4212 16250
rect 4160 16186 4212 16192
rect 3976 16176 4028 16182
rect 3882 16144 3938 16153
rect 3976 16118 4028 16124
rect 3882 16079 3938 16088
rect 4068 16108 4120 16114
rect 3332 15904 3384 15910
rect 3332 15846 3384 15852
rect 3549 15804 3857 15813
rect 3549 15802 3555 15804
rect 3611 15802 3635 15804
rect 3691 15802 3715 15804
rect 3771 15802 3795 15804
rect 3851 15802 3857 15804
rect 3611 15750 3613 15802
rect 3793 15750 3795 15802
rect 3549 15748 3555 15750
rect 3611 15748 3635 15750
rect 3691 15748 3715 15750
rect 3771 15748 3795 15750
rect 3851 15748 3857 15750
rect 3549 15739 3857 15748
rect 3549 14716 3857 14725
rect 3549 14714 3555 14716
rect 3611 14714 3635 14716
rect 3691 14714 3715 14716
rect 3771 14714 3795 14716
rect 3851 14714 3857 14716
rect 3611 14662 3613 14714
rect 3793 14662 3795 14714
rect 3549 14660 3555 14662
rect 3611 14660 3635 14662
rect 3691 14660 3715 14662
rect 3771 14660 3795 14662
rect 3851 14660 3857 14662
rect 3549 14651 3857 14660
rect 3424 14408 3476 14414
rect 3424 14350 3476 14356
rect 3436 12714 3464 14350
rect 3549 13628 3857 13637
rect 3549 13626 3555 13628
rect 3611 13626 3635 13628
rect 3691 13626 3715 13628
rect 3771 13626 3795 13628
rect 3851 13626 3857 13628
rect 3611 13574 3613 13626
rect 3793 13574 3795 13626
rect 3549 13572 3555 13574
rect 3611 13572 3635 13574
rect 3691 13572 3715 13574
rect 3771 13572 3795 13574
rect 3851 13572 3857 13574
rect 3549 13563 3857 13572
rect 3424 12708 3476 12714
rect 3424 12650 3476 12656
rect 3549 12540 3857 12549
rect 3549 12538 3555 12540
rect 3611 12538 3635 12540
rect 3691 12538 3715 12540
rect 3771 12538 3795 12540
rect 3851 12538 3857 12540
rect 3611 12486 3613 12538
rect 3793 12486 3795 12538
rect 3549 12484 3555 12486
rect 3611 12484 3635 12486
rect 3691 12484 3715 12486
rect 3771 12484 3795 12486
rect 3851 12484 3857 12486
rect 3549 12475 3857 12484
rect 3896 12442 3924 16079
rect 4068 16050 4120 16056
rect 3976 13320 4028 13326
rect 3976 13262 4028 13268
rect 3988 12646 4016 13262
rect 3976 12640 4028 12646
rect 3976 12582 4028 12588
rect 3884 12436 3936 12442
rect 4080 12434 4108 16050
rect 4160 14816 4212 14822
rect 4160 14758 4212 14764
rect 4172 14414 4200 14758
rect 4160 14408 4212 14414
rect 4160 14350 4212 14356
rect 4160 13932 4212 13938
rect 4160 13874 4212 13880
rect 3884 12378 3936 12384
rect 3988 12406 4108 12434
rect 3549 11452 3857 11461
rect 3549 11450 3555 11452
rect 3611 11450 3635 11452
rect 3691 11450 3715 11452
rect 3771 11450 3795 11452
rect 3851 11450 3857 11452
rect 3611 11398 3613 11450
rect 3793 11398 3795 11450
rect 3549 11396 3555 11398
rect 3611 11396 3635 11398
rect 3691 11396 3715 11398
rect 3771 11396 3795 11398
rect 3851 11396 3857 11398
rect 3549 11387 3857 11396
rect 3238 11248 3294 11257
rect 3238 11183 3294 11192
rect 3240 11144 3292 11150
rect 3240 11086 3292 11092
rect 3252 9382 3280 11086
rect 3332 11076 3384 11082
rect 3332 11018 3384 11024
rect 3344 10130 3372 11018
rect 3988 10810 4016 12406
rect 4068 11552 4120 11558
rect 4068 11494 4120 11500
rect 3976 10804 4028 10810
rect 3976 10746 4028 10752
rect 3884 10600 3936 10606
rect 3884 10542 3936 10548
rect 3424 10464 3476 10470
rect 3424 10406 3476 10412
rect 3332 10124 3384 10130
rect 3332 10066 3384 10072
rect 3436 9722 3464 10406
rect 3549 10364 3857 10373
rect 3549 10362 3555 10364
rect 3611 10362 3635 10364
rect 3691 10362 3715 10364
rect 3771 10362 3795 10364
rect 3851 10362 3857 10364
rect 3611 10310 3613 10362
rect 3793 10310 3795 10362
rect 3549 10308 3555 10310
rect 3611 10308 3635 10310
rect 3691 10308 3715 10310
rect 3771 10308 3795 10310
rect 3851 10308 3857 10310
rect 3549 10299 3857 10308
rect 3896 10266 3924 10542
rect 3884 10260 3936 10266
rect 3884 10202 3936 10208
rect 3988 10062 4016 10746
rect 3976 10056 4028 10062
rect 3976 9998 4028 10004
rect 3514 9888 3570 9897
rect 3514 9823 3570 9832
rect 3424 9716 3476 9722
rect 3424 9658 3476 9664
rect 3332 9512 3384 9518
rect 3332 9454 3384 9460
rect 3424 9512 3476 9518
rect 3424 9454 3476 9460
rect 3528 9466 3556 9823
rect 3976 9580 4028 9586
rect 3976 9522 4028 9528
rect 3240 9376 3292 9382
rect 3240 9318 3292 9324
rect 3344 8634 3372 9454
rect 3148 8628 3200 8634
rect 3148 8570 3200 8576
rect 3332 8628 3384 8634
rect 3332 8570 3384 8576
rect 3332 8424 3384 8430
rect 3332 8366 3384 8372
rect 3068 7942 3188 7970
rect 3056 7812 3108 7818
rect 3056 7754 3108 7760
rect 2964 6860 3016 6866
rect 2964 6802 3016 6808
rect 2872 6656 2924 6662
rect 2872 6598 2924 6604
rect 2780 6316 2832 6322
rect 2780 6258 2832 6264
rect 2778 5944 2834 5953
rect 2778 5879 2834 5888
rect 2688 5636 2740 5642
rect 2688 5578 2740 5584
rect 2320 5296 2372 5302
rect 2320 5238 2372 5244
rect 2228 5092 2280 5098
rect 2228 5034 2280 5040
rect 2700 4826 2728 5578
rect 2792 5370 2820 5879
rect 2884 5846 2912 6598
rect 3068 6497 3096 7754
rect 3054 6488 3110 6497
rect 3054 6423 3110 6432
rect 2964 6384 3016 6390
rect 2964 6326 3016 6332
rect 2872 5840 2924 5846
rect 2872 5782 2924 5788
rect 2872 5568 2924 5574
rect 2872 5510 2924 5516
rect 2780 5364 2832 5370
rect 2780 5306 2832 5312
rect 2044 4820 2096 4826
rect 2044 4762 2096 4768
rect 2688 4820 2740 4826
rect 2688 4762 2740 4768
rect 1952 4616 2004 4622
rect 1952 4558 2004 4564
rect 1964 4185 1992 4558
rect 1950 4176 2006 4185
rect 1950 4111 2006 4120
rect 2884 4010 2912 5510
rect 2976 5370 3004 6326
rect 2964 5364 3016 5370
rect 2964 5306 3016 5312
rect 2872 4004 2924 4010
rect 2872 3946 2924 3952
rect 1860 3188 1912 3194
rect 1860 3130 1912 3136
rect 2976 3126 3004 5306
rect 3068 3738 3096 6423
rect 3160 6254 3188 7942
rect 3344 6798 3372 8366
rect 3436 8362 3464 9454
rect 3528 9438 3924 9466
rect 3549 9276 3857 9285
rect 3549 9274 3555 9276
rect 3611 9274 3635 9276
rect 3691 9274 3715 9276
rect 3771 9274 3795 9276
rect 3851 9274 3857 9276
rect 3611 9222 3613 9274
rect 3793 9222 3795 9274
rect 3549 9220 3555 9222
rect 3611 9220 3635 9222
rect 3691 9220 3715 9222
rect 3771 9220 3795 9222
rect 3851 9220 3857 9222
rect 3549 9211 3857 9220
rect 3424 8356 3476 8362
rect 3424 8298 3476 8304
rect 3549 8188 3857 8197
rect 3549 8186 3555 8188
rect 3611 8186 3635 8188
rect 3691 8186 3715 8188
rect 3771 8186 3795 8188
rect 3851 8186 3857 8188
rect 3611 8134 3613 8186
rect 3793 8134 3795 8186
rect 3549 8132 3555 8134
rect 3611 8132 3635 8134
rect 3691 8132 3715 8134
rect 3771 8132 3795 8134
rect 3851 8132 3857 8134
rect 3549 8123 3857 8132
rect 3424 7812 3476 7818
rect 3424 7754 3476 7760
rect 3436 7449 3464 7754
rect 3516 7744 3568 7750
rect 3516 7686 3568 7692
rect 3422 7440 3478 7449
rect 3422 7375 3478 7384
rect 3528 7324 3556 7686
rect 3896 7478 3924 9438
rect 3988 8022 4016 9522
rect 4080 9518 4108 11494
rect 4172 10810 4200 13874
rect 4264 11898 4292 19790
rect 4356 19530 4384 20334
rect 4434 19816 4490 19825
rect 4434 19751 4490 19760
rect 4448 19718 4476 19751
rect 4436 19712 4488 19718
rect 4436 19654 4488 19660
rect 4356 19502 4476 19530
rect 4344 19304 4396 19310
rect 4344 19246 4396 19252
rect 4356 17338 4384 19246
rect 4448 18698 4476 19502
rect 4436 18692 4488 18698
rect 4436 18634 4488 18640
rect 4344 17332 4396 17338
rect 4344 17274 4396 17280
rect 4448 15609 4476 18634
rect 4540 18426 4568 20470
rect 4632 19854 4660 22200
rect 4712 20392 4764 20398
rect 4712 20334 4764 20340
rect 4724 19990 4752 20334
rect 4896 20256 4948 20262
rect 4894 20224 4896 20233
rect 4948 20224 4950 20233
rect 4894 20159 4950 20168
rect 4712 19984 4764 19990
rect 4712 19926 4764 19932
rect 5000 19854 5028 22200
rect 5368 20618 5396 22200
rect 5368 20602 5580 20618
rect 5736 20602 5764 22200
rect 6104 20890 6132 22200
rect 6012 20862 6132 20890
rect 6012 20602 6040 20862
rect 6472 20856 6500 22200
rect 6472 20828 6592 20856
rect 6148 20700 6456 20709
rect 6148 20698 6154 20700
rect 6210 20698 6234 20700
rect 6290 20698 6314 20700
rect 6370 20698 6394 20700
rect 6450 20698 6456 20700
rect 6210 20646 6212 20698
rect 6392 20646 6394 20698
rect 6148 20644 6154 20646
rect 6210 20644 6234 20646
rect 6290 20644 6314 20646
rect 6370 20644 6394 20646
rect 6450 20644 6456 20646
rect 6148 20635 6456 20644
rect 5368 20596 5592 20602
rect 5368 20590 5540 20596
rect 5540 20538 5592 20544
rect 5724 20596 5776 20602
rect 5724 20538 5776 20544
rect 6000 20596 6052 20602
rect 6000 20538 6052 20544
rect 5448 20528 5500 20534
rect 5354 20496 5410 20505
rect 5448 20470 5500 20476
rect 5354 20431 5410 20440
rect 5264 20256 5316 20262
rect 5264 20198 5316 20204
rect 4620 19848 4672 19854
rect 4620 19790 4672 19796
rect 4988 19848 5040 19854
rect 4988 19790 5040 19796
rect 4632 18426 4660 19790
rect 4712 19780 4764 19786
rect 4896 19780 4948 19786
rect 4764 19740 4896 19768
rect 4712 19722 4764 19728
rect 4896 19722 4948 19728
rect 5000 19514 5028 19790
rect 5172 19712 5224 19718
rect 5172 19654 5224 19660
rect 4988 19508 5040 19514
rect 4988 19450 5040 19456
rect 5080 19508 5132 19514
rect 5080 19450 5132 19456
rect 5092 19334 5120 19450
rect 5184 19378 5212 19654
rect 4712 19304 4764 19310
rect 4712 19246 4764 19252
rect 4896 19304 4948 19310
rect 4896 19246 4948 19252
rect 5000 19306 5120 19334
rect 5172 19372 5224 19378
rect 5172 19314 5224 19320
rect 4528 18420 4580 18426
rect 4528 18362 4580 18368
rect 4620 18420 4672 18426
rect 4620 18362 4672 18368
rect 4724 18222 4752 19246
rect 4804 19168 4856 19174
rect 4804 19110 4856 19116
rect 4816 18714 4844 19110
rect 4908 18970 4936 19246
rect 4896 18964 4948 18970
rect 4896 18906 4948 18912
rect 5000 18902 5028 19306
rect 4988 18896 5040 18902
rect 4988 18838 5040 18844
rect 4816 18686 4936 18714
rect 4804 18624 4856 18630
rect 4804 18566 4856 18572
rect 4712 18216 4764 18222
rect 4712 18158 4764 18164
rect 4712 17196 4764 17202
rect 4712 17138 4764 17144
rect 4724 16250 4752 17138
rect 4712 16244 4764 16250
rect 4712 16186 4764 16192
rect 4434 15600 4490 15609
rect 4434 15535 4490 15544
rect 4620 15428 4672 15434
rect 4620 15370 4672 15376
rect 4528 15360 4580 15366
rect 4528 15302 4580 15308
rect 4540 15162 4568 15302
rect 4436 15156 4488 15162
rect 4436 15098 4488 15104
rect 4528 15156 4580 15162
rect 4528 15098 4580 15104
rect 4344 15020 4396 15026
rect 4344 14962 4396 14968
rect 4356 14618 4384 14962
rect 4344 14612 4396 14618
rect 4344 14554 4396 14560
rect 4448 13954 4476 15098
rect 4528 14272 4580 14278
rect 4528 14214 4580 14220
rect 4540 14074 4568 14214
rect 4528 14068 4580 14074
rect 4528 14010 4580 14016
rect 4448 13926 4568 13954
rect 4436 13184 4488 13190
rect 4436 13126 4488 13132
rect 4448 12442 4476 13126
rect 4436 12436 4488 12442
rect 4436 12378 4488 12384
rect 4252 11892 4304 11898
rect 4252 11834 4304 11840
rect 4344 11144 4396 11150
rect 4250 11112 4306 11121
rect 4344 11086 4396 11092
rect 4250 11047 4306 11056
rect 4264 11014 4292 11047
rect 4252 11008 4304 11014
rect 4252 10950 4304 10956
rect 4160 10804 4212 10810
rect 4160 10746 4212 10752
rect 4160 10600 4212 10606
rect 4160 10542 4212 10548
rect 4172 10198 4200 10542
rect 4252 10464 4304 10470
rect 4252 10406 4304 10412
rect 4160 10192 4212 10198
rect 4160 10134 4212 10140
rect 4068 9512 4120 9518
rect 4068 9454 4120 9460
rect 4172 9364 4200 10134
rect 4264 9654 4292 10406
rect 4356 9926 4384 11086
rect 4434 10840 4490 10849
rect 4434 10775 4490 10784
rect 4448 10062 4476 10775
rect 4436 10056 4488 10062
rect 4436 9998 4488 10004
rect 4344 9920 4396 9926
rect 4344 9862 4396 9868
rect 4252 9648 4304 9654
rect 4252 9590 4304 9596
rect 4080 9336 4200 9364
rect 4080 8430 4108 9336
rect 4160 8492 4212 8498
rect 4160 8434 4212 8440
rect 4068 8424 4120 8430
rect 4068 8366 4120 8372
rect 4080 8294 4108 8366
rect 4068 8288 4120 8294
rect 4068 8230 4120 8236
rect 3976 8016 4028 8022
rect 3976 7958 4028 7964
rect 3974 7848 4030 7857
rect 3974 7783 4030 7792
rect 3884 7472 3936 7478
rect 3884 7414 3936 7420
rect 3436 7296 3556 7324
rect 3332 6792 3384 6798
rect 3332 6734 3384 6740
rect 3240 6656 3292 6662
rect 3240 6598 3292 6604
rect 3148 6248 3200 6254
rect 3148 6190 3200 6196
rect 3148 6112 3200 6118
rect 3148 6054 3200 6060
rect 3160 5166 3188 6054
rect 3252 5914 3280 6598
rect 3330 6488 3386 6497
rect 3330 6423 3332 6432
rect 3384 6423 3386 6432
rect 3332 6394 3384 6400
rect 3332 6316 3384 6322
rect 3332 6258 3384 6264
rect 3240 5908 3292 5914
rect 3240 5850 3292 5856
rect 3344 5642 3372 6258
rect 3332 5636 3384 5642
rect 3332 5578 3384 5584
rect 3148 5160 3200 5166
rect 3148 5102 3200 5108
rect 3056 3732 3108 3738
rect 3056 3674 3108 3680
rect 3436 3194 3464 7296
rect 3549 7100 3857 7109
rect 3549 7098 3555 7100
rect 3611 7098 3635 7100
rect 3691 7098 3715 7100
rect 3771 7098 3795 7100
rect 3851 7098 3857 7100
rect 3611 7046 3613 7098
rect 3793 7046 3795 7098
rect 3549 7044 3555 7046
rect 3611 7044 3635 7046
rect 3691 7044 3715 7046
rect 3771 7044 3795 7046
rect 3851 7044 3857 7046
rect 3549 7035 3857 7044
rect 3608 6928 3660 6934
rect 3608 6870 3660 6876
rect 3516 6656 3568 6662
rect 3516 6598 3568 6604
rect 3528 6458 3556 6598
rect 3516 6452 3568 6458
rect 3516 6394 3568 6400
rect 3620 6390 3648 6870
rect 3988 6866 4016 7783
rect 4172 7546 4200 8434
rect 4356 7750 4384 9862
rect 4540 8022 4568 13926
rect 4632 13512 4660 15370
rect 4712 14544 4764 14550
rect 4712 14486 4764 14492
rect 4724 13802 4752 14486
rect 4816 13852 4844 18566
rect 4908 16522 4936 18686
rect 4896 16516 4948 16522
rect 4896 16458 4948 16464
rect 4896 14884 4948 14890
rect 4896 14826 4948 14832
rect 4908 14074 4936 14826
rect 4896 14068 4948 14074
rect 4896 14010 4948 14016
rect 5000 14006 5028 18838
rect 5172 18624 5224 18630
rect 5172 18566 5224 18572
rect 5080 17536 5132 17542
rect 5080 17478 5132 17484
rect 5092 17202 5120 17478
rect 5080 17196 5132 17202
rect 5080 17138 5132 17144
rect 5080 15088 5132 15094
rect 5080 15030 5132 15036
rect 4988 14000 5040 14006
rect 4988 13942 5040 13948
rect 4816 13824 5028 13852
rect 4712 13796 4764 13802
rect 4712 13738 4764 13744
rect 4632 13484 4752 13512
rect 4724 10810 4752 13484
rect 4896 12776 4948 12782
rect 4896 12718 4948 12724
rect 4908 12238 4936 12718
rect 4896 12232 4948 12238
rect 4896 12174 4948 12180
rect 4896 12096 4948 12102
rect 4896 12038 4948 12044
rect 4804 11824 4856 11830
rect 4804 11766 4856 11772
rect 4816 11150 4844 11766
rect 4804 11144 4856 11150
rect 4804 11086 4856 11092
rect 4620 10804 4672 10810
rect 4620 10746 4672 10752
rect 4712 10804 4764 10810
rect 4712 10746 4764 10752
rect 4632 9994 4660 10746
rect 4816 10606 4844 11086
rect 4804 10600 4856 10606
rect 4804 10542 4856 10548
rect 4804 10124 4856 10130
rect 4804 10066 4856 10072
rect 4620 9988 4672 9994
rect 4620 9930 4672 9936
rect 4528 8016 4580 8022
rect 4528 7958 4580 7964
rect 4344 7744 4396 7750
rect 4344 7686 4396 7692
rect 4540 7546 4568 7958
rect 4160 7540 4212 7546
rect 4160 7482 4212 7488
rect 4528 7540 4580 7546
rect 4528 7482 4580 7488
rect 4068 7472 4120 7478
rect 4068 7414 4120 7420
rect 4080 6866 4108 7414
rect 4160 7200 4212 7206
rect 4158 7168 4160 7177
rect 4212 7168 4214 7177
rect 4158 7103 4214 7112
rect 3976 6860 4028 6866
rect 3976 6802 4028 6808
rect 4068 6860 4120 6866
rect 4068 6802 4120 6808
rect 4436 6860 4488 6866
rect 4436 6802 4488 6808
rect 3884 6792 3936 6798
rect 3884 6734 3936 6740
rect 3608 6384 3660 6390
rect 3608 6326 3660 6332
rect 3549 6012 3857 6021
rect 3549 6010 3555 6012
rect 3611 6010 3635 6012
rect 3691 6010 3715 6012
rect 3771 6010 3795 6012
rect 3851 6010 3857 6012
rect 3611 5958 3613 6010
rect 3793 5958 3795 6010
rect 3549 5956 3555 5958
rect 3611 5956 3635 5958
rect 3691 5956 3715 5958
rect 3771 5956 3795 5958
rect 3851 5956 3857 5958
rect 3549 5947 3857 5956
rect 3516 5636 3568 5642
rect 3516 5578 3568 5584
rect 3528 5370 3556 5578
rect 3516 5364 3568 5370
rect 3516 5306 3568 5312
rect 3896 5030 3924 6734
rect 3976 6724 4028 6730
rect 3976 6666 4028 6672
rect 4068 6724 4120 6730
rect 4068 6666 4120 6672
rect 3988 5574 4016 6666
rect 4080 6254 4108 6666
rect 4068 6248 4120 6254
rect 4068 6190 4120 6196
rect 3976 5568 4028 5574
rect 3976 5510 4028 5516
rect 3884 5024 3936 5030
rect 3884 4966 3936 4972
rect 3549 4924 3857 4933
rect 3549 4922 3555 4924
rect 3611 4922 3635 4924
rect 3691 4922 3715 4924
rect 3771 4922 3795 4924
rect 3851 4922 3857 4924
rect 3611 4870 3613 4922
rect 3793 4870 3795 4922
rect 3549 4868 3555 4870
rect 3611 4868 3635 4870
rect 3691 4868 3715 4870
rect 3771 4868 3795 4870
rect 3851 4868 3857 4870
rect 3549 4859 3857 4868
rect 4080 4758 4108 6190
rect 4448 5778 4476 6802
rect 4540 6390 4568 7482
rect 4632 6662 4660 9930
rect 4712 9920 4764 9926
rect 4712 9862 4764 9868
rect 4724 9722 4752 9862
rect 4712 9716 4764 9722
rect 4712 9658 4764 9664
rect 4712 7744 4764 7750
rect 4712 7686 4764 7692
rect 4620 6656 4672 6662
rect 4620 6598 4672 6604
rect 4528 6384 4580 6390
rect 4528 6326 4580 6332
rect 4436 5772 4488 5778
rect 4436 5714 4488 5720
rect 4068 4752 4120 4758
rect 4068 4694 4120 4700
rect 3549 3836 3857 3845
rect 3549 3834 3555 3836
rect 3611 3834 3635 3836
rect 3691 3834 3715 3836
rect 3771 3834 3795 3836
rect 3851 3834 3857 3836
rect 3611 3782 3613 3834
rect 3793 3782 3795 3834
rect 3549 3780 3555 3782
rect 3611 3780 3635 3782
rect 3691 3780 3715 3782
rect 3771 3780 3795 3782
rect 3851 3780 3857 3782
rect 3549 3771 3857 3780
rect 3424 3188 3476 3194
rect 3424 3130 3476 3136
rect 2964 3120 3016 3126
rect 2964 3062 3016 3068
rect 1400 3052 1452 3058
rect 1400 2994 1452 3000
rect 1676 3052 1728 3058
rect 1676 2994 1728 3000
rect 1412 2961 1440 2994
rect 1398 2952 1454 2961
rect 1398 2887 1454 2896
rect 1688 2553 1716 2994
rect 2780 2848 2832 2854
rect 2780 2790 2832 2796
rect 1674 2544 1730 2553
rect 1674 2479 1730 2488
rect 2228 2440 2280 2446
rect 2228 2382 2280 2388
rect 2320 2440 2372 2446
rect 2320 2382 2372 2388
rect 2240 2145 2268 2382
rect 2226 2136 2282 2145
rect 2226 2071 2282 2080
rect 2332 1578 2360 2382
rect 2792 1737 2820 2790
rect 3549 2748 3857 2757
rect 3549 2746 3555 2748
rect 3611 2746 3635 2748
rect 3691 2746 3715 2748
rect 3771 2746 3795 2748
rect 3851 2746 3857 2748
rect 3611 2694 3613 2746
rect 3793 2694 3795 2746
rect 3549 2692 3555 2694
rect 3611 2692 3635 2694
rect 3691 2692 3715 2694
rect 3771 2692 3795 2694
rect 3851 2692 3857 2694
rect 3549 2683 3857 2692
rect 4632 2514 4660 6598
rect 4724 6458 4752 7686
rect 4816 7342 4844 10066
rect 4804 7336 4856 7342
rect 4804 7278 4856 7284
rect 4804 6792 4856 6798
rect 4804 6734 4856 6740
rect 4712 6452 4764 6458
rect 4712 6394 4764 6400
rect 4816 6322 4844 6734
rect 4908 6662 4936 12038
rect 5000 6798 5028 13824
rect 5092 12102 5120 15030
rect 5080 12096 5132 12102
rect 5080 12038 5132 12044
rect 5184 11370 5212 18566
rect 5276 11762 5304 20198
rect 5368 19174 5396 20431
rect 5356 19168 5408 19174
rect 5356 19110 5408 19116
rect 5460 18426 5488 20470
rect 5540 20460 5592 20466
rect 5540 20402 5592 20408
rect 5816 20460 5868 20466
rect 5816 20402 5868 20408
rect 6368 20460 6420 20466
rect 6368 20402 6420 20408
rect 5552 19145 5580 20402
rect 5724 20324 5776 20330
rect 5724 20266 5776 20272
rect 5632 19780 5684 19786
rect 5632 19722 5684 19728
rect 5644 19310 5672 19722
rect 5632 19304 5684 19310
rect 5632 19246 5684 19252
rect 5538 19136 5594 19145
rect 5538 19071 5594 19080
rect 5644 18902 5672 19246
rect 5632 18896 5684 18902
rect 5632 18838 5684 18844
rect 5448 18420 5500 18426
rect 5448 18362 5500 18368
rect 5356 17196 5408 17202
rect 5356 17138 5408 17144
rect 5368 16658 5396 17138
rect 5356 16652 5408 16658
rect 5356 16594 5408 16600
rect 5368 16046 5396 16594
rect 5448 16108 5500 16114
rect 5448 16050 5500 16056
rect 5356 16040 5408 16046
rect 5356 15982 5408 15988
rect 5460 15706 5488 16050
rect 5448 15700 5500 15706
rect 5448 15642 5500 15648
rect 5448 15564 5500 15570
rect 5448 15506 5500 15512
rect 5356 14952 5408 14958
rect 5356 14894 5408 14900
rect 5368 14550 5396 14894
rect 5356 14544 5408 14550
rect 5356 14486 5408 14492
rect 5460 14482 5488 15506
rect 5540 14884 5592 14890
rect 5540 14826 5592 14832
rect 5448 14476 5500 14482
rect 5448 14418 5500 14424
rect 5356 14272 5408 14278
rect 5356 14214 5408 14220
rect 5368 14074 5396 14214
rect 5356 14068 5408 14074
rect 5356 14010 5408 14016
rect 5460 13870 5488 14418
rect 5552 14414 5580 14826
rect 5540 14408 5592 14414
rect 5540 14350 5592 14356
rect 5448 13864 5500 13870
rect 5448 13806 5500 13812
rect 5540 13524 5592 13530
rect 5540 13466 5592 13472
rect 5356 13252 5408 13258
rect 5356 13194 5408 13200
rect 5368 12850 5396 13194
rect 5448 13184 5500 13190
rect 5448 13126 5500 13132
rect 5356 12844 5408 12850
rect 5356 12786 5408 12792
rect 5368 12434 5396 12786
rect 5460 12714 5488 13126
rect 5552 12986 5580 13466
rect 5632 13388 5684 13394
rect 5632 13330 5684 13336
rect 5540 12980 5592 12986
rect 5540 12922 5592 12928
rect 5644 12866 5672 13330
rect 5552 12838 5672 12866
rect 5448 12708 5500 12714
rect 5448 12650 5500 12656
rect 5368 12406 5488 12434
rect 5356 12096 5408 12102
rect 5356 12038 5408 12044
rect 5264 11756 5316 11762
rect 5264 11698 5316 11704
rect 5184 11342 5304 11370
rect 5172 11212 5224 11218
rect 5172 11154 5224 11160
rect 5184 11121 5212 11154
rect 5170 11112 5226 11121
rect 5080 11076 5132 11082
rect 5170 11047 5226 11056
rect 5080 11018 5132 11024
rect 5092 10606 5120 11018
rect 5172 10736 5224 10742
rect 5172 10678 5224 10684
rect 5080 10600 5132 10606
rect 5080 10542 5132 10548
rect 5092 9722 5120 10542
rect 5184 10470 5212 10678
rect 5172 10464 5224 10470
rect 5172 10406 5224 10412
rect 5184 10266 5212 10406
rect 5172 10260 5224 10266
rect 5172 10202 5224 10208
rect 5172 10056 5224 10062
rect 5170 10024 5172 10033
rect 5224 10024 5226 10033
rect 5170 9959 5226 9968
rect 5276 9761 5304 11342
rect 5368 9897 5396 12038
rect 5460 11558 5488 12406
rect 5448 11552 5500 11558
rect 5448 11494 5500 11500
rect 5354 9888 5410 9897
rect 5354 9823 5410 9832
rect 5262 9752 5318 9761
rect 5080 9716 5132 9722
rect 5262 9687 5318 9696
rect 5080 9658 5132 9664
rect 5172 8900 5224 8906
rect 5172 8842 5224 8848
rect 5184 8362 5212 8842
rect 5172 8356 5224 8362
rect 5172 8298 5224 8304
rect 5184 7954 5212 8298
rect 5172 7948 5224 7954
rect 5172 7890 5224 7896
rect 5080 7744 5132 7750
rect 5080 7686 5132 7692
rect 5264 7744 5316 7750
rect 5264 7686 5316 7692
rect 5092 7546 5120 7686
rect 5080 7540 5132 7546
rect 5080 7482 5132 7488
rect 5276 7478 5304 7686
rect 5552 7546 5580 12838
rect 5736 12481 5764 20266
rect 5828 18358 5856 20402
rect 6380 19961 6408 20402
rect 6366 19952 6422 19961
rect 6366 19887 6422 19896
rect 6000 19848 6052 19854
rect 6000 19790 6052 19796
rect 5908 19440 5960 19446
rect 5908 19382 5960 19388
rect 5920 18426 5948 19382
rect 6012 19242 6040 19790
rect 6148 19612 6456 19621
rect 6148 19610 6154 19612
rect 6210 19610 6234 19612
rect 6290 19610 6314 19612
rect 6370 19610 6394 19612
rect 6450 19610 6456 19612
rect 6210 19558 6212 19610
rect 6392 19558 6394 19610
rect 6148 19556 6154 19558
rect 6210 19556 6234 19558
rect 6290 19556 6314 19558
rect 6370 19556 6394 19558
rect 6450 19556 6456 19558
rect 6148 19547 6456 19556
rect 6000 19236 6052 19242
rect 6000 19178 6052 19184
rect 5908 18420 5960 18426
rect 5908 18362 5960 18368
rect 5816 18352 5868 18358
rect 5816 18294 5868 18300
rect 5722 12472 5778 12481
rect 5644 12416 5722 12434
rect 5644 12407 5778 12416
rect 5644 12406 5764 12407
rect 5644 11694 5672 12406
rect 5724 12368 5776 12374
rect 5724 12310 5776 12316
rect 5736 11898 5764 12310
rect 5724 11892 5776 11898
rect 5724 11834 5776 11840
rect 5632 11688 5684 11694
rect 5632 11630 5684 11636
rect 5632 11552 5684 11558
rect 5632 11494 5684 11500
rect 5644 8566 5672 11494
rect 5724 10192 5776 10198
rect 5724 10134 5776 10140
rect 5736 8906 5764 10134
rect 5724 8900 5776 8906
rect 5724 8842 5776 8848
rect 5632 8560 5684 8566
rect 5632 8502 5684 8508
rect 5644 8022 5672 8502
rect 5632 8016 5684 8022
rect 5632 7958 5684 7964
rect 5448 7540 5500 7546
rect 5448 7482 5500 7488
rect 5540 7540 5592 7546
rect 5540 7482 5592 7488
rect 5264 7472 5316 7478
rect 5264 7414 5316 7420
rect 5356 7472 5408 7478
rect 5356 7414 5408 7420
rect 5262 6896 5318 6905
rect 5368 6882 5396 7414
rect 5460 7002 5488 7482
rect 5448 6996 5500 7002
rect 5448 6938 5500 6944
rect 5368 6854 5488 6882
rect 5262 6831 5318 6840
rect 5276 6798 5304 6831
rect 4988 6792 5040 6798
rect 4988 6734 5040 6740
rect 5264 6792 5316 6798
rect 5264 6734 5316 6740
rect 4896 6656 4948 6662
rect 4896 6598 4948 6604
rect 5264 6656 5316 6662
rect 5264 6598 5316 6604
rect 4804 6316 4856 6322
rect 4804 6258 4856 6264
rect 5276 5642 5304 6598
rect 5460 6254 5488 6854
rect 5540 6860 5592 6866
rect 5724 6860 5776 6866
rect 5592 6820 5724 6848
rect 5540 6802 5592 6808
rect 5724 6802 5776 6808
rect 5356 6248 5408 6254
rect 5356 6190 5408 6196
rect 5448 6248 5500 6254
rect 5448 6190 5500 6196
rect 5368 5914 5396 6190
rect 5356 5908 5408 5914
rect 5356 5850 5408 5856
rect 5264 5636 5316 5642
rect 5264 5578 5316 5584
rect 5828 2922 5856 18294
rect 6012 18154 6040 19178
rect 6564 19174 6592 20828
rect 6840 20534 6868 22200
rect 6828 20528 6880 20534
rect 6828 20470 6880 20476
rect 7012 20528 7064 20534
rect 7012 20470 7064 20476
rect 6828 20256 6880 20262
rect 6828 20198 6880 20204
rect 6840 19854 6868 20198
rect 6828 19848 6880 19854
rect 6828 19790 6880 19796
rect 7024 19718 7052 20470
rect 7104 20460 7156 20466
rect 7208 20448 7236 22200
rect 7380 20596 7432 20602
rect 7380 20538 7432 20544
rect 7156 20420 7236 20448
rect 7104 20402 7156 20408
rect 7116 20058 7144 20402
rect 7196 20256 7248 20262
rect 7196 20198 7248 20204
rect 7104 20052 7156 20058
rect 7104 19994 7156 20000
rect 7012 19712 7064 19718
rect 7012 19654 7064 19660
rect 7102 19544 7158 19553
rect 7102 19479 7158 19488
rect 7116 19446 7144 19479
rect 7104 19440 7156 19446
rect 7104 19382 7156 19388
rect 6736 19372 6788 19378
rect 6736 19314 6788 19320
rect 6644 19236 6696 19242
rect 6644 19178 6696 19184
rect 6184 19168 6236 19174
rect 6184 19110 6236 19116
rect 6552 19168 6604 19174
rect 6552 19110 6604 19116
rect 6196 18766 6224 19110
rect 6656 18970 6684 19178
rect 6644 18964 6696 18970
rect 6644 18906 6696 18912
rect 6276 18896 6328 18902
rect 6460 18896 6512 18902
rect 6328 18856 6460 18884
rect 6276 18838 6328 18844
rect 6460 18838 6512 18844
rect 6552 18828 6604 18834
rect 6552 18770 6604 18776
rect 6184 18760 6236 18766
rect 6184 18702 6236 18708
rect 6564 18698 6592 18770
rect 6552 18692 6604 18698
rect 6552 18634 6604 18640
rect 6550 18592 6606 18601
rect 6148 18524 6456 18533
rect 6550 18527 6606 18536
rect 6148 18522 6154 18524
rect 6210 18522 6234 18524
rect 6290 18522 6314 18524
rect 6370 18522 6394 18524
rect 6450 18522 6456 18524
rect 6210 18470 6212 18522
rect 6392 18470 6394 18522
rect 6148 18468 6154 18470
rect 6210 18468 6234 18470
rect 6290 18468 6314 18470
rect 6370 18468 6394 18470
rect 6450 18468 6456 18470
rect 6148 18459 6456 18468
rect 6000 18148 6052 18154
rect 6000 18090 6052 18096
rect 6012 17882 6040 18090
rect 6564 18057 6592 18527
rect 6656 18358 6684 18906
rect 6644 18352 6696 18358
rect 6644 18294 6696 18300
rect 6644 18148 6696 18154
rect 6644 18090 6696 18096
rect 6550 18048 6606 18057
rect 6550 17983 6606 17992
rect 6000 17876 6052 17882
rect 6000 17818 6052 17824
rect 6656 17542 6684 18090
rect 6644 17536 6696 17542
rect 6644 17478 6696 17484
rect 6148 17436 6456 17445
rect 6148 17434 6154 17436
rect 6210 17434 6234 17436
rect 6290 17434 6314 17436
rect 6370 17434 6394 17436
rect 6450 17434 6456 17436
rect 6210 17382 6212 17434
rect 6392 17382 6394 17434
rect 6148 17380 6154 17382
rect 6210 17380 6234 17382
rect 6290 17380 6314 17382
rect 6370 17380 6394 17382
rect 6450 17380 6456 17382
rect 6148 17371 6456 17380
rect 6656 17202 6684 17478
rect 6748 17202 6776 19314
rect 6920 17876 6972 17882
rect 6920 17818 6972 17824
rect 6828 17604 6880 17610
rect 6828 17546 6880 17552
rect 6644 17196 6696 17202
rect 6644 17138 6696 17144
rect 6736 17196 6788 17202
rect 6736 17138 6788 17144
rect 6184 16992 6236 16998
rect 6184 16934 6236 16940
rect 6552 16992 6604 16998
rect 6552 16934 6604 16940
rect 6196 16590 6224 16934
rect 6564 16658 6592 16934
rect 6656 16794 6684 17138
rect 6840 16998 6868 17546
rect 6828 16992 6880 16998
rect 6828 16934 6880 16940
rect 6644 16788 6696 16794
rect 6644 16730 6696 16736
rect 6552 16652 6604 16658
rect 6552 16594 6604 16600
rect 6184 16584 6236 16590
rect 6184 16526 6236 16532
rect 6148 16348 6456 16357
rect 6148 16346 6154 16348
rect 6210 16346 6234 16348
rect 6290 16346 6314 16348
rect 6370 16346 6394 16348
rect 6450 16346 6456 16348
rect 6210 16294 6212 16346
rect 6392 16294 6394 16346
rect 6148 16292 6154 16294
rect 6210 16292 6234 16294
rect 6290 16292 6314 16294
rect 6370 16292 6394 16294
rect 6450 16292 6456 16294
rect 6148 16283 6456 16292
rect 6276 16040 6328 16046
rect 6276 15982 6328 15988
rect 6288 15706 6316 15982
rect 6368 15972 6420 15978
rect 6368 15914 6420 15920
rect 6380 15706 6408 15914
rect 6276 15700 6328 15706
rect 6276 15642 6328 15648
rect 6368 15700 6420 15706
rect 6368 15642 6420 15648
rect 6564 15570 6592 16594
rect 6656 16250 6684 16730
rect 6644 16244 6696 16250
rect 6644 16186 6696 16192
rect 6552 15564 6604 15570
rect 6552 15506 6604 15512
rect 6656 15502 6684 16186
rect 6644 15496 6696 15502
rect 6550 15464 6606 15473
rect 6644 15438 6696 15444
rect 6550 15399 6552 15408
rect 6604 15399 6606 15408
rect 6552 15370 6604 15376
rect 6148 15260 6456 15269
rect 6148 15258 6154 15260
rect 6210 15258 6234 15260
rect 6290 15258 6314 15260
rect 6370 15258 6394 15260
rect 6450 15258 6456 15260
rect 6210 15206 6212 15258
rect 6392 15206 6394 15258
rect 6148 15204 6154 15206
rect 6210 15204 6234 15206
rect 6290 15204 6314 15206
rect 6370 15204 6394 15206
rect 6450 15204 6456 15206
rect 6148 15195 6456 15204
rect 6564 15094 6592 15370
rect 6656 15162 6684 15438
rect 6644 15156 6696 15162
rect 6644 15098 6696 15104
rect 6552 15088 6604 15094
rect 6552 15030 6604 15036
rect 6656 14414 6684 15098
rect 6736 14816 6788 14822
rect 6736 14758 6788 14764
rect 6644 14408 6696 14414
rect 6644 14350 6696 14356
rect 6000 14272 6052 14278
rect 6000 14214 6052 14220
rect 6012 13394 6040 14214
rect 6148 14172 6456 14181
rect 6148 14170 6154 14172
rect 6210 14170 6234 14172
rect 6290 14170 6314 14172
rect 6370 14170 6394 14172
rect 6450 14170 6456 14172
rect 6210 14118 6212 14170
rect 6392 14118 6394 14170
rect 6148 14116 6154 14118
rect 6210 14116 6234 14118
rect 6290 14116 6314 14118
rect 6370 14116 6394 14118
rect 6450 14116 6456 14118
rect 6148 14107 6456 14116
rect 6656 14074 6684 14350
rect 6748 14346 6776 14758
rect 6736 14340 6788 14346
rect 6736 14282 6788 14288
rect 6184 14068 6236 14074
rect 6184 14010 6236 14016
rect 6644 14068 6696 14074
rect 6644 14010 6696 14016
rect 6092 13932 6144 13938
rect 6092 13874 6144 13880
rect 6104 13462 6132 13874
rect 6196 13530 6224 14010
rect 6644 13932 6696 13938
rect 6644 13874 6696 13880
rect 6184 13524 6236 13530
rect 6184 13466 6236 13472
rect 6092 13456 6144 13462
rect 6092 13398 6144 13404
rect 6000 13388 6052 13394
rect 6000 13330 6052 13336
rect 6148 13084 6456 13093
rect 6148 13082 6154 13084
rect 6210 13082 6234 13084
rect 6290 13082 6314 13084
rect 6370 13082 6394 13084
rect 6450 13082 6456 13084
rect 6210 13030 6212 13082
rect 6392 13030 6394 13082
rect 6148 13028 6154 13030
rect 6210 13028 6234 13030
rect 6290 13028 6314 13030
rect 6370 13028 6394 13030
rect 6450 13028 6456 13030
rect 6148 13019 6456 13028
rect 6000 12980 6052 12986
rect 6656 12968 6684 13874
rect 6000 12922 6052 12928
rect 6288 12940 6684 12968
rect 6012 12102 6040 12922
rect 6092 12776 6144 12782
rect 6092 12718 6144 12724
rect 6104 12306 6132 12718
rect 6288 12646 6316 12940
rect 6368 12844 6420 12850
rect 6368 12786 6420 12792
rect 6276 12640 6328 12646
rect 6276 12582 6328 12588
rect 6380 12442 6408 12786
rect 6368 12436 6420 12442
rect 6368 12378 6420 12384
rect 6748 12306 6776 14282
rect 6828 13184 6880 13190
rect 6828 13126 6880 13132
rect 6840 12986 6868 13126
rect 6828 12980 6880 12986
rect 6828 12922 6880 12928
rect 6092 12300 6144 12306
rect 6092 12242 6144 12248
rect 6736 12300 6788 12306
rect 6736 12242 6788 12248
rect 6644 12232 6696 12238
rect 6840 12186 6868 12922
rect 6644 12174 6696 12180
rect 6000 12096 6052 12102
rect 6000 12038 6052 12044
rect 6012 11778 6040 12038
rect 6148 11996 6456 12005
rect 6148 11994 6154 11996
rect 6210 11994 6234 11996
rect 6290 11994 6314 11996
rect 6370 11994 6394 11996
rect 6450 11994 6456 11996
rect 6210 11942 6212 11994
rect 6392 11942 6394 11994
rect 6148 11940 6154 11942
rect 6210 11940 6234 11942
rect 6290 11940 6314 11942
rect 6370 11940 6394 11942
rect 6450 11940 6456 11942
rect 6148 11931 6456 11940
rect 6656 11898 6684 12174
rect 6748 12158 6868 12186
rect 6748 12102 6776 12158
rect 6736 12096 6788 12102
rect 6736 12038 6788 12044
rect 6644 11892 6696 11898
rect 6644 11834 6696 11840
rect 6012 11762 6132 11778
rect 6012 11756 6144 11762
rect 6012 11750 6092 11756
rect 6092 11698 6144 11704
rect 6276 11756 6328 11762
rect 6276 11698 6328 11704
rect 6644 11756 6696 11762
rect 6644 11698 6696 11704
rect 5908 11280 5960 11286
rect 5960 11228 6040 11234
rect 5908 11222 6040 11228
rect 5920 11206 6040 11222
rect 5908 9580 5960 9586
rect 6012 9568 6040 11206
rect 6288 11082 6316 11698
rect 6552 11144 6604 11150
rect 6552 11086 6604 11092
rect 6276 11076 6328 11082
rect 6276 11018 6328 11024
rect 6148 10908 6456 10917
rect 6148 10906 6154 10908
rect 6210 10906 6234 10908
rect 6290 10906 6314 10908
rect 6370 10906 6394 10908
rect 6450 10906 6456 10908
rect 6210 10854 6212 10906
rect 6392 10854 6394 10906
rect 6148 10852 6154 10854
rect 6210 10852 6234 10854
rect 6290 10852 6314 10854
rect 6370 10852 6394 10854
rect 6450 10852 6456 10854
rect 6148 10843 6456 10852
rect 6564 10538 6592 11086
rect 6552 10532 6604 10538
rect 6552 10474 6604 10480
rect 6368 10464 6420 10470
rect 6368 10406 6420 10412
rect 6380 9926 6408 10406
rect 6564 10062 6592 10474
rect 6552 10056 6604 10062
rect 6552 9998 6604 10004
rect 6368 9920 6420 9926
rect 6368 9862 6420 9868
rect 6148 9820 6456 9829
rect 6148 9818 6154 9820
rect 6210 9818 6234 9820
rect 6290 9818 6314 9820
rect 6370 9818 6394 9820
rect 6450 9818 6456 9820
rect 6210 9766 6212 9818
rect 6392 9766 6394 9818
rect 6148 9764 6154 9766
rect 6210 9764 6234 9766
rect 6290 9764 6314 9766
rect 6370 9764 6394 9766
rect 6450 9764 6456 9766
rect 6148 9755 6456 9764
rect 6564 9602 6592 9998
rect 5960 9540 6040 9568
rect 5908 9522 5960 9528
rect 6012 9382 6040 9540
rect 6380 9574 6592 9602
rect 6380 9518 6408 9574
rect 6368 9512 6420 9518
rect 6368 9454 6420 9460
rect 6000 9376 6052 9382
rect 6000 9318 6052 9324
rect 6012 7313 6040 9318
rect 6380 8974 6408 9454
rect 6368 8968 6420 8974
rect 6420 8916 6592 8922
rect 6368 8910 6592 8916
rect 6380 8894 6592 8910
rect 6148 8732 6456 8741
rect 6148 8730 6154 8732
rect 6210 8730 6234 8732
rect 6290 8730 6314 8732
rect 6370 8730 6394 8732
rect 6450 8730 6456 8732
rect 6210 8678 6212 8730
rect 6392 8678 6394 8730
rect 6148 8676 6154 8678
rect 6210 8676 6234 8678
rect 6290 8676 6314 8678
rect 6370 8676 6394 8678
rect 6450 8676 6456 8678
rect 6148 8667 6456 8676
rect 6564 8566 6592 8894
rect 6552 8560 6604 8566
rect 6472 8520 6552 8548
rect 6472 7886 6500 8520
rect 6552 8502 6604 8508
rect 6460 7880 6512 7886
rect 6460 7822 6512 7828
rect 6550 7848 6606 7857
rect 6550 7783 6606 7792
rect 6564 7750 6592 7783
rect 6552 7744 6604 7750
rect 6552 7686 6604 7692
rect 6148 7644 6456 7653
rect 6148 7642 6154 7644
rect 6210 7642 6234 7644
rect 6290 7642 6314 7644
rect 6370 7642 6394 7644
rect 6450 7642 6456 7644
rect 6210 7590 6212 7642
rect 6392 7590 6394 7642
rect 6148 7588 6154 7590
rect 6210 7588 6234 7590
rect 6290 7588 6314 7590
rect 6370 7588 6394 7590
rect 6450 7588 6456 7590
rect 6148 7579 6456 7588
rect 6564 7478 6592 7686
rect 6552 7472 6604 7478
rect 6552 7414 6604 7420
rect 5998 7304 6054 7313
rect 5998 7239 6054 7248
rect 5906 7168 5962 7177
rect 5906 7103 5962 7112
rect 5920 6934 5948 7103
rect 5908 6928 5960 6934
rect 5908 6870 5960 6876
rect 5908 6656 5960 6662
rect 5908 6598 5960 6604
rect 5920 6458 5948 6598
rect 6148 6556 6456 6565
rect 6148 6554 6154 6556
rect 6210 6554 6234 6556
rect 6290 6554 6314 6556
rect 6370 6554 6394 6556
rect 6450 6554 6456 6556
rect 6210 6502 6212 6554
rect 6392 6502 6394 6554
rect 6148 6500 6154 6502
rect 6210 6500 6234 6502
rect 6290 6500 6314 6502
rect 6370 6500 6394 6502
rect 6450 6500 6456 6502
rect 6148 6491 6456 6500
rect 5908 6452 5960 6458
rect 5908 6394 5960 6400
rect 5908 6248 5960 6254
rect 5906 6216 5908 6225
rect 5960 6216 5962 6225
rect 5906 6151 5962 6160
rect 6148 5468 6456 5477
rect 6148 5466 6154 5468
rect 6210 5466 6234 5468
rect 6290 5466 6314 5468
rect 6370 5466 6394 5468
rect 6450 5466 6456 5468
rect 6210 5414 6212 5466
rect 6392 5414 6394 5466
rect 6148 5412 6154 5414
rect 6210 5412 6234 5414
rect 6290 5412 6314 5414
rect 6370 5412 6394 5414
rect 6450 5412 6456 5414
rect 6148 5403 6456 5412
rect 6148 4380 6456 4389
rect 6148 4378 6154 4380
rect 6210 4378 6234 4380
rect 6290 4378 6314 4380
rect 6370 4378 6394 4380
rect 6450 4378 6456 4380
rect 6210 4326 6212 4378
rect 6392 4326 6394 4378
rect 6148 4324 6154 4326
rect 6210 4324 6234 4326
rect 6290 4324 6314 4326
rect 6370 4324 6394 4326
rect 6450 4324 6456 4326
rect 6148 4315 6456 4324
rect 5998 3496 6054 3505
rect 5998 3431 6054 3440
rect 6012 3194 6040 3431
rect 6148 3292 6456 3301
rect 6148 3290 6154 3292
rect 6210 3290 6234 3292
rect 6290 3290 6314 3292
rect 6370 3290 6394 3292
rect 6450 3290 6456 3292
rect 6210 3238 6212 3290
rect 6392 3238 6394 3290
rect 6148 3236 6154 3238
rect 6210 3236 6234 3238
rect 6290 3236 6314 3238
rect 6370 3236 6394 3238
rect 6450 3236 6456 3238
rect 6148 3227 6456 3236
rect 6000 3188 6052 3194
rect 6000 3130 6052 3136
rect 5816 2916 5868 2922
rect 5816 2858 5868 2864
rect 6656 2774 6684 11698
rect 6748 11608 6776 12038
rect 6748 11580 6868 11608
rect 6736 9920 6788 9926
rect 6736 9862 6788 9868
rect 6748 9586 6776 9862
rect 6736 9580 6788 9586
rect 6736 9522 6788 9528
rect 6840 7818 6868 11580
rect 6932 11354 6960 17818
rect 7208 16114 7236 20198
rect 7288 19916 7340 19922
rect 7288 19858 7340 19864
rect 7300 19689 7328 19858
rect 7392 19718 7420 20538
rect 7576 20534 7604 22200
rect 7564 20528 7616 20534
rect 7564 20470 7616 20476
rect 7840 20460 7892 20466
rect 7944 20448 7972 22200
rect 8312 20534 8340 22200
rect 8300 20528 8352 20534
rect 8300 20470 8352 20476
rect 7892 20420 7972 20448
rect 8024 20460 8076 20466
rect 7840 20402 7892 20408
rect 8024 20402 8076 20408
rect 7472 20256 7524 20262
rect 7472 20198 7524 20204
rect 7656 20256 7708 20262
rect 7656 20198 7708 20204
rect 7380 19712 7432 19718
rect 7286 19680 7342 19689
rect 7380 19654 7432 19660
rect 7286 19615 7342 19624
rect 7300 19417 7328 19615
rect 7286 19408 7342 19417
rect 7286 19343 7342 19352
rect 7392 17882 7420 19654
rect 7380 17876 7432 17882
rect 7380 17818 7432 17824
rect 7196 16108 7248 16114
rect 7196 16050 7248 16056
rect 7484 14414 7512 20198
rect 7564 19984 7616 19990
rect 7564 19926 7616 19932
rect 7576 19378 7604 19926
rect 7564 19372 7616 19378
rect 7564 19314 7616 19320
rect 7576 18834 7604 19314
rect 7564 18828 7616 18834
rect 7564 18770 7616 18776
rect 7668 17678 7696 20198
rect 7748 19780 7800 19786
rect 7748 19722 7800 19728
rect 7656 17672 7708 17678
rect 7656 17614 7708 17620
rect 7760 17542 7788 19722
rect 7852 17882 7880 20402
rect 7930 19544 7986 19553
rect 7930 19479 7932 19488
rect 7984 19479 7986 19488
rect 7932 19450 7984 19456
rect 7932 19168 7984 19174
rect 7932 19110 7984 19116
rect 7944 18426 7972 19110
rect 7932 18420 7984 18426
rect 7932 18362 7984 18368
rect 7840 17876 7892 17882
rect 7840 17818 7892 17824
rect 8036 17814 8064 20402
rect 8116 20392 8168 20398
rect 8116 20334 8168 20340
rect 8312 20346 8340 20470
rect 8404 20466 8432 22222
rect 8588 22114 8616 22222
rect 8666 22200 8722 23000
rect 9034 22200 9090 23000
rect 9402 22200 9458 23000
rect 9770 22200 9826 23000
rect 10138 22200 10194 23000
rect 10506 22200 10562 23000
rect 10874 22200 10930 23000
rect 11242 22200 11298 23000
rect 11610 22200 11666 23000
rect 11978 22200 12034 23000
rect 12346 22200 12402 23000
rect 12714 22200 12770 23000
rect 13082 22200 13138 23000
rect 13450 22200 13506 23000
rect 13556 22222 13768 22250
rect 8680 22114 8708 22200
rect 8588 22086 8708 22114
rect 8944 20868 8996 20874
rect 8944 20810 8996 20816
rect 8956 20602 8984 20810
rect 9048 20602 9076 22200
rect 8944 20596 8996 20602
rect 8944 20538 8996 20544
rect 9036 20596 9088 20602
rect 9036 20538 9088 20544
rect 9220 20596 9272 20602
rect 9220 20538 9272 20544
rect 8392 20460 8444 20466
rect 8392 20402 8444 20408
rect 8668 20392 8720 20398
rect 8128 19718 8156 20334
rect 8312 20318 8432 20346
rect 8668 20334 8720 20340
rect 8208 20256 8260 20262
rect 8208 20198 8260 20204
rect 8300 20256 8352 20262
rect 8300 20198 8352 20204
rect 8220 20097 8248 20198
rect 8206 20088 8262 20097
rect 8206 20023 8262 20032
rect 8116 19712 8168 19718
rect 8116 19654 8168 19660
rect 8312 19553 8340 20198
rect 8114 19544 8170 19553
rect 8114 19479 8170 19488
rect 8298 19544 8354 19553
rect 8298 19479 8354 19488
rect 8128 19378 8156 19479
rect 8300 19440 8352 19446
rect 8298 19408 8300 19417
rect 8352 19408 8354 19417
rect 8116 19372 8168 19378
rect 8298 19343 8354 19352
rect 8116 19314 8168 19320
rect 8298 19272 8354 19281
rect 8298 19207 8354 19216
rect 8116 19168 8168 19174
rect 8114 19136 8116 19145
rect 8168 19136 8170 19145
rect 8114 19071 8170 19080
rect 8312 18154 8340 19207
rect 8300 18148 8352 18154
rect 8300 18090 8352 18096
rect 8312 18057 8340 18090
rect 8298 18048 8354 18057
rect 8298 17983 8354 17992
rect 8404 17882 8432 20318
rect 8576 20324 8628 20330
rect 8576 20266 8628 20272
rect 8484 20256 8536 20262
rect 8484 20198 8536 20204
rect 8496 19990 8524 20198
rect 8484 19984 8536 19990
rect 8484 19926 8536 19932
rect 8484 19508 8536 19514
rect 8484 19450 8536 19456
rect 8392 17876 8444 17882
rect 8392 17818 8444 17824
rect 8024 17808 8076 17814
rect 8024 17750 8076 17756
rect 8208 17740 8260 17746
rect 8260 17700 8340 17728
rect 8208 17682 8260 17688
rect 8024 17672 8076 17678
rect 8076 17632 8156 17660
rect 8024 17614 8076 17620
rect 7748 17536 7800 17542
rect 7748 17478 7800 17484
rect 7564 17264 7616 17270
rect 7564 17206 7616 17212
rect 7576 15910 7604 17206
rect 7932 16992 7984 16998
rect 7932 16934 7984 16940
rect 7564 15904 7616 15910
rect 7564 15846 7616 15852
rect 7576 15026 7604 15846
rect 7944 15570 7972 16934
rect 8024 16448 8076 16454
rect 8024 16390 8076 16396
rect 7932 15564 7984 15570
rect 7932 15506 7984 15512
rect 7748 15428 7800 15434
rect 7748 15370 7800 15376
rect 7564 15020 7616 15026
rect 7564 14962 7616 14968
rect 7760 14618 7788 15370
rect 8036 15026 8064 16390
rect 8024 15020 8076 15026
rect 8128 15008 8156 17632
rect 8208 17604 8260 17610
rect 8208 17546 8260 17552
rect 8220 17134 8248 17546
rect 8312 17202 8340 17700
rect 8300 17196 8352 17202
rect 8300 17138 8352 17144
rect 8208 17128 8260 17134
rect 8208 17070 8260 17076
rect 8220 16794 8248 17070
rect 8208 16788 8260 16794
rect 8208 16730 8260 16736
rect 8496 16674 8524 19450
rect 8588 18358 8616 20266
rect 8680 20058 8708 20334
rect 9048 20244 9076 20538
rect 9048 20216 9168 20244
rect 8747 20156 9055 20165
rect 8747 20154 8753 20156
rect 8809 20154 8833 20156
rect 8889 20154 8913 20156
rect 8969 20154 8993 20156
rect 9049 20154 9055 20156
rect 8809 20102 8811 20154
rect 8991 20102 8993 20154
rect 8747 20100 8753 20102
rect 8809 20100 8833 20102
rect 8889 20100 8913 20102
rect 8969 20100 8993 20102
rect 9049 20100 9055 20102
rect 8747 20091 9055 20100
rect 8668 20052 8720 20058
rect 8668 19994 8720 20000
rect 8944 19780 8996 19786
rect 8944 19722 8996 19728
rect 8956 19689 8984 19722
rect 9036 19712 9088 19718
rect 8942 19680 8998 19689
rect 9036 19654 9088 19660
rect 8942 19615 8998 19624
rect 9048 19378 9076 19654
rect 8668 19372 8720 19378
rect 8668 19314 8720 19320
rect 9036 19372 9088 19378
rect 9036 19314 9088 19320
rect 8680 18426 8708 19314
rect 8747 19068 9055 19077
rect 8747 19066 8753 19068
rect 8809 19066 8833 19068
rect 8889 19066 8913 19068
rect 8969 19066 8993 19068
rect 9049 19066 9055 19068
rect 8809 19014 8811 19066
rect 8991 19014 8993 19066
rect 8747 19012 8753 19014
rect 8809 19012 8833 19014
rect 8889 19012 8913 19014
rect 8969 19012 8993 19014
rect 9049 19012 9055 19014
rect 8747 19003 9055 19012
rect 8760 18760 8812 18766
rect 8760 18702 8812 18708
rect 8668 18420 8720 18426
rect 8668 18362 8720 18368
rect 8576 18352 8628 18358
rect 8576 18294 8628 18300
rect 8772 18290 8800 18702
rect 9036 18624 9088 18630
rect 9036 18566 9088 18572
rect 8760 18284 8812 18290
rect 8760 18226 8812 18232
rect 9048 18086 9076 18566
rect 9036 18080 9088 18086
rect 9036 18022 9088 18028
rect 8747 17980 9055 17989
rect 8747 17978 8753 17980
rect 8809 17978 8833 17980
rect 8889 17978 8913 17980
rect 8969 17978 8993 17980
rect 9049 17978 9055 17980
rect 8809 17926 8811 17978
rect 8991 17926 8993 17978
rect 8747 17924 8753 17926
rect 8809 17924 8833 17926
rect 8889 17924 8913 17926
rect 8969 17924 8993 17926
rect 9049 17924 9055 17926
rect 8747 17915 9055 17924
rect 9140 17882 9168 20216
rect 9232 19514 9260 20538
rect 9416 20330 9444 22200
rect 9784 20602 9812 22200
rect 9772 20596 9824 20602
rect 9772 20538 9824 20544
rect 9588 20460 9640 20466
rect 9588 20402 9640 20408
rect 9404 20324 9456 20330
rect 9404 20266 9456 20272
rect 9312 20256 9364 20262
rect 9312 20198 9364 20204
rect 9496 20256 9548 20262
rect 9496 20198 9548 20204
rect 9220 19508 9272 19514
rect 9220 19450 9272 19456
rect 9220 18692 9272 18698
rect 9220 18634 9272 18640
rect 8760 17876 8812 17882
rect 8760 17818 8812 17824
rect 9128 17876 9180 17882
rect 9128 17818 9180 17824
rect 8772 17678 8800 17818
rect 8760 17672 8812 17678
rect 8760 17614 8812 17620
rect 8576 17604 8628 17610
rect 8576 17546 8628 17552
rect 8312 16646 8524 16674
rect 8208 16108 8260 16114
rect 8208 16050 8260 16056
rect 8220 15434 8248 16050
rect 8208 15428 8260 15434
rect 8208 15370 8260 15376
rect 8208 15020 8260 15026
rect 8128 14980 8208 15008
rect 8024 14962 8076 14968
rect 8208 14962 8260 14968
rect 7748 14612 7800 14618
rect 7748 14554 7800 14560
rect 7472 14408 7524 14414
rect 7472 14350 7524 14356
rect 7760 13734 7788 14554
rect 7564 13728 7616 13734
rect 7564 13670 7616 13676
rect 7748 13728 7800 13734
rect 7748 13670 7800 13676
rect 7932 13728 7984 13734
rect 7932 13670 7984 13676
rect 7104 13252 7156 13258
rect 7104 13194 7156 13200
rect 7288 13252 7340 13258
rect 7288 13194 7340 13200
rect 7116 13138 7144 13194
rect 7116 13110 7236 13138
rect 7208 12918 7236 13110
rect 7012 12912 7064 12918
rect 7012 12854 7064 12860
rect 7196 12912 7248 12918
rect 7196 12854 7248 12860
rect 7024 11558 7052 12854
rect 7104 12300 7156 12306
rect 7104 12242 7156 12248
rect 7012 11552 7064 11558
rect 7012 11494 7064 11500
rect 6920 11348 6972 11354
rect 6920 11290 6972 11296
rect 6828 7812 6880 7818
rect 6828 7754 6880 7760
rect 6736 7540 6788 7546
rect 6736 7482 6788 7488
rect 6564 2746 6684 2774
rect 6564 2650 6592 2746
rect 6552 2644 6604 2650
rect 6552 2586 6604 2592
rect 4620 2508 4672 2514
rect 4620 2450 4672 2456
rect 6748 2446 6776 7482
rect 7116 6905 7144 12242
rect 7300 11354 7328 13194
rect 7576 13190 7604 13670
rect 7944 13394 7972 13670
rect 7748 13388 7800 13394
rect 7748 13330 7800 13336
rect 7932 13388 7984 13394
rect 7932 13330 7984 13336
rect 7564 13184 7616 13190
rect 7564 13126 7616 13132
rect 7760 12850 7788 13330
rect 7748 12844 7800 12850
rect 7748 12786 7800 12792
rect 7654 12472 7710 12481
rect 7654 12407 7710 12416
rect 7668 12170 7696 12407
rect 7380 12164 7432 12170
rect 7380 12106 7432 12112
rect 7656 12164 7708 12170
rect 7656 12106 7708 12112
rect 7288 11348 7340 11354
rect 7288 11290 7340 11296
rect 7392 10742 7420 12106
rect 7760 11898 7788 12786
rect 7840 12776 7892 12782
rect 7840 12718 7892 12724
rect 7852 12238 7880 12718
rect 8036 12374 8064 14962
rect 8116 14884 8168 14890
rect 8116 14826 8168 14832
rect 8128 13326 8156 14826
rect 8312 14822 8340 16646
rect 8392 16516 8444 16522
rect 8392 16458 8444 16464
rect 8300 14816 8352 14822
rect 8300 14758 8352 14764
rect 8312 14414 8340 14758
rect 8300 14408 8352 14414
rect 8300 14350 8352 14356
rect 8116 13320 8168 13326
rect 8116 13262 8168 13268
rect 8208 13320 8260 13326
rect 8208 13262 8260 13268
rect 8220 12889 8248 13262
rect 8300 13184 8352 13190
rect 8300 13126 8352 13132
rect 8312 12986 8340 13126
rect 8300 12980 8352 12986
rect 8300 12922 8352 12928
rect 8206 12880 8262 12889
rect 8206 12815 8262 12824
rect 8300 12640 8352 12646
rect 8300 12582 8352 12588
rect 8024 12368 8076 12374
rect 8024 12310 8076 12316
rect 7840 12232 7892 12238
rect 7840 12174 7892 12180
rect 7748 11892 7800 11898
rect 7748 11834 7800 11840
rect 8036 11558 8064 12310
rect 8312 12306 8340 12582
rect 8116 12300 8168 12306
rect 8116 12242 8168 12248
rect 8300 12300 8352 12306
rect 8300 12242 8352 12248
rect 8128 11626 8156 12242
rect 8404 12238 8432 16458
rect 8588 15094 8616 17546
rect 8747 16892 9055 16901
rect 8747 16890 8753 16892
rect 8809 16890 8833 16892
rect 8889 16890 8913 16892
rect 8969 16890 8993 16892
rect 9049 16890 9055 16892
rect 8809 16838 8811 16890
rect 8991 16838 8993 16890
rect 8747 16836 8753 16838
rect 8809 16836 8833 16838
rect 8889 16836 8913 16838
rect 8969 16836 8993 16838
rect 9049 16836 9055 16838
rect 8747 16827 9055 16836
rect 9232 16454 9260 18634
rect 9220 16448 9272 16454
rect 9220 16390 9272 16396
rect 9232 16046 9260 16390
rect 9220 16040 9272 16046
rect 9220 15982 9272 15988
rect 8747 15804 9055 15813
rect 8747 15802 8753 15804
rect 8809 15802 8833 15804
rect 8889 15802 8913 15804
rect 8969 15802 8993 15804
rect 9049 15802 9055 15804
rect 8809 15750 8811 15802
rect 8991 15750 8993 15802
rect 8747 15748 8753 15750
rect 8809 15748 8833 15750
rect 8889 15748 8913 15750
rect 8969 15748 8993 15750
rect 9049 15748 9055 15750
rect 8747 15739 9055 15748
rect 9218 15600 9274 15609
rect 9218 15535 9274 15544
rect 9128 15156 9180 15162
rect 9128 15098 9180 15104
rect 8576 15088 8628 15094
rect 8576 15030 8628 15036
rect 8668 14816 8720 14822
rect 8668 14758 8720 14764
rect 8576 14476 8628 14482
rect 8576 14418 8628 14424
rect 8588 13938 8616 14418
rect 8484 13932 8536 13938
rect 8484 13874 8536 13880
rect 8576 13932 8628 13938
rect 8576 13874 8628 13880
rect 8496 13530 8524 13874
rect 8484 13524 8536 13530
rect 8484 13466 8536 13472
rect 8680 12986 8708 14758
rect 8747 14716 9055 14725
rect 8747 14714 8753 14716
rect 8809 14714 8833 14716
rect 8889 14714 8913 14716
rect 8969 14714 8993 14716
rect 9049 14714 9055 14716
rect 8809 14662 8811 14714
rect 8991 14662 8993 14714
rect 8747 14660 8753 14662
rect 8809 14660 8833 14662
rect 8889 14660 8913 14662
rect 8969 14660 8993 14662
rect 9049 14660 9055 14662
rect 8747 14651 9055 14660
rect 9140 14618 9168 15098
rect 9128 14612 9180 14618
rect 9128 14554 9180 14560
rect 8747 13628 9055 13637
rect 8747 13626 8753 13628
rect 8809 13626 8833 13628
rect 8889 13626 8913 13628
rect 8969 13626 8993 13628
rect 9049 13626 9055 13628
rect 8809 13574 8811 13626
rect 8991 13574 8993 13626
rect 8747 13572 8753 13574
rect 8809 13572 8833 13574
rect 8889 13572 8913 13574
rect 8969 13572 8993 13574
rect 9049 13572 9055 13574
rect 8747 13563 9055 13572
rect 8758 13424 8814 13433
rect 8758 13359 8814 13368
rect 8668 12980 8720 12986
rect 8668 12922 8720 12928
rect 8772 12918 8800 13359
rect 8760 12912 8812 12918
rect 8760 12854 8812 12860
rect 8747 12540 9055 12549
rect 8747 12538 8753 12540
rect 8809 12538 8833 12540
rect 8889 12538 8913 12540
rect 8969 12538 8993 12540
rect 9049 12538 9055 12540
rect 8809 12486 8811 12538
rect 8991 12486 8993 12538
rect 8747 12484 8753 12486
rect 8809 12484 8833 12486
rect 8889 12484 8913 12486
rect 8969 12484 8993 12486
rect 9049 12484 9055 12486
rect 8747 12475 9055 12484
rect 9232 12424 9260 15535
rect 9324 15502 9352 20198
rect 9404 19984 9456 19990
rect 9404 19926 9456 19932
rect 9416 19786 9444 19926
rect 9404 19780 9456 19786
rect 9404 19722 9456 19728
rect 9508 19334 9536 20198
rect 9600 19990 9628 20402
rect 9680 20324 9732 20330
rect 9680 20266 9732 20272
rect 9588 19984 9640 19990
rect 9588 19926 9640 19932
rect 9416 19306 9536 19334
rect 9416 19292 9444 19306
rect 9407 19264 9444 19292
rect 9407 18986 9435 19264
rect 9600 19258 9628 19926
rect 9692 19854 9720 20266
rect 9784 20074 9812 20538
rect 9864 20460 9916 20466
rect 9864 20402 9916 20408
rect 9876 20330 9904 20402
rect 9864 20324 9916 20330
rect 9864 20266 9916 20272
rect 9956 20256 10008 20262
rect 9956 20198 10008 20204
rect 9784 20046 9904 20074
rect 9772 19916 9824 19922
rect 9772 19858 9824 19864
rect 9680 19848 9732 19854
rect 9680 19790 9732 19796
rect 9680 19712 9732 19718
rect 9678 19680 9680 19689
rect 9732 19680 9734 19689
rect 9678 19615 9734 19624
rect 9680 19508 9732 19514
rect 9680 19450 9732 19456
rect 9508 19230 9628 19258
rect 9508 19224 9536 19230
rect 9499 19196 9536 19224
rect 9499 18986 9527 19196
rect 9692 19174 9720 19450
rect 9784 19242 9812 19858
rect 9772 19236 9824 19242
rect 9772 19178 9824 19184
rect 9680 19168 9732 19174
rect 9680 19110 9732 19116
rect 9407 18958 9444 18986
rect 9499 18958 9628 18986
rect 9416 17610 9444 18958
rect 9496 18760 9548 18766
rect 9496 18702 9548 18708
rect 9508 18358 9536 18702
rect 9600 18426 9628 18958
rect 9680 18896 9732 18902
rect 9680 18838 9732 18844
rect 9588 18420 9640 18426
rect 9588 18362 9640 18368
rect 9496 18352 9548 18358
rect 9496 18294 9548 18300
rect 9496 18080 9548 18086
rect 9496 18022 9548 18028
rect 9404 17604 9456 17610
rect 9404 17546 9456 17552
rect 9402 17504 9458 17513
rect 9402 17439 9458 17448
rect 9416 17338 9444 17439
rect 9404 17332 9456 17338
rect 9404 17274 9456 17280
rect 9312 15496 9364 15502
rect 9312 15438 9364 15444
rect 9324 12850 9352 15438
rect 9404 14272 9456 14278
rect 9404 14214 9456 14220
rect 9312 12844 9364 12850
rect 9312 12786 9364 12792
rect 9416 12782 9444 14214
rect 9508 12986 9536 18022
rect 9692 17728 9720 18838
rect 9784 18698 9812 19178
rect 9772 18692 9824 18698
rect 9772 18634 9824 18640
rect 9876 17882 9904 20046
rect 9864 17876 9916 17882
rect 9864 17818 9916 17824
rect 9772 17740 9824 17746
rect 9692 17700 9772 17728
rect 9772 17682 9824 17688
rect 9680 17536 9732 17542
rect 9680 17478 9732 17484
rect 9692 17338 9720 17478
rect 9680 17332 9732 17338
rect 9680 17274 9732 17280
rect 9784 17134 9812 17165
rect 9772 17128 9824 17134
rect 9770 17096 9772 17105
rect 9824 17096 9826 17105
rect 9770 17031 9826 17040
rect 9784 13326 9812 17031
rect 9864 15904 9916 15910
rect 9864 15846 9916 15852
rect 9876 15366 9904 15846
rect 9864 15360 9916 15366
rect 9864 15302 9916 15308
rect 9772 13320 9824 13326
rect 9772 13262 9824 13268
rect 9680 13184 9732 13190
rect 9680 13126 9732 13132
rect 9772 13184 9824 13190
rect 9772 13126 9824 13132
rect 9692 12986 9720 13126
rect 9784 12986 9812 13126
rect 9496 12980 9548 12986
rect 9496 12922 9548 12928
rect 9680 12980 9732 12986
rect 9680 12922 9732 12928
rect 9772 12980 9824 12986
rect 9772 12922 9824 12928
rect 9404 12776 9456 12782
rect 9404 12718 9456 12724
rect 9508 12646 9536 12922
rect 9692 12646 9720 12922
rect 9496 12640 9548 12646
rect 9496 12582 9548 12588
rect 9680 12640 9732 12646
rect 9680 12582 9732 12588
rect 9496 12436 9548 12442
rect 9232 12396 9352 12424
rect 9220 12300 9272 12306
rect 9220 12242 9272 12248
rect 8392 12232 8444 12238
rect 8392 12174 8444 12180
rect 8668 12096 8720 12102
rect 8668 12038 8720 12044
rect 8300 11688 8352 11694
rect 8300 11630 8352 11636
rect 8116 11620 8168 11626
rect 8116 11562 8168 11568
rect 8024 11552 8076 11558
rect 8024 11494 8076 11500
rect 8128 11082 8156 11562
rect 8312 11082 8340 11630
rect 8680 11558 8708 12038
rect 9128 11756 9180 11762
rect 9128 11698 9180 11704
rect 8668 11552 8720 11558
rect 8668 11494 8720 11500
rect 8680 11257 8708 11494
rect 8747 11452 9055 11461
rect 8747 11450 8753 11452
rect 8809 11450 8833 11452
rect 8889 11450 8913 11452
rect 8969 11450 8993 11452
rect 9049 11450 9055 11452
rect 8809 11398 8811 11450
rect 8991 11398 8993 11450
rect 8747 11396 8753 11398
rect 8809 11396 8833 11398
rect 8889 11396 8913 11398
rect 8969 11396 8993 11398
rect 9049 11396 9055 11398
rect 8747 11387 9055 11396
rect 9140 11354 9168 11698
rect 9128 11348 9180 11354
rect 9128 11290 9180 11296
rect 8666 11248 8722 11257
rect 8484 11212 8536 11218
rect 8666 11183 8722 11192
rect 8484 11154 8536 11160
rect 8116 11076 8168 11082
rect 8116 11018 8168 11024
rect 8300 11076 8352 11082
rect 8300 11018 8352 11024
rect 7380 10736 7432 10742
rect 7380 10678 7432 10684
rect 7392 9178 7420 10678
rect 8024 9988 8076 9994
rect 8024 9930 8076 9936
rect 8036 9722 8064 9930
rect 8206 9752 8262 9761
rect 8024 9716 8076 9722
rect 8206 9687 8262 9696
rect 8024 9658 8076 9664
rect 7932 9580 7984 9586
rect 7932 9522 7984 9528
rect 7748 9444 7800 9450
rect 7748 9386 7800 9392
rect 7380 9172 7432 9178
rect 7380 9114 7432 9120
rect 7760 8838 7788 9386
rect 7944 9382 7972 9522
rect 7932 9376 7984 9382
rect 7932 9318 7984 9324
rect 7944 9110 7972 9318
rect 7840 9104 7892 9110
rect 7840 9046 7892 9052
rect 7932 9104 7984 9110
rect 7932 9046 7984 9052
rect 7748 8832 7800 8838
rect 7668 8792 7748 8820
rect 7380 8492 7432 8498
rect 7380 8434 7432 8440
rect 7392 8022 7420 8434
rect 7668 8430 7696 8792
rect 7748 8774 7800 8780
rect 7852 8634 7880 9046
rect 8036 9042 8064 9658
rect 8116 9376 8168 9382
rect 8116 9318 8168 9324
rect 8024 9036 8076 9042
rect 8024 8978 8076 8984
rect 8128 8945 8156 9318
rect 8220 8974 8248 9687
rect 8208 8968 8260 8974
rect 8114 8936 8170 8945
rect 8208 8910 8260 8916
rect 8114 8871 8170 8880
rect 8128 8838 8156 8871
rect 8116 8832 8168 8838
rect 8116 8774 8168 8780
rect 7840 8628 7892 8634
rect 7840 8570 7892 8576
rect 7656 8424 7708 8430
rect 7656 8366 7708 8372
rect 8496 8294 8524 11154
rect 9232 11150 9260 12242
rect 9324 12170 9352 12396
rect 9496 12378 9548 12384
rect 9772 12436 9824 12442
rect 9772 12378 9824 12384
rect 9508 12238 9536 12378
rect 9496 12232 9548 12238
rect 9496 12174 9548 12180
rect 9784 12170 9812 12378
rect 9312 12164 9364 12170
rect 9312 12106 9364 12112
rect 9772 12164 9824 12170
rect 9772 12106 9824 12112
rect 9404 11756 9456 11762
rect 9404 11698 9456 11704
rect 9680 11756 9732 11762
rect 9680 11698 9732 11704
rect 9220 11144 9272 11150
rect 9220 11086 9272 11092
rect 9416 11082 9444 11698
rect 9404 11076 9456 11082
rect 9404 11018 9456 11024
rect 8747 10364 9055 10373
rect 8747 10362 8753 10364
rect 8809 10362 8833 10364
rect 8889 10362 8913 10364
rect 8969 10362 8993 10364
rect 9049 10362 9055 10364
rect 8809 10310 8811 10362
rect 8991 10310 8993 10362
rect 8747 10308 8753 10310
rect 8809 10308 8833 10310
rect 8889 10308 8913 10310
rect 8969 10308 8993 10310
rect 9049 10308 9055 10310
rect 8747 10299 9055 10308
rect 8747 9276 9055 9285
rect 8747 9274 8753 9276
rect 8809 9274 8833 9276
rect 8889 9274 8913 9276
rect 8969 9274 8993 9276
rect 9049 9274 9055 9276
rect 8809 9222 8811 9274
rect 8991 9222 8993 9274
rect 8747 9220 8753 9222
rect 8809 9220 8833 9222
rect 8889 9220 8913 9222
rect 8969 9220 8993 9222
rect 9049 9220 9055 9222
rect 8747 9211 9055 9220
rect 8760 9104 8812 9110
rect 8760 9046 8812 9052
rect 8772 8498 8800 9046
rect 8852 8900 8904 8906
rect 8852 8842 8904 8848
rect 8864 8498 8892 8842
rect 9128 8832 9180 8838
rect 9128 8774 9180 8780
rect 8760 8492 8812 8498
rect 8760 8434 8812 8440
rect 8852 8492 8904 8498
rect 8852 8434 8904 8440
rect 8772 8378 8800 8434
rect 8680 8350 8800 8378
rect 8484 8288 8536 8294
rect 8484 8230 8536 8236
rect 7380 8016 7432 8022
rect 7380 7958 7432 7964
rect 7392 7342 7420 7958
rect 8392 7812 8444 7818
rect 8392 7754 8444 7760
rect 8208 7540 8260 7546
rect 8208 7482 8260 7488
rect 7380 7336 7432 7342
rect 7380 7278 7432 7284
rect 8220 7206 8248 7482
rect 8404 7478 8432 7754
rect 8392 7472 8444 7478
rect 8392 7414 8444 7420
rect 8208 7200 8260 7206
rect 8208 7142 8260 7148
rect 7102 6896 7158 6905
rect 7102 6831 7158 6840
rect 8220 6186 8248 7142
rect 8404 6866 8432 7414
rect 8496 7342 8524 8230
rect 8680 7886 8708 8350
rect 8747 8188 9055 8197
rect 8747 8186 8753 8188
rect 8809 8186 8833 8188
rect 8889 8186 8913 8188
rect 8969 8186 8993 8188
rect 9049 8186 9055 8188
rect 8809 8134 8811 8186
rect 8991 8134 8993 8186
rect 8747 8132 8753 8134
rect 8809 8132 8833 8134
rect 8889 8132 8913 8134
rect 8969 8132 8993 8134
rect 9049 8132 9055 8134
rect 8747 8123 9055 8132
rect 8668 7880 8720 7886
rect 8668 7822 8720 7828
rect 9140 7478 9168 8774
rect 9416 7954 9444 11018
rect 9496 9444 9548 9450
rect 9496 9386 9548 9392
rect 9508 9110 9536 9386
rect 9588 9376 9640 9382
rect 9588 9318 9640 9324
rect 9496 9104 9548 9110
rect 9496 9046 9548 9052
rect 9600 8906 9628 9318
rect 9588 8900 9640 8906
rect 9588 8842 9640 8848
rect 9692 8022 9720 11698
rect 9876 10169 9904 15302
rect 9968 12238 9996 20198
rect 10152 19990 10180 22200
rect 10520 20602 10548 22200
rect 10508 20596 10560 20602
rect 10508 20538 10560 20544
rect 10232 20392 10284 20398
rect 10232 20334 10284 20340
rect 10416 20392 10468 20398
rect 10416 20334 10468 20340
rect 10140 19984 10192 19990
rect 10140 19926 10192 19932
rect 10244 19922 10272 20334
rect 10428 20058 10456 20334
rect 10416 20052 10468 20058
rect 10416 19994 10468 20000
rect 10520 19938 10548 20538
rect 10784 20324 10836 20330
rect 10888 20312 10916 22200
rect 11256 20466 11284 22200
rect 11624 20890 11652 22200
rect 11624 20862 11744 20890
rect 11346 20700 11654 20709
rect 11346 20698 11352 20700
rect 11408 20698 11432 20700
rect 11488 20698 11512 20700
rect 11568 20698 11592 20700
rect 11648 20698 11654 20700
rect 11408 20646 11410 20698
rect 11590 20646 11592 20698
rect 11346 20644 11352 20646
rect 11408 20644 11432 20646
rect 11488 20644 11512 20646
rect 11568 20644 11592 20646
rect 11648 20644 11654 20646
rect 11346 20635 11654 20644
rect 11060 20460 11112 20466
rect 11060 20402 11112 20408
rect 11244 20460 11296 20466
rect 11244 20402 11296 20408
rect 10836 20284 10916 20312
rect 10784 20266 10836 20272
rect 10600 20052 10652 20058
rect 10600 19994 10652 20000
rect 10048 19916 10100 19922
rect 10048 19858 10100 19864
rect 10232 19916 10284 19922
rect 10232 19858 10284 19864
rect 10428 19910 10548 19938
rect 10060 19378 10088 19858
rect 10324 19848 10376 19854
rect 10324 19790 10376 19796
rect 10048 19372 10100 19378
rect 10048 19314 10100 19320
rect 10046 18864 10102 18873
rect 10046 18799 10102 18808
rect 10060 18601 10088 18799
rect 10046 18592 10102 18601
rect 10046 18527 10102 18536
rect 10232 18352 10284 18358
rect 10232 18294 10284 18300
rect 10138 17776 10194 17785
rect 10048 17740 10100 17746
rect 10138 17711 10194 17720
rect 10048 17682 10100 17688
rect 10060 17066 10088 17682
rect 10152 17542 10180 17711
rect 10140 17536 10192 17542
rect 10140 17478 10192 17484
rect 10244 17134 10272 18294
rect 10336 17626 10364 19790
rect 10428 17882 10456 19910
rect 10612 18358 10640 19994
rect 10876 19984 10928 19990
rect 10876 19926 10928 19932
rect 10784 19916 10836 19922
rect 10784 19858 10836 19864
rect 10796 19009 10824 19858
rect 10782 19000 10838 19009
rect 10782 18935 10838 18944
rect 10600 18352 10652 18358
rect 10600 18294 10652 18300
rect 10888 18290 10916 19926
rect 10968 19236 11020 19242
rect 10968 19178 11020 19184
rect 10980 18970 11008 19178
rect 10968 18964 11020 18970
rect 10968 18906 11020 18912
rect 10876 18284 10928 18290
rect 10876 18226 10928 18232
rect 10692 18216 10744 18222
rect 10692 18158 10744 18164
rect 10508 18080 10560 18086
rect 10508 18022 10560 18028
rect 10416 17876 10468 17882
rect 10416 17818 10468 17824
rect 10520 17814 10548 18022
rect 10508 17808 10560 17814
rect 10508 17750 10560 17756
rect 10336 17598 10456 17626
rect 10232 17128 10284 17134
rect 10232 17070 10284 17076
rect 10048 17060 10100 17066
rect 10048 17002 10100 17008
rect 10140 16992 10192 16998
rect 10140 16934 10192 16940
rect 10152 16590 10180 16934
rect 10140 16584 10192 16590
rect 10140 16526 10192 16532
rect 10152 16114 10180 16526
rect 10048 16108 10100 16114
rect 10048 16050 10100 16056
rect 10140 16108 10192 16114
rect 10140 16050 10192 16056
rect 10060 15706 10088 16050
rect 10048 15700 10100 15706
rect 10048 15642 10100 15648
rect 10152 15586 10180 16050
rect 10152 15570 10272 15586
rect 10152 15564 10284 15570
rect 10152 15558 10232 15564
rect 10232 15506 10284 15512
rect 10140 15496 10192 15502
rect 10140 15438 10192 15444
rect 10048 14340 10100 14346
rect 10048 14282 10100 14288
rect 9956 12232 10008 12238
rect 9956 12174 10008 12180
rect 9862 10160 9918 10169
rect 9862 10095 9918 10104
rect 9772 9920 9824 9926
rect 9772 9862 9824 9868
rect 9956 9920 10008 9926
rect 9956 9862 10008 9868
rect 9784 9518 9812 9862
rect 9968 9761 9996 9862
rect 9954 9752 10010 9761
rect 9954 9687 10010 9696
rect 9772 9512 9824 9518
rect 9772 9454 9824 9460
rect 10060 8242 10088 14282
rect 10152 12986 10180 15438
rect 10324 15020 10376 15026
rect 10324 14962 10376 14968
rect 10336 13734 10364 14962
rect 10324 13728 10376 13734
rect 10324 13670 10376 13676
rect 10336 13462 10364 13670
rect 10324 13456 10376 13462
rect 10324 13398 10376 13404
rect 10140 12980 10192 12986
rect 10140 12922 10192 12928
rect 10140 12776 10192 12782
rect 10140 12718 10192 12724
rect 10152 10810 10180 12718
rect 10324 12436 10376 12442
rect 10324 12378 10376 12384
rect 10336 12306 10364 12378
rect 10324 12300 10376 12306
rect 10324 12242 10376 12248
rect 10428 11558 10456 17598
rect 10520 12434 10548 17750
rect 10600 17536 10652 17542
rect 10598 17504 10600 17513
rect 10652 17504 10654 17513
rect 10598 17439 10654 17448
rect 10704 17338 10732 18158
rect 10968 17536 11020 17542
rect 10968 17478 11020 17484
rect 10692 17332 10744 17338
rect 10692 17274 10744 17280
rect 10600 17128 10652 17134
rect 10598 17096 10600 17105
rect 10652 17096 10654 17105
rect 10598 17031 10654 17040
rect 10876 16584 10928 16590
rect 10876 16526 10928 16532
rect 10784 16516 10836 16522
rect 10784 16458 10836 16464
rect 10692 16040 10744 16046
rect 10692 15982 10744 15988
rect 10598 15600 10654 15609
rect 10598 15535 10654 15544
rect 10612 15366 10640 15535
rect 10600 15360 10652 15366
rect 10600 15302 10652 15308
rect 10704 14346 10732 15982
rect 10796 15910 10824 16458
rect 10784 15904 10836 15910
rect 10784 15846 10836 15852
rect 10888 15706 10916 16526
rect 10980 16266 11008 17478
rect 11072 16454 11100 20402
rect 11256 19334 11284 20402
rect 11346 19612 11654 19621
rect 11346 19610 11352 19612
rect 11408 19610 11432 19612
rect 11488 19610 11512 19612
rect 11568 19610 11592 19612
rect 11648 19610 11654 19612
rect 11408 19558 11410 19610
rect 11590 19558 11592 19610
rect 11346 19556 11352 19558
rect 11408 19556 11432 19558
rect 11488 19556 11512 19558
rect 11568 19556 11592 19558
rect 11648 19556 11654 19558
rect 11346 19547 11654 19556
rect 11256 19306 11468 19334
rect 11716 19310 11744 20862
rect 11992 20466 12020 22200
rect 11980 20460 12032 20466
rect 11980 20402 12032 20408
rect 12256 20460 12308 20466
rect 12256 20402 12308 20408
rect 12164 20256 12216 20262
rect 12164 20198 12216 20204
rect 12072 19916 12124 19922
rect 12072 19858 12124 19864
rect 11888 19848 11940 19854
rect 11888 19790 11940 19796
rect 11796 19780 11848 19786
rect 11796 19722 11848 19728
rect 11152 19168 11204 19174
rect 11152 19110 11204 19116
rect 11164 17882 11192 19110
rect 11334 19000 11390 19009
rect 11440 18970 11468 19306
rect 11704 19304 11756 19310
rect 11704 19246 11756 19252
rect 11808 19174 11836 19722
rect 11900 19446 11928 19790
rect 11888 19440 11940 19446
rect 11888 19382 11940 19388
rect 11978 19408 12034 19417
rect 11796 19168 11848 19174
rect 11796 19110 11848 19116
rect 11334 18935 11390 18944
rect 11428 18964 11480 18970
rect 11348 18902 11376 18935
rect 11428 18906 11480 18912
rect 11336 18896 11388 18902
rect 11336 18838 11388 18844
rect 11348 18698 11376 18838
rect 11336 18692 11388 18698
rect 11336 18634 11388 18640
rect 11346 18524 11654 18533
rect 11346 18522 11352 18524
rect 11408 18522 11432 18524
rect 11488 18522 11512 18524
rect 11568 18522 11592 18524
rect 11648 18522 11654 18524
rect 11408 18470 11410 18522
rect 11590 18470 11592 18522
rect 11346 18468 11352 18470
rect 11408 18468 11432 18470
rect 11488 18468 11512 18470
rect 11568 18468 11592 18470
rect 11648 18468 11654 18470
rect 11346 18459 11654 18468
rect 11808 18222 11836 19110
rect 11900 18766 11928 19382
rect 12084 19378 12112 19858
rect 11978 19343 11980 19352
rect 12032 19343 12034 19352
rect 12072 19372 12124 19378
rect 11980 19314 12032 19320
rect 12072 19314 12124 19320
rect 11888 18760 11940 18766
rect 11888 18702 11940 18708
rect 12176 18714 12204 20198
rect 12268 19310 12296 20402
rect 12360 20244 12388 22200
rect 12728 20448 12756 22200
rect 13096 20534 13124 22200
rect 13464 22114 13492 22200
rect 13556 22114 13584 22222
rect 13464 22086 13584 22114
rect 13084 20528 13136 20534
rect 13084 20470 13136 20476
rect 12808 20460 12860 20466
rect 12728 20420 12808 20448
rect 12808 20402 12860 20408
rect 13636 20460 13688 20466
rect 13636 20402 13688 20408
rect 12532 20392 12584 20398
rect 12532 20334 12584 20340
rect 12360 20216 12480 20244
rect 12452 19854 12480 20216
rect 12440 19848 12492 19854
rect 12440 19790 12492 19796
rect 12348 19780 12400 19786
rect 12348 19722 12400 19728
rect 12360 19514 12388 19722
rect 12348 19508 12400 19514
rect 12348 19450 12400 19456
rect 12256 19304 12308 19310
rect 12256 19246 12308 19252
rect 12440 18760 12492 18766
rect 11900 18358 11928 18702
rect 12176 18686 12388 18714
rect 12440 18702 12492 18708
rect 11888 18352 11940 18358
rect 11888 18294 11940 18300
rect 11796 18216 11848 18222
rect 11796 18158 11848 18164
rect 11152 17876 11204 17882
rect 11152 17818 11204 17824
rect 11520 17808 11572 17814
rect 11520 17750 11572 17756
rect 11244 17740 11296 17746
rect 11244 17682 11296 17688
rect 11152 16992 11204 16998
rect 11152 16934 11204 16940
rect 11060 16448 11112 16454
rect 11060 16390 11112 16396
rect 10980 16238 11100 16266
rect 11164 16250 11192 16934
rect 11256 16590 11284 17682
rect 11532 17542 11560 17750
rect 11704 17740 11756 17746
rect 11704 17682 11756 17688
rect 11520 17536 11572 17542
rect 11520 17478 11572 17484
rect 11346 17436 11654 17445
rect 11346 17434 11352 17436
rect 11408 17434 11432 17436
rect 11488 17434 11512 17436
rect 11568 17434 11592 17436
rect 11648 17434 11654 17436
rect 11408 17382 11410 17434
rect 11590 17382 11592 17434
rect 11346 17380 11352 17382
rect 11408 17380 11432 17382
rect 11488 17380 11512 17382
rect 11568 17380 11592 17382
rect 11648 17380 11654 17382
rect 11346 17371 11654 17380
rect 11612 17264 11664 17270
rect 11610 17232 11612 17241
rect 11664 17232 11666 17241
rect 11610 17167 11666 17176
rect 11244 16584 11296 16590
rect 11244 16526 11296 16532
rect 11244 16448 11296 16454
rect 11244 16390 11296 16396
rect 11072 15706 11100 16238
rect 11152 16244 11204 16250
rect 11152 16186 11204 16192
rect 11256 16182 11284 16390
rect 11346 16348 11654 16357
rect 11346 16346 11352 16348
rect 11408 16346 11432 16348
rect 11488 16346 11512 16348
rect 11568 16346 11592 16348
rect 11648 16346 11654 16348
rect 11408 16294 11410 16346
rect 11590 16294 11592 16346
rect 11346 16292 11352 16294
rect 11408 16292 11432 16294
rect 11488 16292 11512 16294
rect 11568 16292 11592 16294
rect 11648 16292 11654 16294
rect 11346 16283 11654 16292
rect 11336 16244 11388 16250
rect 11336 16186 11388 16192
rect 11520 16244 11572 16250
rect 11520 16186 11572 16192
rect 11244 16176 11296 16182
rect 11244 16118 11296 16124
rect 10876 15700 10928 15706
rect 10876 15642 10928 15648
rect 11060 15700 11112 15706
rect 11060 15642 11112 15648
rect 11348 15570 11376 16186
rect 11532 15638 11560 16186
rect 11612 15904 11664 15910
rect 11612 15846 11664 15852
rect 11520 15632 11572 15638
rect 11520 15574 11572 15580
rect 11336 15564 11388 15570
rect 11336 15506 11388 15512
rect 11060 15496 11112 15502
rect 11060 15438 11112 15444
rect 11072 14618 11100 15438
rect 11624 15366 11652 15846
rect 11612 15360 11664 15366
rect 11612 15302 11664 15308
rect 11346 15260 11654 15269
rect 11346 15258 11352 15260
rect 11408 15258 11432 15260
rect 11488 15258 11512 15260
rect 11568 15258 11592 15260
rect 11648 15258 11654 15260
rect 11408 15206 11410 15258
rect 11590 15206 11592 15258
rect 11346 15204 11352 15206
rect 11408 15204 11432 15206
rect 11488 15204 11512 15206
rect 11568 15204 11592 15206
rect 11648 15204 11654 15206
rect 11346 15195 11654 15204
rect 11336 15156 11388 15162
rect 11336 15098 11388 15104
rect 11348 14618 11376 15098
rect 11716 14890 11744 17682
rect 11796 17536 11848 17542
rect 11794 17504 11796 17513
rect 11848 17504 11850 17513
rect 11794 17439 11850 17448
rect 11900 17338 11928 18294
rect 12072 17876 12124 17882
rect 12360 17864 12388 18686
rect 12452 18222 12480 18702
rect 12440 18216 12492 18222
rect 12440 18158 12492 18164
rect 12072 17818 12124 17824
rect 12268 17836 12388 17864
rect 11980 17604 12032 17610
rect 11980 17546 12032 17552
rect 11888 17332 11940 17338
rect 11888 17274 11940 17280
rect 11796 17196 11848 17202
rect 11796 17138 11848 17144
rect 11808 16590 11836 17138
rect 11900 16794 11928 17274
rect 11992 17202 12020 17546
rect 12084 17542 12112 17818
rect 12164 17740 12216 17746
rect 12164 17682 12216 17688
rect 12176 17649 12204 17682
rect 12162 17640 12218 17649
rect 12162 17575 12218 17584
rect 12072 17536 12124 17542
rect 12072 17478 12124 17484
rect 12084 17270 12112 17478
rect 12072 17264 12124 17270
rect 12072 17206 12124 17212
rect 11980 17196 12032 17202
rect 11980 17138 12032 17144
rect 12164 17128 12216 17134
rect 12164 17070 12216 17076
rect 12268 17082 12296 17836
rect 12452 17202 12480 18158
rect 12440 17196 12492 17202
rect 12440 17138 12492 17144
rect 11888 16788 11940 16794
rect 11888 16730 11940 16736
rect 11886 16688 11942 16697
rect 11886 16623 11942 16632
rect 11796 16584 11848 16590
rect 11796 16526 11848 16532
rect 11900 16402 11928 16623
rect 11808 16374 11928 16402
rect 11704 14884 11756 14890
rect 11704 14826 11756 14832
rect 11520 14816 11572 14822
rect 11520 14758 11572 14764
rect 11060 14612 11112 14618
rect 11060 14554 11112 14560
rect 11336 14612 11388 14618
rect 11336 14554 11388 14560
rect 10692 14340 10744 14346
rect 10692 14282 10744 14288
rect 11072 14006 11100 14554
rect 11532 14346 11560 14758
rect 11520 14340 11572 14346
rect 11520 14282 11572 14288
rect 11346 14172 11654 14181
rect 11346 14170 11352 14172
rect 11408 14170 11432 14172
rect 11488 14170 11512 14172
rect 11568 14170 11592 14172
rect 11648 14170 11654 14172
rect 11408 14118 11410 14170
rect 11590 14118 11592 14170
rect 11346 14116 11352 14118
rect 11408 14116 11432 14118
rect 11488 14116 11512 14118
rect 11568 14116 11592 14118
rect 11648 14116 11654 14118
rect 11346 14107 11654 14116
rect 11060 14000 11112 14006
rect 11060 13942 11112 13948
rect 11704 13728 11756 13734
rect 11704 13670 11756 13676
rect 11716 13258 11744 13670
rect 11704 13252 11756 13258
rect 11704 13194 11756 13200
rect 11244 13184 11296 13190
rect 11244 13126 11296 13132
rect 11256 12986 11284 13126
rect 11346 13084 11654 13093
rect 11346 13082 11352 13084
rect 11408 13082 11432 13084
rect 11488 13082 11512 13084
rect 11568 13082 11592 13084
rect 11648 13082 11654 13084
rect 11408 13030 11410 13082
rect 11590 13030 11592 13082
rect 11346 13028 11352 13030
rect 11408 13028 11432 13030
rect 11488 13028 11512 13030
rect 11568 13028 11592 13030
rect 11648 13028 11654 13030
rect 11346 13019 11654 13028
rect 11244 12980 11296 12986
rect 11244 12922 11296 12928
rect 11716 12782 11744 13194
rect 11704 12776 11756 12782
rect 11704 12718 11756 12724
rect 10968 12640 11020 12646
rect 10968 12582 11020 12588
rect 10520 12406 10732 12434
rect 10508 12300 10560 12306
rect 10508 12242 10560 12248
rect 10520 11830 10548 12242
rect 10600 12096 10652 12102
rect 10600 12038 10652 12044
rect 10612 11830 10640 12038
rect 10508 11824 10560 11830
rect 10508 11766 10560 11772
rect 10600 11824 10652 11830
rect 10600 11766 10652 11772
rect 10416 11552 10468 11558
rect 10416 11494 10468 11500
rect 10428 10810 10456 11494
rect 10140 10804 10192 10810
rect 10140 10746 10192 10752
rect 10416 10804 10468 10810
rect 10416 10746 10468 10752
rect 10152 9654 10180 10746
rect 10230 10704 10286 10713
rect 10230 10639 10286 10648
rect 10244 10266 10272 10639
rect 10232 10260 10284 10266
rect 10232 10202 10284 10208
rect 10140 9648 10192 9654
rect 10140 9590 10192 9596
rect 10508 9376 10560 9382
rect 10508 9318 10560 9324
rect 10520 8974 10548 9318
rect 10704 8974 10732 12406
rect 10784 12232 10836 12238
rect 10784 12174 10836 12180
rect 10796 11694 10824 12174
rect 10876 12096 10928 12102
rect 10876 12038 10928 12044
rect 10888 11898 10916 12038
rect 10876 11892 10928 11898
rect 10876 11834 10928 11840
rect 10784 11688 10836 11694
rect 10784 11630 10836 11636
rect 10784 11144 10836 11150
rect 10784 11086 10836 11092
rect 10796 10674 10824 11086
rect 10784 10668 10836 10674
rect 10784 10610 10836 10616
rect 10980 9081 11008 12582
rect 11704 12164 11756 12170
rect 11704 12106 11756 12112
rect 11060 12096 11112 12102
rect 11060 12038 11112 12044
rect 10966 9072 11022 9081
rect 10966 9007 11022 9016
rect 10508 8968 10560 8974
rect 10508 8910 10560 8916
rect 10692 8968 10744 8974
rect 10692 8910 10744 8916
rect 10140 8900 10192 8906
rect 10140 8842 10192 8848
rect 10152 8362 10180 8842
rect 10520 8362 10548 8910
rect 11072 8634 11100 12038
rect 11346 11996 11654 12005
rect 11346 11994 11352 11996
rect 11408 11994 11432 11996
rect 11488 11994 11512 11996
rect 11568 11994 11592 11996
rect 11648 11994 11654 11996
rect 11408 11942 11410 11994
rect 11590 11942 11592 11994
rect 11346 11940 11352 11942
rect 11408 11940 11432 11942
rect 11488 11940 11512 11942
rect 11568 11940 11592 11942
rect 11648 11940 11654 11942
rect 11346 11931 11654 11940
rect 11150 11792 11206 11801
rect 11150 11727 11206 11736
rect 11060 8628 11112 8634
rect 11060 8570 11112 8576
rect 11164 8566 11192 11727
rect 11612 11552 11664 11558
rect 11612 11494 11664 11500
rect 11624 11354 11652 11494
rect 11612 11348 11664 11354
rect 11612 11290 11664 11296
rect 11716 11150 11744 12106
rect 11704 11144 11756 11150
rect 11704 11086 11756 11092
rect 11346 10908 11654 10917
rect 11346 10906 11352 10908
rect 11408 10906 11432 10908
rect 11488 10906 11512 10908
rect 11568 10906 11592 10908
rect 11648 10906 11654 10908
rect 11408 10854 11410 10906
rect 11590 10854 11592 10906
rect 11346 10852 11352 10854
rect 11408 10852 11432 10854
rect 11488 10852 11512 10854
rect 11568 10852 11592 10854
rect 11648 10852 11654 10854
rect 11346 10843 11654 10852
rect 11346 9820 11654 9829
rect 11346 9818 11352 9820
rect 11408 9818 11432 9820
rect 11488 9818 11512 9820
rect 11568 9818 11592 9820
rect 11648 9818 11654 9820
rect 11408 9766 11410 9818
rect 11590 9766 11592 9818
rect 11346 9764 11352 9766
rect 11408 9764 11432 9766
rect 11488 9764 11512 9766
rect 11568 9764 11592 9766
rect 11648 9764 11654 9766
rect 11346 9755 11654 9764
rect 11716 9382 11744 11086
rect 11704 9376 11756 9382
rect 11704 9318 11756 9324
rect 11346 8732 11654 8741
rect 11346 8730 11352 8732
rect 11408 8730 11432 8732
rect 11488 8730 11512 8732
rect 11568 8730 11592 8732
rect 11648 8730 11654 8732
rect 11408 8678 11410 8730
rect 11590 8678 11592 8730
rect 11346 8676 11352 8678
rect 11408 8676 11432 8678
rect 11488 8676 11512 8678
rect 11568 8676 11592 8678
rect 11648 8676 11654 8678
rect 11346 8667 11654 8676
rect 11428 8628 11480 8634
rect 11428 8570 11480 8576
rect 11152 8560 11204 8566
rect 11152 8502 11204 8508
rect 10968 8492 11020 8498
rect 10968 8434 11020 8440
rect 10140 8356 10192 8362
rect 10140 8298 10192 8304
rect 10508 8356 10560 8362
rect 10508 8298 10560 8304
rect 10876 8288 10928 8294
rect 10060 8214 10548 8242
rect 10876 8230 10928 8236
rect 10520 8090 10548 8214
rect 10508 8084 10560 8090
rect 10508 8026 10560 8032
rect 9680 8016 9732 8022
rect 9680 7958 9732 7964
rect 9404 7948 9456 7954
rect 9404 7890 9456 7896
rect 9680 7880 9732 7886
rect 9680 7822 9732 7828
rect 9404 7744 9456 7750
rect 9404 7686 9456 7692
rect 9416 7546 9444 7686
rect 9404 7540 9456 7546
rect 9404 7482 9456 7488
rect 9128 7472 9180 7478
rect 9128 7414 9180 7420
rect 8484 7336 8536 7342
rect 8484 7278 8536 7284
rect 8496 6866 8524 7278
rect 8852 7268 8904 7274
rect 9036 7268 9088 7274
rect 8904 7228 9036 7256
rect 8852 7210 8904 7216
rect 9036 7210 9088 7216
rect 8747 7100 9055 7109
rect 8747 7098 8753 7100
rect 8809 7098 8833 7100
rect 8889 7098 8913 7100
rect 8969 7098 8993 7100
rect 9049 7098 9055 7100
rect 8809 7046 8811 7098
rect 8991 7046 8993 7098
rect 8747 7044 8753 7046
rect 8809 7044 8833 7046
rect 8889 7044 8913 7046
rect 8969 7044 8993 7046
rect 9049 7044 9055 7046
rect 8747 7035 9055 7044
rect 9692 7002 9720 7822
rect 9864 7404 9916 7410
rect 9864 7346 9916 7352
rect 9772 7200 9824 7206
rect 9772 7142 9824 7148
rect 9784 7002 9812 7142
rect 9680 6996 9732 7002
rect 9680 6938 9732 6944
rect 9772 6996 9824 7002
rect 9772 6938 9824 6944
rect 9876 6866 9904 7346
rect 8392 6860 8444 6866
rect 8392 6802 8444 6808
rect 8484 6860 8536 6866
rect 8484 6802 8536 6808
rect 9864 6860 9916 6866
rect 9864 6802 9916 6808
rect 9220 6656 9272 6662
rect 9220 6598 9272 6604
rect 9312 6656 9364 6662
rect 9312 6598 9364 6604
rect 9232 6390 9260 6598
rect 9220 6384 9272 6390
rect 9220 6326 9272 6332
rect 8208 6180 8260 6186
rect 8208 6122 8260 6128
rect 8747 6012 9055 6021
rect 8747 6010 8753 6012
rect 8809 6010 8833 6012
rect 8889 6010 8913 6012
rect 8969 6010 8993 6012
rect 9049 6010 9055 6012
rect 8809 5958 8811 6010
rect 8991 5958 8993 6010
rect 8747 5956 8753 5958
rect 8809 5956 8833 5958
rect 8889 5956 8913 5958
rect 8969 5956 8993 5958
rect 9049 5956 9055 5958
rect 8747 5947 9055 5956
rect 9324 5817 9352 6598
rect 10520 6322 10548 8026
rect 10598 7984 10654 7993
rect 10598 7919 10654 7928
rect 10612 7886 10640 7919
rect 10600 7880 10652 7886
rect 10600 7822 10652 7828
rect 10612 7478 10640 7822
rect 10600 7472 10652 7478
rect 10600 7414 10652 7420
rect 10888 7342 10916 8230
rect 10876 7336 10928 7342
rect 10876 7278 10928 7284
rect 10508 6316 10560 6322
rect 10508 6258 10560 6264
rect 9310 5808 9366 5817
rect 9310 5743 9366 5752
rect 10980 5642 11008 8434
rect 11440 7954 11468 8570
rect 11428 7948 11480 7954
rect 11428 7890 11480 7896
rect 11808 7886 11836 16374
rect 12072 16108 12124 16114
rect 12072 16050 12124 16056
rect 11980 16040 12032 16046
rect 12084 16017 12112 16050
rect 11980 15982 12032 15988
rect 12070 16008 12126 16017
rect 11992 15706 12020 15982
rect 12070 15943 12126 15952
rect 12084 15910 12112 15943
rect 12072 15904 12124 15910
rect 12072 15846 12124 15852
rect 11980 15700 12032 15706
rect 11980 15642 12032 15648
rect 12176 15570 12204 17070
rect 12268 17054 12388 17082
rect 12360 16697 12388 17054
rect 12346 16688 12402 16697
rect 12346 16623 12402 16632
rect 12348 16516 12400 16522
rect 12348 16458 12400 16464
rect 12164 15564 12216 15570
rect 12164 15506 12216 15512
rect 12360 15502 12388 16458
rect 12348 15496 12400 15502
rect 12348 15438 12400 15444
rect 12072 15428 12124 15434
rect 12072 15370 12124 15376
rect 11888 15360 11940 15366
rect 11888 15302 11940 15308
rect 11900 12986 11928 15302
rect 11888 12980 11940 12986
rect 11888 12922 11940 12928
rect 11888 12776 11940 12782
rect 11888 12718 11940 12724
rect 11900 11694 11928 12718
rect 11888 11688 11940 11694
rect 11888 11630 11940 11636
rect 11980 9988 12032 9994
rect 11980 9930 12032 9936
rect 11992 9110 12020 9930
rect 11980 9104 12032 9110
rect 11980 9046 12032 9052
rect 11980 8288 12032 8294
rect 11980 8230 12032 8236
rect 11992 7886 12020 8230
rect 11060 7880 11112 7886
rect 11060 7822 11112 7828
rect 11796 7880 11848 7886
rect 11796 7822 11848 7828
rect 11980 7880 12032 7886
rect 11980 7822 12032 7828
rect 11072 7546 11100 7822
rect 11346 7644 11654 7653
rect 11346 7642 11352 7644
rect 11408 7642 11432 7644
rect 11488 7642 11512 7644
rect 11568 7642 11592 7644
rect 11648 7642 11654 7644
rect 11408 7590 11410 7642
rect 11590 7590 11592 7642
rect 11346 7588 11352 7590
rect 11408 7588 11432 7590
rect 11488 7588 11512 7590
rect 11568 7588 11592 7590
rect 11648 7588 11654 7590
rect 11346 7579 11654 7588
rect 11992 7546 12020 7822
rect 11060 7540 11112 7546
rect 11060 7482 11112 7488
rect 11980 7540 12032 7546
rect 11980 7482 12032 7488
rect 11346 6556 11654 6565
rect 11346 6554 11352 6556
rect 11408 6554 11432 6556
rect 11488 6554 11512 6556
rect 11568 6554 11592 6556
rect 11648 6554 11654 6556
rect 11408 6502 11410 6554
rect 11590 6502 11592 6554
rect 11346 6500 11352 6502
rect 11408 6500 11432 6502
rect 11488 6500 11512 6502
rect 11568 6500 11592 6502
rect 11648 6500 11654 6502
rect 11346 6491 11654 6500
rect 11980 6452 12032 6458
rect 12084 6440 12112 15370
rect 12440 13728 12492 13734
rect 12440 13670 12492 13676
rect 12348 13252 12400 13258
rect 12348 13194 12400 13200
rect 12256 13184 12308 13190
rect 12256 13126 12308 13132
rect 12268 12986 12296 13126
rect 12256 12980 12308 12986
rect 12256 12922 12308 12928
rect 12164 12844 12216 12850
rect 12164 12786 12216 12792
rect 12176 12646 12204 12786
rect 12164 12640 12216 12646
rect 12164 12582 12216 12588
rect 12360 12306 12388 13194
rect 12452 12918 12480 13670
rect 12440 12912 12492 12918
rect 12440 12854 12492 12860
rect 12544 12424 12572 20334
rect 12624 19848 12676 19854
rect 12624 19790 12676 19796
rect 12716 19848 12768 19854
rect 12716 19790 12768 19796
rect 12636 19514 12664 19790
rect 12624 19508 12676 19514
rect 12624 19450 12676 19456
rect 12624 17876 12676 17882
rect 12624 17818 12676 17824
rect 12636 17610 12664 17818
rect 12624 17604 12676 17610
rect 12624 17546 12676 17552
rect 12728 16250 12756 19790
rect 12820 19514 12848 20402
rect 12992 20392 13044 20398
rect 12992 20334 13044 20340
rect 12808 19508 12860 19514
rect 12808 19450 12860 19456
rect 12808 18080 12860 18086
rect 12808 18022 12860 18028
rect 12716 16244 12768 16250
rect 12716 16186 12768 16192
rect 12820 15026 12848 18022
rect 12900 15904 12952 15910
rect 12900 15846 12952 15852
rect 12808 15020 12860 15026
rect 12808 14962 12860 14968
rect 12806 14920 12862 14929
rect 12806 14855 12862 14864
rect 12820 13841 12848 14855
rect 12806 13832 12862 13841
rect 12806 13767 12862 13776
rect 12716 13320 12768 13326
rect 12716 13262 12768 13268
rect 12624 12980 12676 12986
rect 12624 12922 12676 12928
rect 12636 12714 12664 12922
rect 12728 12850 12756 13262
rect 12820 12889 12848 13767
rect 12806 12880 12862 12889
rect 12716 12844 12768 12850
rect 12806 12815 12862 12824
rect 12716 12786 12768 12792
rect 12624 12708 12676 12714
rect 12624 12650 12676 12656
rect 12912 12646 12940 15846
rect 13004 14929 13032 20334
rect 13360 19916 13412 19922
rect 13360 19858 13412 19864
rect 13176 19712 13228 19718
rect 13176 19654 13228 19660
rect 13188 18290 13216 19654
rect 13372 19514 13400 19858
rect 13452 19848 13504 19854
rect 13452 19790 13504 19796
rect 13544 19848 13596 19854
rect 13544 19790 13596 19796
rect 13360 19508 13412 19514
rect 13360 19450 13412 19456
rect 13464 18970 13492 19790
rect 13452 18964 13504 18970
rect 13452 18906 13504 18912
rect 13268 18760 13320 18766
rect 13268 18702 13320 18708
rect 13176 18284 13228 18290
rect 13176 18226 13228 18232
rect 13082 17640 13138 17649
rect 13082 17575 13138 17584
rect 13096 17202 13124 17575
rect 13176 17536 13228 17542
rect 13174 17504 13176 17513
rect 13228 17504 13230 17513
rect 13174 17439 13230 17448
rect 13084 17196 13136 17202
rect 13084 17138 13136 17144
rect 13096 16561 13124 17138
rect 13082 16552 13138 16561
rect 13082 16487 13138 16496
rect 13084 15564 13136 15570
rect 13084 15506 13136 15512
rect 12990 14920 13046 14929
rect 12990 14855 13046 14864
rect 12992 14816 13044 14822
rect 12992 14758 13044 14764
rect 13004 12850 13032 14758
rect 12992 12844 13044 12850
rect 12992 12786 13044 12792
rect 12900 12640 12952 12646
rect 12900 12582 12952 12588
rect 12452 12396 12572 12424
rect 12348 12300 12400 12306
rect 12348 12242 12400 12248
rect 12164 12096 12216 12102
rect 12164 12038 12216 12044
rect 12256 12096 12308 12102
rect 12256 12038 12308 12044
rect 12176 11830 12204 12038
rect 12164 11824 12216 11830
rect 12268 11801 12296 12038
rect 12164 11766 12216 11772
rect 12254 11792 12310 11801
rect 12254 11727 12310 11736
rect 12452 11257 12480 12396
rect 12808 12368 12860 12374
rect 12544 12316 12808 12322
rect 12544 12310 12860 12316
rect 12544 12294 12848 12310
rect 12544 12170 12572 12294
rect 12532 12164 12584 12170
rect 12532 12106 12584 12112
rect 12438 11248 12494 11257
rect 12256 11212 12308 11218
rect 12438 11183 12494 11192
rect 12256 11154 12308 11160
rect 12268 10810 12296 11154
rect 12256 10804 12308 10810
rect 12256 10746 12308 10752
rect 12164 10736 12216 10742
rect 12164 10678 12216 10684
rect 12176 9994 12204 10678
rect 12268 10062 12296 10746
rect 12912 10577 12940 12582
rect 13004 12442 13032 12786
rect 12992 12436 13044 12442
rect 12992 12378 13044 12384
rect 12992 11552 13044 11558
rect 13096 11540 13124 15506
rect 13176 13796 13228 13802
rect 13176 13738 13228 13744
rect 13188 13530 13216 13738
rect 13176 13524 13228 13530
rect 13176 13466 13228 13472
rect 13176 13184 13228 13190
rect 13176 13126 13228 13132
rect 13188 12442 13216 13126
rect 13176 12436 13228 12442
rect 13176 12378 13228 12384
rect 13280 11762 13308 18702
rect 13452 18624 13504 18630
rect 13452 18566 13504 18572
rect 13360 16584 13412 16590
rect 13360 16526 13412 16532
rect 13372 14074 13400 16526
rect 13360 14068 13412 14074
rect 13360 14010 13412 14016
rect 13360 12844 13412 12850
rect 13360 12786 13412 12792
rect 13268 11756 13320 11762
rect 13268 11698 13320 11704
rect 13372 11558 13400 12786
rect 13464 12753 13492 18566
rect 13556 16726 13584 19790
rect 13648 18970 13676 20402
rect 13740 19938 13768 22222
rect 13818 22200 13874 23000
rect 14186 22200 14242 23000
rect 14554 22200 14610 23000
rect 14922 22200 14978 23000
rect 15290 22200 15346 23000
rect 15658 22200 15714 23000
rect 16026 22200 16082 23000
rect 16394 22200 16450 23000
rect 16762 22200 16818 23000
rect 17130 22200 17186 23000
rect 17498 22200 17554 23000
rect 17866 22200 17922 23000
rect 18234 22200 18290 23000
rect 18602 22200 18658 23000
rect 18970 22200 19026 23000
rect 19076 22222 19288 22250
rect 13832 20330 13860 22200
rect 13912 20392 13964 20398
rect 13912 20334 13964 20340
rect 13820 20324 13872 20330
rect 13820 20266 13872 20272
rect 13924 20262 13952 20334
rect 14200 20262 14228 22200
rect 14280 20460 14332 20466
rect 14280 20402 14332 20408
rect 13912 20256 13964 20262
rect 13912 20198 13964 20204
rect 14188 20256 14240 20262
rect 14188 20198 14240 20204
rect 13945 20156 14253 20165
rect 13945 20154 13951 20156
rect 14007 20154 14031 20156
rect 14087 20154 14111 20156
rect 14167 20154 14191 20156
rect 14247 20154 14253 20156
rect 14007 20102 14009 20154
rect 14189 20102 14191 20154
rect 13945 20100 13951 20102
rect 14007 20100 14031 20102
rect 14087 20100 14111 20102
rect 14167 20100 14191 20102
rect 14247 20100 14253 20102
rect 13945 20091 14253 20100
rect 14292 20058 14320 20402
rect 14464 20392 14516 20398
rect 14464 20334 14516 20340
rect 14280 20052 14332 20058
rect 14280 19994 14332 20000
rect 14476 19938 14504 20334
rect 14568 20058 14596 22200
rect 14936 20618 14964 22200
rect 14936 20590 15240 20618
rect 15108 20528 15160 20534
rect 15108 20470 15160 20476
rect 14740 20392 14792 20398
rect 14740 20334 14792 20340
rect 14832 20392 14884 20398
rect 14832 20334 14884 20340
rect 15120 20346 15148 20470
rect 15212 20466 15240 20590
rect 15200 20460 15252 20466
rect 15200 20402 15252 20408
rect 14556 20052 14608 20058
rect 14556 19994 14608 20000
rect 13740 19910 13860 19938
rect 14476 19910 14688 19938
rect 13832 19854 13860 19910
rect 13820 19848 13872 19854
rect 13820 19790 13872 19796
rect 14556 19712 14608 19718
rect 14556 19654 14608 19660
rect 14464 19372 14516 19378
rect 14464 19314 14516 19320
rect 14372 19168 14424 19174
rect 14372 19110 14424 19116
rect 13945 19068 14253 19077
rect 13945 19066 13951 19068
rect 14007 19066 14031 19068
rect 14087 19066 14111 19068
rect 14167 19066 14191 19068
rect 14247 19066 14253 19068
rect 14007 19014 14009 19066
rect 14189 19014 14191 19066
rect 13945 19012 13951 19014
rect 14007 19012 14031 19014
rect 14087 19012 14111 19014
rect 14167 19012 14191 19014
rect 14247 19012 14253 19014
rect 13945 19003 14253 19012
rect 14384 18970 14412 19110
rect 14476 18970 14504 19314
rect 13636 18964 13688 18970
rect 13636 18906 13688 18912
rect 14096 18964 14148 18970
rect 14096 18906 14148 18912
rect 14372 18964 14424 18970
rect 14372 18906 14424 18912
rect 14464 18964 14516 18970
rect 14464 18906 14516 18912
rect 14108 18766 14136 18906
rect 14096 18760 14148 18766
rect 14096 18702 14148 18708
rect 14384 18358 14412 18906
rect 14372 18352 14424 18358
rect 14372 18294 14424 18300
rect 13945 17980 14253 17989
rect 13945 17978 13951 17980
rect 14007 17978 14031 17980
rect 14087 17978 14111 17980
rect 14167 17978 14191 17980
rect 14247 17978 14253 17980
rect 14007 17926 14009 17978
rect 14189 17926 14191 17978
rect 13945 17924 13951 17926
rect 14007 17924 14031 17926
rect 14087 17924 14111 17926
rect 14167 17924 14191 17926
rect 14247 17924 14253 17926
rect 13945 17915 14253 17924
rect 14568 17814 14596 19654
rect 14556 17808 14608 17814
rect 14556 17750 14608 17756
rect 14004 17740 14056 17746
rect 14004 17682 14056 17688
rect 13728 17672 13780 17678
rect 13728 17614 13780 17620
rect 13636 16992 13688 16998
rect 13636 16934 13688 16940
rect 13648 16794 13676 16934
rect 13740 16794 13768 17614
rect 14016 17066 14044 17682
rect 14372 17536 14424 17542
rect 14372 17478 14424 17484
rect 14384 17241 14412 17478
rect 14556 17332 14608 17338
rect 14556 17274 14608 17280
rect 14370 17232 14426 17241
rect 14370 17167 14426 17176
rect 14004 17060 14056 17066
rect 14004 17002 14056 17008
rect 14568 16998 14596 17274
rect 14556 16992 14608 16998
rect 14556 16934 14608 16940
rect 13945 16892 14253 16901
rect 13945 16890 13951 16892
rect 14007 16890 14031 16892
rect 14087 16890 14111 16892
rect 14167 16890 14191 16892
rect 14247 16890 14253 16892
rect 14007 16838 14009 16890
rect 14189 16838 14191 16890
rect 13945 16836 13951 16838
rect 14007 16836 14031 16838
rect 14087 16836 14111 16838
rect 14167 16836 14191 16838
rect 14247 16836 14253 16838
rect 13945 16827 14253 16836
rect 13636 16788 13688 16794
rect 13636 16730 13688 16736
rect 13728 16788 13780 16794
rect 13728 16730 13780 16736
rect 13544 16720 13596 16726
rect 13544 16662 13596 16668
rect 13648 16590 13676 16730
rect 13636 16584 13688 16590
rect 13636 16526 13688 16532
rect 13740 16250 13768 16730
rect 14660 16250 14688 19910
rect 13728 16244 13780 16250
rect 13728 16186 13780 16192
rect 14648 16244 14700 16250
rect 14648 16186 14700 16192
rect 13740 16114 13768 16186
rect 13728 16108 13780 16114
rect 13912 16108 13964 16114
rect 13728 16050 13780 16056
rect 13832 16068 13912 16096
rect 13544 15904 13596 15910
rect 13544 15846 13596 15852
rect 13450 12744 13506 12753
rect 13450 12679 13506 12688
rect 13044 11512 13124 11540
rect 13360 11552 13412 11558
rect 12992 11494 13044 11500
rect 13360 11494 13412 11500
rect 12898 10568 12954 10577
rect 12898 10503 12954 10512
rect 12256 10056 12308 10062
rect 12256 9998 12308 10004
rect 12164 9988 12216 9994
rect 12164 9930 12216 9936
rect 12164 9648 12216 9654
rect 12164 9590 12216 9596
rect 12176 9178 12204 9590
rect 12164 9172 12216 9178
rect 12164 9114 12216 9120
rect 12532 8832 12584 8838
rect 12532 8774 12584 8780
rect 12544 8566 12572 8774
rect 12532 8560 12584 8566
rect 12532 8502 12584 8508
rect 12544 6866 12572 8502
rect 13004 7818 13032 11494
rect 13084 11076 13136 11082
rect 13084 11018 13136 11024
rect 13096 10198 13124 11018
rect 13084 10192 13136 10198
rect 13084 10134 13136 10140
rect 13556 9382 13584 15846
rect 13740 15706 13768 16050
rect 13728 15700 13780 15706
rect 13728 15642 13780 15648
rect 13740 15162 13768 15642
rect 13728 15156 13780 15162
rect 13728 15098 13780 15104
rect 13740 15026 13768 15098
rect 13728 15020 13780 15026
rect 13728 14962 13780 14968
rect 13740 14618 13768 14962
rect 13728 14612 13780 14618
rect 13728 14554 13780 14560
rect 13740 14074 13768 14554
rect 13832 14498 13860 16068
rect 13912 16050 13964 16056
rect 13945 15804 14253 15813
rect 13945 15802 13951 15804
rect 14007 15802 14031 15804
rect 14087 15802 14111 15804
rect 14167 15802 14191 15804
rect 14247 15802 14253 15804
rect 14007 15750 14009 15802
rect 14189 15750 14191 15802
rect 13945 15748 13951 15750
rect 14007 15748 14031 15750
rect 14087 15748 14111 15750
rect 14167 15748 14191 15750
rect 14247 15748 14253 15750
rect 13945 15739 14253 15748
rect 14372 15428 14424 15434
rect 14372 15370 14424 15376
rect 13945 14716 14253 14725
rect 13945 14714 13951 14716
rect 14007 14714 14031 14716
rect 14087 14714 14111 14716
rect 14167 14714 14191 14716
rect 14247 14714 14253 14716
rect 14007 14662 14009 14714
rect 14189 14662 14191 14714
rect 13945 14660 13951 14662
rect 14007 14660 14031 14662
rect 14087 14660 14111 14662
rect 14167 14660 14191 14662
rect 14247 14660 14253 14662
rect 13945 14651 14253 14660
rect 14384 14618 14412 15370
rect 14372 14612 14424 14618
rect 14372 14554 14424 14560
rect 13912 14544 13964 14550
rect 13832 14492 13912 14498
rect 13832 14486 13964 14492
rect 13832 14470 13952 14486
rect 13728 14068 13780 14074
rect 13728 14010 13780 14016
rect 13832 14006 13860 14470
rect 14280 14068 14332 14074
rect 14280 14010 14332 14016
rect 13820 14000 13872 14006
rect 13820 13942 13872 13948
rect 13912 13932 13964 13938
rect 13912 13874 13964 13880
rect 13924 13818 13952 13874
rect 14292 13818 14320 14010
rect 13924 13790 14320 13818
rect 13945 13628 14253 13637
rect 13945 13626 13951 13628
rect 14007 13626 14031 13628
rect 14087 13626 14111 13628
rect 14167 13626 14191 13628
rect 14247 13626 14253 13628
rect 14007 13574 14009 13626
rect 14189 13574 14191 13626
rect 13945 13572 13951 13574
rect 14007 13572 14031 13574
rect 14087 13572 14111 13574
rect 14167 13572 14191 13574
rect 14247 13572 14253 13574
rect 13945 13563 14253 13572
rect 13636 12640 13688 12646
rect 13636 12582 13688 12588
rect 13648 9722 13676 12582
rect 13945 12540 14253 12549
rect 13945 12538 13951 12540
rect 14007 12538 14031 12540
rect 14087 12538 14111 12540
rect 14167 12538 14191 12540
rect 14247 12538 14253 12540
rect 14007 12486 14009 12538
rect 14189 12486 14191 12538
rect 13945 12484 13951 12486
rect 14007 12484 14031 12486
rect 14087 12484 14111 12486
rect 14167 12484 14191 12486
rect 14247 12484 14253 12486
rect 13945 12475 14253 12484
rect 14004 12164 14056 12170
rect 14004 12106 14056 12112
rect 14016 11642 14044 12106
rect 14188 12096 14240 12102
rect 14188 12038 14240 12044
rect 14200 11778 14228 12038
rect 14292 11898 14320 13790
rect 14384 13394 14412 14554
rect 14464 13932 14516 13938
rect 14464 13874 14516 13880
rect 14372 13388 14424 13394
rect 14372 13330 14424 13336
rect 14476 12646 14504 13874
rect 14464 12640 14516 12646
rect 14464 12582 14516 12588
rect 14280 11892 14332 11898
rect 14280 11834 14332 11840
rect 14200 11750 14320 11778
rect 13832 11614 14044 11642
rect 14292 11626 14320 11750
rect 14280 11620 14332 11626
rect 13832 11286 13860 11614
rect 14280 11562 14332 11568
rect 13945 11452 14253 11461
rect 13945 11450 13951 11452
rect 14007 11450 14031 11452
rect 14087 11450 14111 11452
rect 14167 11450 14191 11452
rect 14247 11450 14253 11452
rect 14007 11398 14009 11450
rect 14189 11398 14191 11450
rect 13945 11396 13951 11398
rect 14007 11396 14031 11398
rect 14087 11396 14111 11398
rect 14167 11396 14191 11398
rect 14247 11396 14253 11398
rect 13945 11387 14253 11396
rect 13820 11280 13872 11286
rect 13820 11222 13872 11228
rect 14096 11144 14148 11150
rect 14292 11098 14320 11562
rect 14752 11354 14780 20334
rect 14844 19854 14872 20334
rect 15120 20318 15240 20346
rect 15304 20330 15332 22200
rect 15568 20868 15620 20874
rect 15568 20810 15620 20816
rect 15580 20534 15608 20810
rect 15672 20618 15700 22200
rect 15672 20590 15792 20618
rect 16040 20602 16068 22200
rect 15568 20528 15620 20534
rect 15568 20470 15620 20476
rect 15660 20460 15712 20466
rect 15660 20402 15712 20408
rect 15212 19990 15240 20318
rect 15292 20324 15344 20330
rect 15292 20266 15344 20272
rect 15200 19984 15252 19990
rect 15200 19926 15252 19932
rect 15016 19916 15068 19922
rect 15016 19858 15068 19864
rect 14832 19848 14884 19854
rect 14832 19790 14884 19796
rect 14832 19712 14884 19718
rect 14832 19654 14884 19660
rect 14924 19712 14976 19718
rect 14924 19654 14976 19660
rect 14844 19242 14872 19654
rect 14936 19378 14964 19654
rect 15028 19514 15056 19858
rect 15292 19848 15344 19854
rect 15292 19790 15344 19796
rect 15016 19508 15068 19514
rect 15016 19450 15068 19456
rect 14924 19372 14976 19378
rect 14924 19314 14976 19320
rect 15200 19372 15252 19378
rect 15200 19314 15252 19320
rect 14832 19236 14884 19242
rect 14832 19178 14884 19184
rect 14832 18284 14884 18290
rect 14832 18226 14884 18232
rect 14844 17338 14872 18226
rect 15212 17354 15240 19314
rect 14832 17332 14884 17338
rect 14832 17274 14884 17280
rect 15120 17326 15240 17354
rect 15120 16454 15148 17326
rect 15200 17196 15252 17202
rect 15200 17138 15252 17144
rect 15108 16448 15160 16454
rect 15108 16390 15160 16396
rect 15108 16244 15160 16250
rect 15108 16186 15160 16192
rect 15016 14068 15068 14074
rect 15016 14010 15068 14016
rect 15028 13938 15056 14010
rect 15016 13932 15068 13938
rect 15016 13874 15068 13880
rect 15120 13433 15148 16186
rect 15212 15910 15240 17138
rect 15200 15904 15252 15910
rect 15200 15846 15252 15852
rect 15106 13424 15162 13433
rect 15106 13359 15162 13368
rect 14924 13184 14976 13190
rect 15304 13172 15332 19790
rect 15672 19514 15700 20402
rect 15764 20058 15792 20590
rect 16028 20596 16080 20602
rect 16028 20538 16080 20544
rect 15842 20496 15898 20505
rect 16408 20482 16436 22200
rect 16776 20890 16804 22200
rect 16776 20862 16988 20890
rect 16544 20700 16852 20709
rect 16544 20698 16550 20700
rect 16606 20698 16630 20700
rect 16686 20698 16710 20700
rect 16766 20698 16790 20700
rect 16846 20698 16852 20700
rect 16606 20646 16608 20698
rect 16788 20646 16790 20698
rect 16544 20644 16550 20646
rect 16606 20644 16630 20646
rect 16686 20644 16710 20646
rect 16766 20644 16790 20646
rect 16846 20644 16852 20646
rect 16544 20635 16852 20644
rect 16960 20602 16988 20862
rect 16948 20596 17000 20602
rect 16948 20538 17000 20544
rect 15842 20431 15898 20440
rect 16120 20460 16172 20466
rect 15752 20052 15804 20058
rect 15752 19994 15804 20000
rect 15752 19712 15804 19718
rect 15752 19654 15804 19660
rect 15660 19508 15712 19514
rect 15660 19450 15712 19456
rect 15660 19372 15712 19378
rect 15764 19360 15792 19654
rect 15856 19378 15884 20431
rect 16120 20402 16172 20408
rect 16212 20460 16264 20466
rect 16408 20454 16620 20482
rect 16212 20402 16264 20408
rect 16132 19922 16160 20402
rect 16120 19916 16172 19922
rect 16120 19858 16172 19864
rect 16224 19514 16252 20402
rect 16592 20330 16620 20454
rect 16856 20460 16908 20466
rect 16856 20402 16908 20408
rect 16580 20324 16632 20330
rect 16580 20266 16632 20272
rect 16868 20058 16896 20402
rect 17144 20262 17172 22200
rect 17408 20460 17460 20466
rect 17408 20402 17460 20408
rect 17132 20256 17184 20262
rect 17132 20198 17184 20204
rect 17420 20058 17448 20402
rect 17512 20330 17540 22200
rect 17880 20618 17908 22200
rect 17880 20602 18000 20618
rect 17880 20596 18012 20602
rect 17880 20590 17960 20596
rect 17960 20538 18012 20544
rect 17776 20460 17828 20466
rect 17776 20402 17828 20408
rect 18144 20460 18196 20466
rect 18144 20402 18196 20408
rect 17500 20324 17552 20330
rect 17500 20266 17552 20272
rect 17788 20058 17816 20402
rect 16856 20052 16908 20058
rect 16856 19994 16908 20000
rect 17408 20052 17460 20058
rect 17408 19994 17460 20000
rect 17776 20052 17828 20058
rect 17776 19994 17828 20000
rect 16304 19848 16356 19854
rect 16304 19790 16356 19796
rect 16396 19848 16448 19854
rect 16396 19790 16448 19796
rect 16948 19848 17000 19854
rect 16948 19790 17000 19796
rect 17224 19848 17276 19854
rect 17224 19790 17276 19796
rect 18052 19848 18104 19854
rect 18052 19790 18104 19796
rect 16212 19508 16264 19514
rect 16212 19450 16264 19456
rect 15712 19332 15792 19360
rect 15844 19372 15896 19378
rect 15660 19314 15712 19320
rect 15844 19314 15896 19320
rect 16028 19236 16080 19242
rect 16028 19178 16080 19184
rect 15752 18284 15804 18290
rect 15752 18226 15804 18232
rect 15568 18216 15620 18222
rect 15568 18158 15620 18164
rect 15580 17882 15608 18158
rect 15764 17882 15792 18226
rect 15568 17876 15620 17882
rect 15568 17818 15620 17824
rect 15752 17876 15804 17882
rect 15752 17818 15804 17824
rect 15844 17740 15896 17746
rect 15844 17682 15896 17688
rect 15752 17672 15804 17678
rect 15752 17614 15804 17620
rect 15476 17604 15528 17610
rect 15476 17546 15528 17552
rect 15384 17128 15436 17134
rect 15384 17070 15436 17076
rect 15396 16454 15424 17070
rect 15384 16448 15436 16454
rect 15384 16390 15436 16396
rect 15396 14958 15424 16390
rect 15488 16114 15516 17546
rect 15764 17202 15792 17614
rect 15856 17338 15884 17682
rect 15844 17332 15896 17338
rect 15844 17274 15896 17280
rect 15752 17196 15804 17202
rect 15752 17138 15804 17144
rect 16040 17116 16068 19178
rect 16316 18426 16344 19790
rect 16408 19310 16436 19790
rect 16544 19612 16852 19621
rect 16544 19610 16550 19612
rect 16606 19610 16630 19612
rect 16686 19610 16710 19612
rect 16766 19610 16790 19612
rect 16846 19610 16852 19612
rect 16606 19558 16608 19610
rect 16788 19558 16790 19610
rect 16544 19556 16550 19558
rect 16606 19556 16630 19558
rect 16686 19556 16710 19558
rect 16766 19556 16790 19558
rect 16846 19556 16852 19558
rect 16544 19547 16852 19556
rect 16396 19304 16448 19310
rect 16856 19304 16908 19310
rect 16396 19246 16448 19252
rect 16578 19272 16634 19281
rect 16856 19246 16908 19252
rect 16578 19207 16634 19216
rect 16592 18902 16620 19207
rect 16868 18970 16896 19246
rect 16856 18964 16908 18970
rect 16856 18906 16908 18912
rect 16580 18896 16632 18902
rect 16580 18838 16632 18844
rect 16592 18698 16620 18838
rect 16580 18692 16632 18698
rect 16580 18634 16632 18640
rect 16544 18524 16852 18533
rect 16544 18522 16550 18524
rect 16606 18522 16630 18524
rect 16686 18522 16710 18524
rect 16766 18522 16790 18524
rect 16846 18522 16852 18524
rect 16606 18470 16608 18522
rect 16788 18470 16790 18522
rect 16544 18468 16550 18470
rect 16606 18468 16630 18470
rect 16686 18468 16710 18470
rect 16766 18468 16790 18470
rect 16846 18468 16852 18470
rect 16544 18459 16852 18468
rect 16304 18420 16356 18426
rect 16304 18362 16356 18368
rect 16960 17814 16988 19790
rect 17236 19514 17264 19790
rect 17224 19508 17276 19514
rect 17224 19450 17276 19456
rect 17960 19440 18012 19446
rect 17960 19382 18012 19388
rect 17132 19372 17184 19378
rect 17132 19314 17184 19320
rect 17040 19304 17092 19310
rect 17040 19246 17092 19252
rect 17052 18970 17080 19246
rect 17040 18964 17092 18970
rect 17040 18906 17092 18912
rect 17144 18902 17172 19314
rect 17132 18896 17184 18902
rect 17132 18838 17184 18844
rect 17222 18864 17278 18873
rect 17222 18799 17278 18808
rect 17236 18698 17264 18799
rect 17972 18766 18000 19382
rect 17960 18760 18012 18766
rect 17960 18702 18012 18708
rect 17224 18692 17276 18698
rect 17224 18634 17276 18640
rect 18064 18358 18092 19790
rect 18156 19514 18184 20402
rect 18248 20058 18276 22200
rect 18616 20618 18644 22200
rect 18984 22114 19012 22200
rect 19076 22114 19104 22222
rect 18984 22086 19104 22114
rect 18616 20602 18736 20618
rect 18616 20596 18748 20602
rect 18616 20590 18696 20596
rect 18696 20538 18748 20544
rect 19064 20528 19116 20534
rect 19064 20470 19116 20476
rect 18880 20460 18932 20466
rect 18880 20402 18932 20408
rect 18972 20460 19024 20466
rect 18972 20402 19024 20408
rect 18696 20256 18748 20262
rect 18696 20198 18748 20204
rect 18236 20052 18288 20058
rect 18236 19994 18288 20000
rect 18604 19848 18656 19854
rect 18604 19790 18656 19796
rect 18616 19514 18644 19790
rect 18144 19508 18196 19514
rect 18144 19450 18196 19456
rect 18604 19508 18656 19514
rect 18604 19450 18656 19456
rect 18420 19372 18472 19378
rect 18420 19314 18472 19320
rect 18236 19304 18288 19310
rect 18288 19264 18368 19292
rect 18236 19246 18288 19252
rect 18144 19236 18196 19242
rect 18144 19178 18196 19184
rect 18052 18352 18104 18358
rect 18052 18294 18104 18300
rect 17408 18284 17460 18290
rect 17408 18226 17460 18232
rect 16948 17808 17000 17814
rect 17420 17785 17448 18226
rect 18156 18170 18184 19178
rect 18340 18630 18368 19264
rect 18328 18624 18380 18630
rect 18328 18566 18380 18572
rect 18064 18142 18184 18170
rect 18340 18154 18368 18566
rect 18432 18426 18460 19314
rect 18420 18420 18472 18426
rect 18420 18362 18472 18368
rect 18708 18329 18736 20198
rect 18892 20058 18920 20402
rect 18880 20052 18932 20058
rect 18880 19994 18932 20000
rect 18788 19848 18840 19854
rect 18788 19790 18840 19796
rect 18800 18737 18828 19790
rect 18984 19514 19012 20402
rect 19076 19514 19104 20470
rect 19260 20346 19288 22222
rect 19338 22200 19394 23000
rect 19706 22200 19762 23000
rect 20074 22200 20130 23000
rect 20442 22200 20498 23000
rect 20810 22200 20866 23000
rect 21178 22200 21234 23000
rect 19352 20448 19380 22200
rect 19616 20460 19668 20466
rect 19352 20420 19472 20448
rect 19260 20330 19380 20346
rect 19260 20324 19392 20330
rect 19260 20318 19340 20324
rect 19340 20266 19392 20272
rect 19444 20262 19472 20420
rect 19616 20402 19668 20408
rect 19628 20369 19656 20402
rect 19720 20398 19748 22200
rect 20088 20602 20116 22200
rect 20076 20596 20128 20602
rect 20076 20538 20128 20544
rect 19890 20496 19946 20505
rect 19890 20431 19946 20440
rect 19984 20460 20036 20466
rect 19708 20392 19760 20398
rect 19614 20360 19670 20369
rect 19708 20334 19760 20340
rect 19614 20295 19670 20304
rect 19432 20256 19484 20262
rect 19432 20198 19484 20204
rect 19143 20156 19451 20165
rect 19143 20154 19149 20156
rect 19205 20154 19229 20156
rect 19285 20154 19309 20156
rect 19365 20154 19389 20156
rect 19445 20154 19451 20156
rect 19205 20102 19207 20154
rect 19387 20102 19389 20154
rect 19143 20100 19149 20102
rect 19205 20100 19229 20102
rect 19285 20100 19309 20102
rect 19365 20100 19389 20102
rect 19445 20100 19451 20102
rect 19143 20091 19451 20100
rect 19904 20058 19932 20431
rect 19984 20402 20036 20408
rect 20352 20460 20404 20466
rect 20352 20402 20404 20408
rect 19892 20052 19944 20058
rect 19892 19994 19944 20000
rect 19708 19848 19760 19854
rect 19996 19825 20024 20402
rect 20258 20088 20314 20097
rect 20258 20023 20260 20032
rect 20312 20023 20314 20032
rect 20260 19994 20312 20000
rect 20364 19961 20392 20402
rect 20456 20262 20484 22200
rect 20444 20256 20496 20262
rect 20444 20198 20496 20204
rect 20824 20058 20852 22200
rect 20902 20904 20958 20913
rect 20902 20839 20958 20848
rect 20812 20052 20864 20058
rect 20812 19994 20864 20000
rect 20350 19952 20406 19961
rect 20350 19887 20406 19896
rect 20260 19848 20312 19854
rect 19708 19790 19760 19796
rect 19982 19816 20038 19825
rect 18972 19508 19024 19514
rect 18972 19450 19024 19456
rect 19064 19508 19116 19514
rect 19064 19450 19116 19456
rect 18880 19372 18932 19378
rect 18880 19314 18932 19320
rect 19524 19372 19576 19378
rect 19524 19314 19576 19320
rect 18786 18728 18842 18737
rect 18786 18663 18842 18672
rect 18694 18320 18750 18329
rect 18694 18255 18750 18264
rect 18420 18216 18472 18222
rect 18420 18158 18472 18164
rect 18328 18148 18380 18154
rect 18064 18086 18092 18142
rect 18328 18090 18380 18096
rect 18052 18080 18104 18086
rect 18052 18022 18104 18028
rect 17500 17808 17552 17814
rect 16948 17750 17000 17756
rect 17406 17776 17462 17785
rect 17500 17750 17552 17756
rect 17406 17711 17462 17720
rect 16304 17672 16356 17678
rect 16304 17614 16356 17620
rect 16316 17338 16344 17614
rect 16948 17536 17000 17542
rect 16948 17478 17000 17484
rect 17224 17536 17276 17542
rect 17224 17478 17276 17484
rect 17408 17536 17460 17542
rect 17408 17478 17460 17484
rect 16544 17436 16852 17445
rect 16544 17434 16550 17436
rect 16606 17434 16630 17436
rect 16686 17434 16710 17436
rect 16766 17434 16790 17436
rect 16846 17434 16852 17436
rect 16606 17382 16608 17434
rect 16788 17382 16790 17434
rect 16544 17380 16550 17382
rect 16606 17380 16630 17382
rect 16686 17380 16710 17382
rect 16766 17380 16790 17382
rect 16846 17380 16852 17382
rect 16544 17371 16852 17380
rect 16304 17332 16356 17338
rect 16304 17274 16356 17280
rect 15948 17088 16068 17116
rect 15476 16108 15528 16114
rect 15476 16050 15528 16056
rect 15488 15706 15516 16050
rect 15752 15904 15804 15910
rect 15752 15846 15804 15852
rect 15476 15700 15528 15706
rect 15476 15642 15528 15648
rect 15476 15156 15528 15162
rect 15476 15098 15528 15104
rect 15384 14952 15436 14958
rect 15384 14894 15436 14900
rect 15488 14482 15516 15098
rect 15764 14958 15792 15846
rect 15752 14952 15804 14958
rect 15752 14894 15804 14900
rect 15476 14476 15528 14482
rect 15476 14418 15528 14424
rect 15568 14408 15620 14414
rect 15568 14350 15620 14356
rect 15476 13728 15528 13734
rect 15476 13670 15528 13676
rect 15488 13394 15516 13670
rect 15580 13394 15608 14350
rect 15844 13864 15896 13870
rect 15844 13806 15896 13812
rect 15752 13796 15804 13802
rect 15752 13738 15804 13744
rect 15476 13388 15528 13394
rect 15476 13330 15528 13336
rect 15568 13388 15620 13394
rect 15568 13330 15620 13336
rect 14976 13144 15332 13172
rect 15568 13184 15620 13190
rect 14924 13126 14976 13132
rect 15568 13126 15620 13132
rect 15580 12434 15608 13126
rect 15764 12850 15792 13738
rect 15856 13326 15884 13806
rect 15948 13433 15976 17088
rect 16960 16726 16988 17478
rect 17040 17196 17092 17202
rect 17040 17138 17092 17144
rect 16948 16720 17000 16726
rect 16948 16662 17000 16668
rect 16316 16510 16528 16538
rect 16316 16250 16344 16510
rect 16500 16454 16528 16510
rect 16396 16448 16448 16454
rect 16396 16390 16448 16396
rect 16488 16448 16540 16454
rect 16488 16390 16540 16396
rect 16408 16250 16436 16390
rect 16544 16348 16852 16357
rect 16544 16346 16550 16348
rect 16606 16346 16630 16348
rect 16686 16346 16710 16348
rect 16766 16346 16790 16348
rect 16846 16346 16852 16348
rect 16606 16294 16608 16346
rect 16788 16294 16790 16346
rect 16544 16292 16550 16294
rect 16606 16292 16630 16294
rect 16686 16292 16710 16294
rect 16766 16292 16790 16294
rect 16846 16292 16852 16294
rect 16544 16283 16852 16292
rect 16304 16244 16356 16250
rect 16304 16186 16356 16192
rect 16396 16244 16448 16250
rect 16396 16186 16448 16192
rect 16212 16176 16264 16182
rect 16212 16118 16264 16124
rect 16118 15600 16174 15609
rect 16118 15535 16174 15544
rect 16028 14340 16080 14346
rect 16028 14282 16080 14288
rect 16040 13734 16068 14282
rect 16028 13728 16080 13734
rect 16028 13670 16080 13676
rect 15934 13424 15990 13433
rect 15934 13359 15990 13368
rect 15844 13320 15896 13326
rect 15844 13262 15896 13268
rect 16040 13190 16068 13670
rect 16028 13184 16080 13190
rect 16028 13126 16080 13132
rect 15752 12844 15804 12850
rect 15752 12786 15804 12792
rect 15304 12406 15608 12434
rect 14740 11348 14792 11354
rect 14740 11290 14792 11296
rect 14148 11092 14320 11098
rect 14096 11086 14320 11092
rect 14108 11070 14320 11086
rect 14464 11076 14516 11082
rect 14108 10810 14136 11070
rect 14464 11018 14516 11024
rect 14096 10804 14148 10810
rect 14096 10746 14148 10752
rect 14476 10470 14504 11018
rect 14648 10600 14700 10606
rect 14752 10588 14780 11290
rect 14700 10560 14780 10588
rect 14648 10542 14700 10548
rect 14464 10464 14516 10470
rect 14464 10406 14516 10412
rect 13945 10364 14253 10373
rect 13945 10362 13951 10364
rect 14007 10362 14031 10364
rect 14087 10362 14111 10364
rect 14167 10362 14191 10364
rect 14247 10362 14253 10364
rect 14007 10310 14009 10362
rect 14189 10310 14191 10362
rect 13945 10308 13951 10310
rect 14007 10308 14031 10310
rect 14087 10308 14111 10310
rect 14167 10308 14191 10310
rect 14247 10308 14253 10310
rect 13945 10299 14253 10308
rect 13636 9716 13688 9722
rect 13636 9658 13688 9664
rect 13544 9376 13596 9382
rect 13544 9318 13596 9324
rect 13820 9376 13872 9382
rect 13820 9318 13872 9324
rect 13360 8968 13412 8974
rect 13360 8910 13412 8916
rect 12992 7812 13044 7818
rect 12992 7754 13044 7760
rect 12532 6860 12584 6866
rect 12532 6802 12584 6808
rect 12716 6656 12768 6662
rect 12716 6598 12768 6604
rect 12728 6458 12756 6598
rect 12032 6412 12112 6440
rect 12716 6452 12768 6458
rect 11980 6394 12032 6400
rect 12716 6394 12768 6400
rect 13084 6316 13136 6322
rect 13084 6258 13136 6264
rect 13096 5681 13124 6258
rect 13372 6254 13400 8910
rect 13832 8838 13860 9318
rect 13945 9276 14253 9285
rect 13945 9274 13951 9276
rect 14007 9274 14031 9276
rect 14087 9274 14111 9276
rect 14167 9274 14191 9276
rect 14247 9274 14253 9276
rect 14007 9222 14009 9274
rect 14189 9222 14191 9274
rect 13945 9220 13951 9222
rect 14007 9220 14031 9222
rect 14087 9220 14111 9222
rect 14167 9220 14191 9222
rect 14247 9220 14253 9222
rect 13945 9211 14253 9220
rect 13912 9172 13964 9178
rect 13912 9114 13964 9120
rect 13924 8838 13952 9114
rect 14476 8906 14504 10406
rect 15304 9625 15332 12406
rect 15384 12368 15436 12374
rect 15384 12310 15436 12316
rect 15396 10742 15424 12310
rect 16132 11830 16160 15535
rect 16224 12918 16252 16118
rect 17052 15978 17080 17138
rect 17132 17128 17184 17134
rect 17132 17070 17184 17076
rect 17040 15972 17092 15978
rect 17040 15914 17092 15920
rect 17144 15706 17172 17070
rect 17236 16250 17264 17478
rect 17420 17270 17448 17478
rect 17408 17264 17460 17270
rect 17314 17232 17370 17241
rect 17408 17206 17460 17212
rect 17314 17167 17370 17176
rect 17328 17134 17356 17167
rect 17316 17128 17368 17134
rect 17316 17070 17368 17076
rect 17512 16590 17540 17750
rect 17592 17740 17644 17746
rect 17592 17682 17644 17688
rect 17604 17116 17632 17682
rect 18064 17678 18092 18022
rect 18052 17672 18104 17678
rect 18052 17614 18104 17620
rect 17684 17604 17736 17610
rect 17684 17546 17736 17552
rect 17696 17338 17724 17546
rect 17684 17332 17736 17338
rect 17684 17274 17736 17280
rect 17776 17264 17828 17270
rect 17776 17206 17828 17212
rect 17684 17128 17736 17134
rect 17604 17088 17684 17116
rect 17684 17070 17736 17076
rect 17500 16584 17552 16590
rect 17500 16526 17552 16532
rect 17696 16522 17724 17070
rect 17684 16516 17736 16522
rect 17684 16458 17736 16464
rect 17788 16454 17816 17206
rect 17868 17196 17920 17202
rect 17868 17138 17920 17144
rect 17880 16794 17908 17138
rect 18064 17105 18092 17614
rect 18144 17536 18196 17542
rect 18144 17478 18196 17484
rect 18050 17096 18106 17105
rect 18050 17031 18106 17040
rect 18156 16794 18184 17478
rect 18236 17196 18288 17202
rect 18236 17138 18288 17144
rect 17868 16788 17920 16794
rect 17868 16730 17920 16736
rect 18144 16788 18196 16794
rect 18144 16730 18196 16736
rect 18052 16652 18104 16658
rect 18052 16594 18104 16600
rect 17316 16448 17368 16454
rect 17316 16390 17368 16396
rect 17776 16448 17828 16454
rect 17776 16390 17828 16396
rect 17224 16244 17276 16250
rect 17224 16186 17276 16192
rect 17132 15700 17184 15706
rect 17132 15642 17184 15648
rect 16948 15496 17000 15502
rect 16948 15438 17000 15444
rect 16544 15260 16852 15269
rect 16544 15258 16550 15260
rect 16606 15258 16630 15260
rect 16686 15258 16710 15260
rect 16766 15258 16790 15260
rect 16846 15258 16852 15260
rect 16606 15206 16608 15258
rect 16788 15206 16790 15258
rect 16544 15204 16550 15206
rect 16606 15204 16630 15206
rect 16686 15204 16710 15206
rect 16766 15204 16790 15206
rect 16846 15204 16852 15206
rect 16544 15195 16852 15204
rect 16960 15162 16988 15438
rect 16948 15156 17000 15162
rect 16948 15098 17000 15104
rect 17224 14952 17276 14958
rect 17224 14894 17276 14900
rect 17236 14618 17264 14894
rect 17224 14612 17276 14618
rect 17224 14554 17276 14560
rect 16396 14408 16448 14414
rect 16396 14350 16448 14356
rect 16408 14074 16436 14350
rect 16544 14172 16852 14181
rect 16544 14170 16550 14172
rect 16606 14170 16630 14172
rect 16686 14170 16710 14172
rect 16766 14170 16790 14172
rect 16846 14170 16852 14172
rect 16606 14118 16608 14170
rect 16788 14118 16790 14170
rect 16544 14116 16550 14118
rect 16606 14116 16630 14118
rect 16686 14116 16710 14118
rect 16766 14116 16790 14118
rect 16846 14116 16852 14118
rect 16544 14107 16852 14116
rect 16396 14068 16448 14074
rect 16396 14010 16448 14016
rect 16580 14000 16632 14006
rect 16580 13942 16632 13948
rect 16592 13462 16620 13942
rect 16948 13932 17000 13938
rect 16948 13874 17000 13880
rect 16580 13456 16632 13462
rect 16580 13398 16632 13404
rect 16544 13084 16852 13093
rect 16544 13082 16550 13084
rect 16606 13082 16630 13084
rect 16686 13082 16710 13084
rect 16766 13082 16790 13084
rect 16846 13082 16852 13084
rect 16606 13030 16608 13082
rect 16788 13030 16790 13082
rect 16544 13028 16550 13030
rect 16606 13028 16630 13030
rect 16686 13028 16710 13030
rect 16766 13028 16790 13030
rect 16846 13028 16852 13030
rect 16544 13019 16852 13028
rect 16212 12912 16264 12918
rect 16212 12854 16264 12860
rect 16764 12776 16816 12782
rect 16764 12718 16816 12724
rect 16776 12442 16804 12718
rect 16764 12436 16816 12442
rect 16764 12378 16816 12384
rect 16544 11996 16852 12005
rect 16544 11994 16550 11996
rect 16606 11994 16630 11996
rect 16686 11994 16710 11996
rect 16766 11994 16790 11996
rect 16846 11994 16852 11996
rect 16606 11942 16608 11994
rect 16788 11942 16790 11994
rect 16544 11940 16550 11942
rect 16606 11940 16630 11942
rect 16686 11940 16710 11942
rect 16766 11940 16790 11942
rect 16846 11940 16852 11942
rect 16544 11931 16852 11940
rect 16120 11824 16172 11830
rect 16120 11766 16172 11772
rect 15568 11756 15620 11762
rect 15568 11698 15620 11704
rect 15580 11286 15608 11698
rect 15660 11688 15712 11694
rect 15660 11630 15712 11636
rect 15568 11280 15620 11286
rect 15568 11222 15620 11228
rect 15672 10810 15700 11630
rect 16580 11552 16632 11558
rect 16580 11494 16632 11500
rect 16960 11506 16988 13874
rect 17132 13864 17184 13870
rect 17130 13832 17132 13841
rect 17184 13832 17186 13841
rect 17130 13767 17186 13776
rect 17040 13184 17092 13190
rect 17040 13126 17092 13132
rect 17132 13184 17184 13190
rect 17132 13126 17184 13132
rect 17052 12986 17080 13126
rect 17040 12980 17092 12986
rect 17040 12922 17092 12928
rect 17040 12708 17092 12714
rect 17040 12650 17092 12656
rect 17052 12306 17080 12650
rect 17040 12300 17092 12306
rect 17040 12242 17092 12248
rect 17052 11801 17080 12242
rect 17144 12102 17172 13126
rect 17132 12096 17184 12102
rect 17132 12038 17184 12044
rect 17224 12096 17276 12102
rect 17224 12038 17276 12044
rect 17038 11792 17094 11801
rect 17038 11727 17094 11736
rect 17132 11756 17184 11762
rect 17132 11698 17184 11704
rect 15750 11248 15806 11257
rect 16592 11218 16620 11494
rect 16960 11478 17080 11506
rect 16948 11348 17000 11354
rect 16948 11290 17000 11296
rect 15750 11183 15806 11192
rect 16212 11212 16264 11218
rect 15660 10804 15712 10810
rect 15660 10746 15712 10752
rect 15384 10736 15436 10742
rect 15384 10678 15436 10684
rect 15672 10606 15700 10746
rect 15660 10600 15712 10606
rect 15660 10542 15712 10548
rect 15672 10130 15700 10542
rect 15660 10124 15712 10130
rect 15660 10066 15712 10072
rect 15384 9988 15436 9994
rect 15436 9948 15516 9976
rect 15384 9930 15436 9936
rect 14554 9616 14610 9625
rect 15290 9616 15346 9625
rect 14554 9551 14556 9560
rect 14608 9551 14610 9560
rect 15016 9580 15068 9586
rect 14556 9522 14608 9528
rect 15290 9551 15346 9560
rect 15016 9522 15068 9528
rect 15028 9178 15056 9522
rect 15488 9382 15516 9948
rect 15764 9518 15792 11183
rect 16212 11154 16264 11160
rect 16580 11212 16632 11218
rect 16580 11154 16632 11160
rect 16224 11082 16252 11154
rect 16212 11076 16264 11082
rect 16212 11018 16264 11024
rect 16396 11008 16448 11014
rect 16396 10950 16448 10956
rect 16408 10606 16436 10950
rect 16544 10908 16852 10917
rect 16544 10906 16550 10908
rect 16606 10906 16630 10908
rect 16686 10906 16710 10908
rect 16766 10906 16790 10908
rect 16846 10906 16852 10908
rect 16606 10854 16608 10906
rect 16788 10854 16790 10906
rect 16544 10852 16550 10854
rect 16606 10852 16630 10854
rect 16686 10852 16710 10854
rect 16766 10852 16790 10854
rect 16846 10852 16852 10854
rect 16544 10843 16852 10852
rect 16764 10804 16816 10810
rect 16764 10746 16816 10752
rect 16396 10600 16448 10606
rect 16396 10542 16448 10548
rect 16396 10464 16448 10470
rect 16396 10406 16448 10412
rect 16408 9625 16436 10406
rect 16578 10160 16634 10169
rect 16578 10095 16580 10104
rect 16632 10095 16634 10104
rect 16580 10066 16632 10072
rect 16776 9926 16804 10746
rect 16960 10690 16988 11290
rect 17052 10810 17080 11478
rect 17144 11354 17172 11698
rect 17132 11348 17184 11354
rect 17132 11290 17184 11296
rect 17040 10804 17092 10810
rect 17040 10746 17092 10752
rect 17236 10690 17264 12038
rect 17328 11914 17356 16390
rect 17960 16244 18012 16250
rect 17960 16186 18012 16192
rect 17972 16153 18000 16186
rect 17958 16144 18014 16153
rect 17958 16079 18014 16088
rect 17592 16040 17644 16046
rect 17592 15982 17644 15988
rect 17604 15570 17632 15982
rect 17592 15564 17644 15570
rect 17592 15506 17644 15512
rect 17960 15496 18012 15502
rect 17960 15438 18012 15444
rect 17972 14890 18000 15438
rect 17960 14884 18012 14890
rect 17960 14826 18012 14832
rect 17868 14272 17920 14278
rect 17868 14214 17920 14220
rect 17684 13796 17736 13802
rect 17684 13738 17736 13744
rect 17592 13388 17644 13394
rect 17592 13330 17644 13336
rect 17500 12844 17552 12850
rect 17500 12786 17552 12792
rect 17512 12306 17540 12786
rect 17604 12646 17632 13330
rect 17592 12640 17644 12646
rect 17592 12582 17644 12588
rect 17500 12300 17552 12306
rect 17500 12242 17552 12248
rect 17328 11886 17540 11914
rect 17316 11824 17368 11830
rect 17316 11766 17368 11772
rect 17328 11354 17356 11766
rect 17512 11540 17540 11886
rect 17604 11694 17632 12582
rect 17592 11688 17644 11694
rect 17592 11630 17644 11636
rect 17512 11512 17632 11540
rect 17316 11348 17368 11354
rect 17316 11290 17368 11296
rect 16960 10662 17172 10690
rect 17236 10662 17356 10690
rect 17040 10600 17092 10606
rect 17040 10542 17092 10548
rect 17052 10130 17080 10542
rect 16856 10124 16908 10130
rect 16856 10066 16908 10072
rect 17040 10124 17092 10130
rect 17040 10066 17092 10072
rect 16868 9976 16896 10066
rect 16868 9948 16988 9976
rect 16764 9920 16816 9926
rect 16764 9862 16816 9868
rect 16544 9820 16852 9829
rect 16544 9818 16550 9820
rect 16606 9818 16630 9820
rect 16686 9818 16710 9820
rect 16766 9818 16790 9820
rect 16846 9818 16852 9820
rect 16606 9766 16608 9818
rect 16788 9766 16790 9818
rect 16544 9764 16550 9766
rect 16606 9764 16630 9766
rect 16686 9764 16710 9766
rect 16766 9764 16790 9766
rect 16846 9764 16852 9766
rect 16544 9755 16852 9764
rect 16394 9616 16450 9625
rect 16394 9551 16450 9560
rect 15752 9512 15804 9518
rect 15752 9454 15804 9460
rect 16396 9444 16448 9450
rect 16396 9386 16448 9392
rect 15476 9376 15528 9382
rect 15476 9318 15528 9324
rect 15016 9172 15068 9178
rect 15016 9114 15068 9120
rect 15660 8968 15712 8974
rect 15660 8910 15712 8916
rect 14464 8900 14516 8906
rect 14464 8842 14516 8848
rect 13820 8832 13872 8838
rect 13820 8774 13872 8780
rect 13912 8832 13964 8838
rect 13912 8774 13964 8780
rect 13832 8566 13860 8774
rect 13820 8560 13872 8566
rect 13820 8502 13872 8508
rect 13832 7886 13860 8502
rect 13924 8362 13952 8774
rect 15672 8634 15700 8910
rect 15660 8628 15712 8634
rect 15660 8570 15712 8576
rect 16408 8566 16436 9386
rect 16960 8906 16988 9948
rect 17144 9722 17172 10662
rect 17224 10600 17276 10606
rect 17224 10542 17276 10548
rect 17236 10266 17264 10542
rect 17224 10260 17276 10266
rect 17224 10202 17276 10208
rect 17224 9920 17276 9926
rect 17224 9862 17276 9868
rect 17132 9716 17184 9722
rect 17132 9658 17184 9664
rect 16948 8900 17000 8906
rect 16948 8842 17000 8848
rect 17040 8832 17092 8838
rect 17040 8774 17092 8780
rect 16544 8732 16852 8741
rect 16544 8730 16550 8732
rect 16606 8730 16630 8732
rect 16686 8730 16710 8732
rect 16766 8730 16790 8732
rect 16846 8730 16852 8732
rect 16606 8678 16608 8730
rect 16788 8678 16790 8730
rect 16544 8676 16550 8678
rect 16606 8676 16630 8678
rect 16686 8676 16710 8678
rect 16766 8676 16790 8678
rect 16846 8676 16852 8678
rect 16544 8667 16852 8676
rect 17052 8650 17080 8774
rect 17144 8673 17172 9658
rect 16580 8628 16632 8634
rect 16580 8570 16632 8576
rect 16960 8622 17080 8650
rect 17130 8664 17186 8673
rect 16396 8560 16448 8566
rect 16396 8502 16448 8508
rect 14280 8492 14332 8498
rect 14280 8434 14332 8440
rect 13912 8356 13964 8362
rect 13912 8298 13964 8304
rect 13945 8188 14253 8197
rect 13945 8186 13951 8188
rect 14007 8186 14031 8188
rect 14087 8186 14111 8188
rect 14167 8186 14191 8188
rect 14247 8186 14253 8188
rect 14007 8134 14009 8186
rect 14189 8134 14191 8186
rect 13945 8132 13951 8134
rect 14007 8132 14031 8134
rect 14087 8132 14111 8134
rect 14167 8132 14191 8134
rect 14247 8132 14253 8134
rect 13945 8123 14253 8132
rect 14292 8022 14320 8434
rect 16592 8362 16620 8570
rect 16960 8514 16988 8622
rect 17130 8599 17186 8608
rect 16684 8486 16988 8514
rect 17040 8492 17092 8498
rect 15200 8356 15252 8362
rect 15200 8298 15252 8304
rect 16580 8356 16632 8362
rect 16580 8298 16632 8304
rect 14280 8016 14332 8022
rect 14280 7958 14332 7964
rect 13820 7880 13872 7886
rect 13820 7822 13872 7828
rect 15212 7818 15240 8298
rect 16592 7970 16620 8298
rect 16500 7954 16620 7970
rect 16488 7948 16620 7954
rect 16540 7942 16620 7948
rect 16488 7890 16540 7896
rect 16684 7886 16712 8486
rect 17040 8434 17092 8440
rect 16948 8424 17000 8430
rect 16948 8366 17000 8372
rect 16960 8090 16988 8366
rect 16948 8084 17000 8090
rect 16948 8026 17000 8032
rect 16672 7880 16724 7886
rect 16672 7822 16724 7828
rect 13728 7812 13780 7818
rect 13728 7754 13780 7760
rect 15200 7812 15252 7818
rect 15200 7754 15252 7760
rect 16396 7812 16448 7818
rect 16396 7754 16448 7760
rect 13740 6322 13768 7754
rect 16408 7342 16436 7754
rect 16544 7644 16852 7653
rect 16544 7642 16550 7644
rect 16606 7642 16630 7644
rect 16686 7642 16710 7644
rect 16766 7642 16790 7644
rect 16846 7642 16852 7644
rect 16606 7590 16608 7642
rect 16788 7590 16790 7642
rect 16544 7588 16550 7590
rect 16606 7588 16630 7590
rect 16686 7588 16710 7590
rect 16766 7588 16790 7590
rect 16846 7588 16852 7590
rect 16544 7579 16852 7588
rect 17052 7546 17080 8434
rect 17236 7993 17264 9862
rect 17328 8566 17356 10662
rect 17408 10668 17460 10674
rect 17408 10610 17460 10616
rect 17420 10266 17448 10610
rect 17408 10260 17460 10266
rect 17408 10202 17460 10208
rect 17500 9716 17552 9722
rect 17500 9658 17552 9664
rect 17408 8968 17460 8974
rect 17512 8945 17540 9658
rect 17408 8910 17460 8916
rect 17498 8936 17554 8945
rect 17420 8634 17448 8910
rect 17498 8871 17500 8880
rect 17552 8871 17554 8880
rect 17500 8842 17552 8848
rect 17604 8838 17632 11512
rect 17696 11286 17724 13738
rect 17880 13326 17908 14214
rect 17868 13320 17920 13326
rect 17868 13262 17920 13268
rect 17776 13184 17828 13190
rect 17776 13126 17828 13132
rect 17788 11898 17816 13126
rect 17868 12232 17920 12238
rect 17868 12174 17920 12180
rect 17880 12102 17908 12174
rect 17868 12096 17920 12102
rect 17868 12038 17920 12044
rect 17776 11892 17828 11898
rect 17776 11834 17828 11840
rect 17774 11792 17830 11801
rect 17774 11727 17830 11736
rect 17788 11558 17816 11727
rect 17776 11552 17828 11558
rect 17776 11494 17828 11500
rect 17684 11280 17736 11286
rect 17684 11222 17736 11228
rect 17684 9104 17736 9110
rect 17684 9046 17736 9052
rect 17592 8832 17644 8838
rect 17590 8800 17592 8809
rect 17644 8800 17646 8809
rect 17590 8735 17646 8744
rect 17408 8628 17460 8634
rect 17408 8570 17460 8576
rect 17316 8560 17368 8566
rect 17316 8502 17368 8508
rect 17696 8294 17724 9046
rect 17500 8288 17552 8294
rect 17500 8230 17552 8236
rect 17684 8288 17736 8294
rect 17684 8230 17736 8236
rect 17222 7984 17278 7993
rect 17222 7919 17278 7928
rect 17512 7546 17540 8230
rect 17788 7886 17816 11494
rect 17880 10713 17908 12038
rect 17960 11688 18012 11694
rect 17960 11630 18012 11636
rect 17972 11218 18000 11630
rect 17960 11212 18012 11218
rect 17960 11154 18012 11160
rect 17960 11076 18012 11082
rect 17960 11018 18012 11024
rect 17866 10704 17922 10713
rect 17866 10639 17922 10648
rect 17972 9926 18000 11018
rect 17960 9920 18012 9926
rect 17960 9862 18012 9868
rect 17958 9480 18014 9489
rect 17958 9415 18014 9424
rect 17972 9110 18000 9415
rect 17960 9104 18012 9110
rect 17960 9046 18012 9052
rect 17972 8634 18000 9046
rect 17960 8628 18012 8634
rect 17960 8570 18012 8576
rect 18064 7886 18092 16594
rect 18144 16584 18196 16590
rect 18142 16552 18144 16561
rect 18196 16552 18198 16561
rect 18142 16487 18198 16496
rect 18156 16046 18184 16487
rect 18144 16040 18196 16046
rect 18144 15982 18196 15988
rect 18144 15700 18196 15706
rect 18144 15642 18196 15648
rect 18156 15434 18184 15642
rect 18144 15428 18196 15434
rect 18144 15370 18196 15376
rect 18156 15094 18184 15370
rect 18144 15088 18196 15094
rect 18144 15030 18196 15036
rect 18248 14074 18276 17138
rect 18236 14068 18288 14074
rect 18236 14010 18288 14016
rect 18236 13932 18288 13938
rect 18236 13874 18288 13880
rect 18144 13864 18196 13870
rect 18144 13806 18196 13812
rect 18156 12186 18184 13806
rect 18248 13530 18276 13874
rect 18236 13524 18288 13530
rect 18236 13466 18288 13472
rect 18340 12209 18368 18090
rect 18432 17678 18460 18158
rect 18788 17740 18840 17746
rect 18788 17682 18840 17688
rect 18420 17672 18472 17678
rect 18420 17614 18472 17620
rect 18800 16726 18828 17682
rect 18788 16720 18840 16726
rect 18788 16662 18840 16668
rect 18604 16448 18656 16454
rect 18604 16390 18656 16396
rect 18616 15978 18644 16390
rect 18788 16108 18840 16114
rect 18788 16050 18840 16056
rect 18604 15972 18656 15978
rect 18604 15914 18656 15920
rect 18418 15464 18474 15473
rect 18418 15399 18474 15408
rect 18432 15366 18460 15399
rect 18420 15360 18472 15366
rect 18420 15302 18472 15308
rect 18696 14884 18748 14890
rect 18696 14826 18748 14832
rect 18708 14482 18736 14826
rect 18696 14476 18748 14482
rect 18696 14418 18748 14424
rect 18512 14340 18564 14346
rect 18512 14282 18564 14288
rect 18420 12776 18472 12782
rect 18420 12718 18472 12724
rect 18432 12306 18460 12718
rect 18420 12300 18472 12306
rect 18420 12242 18472 12248
rect 18326 12200 18382 12209
rect 18156 12158 18276 12186
rect 18144 12096 18196 12102
rect 18144 12038 18196 12044
rect 18156 10810 18184 12038
rect 18248 11626 18276 12158
rect 18326 12135 18382 12144
rect 18328 12096 18380 12102
rect 18328 12038 18380 12044
rect 18340 11898 18368 12038
rect 18328 11892 18380 11898
rect 18328 11834 18380 11840
rect 18236 11620 18288 11626
rect 18236 11562 18288 11568
rect 18328 11620 18380 11626
rect 18328 11562 18380 11568
rect 18340 11082 18368 11562
rect 18432 11150 18460 12242
rect 18420 11144 18472 11150
rect 18420 11086 18472 11092
rect 18328 11076 18380 11082
rect 18328 11018 18380 11024
rect 18144 10804 18196 10810
rect 18340 10792 18368 11018
rect 18340 10764 18460 10792
rect 18144 10746 18196 10752
rect 18234 10704 18290 10713
rect 18234 10639 18290 10648
rect 18328 10668 18380 10674
rect 18144 9648 18196 9654
rect 18142 9616 18144 9625
rect 18196 9616 18198 9625
rect 18142 9551 18198 9560
rect 18144 9512 18196 9518
rect 18144 9454 18196 9460
rect 18156 9178 18184 9454
rect 18144 9172 18196 9178
rect 18144 9114 18196 9120
rect 18156 8906 18184 9114
rect 18144 8900 18196 8906
rect 18144 8842 18196 8848
rect 17776 7880 17828 7886
rect 17776 7822 17828 7828
rect 18052 7880 18104 7886
rect 18052 7822 18104 7828
rect 17868 7812 17920 7818
rect 17868 7754 17920 7760
rect 17776 7744 17828 7750
rect 17776 7686 17828 7692
rect 17788 7546 17816 7686
rect 17040 7540 17092 7546
rect 17040 7482 17092 7488
rect 17500 7540 17552 7546
rect 17500 7482 17552 7488
rect 17776 7540 17828 7546
rect 17776 7482 17828 7488
rect 17880 7426 17908 7754
rect 17960 7744 18012 7750
rect 17960 7686 18012 7692
rect 17972 7478 18000 7686
rect 18064 7478 18092 7822
rect 17788 7398 17908 7426
rect 17960 7472 18012 7478
rect 17960 7414 18012 7420
rect 18052 7472 18104 7478
rect 18052 7414 18104 7420
rect 16396 7336 16448 7342
rect 16396 7278 16448 7284
rect 17788 7206 17816 7398
rect 17776 7200 17828 7206
rect 17776 7142 17828 7148
rect 13945 7100 14253 7109
rect 13945 7098 13951 7100
rect 14007 7098 14031 7100
rect 14087 7098 14111 7100
rect 14167 7098 14191 7100
rect 14247 7098 14253 7100
rect 14007 7046 14009 7098
rect 14189 7046 14191 7098
rect 13945 7044 13951 7046
rect 14007 7044 14031 7046
rect 14087 7044 14111 7046
rect 14167 7044 14191 7046
rect 14247 7044 14253 7046
rect 13945 7035 14253 7044
rect 17788 7002 17816 7142
rect 17776 6996 17828 7002
rect 17776 6938 17828 6944
rect 18248 6866 18276 10639
rect 18328 10610 18380 10616
rect 18340 10266 18368 10610
rect 18328 10260 18380 10266
rect 18328 10202 18380 10208
rect 18328 8832 18380 8838
rect 18328 8774 18380 8780
rect 15384 6860 15436 6866
rect 15384 6802 15436 6808
rect 18236 6860 18288 6866
rect 18236 6802 18288 6808
rect 14648 6724 14700 6730
rect 14648 6666 14700 6672
rect 14660 6458 14688 6666
rect 14648 6452 14700 6458
rect 14648 6394 14700 6400
rect 14094 6352 14150 6361
rect 13728 6316 13780 6322
rect 14094 6287 14150 6296
rect 14556 6316 14608 6322
rect 13728 6258 13780 6264
rect 14108 6254 14136 6287
rect 14556 6258 14608 6264
rect 13176 6248 13228 6254
rect 13176 6190 13228 6196
rect 13360 6248 13412 6254
rect 13360 6190 13412 6196
rect 14096 6248 14148 6254
rect 14096 6190 14148 6196
rect 13188 5914 13216 6190
rect 13945 6012 14253 6021
rect 13945 6010 13951 6012
rect 14007 6010 14031 6012
rect 14087 6010 14111 6012
rect 14167 6010 14191 6012
rect 14247 6010 14253 6012
rect 14007 5958 14009 6010
rect 14189 5958 14191 6010
rect 13945 5956 13951 5958
rect 14007 5956 14031 5958
rect 14087 5956 14111 5958
rect 14167 5956 14191 5958
rect 14247 5956 14253 5958
rect 13945 5947 14253 5956
rect 13176 5908 13228 5914
rect 13176 5850 13228 5856
rect 14568 5778 14596 6258
rect 14660 6254 14688 6394
rect 15396 6390 15424 6802
rect 16948 6792 17000 6798
rect 16948 6734 17000 6740
rect 16544 6556 16852 6565
rect 16544 6554 16550 6556
rect 16606 6554 16630 6556
rect 16686 6554 16710 6556
rect 16766 6554 16790 6556
rect 16846 6554 16852 6556
rect 16606 6502 16608 6554
rect 16788 6502 16790 6554
rect 16544 6500 16550 6502
rect 16606 6500 16630 6502
rect 16686 6500 16710 6502
rect 16766 6500 16790 6502
rect 16846 6500 16852 6502
rect 16544 6491 16852 6500
rect 15384 6384 15436 6390
rect 15384 6326 15436 6332
rect 16960 6322 16988 6734
rect 16948 6316 17000 6322
rect 16948 6258 17000 6264
rect 14648 6248 14700 6254
rect 14648 6190 14700 6196
rect 14556 5772 14608 5778
rect 14556 5714 14608 5720
rect 13082 5672 13138 5681
rect 10968 5636 11020 5642
rect 13082 5607 13138 5616
rect 10968 5578 11020 5584
rect 11346 5468 11654 5477
rect 11346 5466 11352 5468
rect 11408 5466 11432 5468
rect 11488 5466 11512 5468
rect 11568 5466 11592 5468
rect 11648 5466 11654 5468
rect 11408 5414 11410 5466
rect 11590 5414 11592 5466
rect 11346 5412 11352 5414
rect 11408 5412 11432 5414
rect 11488 5412 11512 5414
rect 11568 5412 11592 5414
rect 11648 5412 11654 5414
rect 11346 5403 11654 5412
rect 16544 5468 16852 5477
rect 16544 5466 16550 5468
rect 16606 5466 16630 5468
rect 16686 5466 16710 5468
rect 16766 5466 16790 5468
rect 16846 5466 16852 5468
rect 16606 5414 16608 5466
rect 16788 5414 16790 5466
rect 16544 5412 16550 5414
rect 16606 5412 16630 5414
rect 16686 5412 16710 5414
rect 16766 5412 16790 5414
rect 16846 5412 16852 5414
rect 16544 5403 16852 5412
rect 8747 4924 9055 4933
rect 8747 4922 8753 4924
rect 8809 4922 8833 4924
rect 8889 4922 8913 4924
rect 8969 4922 8993 4924
rect 9049 4922 9055 4924
rect 8809 4870 8811 4922
rect 8991 4870 8993 4922
rect 8747 4868 8753 4870
rect 8809 4868 8833 4870
rect 8889 4868 8913 4870
rect 8969 4868 8993 4870
rect 9049 4868 9055 4870
rect 8747 4859 9055 4868
rect 13945 4924 14253 4933
rect 13945 4922 13951 4924
rect 14007 4922 14031 4924
rect 14087 4922 14111 4924
rect 14167 4922 14191 4924
rect 14247 4922 14253 4924
rect 14007 4870 14009 4922
rect 14189 4870 14191 4922
rect 13945 4868 13951 4870
rect 14007 4868 14031 4870
rect 14087 4868 14111 4870
rect 14167 4868 14191 4870
rect 14247 4868 14253 4870
rect 13945 4859 14253 4868
rect 11346 4380 11654 4389
rect 11346 4378 11352 4380
rect 11408 4378 11432 4380
rect 11488 4378 11512 4380
rect 11568 4378 11592 4380
rect 11648 4378 11654 4380
rect 11408 4326 11410 4378
rect 11590 4326 11592 4378
rect 11346 4324 11352 4326
rect 11408 4324 11432 4326
rect 11488 4324 11512 4326
rect 11568 4324 11592 4326
rect 11648 4324 11654 4326
rect 11346 4315 11654 4324
rect 16544 4380 16852 4389
rect 16544 4378 16550 4380
rect 16606 4378 16630 4380
rect 16686 4378 16710 4380
rect 16766 4378 16790 4380
rect 16846 4378 16852 4380
rect 16606 4326 16608 4378
rect 16788 4326 16790 4378
rect 16544 4324 16550 4326
rect 16606 4324 16630 4326
rect 16686 4324 16710 4326
rect 16766 4324 16790 4326
rect 16846 4324 16852 4326
rect 16544 4315 16852 4324
rect 18340 4010 18368 8774
rect 18432 7834 18460 10764
rect 18524 10062 18552 14282
rect 18604 13864 18656 13870
rect 18604 13806 18656 13812
rect 18616 12986 18644 13806
rect 18696 13320 18748 13326
rect 18696 13262 18748 13268
rect 18604 12980 18656 12986
rect 18604 12922 18656 12928
rect 18708 12442 18736 13262
rect 18696 12436 18748 12442
rect 18696 12378 18748 12384
rect 18696 11756 18748 11762
rect 18696 11698 18748 11704
rect 18602 11656 18658 11665
rect 18602 11591 18658 11600
rect 18616 11257 18644 11591
rect 18708 11354 18736 11698
rect 18696 11348 18748 11354
rect 18696 11290 18748 11296
rect 18800 11286 18828 16050
rect 18892 15434 18920 19314
rect 19536 19242 19564 19314
rect 19524 19236 19576 19242
rect 19524 19178 19576 19184
rect 19143 19068 19451 19077
rect 19143 19066 19149 19068
rect 19205 19066 19229 19068
rect 19285 19066 19309 19068
rect 19365 19066 19389 19068
rect 19445 19066 19451 19068
rect 19205 19014 19207 19066
rect 19387 19014 19389 19066
rect 19143 19012 19149 19014
rect 19205 19012 19229 19014
rect 19285 19012 19309 19014
rect 19365 19012 19389 19014
rect 19445 19012 19451 19014
rect 19143 19003 19451 19012
rect 19143 17980 19451 17989
rect 19143 17978 19149 17980
rect 19205 17978 19229 17980
rect 19285 17978 19309 17980
rect 19365 17978 19389 17980
rect 19445 17978 19451 17980
rect 19205 17926 19207 17978
rect 19387 17926 19389 17978
rect 19143 17924 19149 17926
rect 19205 17924 19229 17926
rect 19285 17924 19309 17926
rect 19365 17924 19389 17926
rect 19445 17924 19451 17926
rect 19143 17915 19451 17924
rect 19143 16892 19451 16901
rect 19143 16890 19149 16892
rect 19205 16890 19229 16892
rect 19285 16890 19309 16892
rect 19365 16890 19389 16892
rect 19445 16890 19451 16892
rect 19205 16838 19207 16890
rect 19387 16838 19389 16890
rect 19143 16836 19149 16838
rect 19205 16836 19229 16838
rect 19285 16836 19309 16838
rect 19365 16836 19389 16838
rect 19445 16836 19451 16838
rect 19143 16827 19451 16836
rect 19616 16652 19668 16658
rect 19616 16594 19668 16600
rect 19143 15804 19451 15813
rect 19143 15802 19149 15804
rect 19205 15802 19229 15804
rect 19285 15802 19309 15804
rect 19365 15802 19389 15804
rect 19445 15802 19451 15804
rect 19205 15750 19207 15802
rect 19387 15750 19389 15802
rect 19143 15748 19149 15750
rect 19205 15748 19229 15750
rect 19285 15748 19309 15750
rect 19365 15748 19389 15750
rect 19445 15748 19451 15750
rect 19143 15739 19451 15748
rect 18880 15428 18932 15434
rect 18880 15370 18932 15376
rect 18972 15020 19024 15026
rect 18972 14962 19024 14968
rect 19524 15020 19576 15026
rect 19524 14962 19576 14968
rect 18880 14068 18932 14074
rect 18880 14010 18932 14016
rect 18892 12442 18920 14010
rect 18984 14006 19012 14962
rect 19064 14952 19116 14958
rect 19064 14894 19116 14900
rect 19076 14618 19104 14894
rect 19143 14716 19451 14725
rect 19143 14714 19149 14716
rect 19205 14714 19229 14716
rect 19285 14714 19309 14716
rect 19365 14714 19389 14716
rect 19445 14714 19451 14716
rect 19205 14662 19207 14714
rect 19387 14662 19389 14714
rect 19143 14660 19149 14662
rect 19205 14660 19229 14662
rect 19285 14660 19309 14662
rect 19365 14660 19389 14662
rect 19445 14660 19451 14662
rect 19143 14651 19451 14660
rect 19064 14612 19116 14618
rect 19064 14554 19116 14560
rect 19064 14408 19116 14414
rect 19064 14350 19116 14356
rect 19076 14074 19104 14350
rect 19536 14278 19564 14962
rect 19524 14272 19576 14278
rect 19524 14214 19576 14220
rect 19064 14068 19116 14074
rect 19064 14010 19116 14016
rect 18972 14000 19024 14006
rect 18972 13942 19024 13948
rect 18972 13796 19024 13802
rect 18972 13738 19024 13744
rect 18984 13394 19012 13738
rect 19143 13628 19451 13637
rect 19143 13626 19149 13628
rect 19205 13626 19229 13628
rect 19285 13626 19309 13628
rect 19365 13626 19389 13628
rect 19445 13626 19451 13628
rect 19205 13574 19207 13626
rect 19387 13574 19389 13626
rect 19143 13572 19149 13574
rect 19205 13572 19229 13574
rect 19285 13572 19309 13574
rect 19365 13572 19389 13574
rect 19445 13572 19451 13574
rect 19143 13563 19451 13572
rect 18972 13388 19024 13394
rect 18972 13330 19024 13336
rect 18984 13297 19012 13330
rect 18970 13288 19026 13297
rect 18970 13223 19026 13232
rect 18972 12844 19024 12850
rect 18972 12786 19024 12792
rect 19524 12844 19576 12850
rect 19524 12786 19576 12792
rect 18880 12436 18932 12442
rect 18880 12378 18932 12384
rect 18880 12164 18932 12170
rect 18880 12106 18932 12112
rect 18892 11694 18920 12106
rect 18880 11688 18932 11694
rect 18880 11630 18932 11636
rect 18788 11280 18840 11286
rect 18602 11248 18658 11257
rect 18788 11222 18840 11228
rect 18602 11183 18658 11192
rect 18696 11212 18748 11218
rect 18616 11150 18644 11183
rect 18696 11154 18748 11160
rect 18604 11144 18656 11150
rect 18604 11086 18656 11092
rect 18708 10962 18736 11154
rect 18616 10934 18736 10962
rect 18512 10056 18564 10062
rect 18512 9998 18564 10004
rect 18512 9376 18564 9382
rect 18512 9318 18564 9324
rect 18524 8362 18552 9318
rect 18616 8838 18644 10934
rect 18892 10606 18920 11630
rect 18880 10600 18932 10606
rect 18880 10542 18932 10548
rect 18696 10532 18748 10538
rect 18696 10474 18748 10480
rect 18708 8838 18736 10474
rect 18880 10464 18932 10470
rect 18880 10406 18932 10412
rect 18788 10056 18840 10062
rect 18788 9998 18840 10004
rect 18604 8832 18656 8838
rect 18604 8774 18656 8780
rect 18696 8832 18748 8838
rect 18696 8774 18748 8780
rect 18708 8378 18736 8774
rect 18512 8356 18564 8362
rect 18512 8298 18564 8304
rect 18616 8350 18736 8378
rect 18432 7806 18552 7834
rect 18420 7744 18472 7750
rect 18420 7686 18472 7692
rect 18432 5370 18460 7686
rect 18524 6730 18552 7806
rect 18616 7750 18644 8350
rect 18696 8288 18748 8294
rect 18696 8230 18748 8236
rect 18708 7954 18736 8230
rect 18696 7948 18748 7954
rect 18696 7890 18748 7896
rect 18604 7744 18656 7750
rect 18604 7686 18656 7692
rect 18708 7342 18736 7890
rect 18800 7818 18828 9998
rect 18788 7812 18840 7818
rect 18788 7754 18840 7760
rect 18696 7336 18748 7342
rect 18696 7278 18748 7284
rect 18892 6769 18920 10406
rect 18984 9058 19012 12786
rect 19143 12540 19451 12549
rect 19143 12538 19149 12540
rect 19205 12538 19229 12540
rect 19285 12538 19309 12540
rect 19365 12538 19389 12540
rect 19445 12538 19451 12540
rect 19205 12486 19207 12538
rect 19387 12486 19389 12538
rect 19143 12484 19149 12486
rect 19205 12484 19229 12486
rect 19285 12484 19309 12486
rect 19365 12484 19389 12486
rect 19445 12484 19451 12486
rect 19143 12475 19451 12484
rect 19248 11824 19300 11830
rect 19248 11766 19300 11772
rect 19064 11688 19116 11694
rect 19064 11630 19116 11636
rect 19076 11218 19104 11630
rect 19260 11626 19288 11766
rect 19248 11620 19300 11626
rect 19248 11562 19300 11568
rect 19143 11452 19451 11461
rect 19143 11450 19149 11452
rect 19205 11450 19229 11452
rect 19285 11450 19309 11452
rect 19365 11450 19389 11452
rect 19445 11450 19451 11452
rect 19205 11398 19207 11450
rect 19387 11398 19389 11450
rect 19143 11396 19149 11398
rect 19205 11396 19229 11398
rect 19285 11396 19309 11398
rect 19365 11396 19389 11398
rect 19445 11396 19451 11398
rect 19143 11387 19451 11396
rect 19246 11248 19302 11257
rect 19064 11212 19116 11218
rect 19246 11183 19302 11192
rect 19064 11154 19116 11160
rect 19260 11082 19288 11183
rect 19248 11076 19300 11082
rect 19248 11018 19300 11024
rect 19432 11008 19484 11014
rect 19432 10950 19484 10956
rect 19444 10674 19472 10950
rect 19432 10668 19484 10674
rect 19432 10610 19484 10616
rect 19143 10364 19451 10373
rect 19143 10362 19149 10364
rect 19205 10362 19229 10364
rect 19285 10362 19309 10364
rect 19365 10362 19389 10364
rect 19445 10362 19451 10364
rect 19205 10310 19207 10362
rect 19387 10310 19389 10362
rect 19143 10308 19149 10310
rect 19205 10308 19229 10310
rect 19285 10308 19309 10310
rect 19365 10308 19389 10310
rect 19445 10308 19451 10310
rect 19143 10299 19451 10308
rect 19156 10260 19208 10266
rect 19156 10202 19208 10208
rect 19168 10146 19196 10202
rect 19432 10192 19484 10198
rect 19168 10140 19432 10146
rect 19168 10134 19484 10140
rect 19536 10146 19564 12786
rect 19628 12434 19656 16594
rect 19720 13734 19748 19790
rect 20260 19790 20312 19796
rect 19982 19751 20038 19760
rect 19800 19712 19852 19718
rect 19800 19654 19852 19660
rect 20168 19712 20220 19718
rect 20168 19654 20220 19660
rect 19812 19446 19840 19654
rect 19984 19508 20036 19514
rect 19984 19450 20036 19456
rect 19800 19440 19852 19446
rect 19800 19382 19852 19388
rect 19996 19378 20024 19450
rect 19984 19372 20036 19378
rect 19984 19314 20036 19320
rect 19892 18216 19944 18222
rect 19892 18158 19944 18164
rect 19800 17672 19852 17678
rect 19800 17614 19852 17620
rect 19812 16998 19840 17614
rect 19904 17338 19932 18158
rect 19892 17332 19944 17338
rect 19892 17274 19944 17280
rect 19800 16992 19852 16998
rect 19800 16934 19852 16940
rect 19800 14476 19852 14482
rect 19800 14418 19852 14424
rect 19812 13938 19840 14418
rect 19800 13932 19852 13938
rect 19800 13874 19852 13880
rect 19708 13728 19760 13734
rect 19708 13670 19760 13676
rect 19996 12434 20024 19314
rect 20180 19174 20208 19654
rect 20272 19514 20300 19790
rect 20720 19780 20772 19786
rect 20720 19722 20772 19728
rect 20260 19508 20312 19514
rect 20260 19450 20312 19456
rect 20168 19168 20220 19174
rect 20168 19110 20220 19116
rect 20628 18760 20680 18766
rect 20626 18728 20628 18737
rect 20680 18728 20682 18737
rect 20626 18663 20682 18672
rect 20352 18624 20404 18630
rect 20352 18566 20404 18572
rect 20260 16108 20312 16114
rect 20260 16050 20312 16056
rect 20168 15904 20220 15910
rect 20168 15846 20220 15852
rect 20180 15609 20208 15846
rect 20272 15706 20300 16050
rect 20260 15700 20312 15706
rect 20260 15642 20312 15648
rect 20166 15600 20222 15609
rect 20166 15535 20222 15544
rect 20076 14272 20128 14278
rect 20076 14214 20128 14220
rect 20088 14074 20116 14214
rect 20076 14068 20128 14074
rect 20076 14010 20128 14016
rect 20260 12776 20312 12782
rect 20260 12718 20312 12724
rect 19628 12406 19932 12434
rect 19996 12406 20116 12434
rect 19616 12368 19668 12374
rect 19616 12310 19668 12316
rect 19628 10742 19656 12310
rect 19708 12096 19760 12102
rect 19708 12038 19760 12044
rect 19720 10810 19748 12038
rect 19800 11688 19852 11694
rect 19800 11630 19852 11636
rect 19812 11218 19840 11630
rect 19800 11212 19852 11218
rect 19800 11154 19852 11160
rect 19708 10804 19760 10810
rect 19708 10746 19760 10752
rect 19616 10736 19668 10742
rect 19616 10678 19668 10684
rect 19812 10266 19840 11154
rect 19904 11014 19932 12406
rect 19984 11688 20036 11694
rect 19984 11630 20036 11636
rect 19996 11150 20024 11630
rect 19984 11144 20036 11150
rect 19984 11086 20036 11092
rect 19892 11008 19944 11014
rect 19892 10950 19944 10956
rect 19892 10804 19944 10810
rect 19892 10746 19944 10752
rect 19800 10260 19852 10266
rect 19800 10202 19852 10208
rect 19168 10118 19472 10134
rect 19536 10118 19840 10146
rect 19524 10056 19576 10062
rect 19524 9998 19576 10004
rect 19708 10056 19760 10062
rect 19708 9998 19760 10004
rect 19536 9722 19564 9998
rect 19616 9920 19668 9926
rect 19616 9862 19668 9868
rect 19524 9716 19576 9722
rect 19524 9658 19576 9664
rect 19628 9450 19656 9862
rect 19616 9444 19668 9450
rect 19616 9386 19668 9392
rect 19143 9276 19451 9285
rect 19143 9274 19149 9276
rect 19205 9274 19229 9276
rect 19285 9274 19309 9276
rect 19365 9274 19389 9276
rect 19445 9274 19451 9276
rect 19205 9222 19207 9274
rect 19387 9222 19389 9274
rect 19143 9220 19149 9222
rect 19205 9220 19229 9222
rect 19285 9220 19309 9222
rect 19365 9220 19389 9222
rect 19445 9220 19451 9222
rect 19143 9211 19451 9220
rect 19156 9172 19208 9178
rect 19156 9114 19208 9120
rect 19340 9172 19392 9178
rect 19340 9114 19392 9120
rect 19168 9058 19196 9114
rect 18984 9030 19196 9058
rect 19248 9036 19300 9042
rect 19248 8978 19300 8984
rect 18972 8832 19024 8838
rect 18972 8774 19024 8780
rect 18984 8566 19012 8774
rect 19260 8673 19288 8978
rect 19352 8974 19380 9114
rect 19720 9058 19748 9998
rect 19444 9030 19748 9058
rect 19340 8968 19392 8974
rect 19340 8910 19392 8916
rect 19444 8906 19472 9030
rect 19432 8900 19484 8906
rect 19432 8842 19484 8848
rect 19246 8664 19302 8673
rect 19246 8599 19302 8608
rect 18972 8560 19024 8566
rect 18972 8502 19024 8508
rect 19248 8492 19300 8498
rect 19248 8434 19300 8440
rect 19260 8401 19288 8434
rect 19246 8392 19302 8401
rect 19444 8362 19472 8842
rect 19524 8832 19576 8838
rect 19524 8774 19576 8780
rect 19536 8498 19564 8774
rect 19524 8492 19576 8498
rect 19524 8434 19576 8440
rect 19616 8424 19668 8430
rect 19616 8366 19668 8372
rect 19246 8327 19302 8336
rect 19432 8356 19484 8362
rect 19432 8298 19484 8304
rect 19143 8188 19451 8197
rect 19143 8186 19149 8188
rect 19205 8186 19229 8188
rect 19285 8186 19309 8188
rect 19365 8186 19389 8188
rect 19445 8186 19451 8188
rect 19205 8134 19207 8186
rect 19387 8134 19389 8186
rect 19143 8132 19149 8134
rect 19205 8132 19229 8134
rect 19285 8132 19309 8134
rect 19365 8132 19389 8134
rect 19445 8132 19451 8134
rect 19143 8123 19451 8132
rect 19628 8090 19656 8366
rect 19616 8084 19668 8090
rect 19616 8026 19668 8032
rect 19143 7100 19451 7109
rect 19143 7098 19149 7100
rect 19205 7098 19229 7100
rect 19285 7098 19309 7100
rect 19365 7098 19389 7100
rect 19445 7098 19451 7100
rect 19205 7046 19207 7098
rect 19387 7046 19389 7098
rect 19143 7044 19149 7046
rect 19205 7044 19229 7046
rect 19285 7044 19309 7046
rect 19365 7044 19389 7046
rect 19445 7044 19451 7046
rect 19143 7035 19451 7044
rect 18878 6760 18934 6769
rect 18512 6724 18564 6730
rect 18878 6695 18934 6704
rect 18512 6666 18564 6672
rect 19812 6662 19840 10118
rect 19904 9042 19932 10746
rect 20088 10674 20116 12406
rect 20272 12238 20300 12718
rect 20260 12232 20312 12238
rect 20260 12174 20312 12180
rect 20168 11552 20220 11558
rect 20168 11494 20220 11500
rect 20180 11354 20208 11494
rect 20168 11348 20220 11354
rect 20168 11290 20220 11296
rect 20364 11082 20392 18566
rect 20536 18284 20588 18290
rect 20536 18226 20588 18232
rect 20548 17882 20576 18226
rect 20732 18154 20760 19722
rect 20916 19514 20944 20839
rect 21192 19990 21220 22200
rect 21546 21312 21602 21321
rect 21546 21247 21602 21256
rect 21364 20460 21416 20466
rect 21364 20402 21416 20408
rect 21180 19984 21232 19990
rect 21180 19926 21232 19932
rect 20996 19848 21048 19854
rect 20996 19790 21048 19796
rect 20904 19508 20956 19514
rect 20904 19450 20956 19456
rect 20904 19372 20956 19378
rect 20904 19314 20956 19320
rect 20812 19236 20864 19242
rect 20812 19178 20864 19184
rect 20824 18766 20852 19178
rect 20916 18970 20944 19314
rect 20904 18964 20956 18970
rect 20904 18906 20956 18912
rect 20812 18760 20864 18766
rect 20812 18702 20864 18708
rect 20720 18148 20772 18154
rect 20720 18090 20772 18096
rect 20536 17876 20588 17882
rect 20536 17818 20588 17824
rect 20628 17672 20680 17678
rect 20628 17614 20680 17620
rect 20536 17196 20588 17202
rect 20536 17138 20588 17144
rect 20548 16250 20576 17138
rect 20640 16794 20668 17614
rect 20628 16788 20680 16794
rect 20628 16730 20680 16736
rect 20812 16584 20864 16590
rect 20812 16526 20864 16532
rect 20536 16244 20588 16250
rect 20536 16186 20588 16192
rect 20720 15428 20772 15434
rect 20720 15370 20772 15376
rect 20732 15162 20760 15370
rect 20720 15156 20772 15162
rect 20720 15098 20772 15104
rect 20628 14408 20680 14414
rect 20628 14350 20680 14356
rect 20534 12200 20590 12209
rect 20534 12135 20536 12144
rect 20588 12135 20590 12144
rect 20536 12106 20588 12112
rect 20548 11898 20576 12106
rect 20536 11892 20588 11898
rect 20536 11834 20588 11840
rect 20352 11076 20404 11082
rect 20352 11018 20404 11024
rect 20536 11076 20588 11082
rect 20536 11018 20588 11024
rect 19984 10668 20036 10674
rect 19984 10610 20036 10616
rect 20076 10668 20128 10674
rect 20076 10610 20128 10616
rect 19996 10266 20024 10610
rect 19984 10260 20036 10266
rect 19984 10202 20036 10208
rect 20548 10169 20576 11018
rect 20640 10810 20668 14350
rect 20824 13274 20852 16526
rect 21008 16454 21036 19790
rect 21088 19508 21140 19514
rect 21088 19450 21140 19456
rect 21100 19281 21128 19450
rect 21272 19372 21324 19378
rect 21272 19314 21324 19320
rect 21086 19272 21142 19281
rect 21086 19207 21142 19216
rect 21284 18902 21312 19314
rect 21272 18896 21324 18902
rect 21272 18838 21324 18844
rect 21272 18760 21324 18766
rect 21272 18702 21324 18708
rect 21284 18426 21312 18702
rect 21272 18420 21324 18426
rect 21272 18362 21324 18368
rect 21180 18284 21232 18290
rect 21180 18226 21232 18232
rect 21086 17640 21142 17649
rect 21086 17575 21142 17584
rect 21100 17542 21128 17575
rect 21088 17536 21140 17542
rect 21088 17478 21140 17484
rect 20996 16448 21048 16454
rect 20996 16390 21048 16396
rect 21192 16250 21220 18226
rect 21376 18193 21404 20402
rect 21454 19816 21510 19825
rect 21454 19751 21510 19760
rect 21468 19718 21496 19751
rect 21456 19712 21508 19718
rect 21456 19654 21508 19660
rect 21456 19168 21508 19174
rect 21456 19110 21508 19116
rect 21468 18873 21496 19110
rect 21560 18970 21588 21247
rect 21742 20700 22050 20709
rect 21742 20698 21748 20700
rect 21804 20698 21828 20700
rect 21884 20698 21908 20700
rect 21964 20698 21988 20700
rect 22044 20698 22050 20700
rect 21804 20646 21806 20698
rect 21986 20646 21988 20698
rect 21742 20644 21748 20646
rect 21804 20644 21828 20646
rect 21884 20644 21908 20646
rect 21964 20644 21988 20646
rect 22044 20644 22050 20646
rect 21742 20635 22050 20644
rect 21742 19612 22050 19621
rect 21742 19610 21748 19612
rect 21804 19610 21828 19612
rect 21884 19610 21908 19612
rect 21964 19610 21988 19612
rect 22044 19610 22050 19612
rect 21804 19558 21806 19610
rect 21986 19558 21988 19610
rect 21742 19556 21748 19558
rect 21804 19556 21828 19558
rect 21884 19556 21908 19558
rect 21964 19556 21988 19558
rect 22044 19556 22050 19558
rect 21742 19547 22050 19556
rect 21548 18964 21600 18970
rect 21548 18906 21600 18912
rect 21454 18864 21510 18873
rect 21454 18799 21510 18808
rect 22284 18828 22336 18834
rect 22284 18770 22336 18776
rect 21456 18624 21508 18630
rect 21456 18566 21508 18572
rect 21468 18329 21496 18566
rect 21742 18524 22050 18533
rect 21742 18522 21748 18524
rect 21804 18522 21828 18524
rect 21884 18522 21908 18524
rect 21964 18522 21988 18524
rect 22044 18522 22050 18524
rect 21804 18470 21806 18522
rect 21986 18470 21988 18522
rect 21742 18468 21748 18470
rect 21804 18468 21828 18470
rect 21884 18468 21908 18470
rect 21964 18468 21988 18470
rect 22044 18468 22050 18470
rect 21742 18459 22050 18468
rect 21454 18320 21510 18329
rect 21454 18255 21510 18264
rect 21362 18184 21418 18193
rect 21362 18119 21418 18128
rect 21456 18080 21508 18086
rect 21454 18048 21456 18057
rect 21508 18048 21510 18057
rect 21454 17983 21510 17992
rect 21272 17672 21324 17678
rect 21272 17614 21324 17620
rect 21180 16244 21232 16250
rect 21180 16186 21232 16192
rect 20904 16108 20956 16114
rect 20904 16050 20956 16056
rect 20916 15162 20944 16050
rect 21086 16008 21142 16017
rect 21086 15943 21088 15952
rect 21140 15943 21142 15952
rect 21088 15914 21140 15920
rect 21284 15706 21312 17614
rect 21456 17536 21508 17542
rect 21456 17478 21508 17484
rect 21468 17241 21496 17478
rect 21742 17436 22050 17445
rect 21742 17434 21748 17436
rect 21804 17434 21828 17436
rect 21884 17434 21908 17436
rect 21964 17434 21988 17436
rect 22044 17434 22050 17436
rect 21804 17382 21806 17434
rect 21986 17382 21988 17434
rect 21742 17380 21748 17382
rect 21804 17380 21828 17382
rect 21884 17380 21908 17382
rect 21964 17380 21988 17382
rect 22044 17380 22050 17382
rect 21742 17371 22050 17380
rect 21454 17232 21510 17241
rect 21454 17167 21510 17176
rect 21456 16992 21508 16998
rect 21456 16934 21508 16940
rect 21468 16833 21496 16934
rect 21454 16824 21510 16833
rect 21454 16759 21510 16768
rect 21454 16552 21510 16561
rect 21454 16487 21510 16496
rect 21468 16454 21496 16487
rect 21456 16448 21508 16454
rect 21456 16390 21508 16396
rect 21742 16348 22050 16357
rect 21742 16346 21748 16348
rect 21804 16346 21828 16348
rect 21884 16346 21908 16348
rect 21964 16346 21988 16348
rect 22044 16346 22050 16348
rect 21804 16294 21806 16346
rect 21986 16294 21988 16346
rect 21742 16292 21748 16294
rect 21804 16292 21828 16294
rect 21884 16292 21908 16294
rect 21964 16292 21988 16294
rect 22044 16292 22050 16294
rect 21742 16283 22050 16292
rect 21364 16108 21416 16114
rect 21364 16050 21416 16056
rect 21272 15700 21324 15706
rect 21272 15642 21324 15648
rect 20996 15496 21048 15502
rect 20996 15438 21048 15444
rect 20904 15156 20956 15162
rect 20904 15098 20956 15104
rect 20904 15020 20956 15026
rect 20904 14962 20956 14968
rect 20732 13246 20852 13274
rect 20732 12986 20760 13246
rect 20812 13184 20864 13190
rect 20812 13126 20864 13132
rect 20720 12980 20772 12986
rect 20720 12922 20772 12928
rect 20718 12744 20774 12753
rect 20718 12679 20720 12688
rect 20772 12679 20774 12688
rect 20720 12650 20772 12656
rect 20824 11830 20852 13126
rect 20812 11824 20864 11830
rect 20812 11766 20864 11772
rect 20812 11348 20864 11354
rect 20812 11290 20864 11296
rect 20824 10810 20852 11290
rect 20628 10804 20680 10810
rect 20628 10746 20680 10752
rect 20812 10804 20864 10810
rect 20812 10746 20864 10752
rect 20812 10600 20864 10606
rect 20812 10542 20864 10548
rect 20720 10532 20772 10538
rect 20720 10474 20772 10480
rect 20628 10464 20680 10470
rect 20628 10406 20680 10412
rect 20534 10160 20590 10169
rect 20640 10130 20668 10406
rect 20534 10095 20590 10104
rect 20628 10124 20680 10130
rect 20628 10066 20680 10072
rect 20732 10033 20760 10474
rect 20718 10024 20774 10033
rect 20444 9988 20496 9994
rect 20444 9930 20496 9936
rect 20628 9988 20680 9994
rect 20718 9959 20774 9968
rect 20628 9930 20680 9936
rect 20168 9920 20220 9926
rect 20168 9862 20220 9868
rect 20180 9722 20208 9862
rect 20168 9716 20220 9722
rect 20168 9658 20220 9664
rect 19984 9172 20036 9178
rect 19984 9114 20036 9120
rect 19892 9036 19944 9042
rect 19892 8978 19944 8984
rect 19996 8974 20024 9114
rect 20168 9104 20220 9110
rect 20168 9046 20220 9052
rect 19984 8968 20036 8974
rect 19984 8910 20036 8916
rect 20074 8936 20130 8945
rect 20074 8871 20130 8880
rect 20088 8838 20116 8871
rect 20076 8832 20128 8838
rect 19982 8800 20038 8809
rect 20076 8774 20128 8780
rect 19982 8735 20038 8744
rect 19996 7750 20024 8735
rect 19984 7744 20036 7750
rect 19984 7686 20036 7692
rect 19800 6656 19852 6662
rect 19800 6598 19852 6604
rect 19143 6012 19451 6021
rect 19143 6010 19149 6012
rect 19205 6010 19229 6012
rect 19285 6010 19309 6012
rect 19365 6010 19389 6012
rect 19445 6010 19451 6012
rect 19205 5958 19207 6010
rect 19387 5958 19389 6010
rect 19143 5956 19149 5958
rect 19205 5956 19229 5958
rect 19285 5956 19309 5958
rect 19365 5956 19389 5958
rect 19445 5956 19451 5958
rect 19143 5947 19451 5956
rect 18420 5364 18472 5370
rect 18420 5306 18472 5312
rect 19143 4924 19451 4933
rect 19143 4922 19149 4924
rect 19205 4922 19229 4924
rect 19285 4922 19309 4924
rect 19365 4922 19389 4924
rect 19445 4922 19451 4924
rect 19205 4870 19207 4922
rect 19387 4870 19389 4922
rect 19143 4868 19149 4870
rect 19205 4868 19229 4870
rect 19285 4868 19309 4870
rect 19365 4868 19389 4870
rect 19445 4868 19451 4870
rect 19143 4859 19451 4868
rect 18328 4004 18380 4010
rect 18328 3946 18380 3952
rect 8747 3836 9055 3845
rect 8747 3834 8753 3836
rect 8809 3834 8833 3836
rect 8889 3834 8913 3836
rect 8969 3834 8993 3836
rect 9049 3834 9055 3836
rect 8809 3782 8811 3834
rect 8991 3782 8993 3834
rect 8747 3780 8753 3782
rect 8809 3780 8833 3782
rect 8889 3780 8913 3782
rect 8969 3780 8993 3782
rect 9049 3780 9055 3782
rect 8747 3771 9055 3780
rect 13945 3836 14253 3845
rect 13945 3834 13951 3836
rect 14007 3834 14031 3836
rect 14087 3834 14111 3836
rect 14167 3834 14191 3836
rect 14247 3834 14253 3836
rect 14007 3782 14009 3834
rect 14189 3782 14191 3834
rect 13945 3780 13951 3782
rect 14007 3780 14031 3782
rect 14087 3780 14111 3782
rect 14167 3780 14191 3782
rect 14247 3780 14253 3782
rect 13945 3771 14253 3780
rect 19143 3836 19451 3845
rect 19143 3834 19149 3836
rect 19205 3834 19229 3836
rect 19285 3834 19309 3836
rect 19365 3834 19389 3836
rect 19445 3834 19451 3836
rect 19205 3782 19207 3834
rect 19387 3782 19389 3834
rect 19143 3780 19149 3782
rect 19205 3780 19229 3782
rect 19285 3780 19309 3782
rect 19365 3780 19389 3782
rect 19445 3780 19451 3782
rect 19143 3771 19451 3780
rect 11346 3292 11654 3301
rect 11346 3290 11352 3292
rect 11408 3290 11432 3292
rect 11488 3290 11512 3292
rect 11568 3290 11592 3292
rect 11648 3290 11654 3292
rect 11408 3238 11410 3290
rect 11590 3238 11592 3290
rect 11346 3236 11352 3238
rect 11408 3236 11432 3238
rect 11488 3236 11512 3238
rect 11568 3236 11592 3238
rect 11648 3236 11654 3238
rect 11346 3227 11654 3236
rect 16544 3292 16852 3301
rect 16544 3290 16550 3292
rect 16606 3290 16630 3292
rect 16686 3290 16710 3292
rect 16766 3290 16790 3292
rect 16846 3290 16852 3292
rect 16606 3238 16608 3290
rect 16788 3238 16790 3290
rect 16544 3236 16550 3238
rect 16606 3236 16630 3238
rect 16686 3236 16710 3238
rect 16766 3236 16790 3238
rect 16846 3236 16852 3238
rect 16544 3227 16852 3236
rect 8668 3052 8720 3058
rect 8668 2994 8720 3000
rect 16120 3052 16172 3058
rect 16120 2994 16172 3000
rect 8680 2650 8708 2994
rect 8747 2748 9055 2757
rect 8747 2746 8753 2748
rect 8809 2746 8833 2748
rect 8889 2746 8913 2748
rect 8969 2746 8993 2748
rect 9049 2746 9055 2748
rect 8809 2694 8811 2746
rect 8991 2694 8993 2746
rect 8747 2692 8753 2694
rect 8809 2692 8833 2694
rect 8889 2692 8913 2694
rect 8969 2692 8993 2694
rect 9049 2692 9055 2694
rect 8747 2683 9055 2692
rect 13945 2748 14253 2757
rect 13945 2746 13951 2748
rect 14007 2746 14031 2748
rect 14087 2746 14111 2748
rect 14167 2746 14191 2748
rect 14247 2746 14253 2748
rect 14007 2694 14009 2746
rect 14189 2694 14191 2746
rect 13945 2692 13951 2694
rect 14007 2692 14031 2694
rect 14087 2692 14111 2694
rect 14167 2692 14191 2694
rect 14247 2692 14253 2694
rect 13945 2683 14253 2692
rect 16132 2650 16160 2994
rect 16854 2952 16910 2961
rect 19996 2922 20024 7686
rect 16854 2887 16856 2896
rect 16908 2887 16910 2896
rect 19984 2916 20036 2922
rect 16856 2858 16908 2864
rect 19984 2858 20036 2864
rect 20088 2774 20116 8774
rect 20180 7954 20208 9046
rect 20352 8492 20404 8498
rect 20352 8434 20404 8440
rect 20258 7984 20314 7993
rect 20168 7948 20220 7954
rect 20258 7919 20314 7928
rect 20168 7890 20220 7896
rect 20272 7750 20300 7919
rect 20260 7744 20312 7750
rect 20260 7686 20312 7692
rect 20272 2854 20300 7686
rect 20364 7478 20392 8434
rect 20456 8430 20484 9930
rect 20536 9920 20588 9926
rect 20536 9862 20588 9868
rect 20548 9722 20576 9862
rect 20536 9716 20588 9722
rect 20536 9658 20588 9664
rect 20640 9178 20668 9930
rect 20824 9674 20852 10542
rect 20732 9646 20852 9674
rect 20628 9172 20680 9178
rect 20628 9114 20680 9120
rect 20732 9110 20760 9646
rect 20812 9444 20864 9450
rect 20812 9386 20864 9392
rect 20720 9104 20772 9110
rect 20720 9046 20772 9052
rect 20628 8968 20680 8974
rect 20628 8910 20680 8916
rect 20536 8900 20588 8906
rect 20536 8842 20588 8848
rect 20548 8430 20576 8842
rect 20640 8537 20668 8910
rect 20824 8634 20852 9386
rect 20812 8628 20864 8634
rect 20812 8570 20864 8576
rect 20626 8528 20682 8537
rect 20626 8463 20682 8472
rect 20444 8424 20496 8430
rect 20444 8366 20496 8372
rect 20536 8424 20588 8430
rect 20536 8366 20588 8372
rect 20352 7472 20404 7478
rect 20352 7414 20404 7420
rect 20364 3738 20392 7414
rect 20352 3732 20404 3738
rect 20352 3674 20404 3680
rect 20456 3194 20484 8366
rect 20640 8090 20668 8463
rect 20628 8084 20680 8090
rect 20628 8026 20680 8032
rect 20916 7546 20944 14962
rect 21008 14618 21036 15438
rect 21180 14816 21232 14822
rect 21180 14758 21232 14764
rect 20996 14612 21048 14618
rect 20996 14554 21048 14560
rect 20996 14408 21048 14414
rect 20996 14350 21048 14356
rect 21086 14376 21142 14385
rect 21008 13530 21036 14350
rect 21086 14311 21142 14320
rect 21100 14278 21128 14311
rect 21088 14272 21140 14278
rect 21088 14214 21140 14220
rect 20996 13524 21048 13530
rect 20996 13466 21048 13472
rect 20994 13424 21050 13433
rect 20994 13359 21050 13368
rect 21008 12986 21036 13359
rect 20996 12980 21048 12986
rect 20996 12922 21048 12928
rect 21088 12844 21140 12850
rect 21088 12786 21140 12792
rect 21100 12345 21128 12786
rect 21086 12336 21142 12345
rect 21086 12271 21142 12280
rect 21088 11552 21140 11558
rect 21088 11494 21140 11500
rect 20996 11144 21048 11150
rect 20994 11112 20996 11121
rect 21048 11112 21050 11121
rect 21100 11082 21128 11494
rect 21192 11354 21220 14758
rect 21272 13932 21324 13938
rect 21272 13874 21324 13880
rect 21180 11348 21232 11354
rect 21180 11290 21232 11296
rect 21180 11212 21232 11218
rect 21180 11154 21232 11160
rect 20994 11047 21050 11056
rect 21088 11076 21140 11082
rect 21088 11018 21140 11024
rect 21100 10713 21128 11018
rect 21086 10704 21142 10713
rect 21086 10639 21142 10648
rect 20994 9072 21050 9081
rect 20994 9007 20996 9016
rect 21048 9007 21050 9016
rect 20996 8978 21048 8984
rect 20996 7880 21048 7886
rect 20996 7822 21048 7828
rect 20904 7540 20956 7546
rect 20904 7482 20956 7488
rect 20626 7440 20682 7449
rect 20536 7404 20588 7410
rect 20626 7375 20682 7384
rect 20536 7346 20588 7352
rect 20548 6390 20576 7346
rect 20640 6866 20668 7375
rect 20720 7336 20772 7342
rect 20720 7278 20772 7284
rect 20732 7041 20760 7278
rect 20718 7032 20774 7041
rect 20718 6967 20774 6976
rect 20628 6860 20680 6866
rect 20628 6802 20680 6808
rect 20812 6792 20864 6798
rect 20810 6760 20812 6769
rect 20864 6760 20866 6769
rect 20810 6695 20866 6704
rect 20628 6656 20680 6662
rect 20628 6598 20680 6604
rect 20640 6458 20668 6598
rect 20628 6452 20680 6458
rect 20628 6394 20680 6400
rect 20536 6384 20588 6390
rect 20536 6326 20588 6332
rect 20720 6248 20772 6254
rect 20718 6216 20720 6225
rect 20772 6216 20774 6225
rect 20718 6151 20774 6160
rect 21008 4690 21036 7822
rect 21088 7812 21140 7818
rect 21088 7754 21140 7760
rect 20996 4684 21048 4690
rect 20996 4626 21048 4632
rect 20720 4616 20772 4622
rect 20720 4558 20772 4564
rect 20732 4185 20760 4558
rect 21100 4282 21128 7754
rect 21192 6361 21220 11154
rect 21284 10266 21312 13874
rect 21376 13530 21404 16050
rect 21456 15904 21508 15910
rect 21456 15846 21508 15852
rect 21468 15609 21496 15846
rect 21548 15700 21600 15706
rect 21548 15642 21600 15648
rect 21454 15600 21510 15609
rect 21454 15535 21510 15544
rect 21560 15065 21588 15642
rect 21640 15632 21692 15638
rect 21640 15574 21692 15580
rect 21546 15056 21602 15065
rect 21546 14991 21602 15000
rect 21456 14816 21508 14822
rect 21454 14784 21456 14793
rect 21508 14784 21510 14793
rect 21454 14719 21510 14728
rect 21456 14272 21508 14278
rect 21456 14214 21508 14220
rect 21468 13977 21496 14214
rect 21454 13968 21510 13977
rect 21454 13903 21510 13912
rect 21548 13796 21600 13802
rect 21548 13738 21600 13744
rect 21456 13728 21508 13734
rect 21456 13670 21508 13676
rect 21468 13569 21496 13670
rect 21454 13560 21510 13569
rect 21364 13524 21416 13530
rect 21454 13495 21510 13504
rect 21364 13466 21416 13472
rect 21364 13388 21416 13394
rect 21364 13330 21416 13336
rect 21376 11898 21404 13330
rect 21560 13326 21588 13738
rect 21548 13320 21600 13326
rect 21546 13288 21548 13297
rect 21600 13288 21602 13297
rect 21546 13223 21602 13232
rect 21652 13190 21680 15574
rect 22100 15428 22152 15434
rect 22100 15370 22152 15376
rect 21742 15260 22050 15269
rect 21742 15258 21748 15260
rect 21804 15258 21828 15260
rect 21884 15258 21908 15260
rect 21964 15258 21988 15260
rect 22044 15258 22050 15260
rect 21804 15206 21806 15258
rect 21986 15206 21988 15258
rect 21742 15204 21748 15206
rect 21804 15204 21828 15206
rect 21884 15204 21908 15206
rect 21964 15204 21988 15206
rect 22044 15204 22050 15206
rect 21742 15195 22050 15204
rect 21742 14172 22050 14181
rect 21742 14170 21748 14172
rect 21804 14170 21828 14172
rect 21884 14170 21908 14172
rect 21964 14170 21988 14172
rect 22044 14170 22050 14172
rect 21804 14118 21806 14170
rect 21986 14118 21988 14170
rect 21742 14116 21748 14118
rect 21804 14116 21828 14118
rect 21884 14116 21908 14118
rect 21964 14116 21988 14118
rect 22044 14116 22050 14118
rect 21742 14107 22050 14116
rect 21640 13184 21692 13190
rect 21640 13126 21692 13132
rect 21742 13084 22050 13093
rect 21742 13082 21748 13084
rect 21804 13082 21828 13084
rect 21884 13082 21908 13084
rect 21964 13082 21988 13084
rect 22044 13082 22050 13084
rect 21804 13030 21806 13082
rect 21986 13030 21988 13082
rect 21742 13028 21748 13030
rect 21804 13028 21828 13030
rect 21884 13028 21908 13030
rect 21964 13028 21988 13030
rect 22044 13028 22050 13030
rect 21742 13019 22050 13028
rect 22112 12968 22140 15370
rect 21652 12940 22140 12968
rect 21456 12844 21508 12850
rect 21456 12786 21508 12792
rect 21468 12753 21496 12786
rect 21454 12744 21510 12753
rect 21454 12679 21510 12688
rect 21468 12374 21496 12679
rect 21456 12368 21508 12374
rect 21456 12310 21508 12316
rect 21456 12164 21508 12170
rect 21456 12106 21508 12112
rect 21364 11892 21416 11898
rect 21364 11834 21416 11840
rect 21468 11801 21496 12106
rect 21454 11792 21510 11801
rect 21454 11727 21510 11736
rect 21548 11756 21600 11762
rect 21548 11698 21600 11704
rect 21364 11688 21416 11694
rect 21364 11630 21416 11636
rect 21376 10962 21404 11630
rect 21456 11620 21508 11626
rect 21456 11562 21508 11568
rect 21468 11150 21496 11562
rect 21560 11529 21588 11698
rect 21546 11520 21602 11529
rect 21546 11455 21602 11464
rect 21456 11144 21508 11150
rect 21454 11112 21456 11121
rect 21508 11112 21510 11121
rect 21454 11047 21510 11056
rect 21376 10934 21496 10962
rect 21468 10674 21496 10934
rect 21456 10668 21508 10674
rect 21456 10610 21508 10616
rect 21362 10568 21418 10577
rect 21362 10503 21418 10512
rect 21376 10266 21404 10503
rect 21468 10305 21496 10610
rect 21454 10296 21510 10305
rect 21272 10260 21324 10266
rect 21272 10202 21324 10208
rect 21364 10260 21416 10266
rect 21454 10231 21510 10240
rect 21364 10202 21416 10208
rect 21456 10056 21508 10062
rect 21456 9998 21508 10004
rect 21468 9489 21496 9998
rect 21652 9586 21680 12940
rect 22296 12730 22324 18770
rect 22376 16176 22428 16182
rect 22376 16118 22428 16124
rect 22112 12702 22324 12730
rect 22112 12442 22140 12702
rect 22100 12436 22152 12442
rect 22100 12378 22152 12384
rect 21742 11996 22050 12005
rect 21742 11994 21748 11996
rect 21804 11994 21828 11996
rect 21884 11994 21908 11996
rect 21964 11994 21988 11996
rect 22044 11994 22050 11996
rect 21804 11942 21806 11994
rect 21986 11942 21988 11994
rect 21742 11940 21748 11942
rect 21804 11940 21828 11942
rect 21884 11940 21908 11942
rect 21964 11940 21988 11942
rect 22044 11940 22050 11942
rect 21742 11931 22050 11940
rect 21742 10908 22050 10917
rect 21742 10906 21748 10908
rect 21804 10906 21828 10908
rect 21884 10906 21908 10908
rect 21964 10906 21988 10908
rect 22044 10906 22050 10908
rect 21804 10854 21806 10906
rect 21986 10854 21988 10906
rect 21742 10852 21748 10854
rect 21804 10852 21828 10854
rect 21884 10852 21908 10854
rect 21964 10852 21988 10854
rect 22044 10852 22050 10854
rect 21742 10843 22050 10852
rect 21742 9820 22050 9829
rect 21742 9818 21748 9820
rect 21804 9818 21828 9820
rect 21884 9818 21908 9820
rect 21964 9818 21988 9820
rect 22044 9818 22050 9820
rect 21804 9766 21806 9818
rect 21986 9766 21988 9818
rect 21742 9764 21748 9766
rect 21804 9764 21828 9766
rect 21884 9764 21908 9766
rect 21964 9764 21988 9766
rect 22044 9764 22050 9766
rect 21742 9755 22050 9764
rect 21640 9580 21692 9586
rect 21640 9522 21692 9528
rect 21548 9512 21600 9518
rect 21454 9480 21510 9489
rect 21548 9454 21600 9460
rect 21454 9415 21510 9424
rect 21560 9081 21588 9454
rect 21546 9072 21602 9081
rect 21546 9007 21602 9016
rect 21272 8424 21324 8430
rect 21272 8366 21324 8372
rect 21284 8090 21312 8366
rect 21560 8090 21588 9007
rect 21742 8732 22050 8741
rect 21742 8730 21748 8732
rect 21804 8730 21828 8732
rect 21884 8730 21908 8732
rect 21964 8730 21988 8732
rect 22044 8730 22050 8732
rect 21804 8678 21806 8730
rect 21986 8678 21988 8730
rect 21742 8676 21748 8678
rect 21804 8676 21828 8678
rect 21884 8676 21908 8678
rect 21964 8676 21988 8678
rect 22044 8676 22050 8678
rect 21742 8667 22050 8676
rect 21272 8084 21324 8090
rect 21272 8026 21324 8032
rect 21548 8084 21600 8090
rect 21548 8026 21600 8032
rect 21454 7848 21510 7857
rect 21454 7783 21510 7792
rect 21468 6798 21496 7783
rect 21742 7644 22050 7653
rect 21742 7642 21748 7644
rect 21804 7642 21828 7644
rect 21884 7642 21908 7644
rect 21964 7642 21988 7644
rect 22044 7642 22050 7644
rect 21804 7590 21806 7642
rect 21986 7590 21988 7642
rect 21742 7588 21748 7590
rect 21804 7588 21828 7590
rect 21884 7588 21908 7590
rect 21964 7588 21988 7590
rect 22044 7588 22050 7590
rect 21742 7579 22050 7588
rect 22388 6866 22416 16118
rect 22376 6860 22428 6866
rect 22376 6802 22428 6808
rect 21456 6792 21508 6798
rect 21456 6734 21508 6740
rect 21742 6556 22050 6565
rect 21742 6554 21748 6556
rect 21804 6554 21828 6556
rect 21884 6554 21908 6556
rect 21964 6554 21988 6556
rect 22044 6554 22050 6556
rect 21804 6502 21806 6554
rect 21986 6502 21988 6554
rect 21742 6500 21748 6502
rect 21804 6500 21828 6502
rect 21884 6500 21908 6502
rect 21964 6500 21988 6502
rect 22044 6500 22050 6502
rect 21742 6491 22050 6500
rect 21178 6352 21234 6361
rect 21178 6287 21234 6296
rect 21546 5808 21602 5817
rect 21546 5743 21602 5752
rect 21560 5710 21588 5743
rect 21272 5704 21324 5710
rect 21272 5646 21324 5652
rect 21548 5704 21600 5710
rect 21548 5646 21600 5652
rect 21284 5273 21312 5646
rect 21742 5468 22050 5477
rect 21742 5466 21748 5468
rect 21804 5466 21828 5468
rect 21884 5466 21908 5468
rect 21964 5466 21988 5468
rect 22044 5466 22050 5468
rect 21804 5414 21806 5466
rect 21986 5414 21988 5466
rect 21742 5412 21748 5414
rect 21804 5412 21828 5414
rect 21884 5412 21908 5414
rect 21964 5412 21988 5414
rect 22044 5412 22050 5414
rect 21742 5403 22050 5412
rect 21270 5264 21326 5273
rect 21270 5199 21326 5208
rect 21548 5228 21600 5234
rect 21548 5170 21600 5176
rect 21560 5001 21588 5170
rect 21546 4992 21602 5001
rect 21546 4927 21602 4936
rect 21546 4584 21602 4593
rect 21546 4519 21602 4528
rect 21088 4276 21140 4282
rect 21088 4218 21140 4224
rect 20718 4176 20774 4185
rect 21560 4146 21588 4519
rect 21742 4380 22050 4389
rect 21742 4378 21748 4380
rect 21804 4378 21828 4380
rect 21884 4378 21908 4380
rect 21964 4378 21988 4380
rect 22044 4378 22050 4380
rect 21804 4326 21806 4378
rect 21986 4326 21988 4378
rect 21742 4324 21748 4326
rect 21804 4324 21828 4326
rect 21884 4324 21908 4326
rect 21964 4324 21988 4326
rect 22044 4324 22050 4326
rect 21742 4315 22050 4324
rect 20718 4111 20774 4120
rect 21272 4140 21324 4146
rect 21272 4082 21324 4088
rect 21548 4140 21600 4146
rect 21548 4082 21600 4088
rect 21284 3777 21312 4082
rect 21270 3768 21326 3777
rect 21270 3703 21326 3712
rect 21548 3528 21600 3534
rect 21546 3496 21548 3505
rect 21600 3496 21602 3505
rect 21546 3431 21602 3440
rect 21742 3292 22050 3301
rect 21742 3290 21748 3292
rect 21804 3290 21828 3292
rect 21884 3290 21908 3292
rect 21964 3290 21988 3292
rect 22044 3290 22050 3292
rect 21804 3238 21806 3290
rect 21986 3238 21988 3290
rect 21742 3236 21748 3238
rect 21804 3236 21828 3238
rect 21884 3236 21908 3238
rect 21964 3236 21988 3238
rect 22044 3236 22050 3238
rect 21742 3227 22050 3236
rect 20444 3188 20496 3194
rect 20444 3130 20496 3136
rect 20628 3052 20680 3058
rect 20628 2994 20680 3000
rect 21272 3052 21324 3058
rect 21272 2994 21324 3000
rect 21548 3052 21600 3058
rect 21548 2994 21600 3000
rect 20260 2848 20312 2854
rect 20260 2790 20312 2796
rect 19143 2748 19451 2757
rect 19143 2746 19149 2748
rect 19205 2746 19229 2748
rect 19285 2746 19309 2748
rect 19365 2746 19389 2748
rect 19445 2746 19451 2748
rect 20088 2746 20208 2774
rect 19205 2694 19207 2746
rect 19387 2694 19389 2746
rect 19143 2692 19149 2694
rect 19205 2692 19229 2694
rect 19285 2692 19309 2694
rect 19365 2692 19389 2694
rect 19445 2692 19451 2694
rect 19143 2683 19451 2692
rect 8668 2644 8720 2650
rect 8668 2586 8720 2592
rect 16120 2644 16172 2650
rect 16120 2586 16172 2592
rect 6736 2440 6788 2446
rect 6736 2382 6788 2388
rect 20180 2378 20208 2746
rect 20640 2650 20668 2994
rect 20720 2848 20772 2854
rect 20720 2790 20772 2796
rect 20628 2644 20680 2650
rect 20732 2632 20760 2790
rect 20812 2644 20864 2650
rect 20732 2604 20812 2632
rect 20628 2586 20680 2592
rect 20812 2586 20864 2592
rect 21284 2553 21312 2994
rect 21560 2961 21588 2994
rect 21546 2952 21602 2961
rect 21546 2887 21602 2896
rect 21270 2544 21326 2553
rect 21270 2479 21326 2488
rect 20628 2440 20680 2446
rect 20628 2382 20680 2388
rect 21272 2440 21324 2446
rect 21272 2382 21324 2388
rect 21548 2440 21600 2446
rect 21548 2382 21600 2388
rect 20168 2372 20220 2378
rect 20168 2314 20220 2320
rect 20640 2310 20668 2382
rect 6828 2304 6880 2310
rect 6828 2246 6880 2252
rect 11704 2304 11756 2310
rect 11704 2246 11756 2252
rect 16028 2304 16080 2310
rect 16028 2246 16080 2252
rect 20628 2304 20680 2310
rect 20628 2246 20680 2252
rect 6148 2204 6456 2213
rect 6148 2202 6154 2204
rect 6210 2202 6234 2204
rect 6290 2202 6314 2204
rect 6370 2202 6394 2204
rect 6450 2202 6456 2204
rect 6210 2150 6212 2202
rect 6392 2150 6394 2202
rect 6148 2148 6154 2150
rect 6210 2148 6234 2150
rect 6290 2148 6314 2150
rect 6370 2148 6394 2150
rect 6450 2148 6456 2150
rect 6148 2139 6456 2148
rect 2778 1728 2834 1737
rect 2778 1663 2834 1672
rect 2240 1550 2360 1578
rect 2240 800 2268 1550
rect 6840 800 6868 2246
rect 11346 2204 11654 2213
rect 11346 2202 11352 2204
rect 11408 2202 11432 2204
rect 11488 2202 11512 2204
rect 11568 2202 11592 2204
rect 11648 2202 11654 2204
rect 11408 2150 11410 2202
rect 11590 2150 11592 2202
rect 11346 2148 11352 2150
rect 11408 2148 11432 2150
rect 11488 2148 11512 2150
rect 11568 2148 11592 2150
rect 11648 2148 11654 2150
rect 11346 2139 11654 2148
rect 11440 870 11560 898
rect 11440 800 11468 870
rect 2226 0 2282 800
rect 6826 0 6882 800
rect 11426 0 11482 800
rect 11532 762 11560 870
rect 11716 762 11744 2246
rect 16040 800 16068 2246
rect 16544 2204 16852 2213
rect 16544 2202 16550 2204
rect 16606 2202 16630 2204
rect 16686 2202 16710 2204
rect 16766 2202 16790 2204
rect 16846 2202 16852 2204
rect 16606 2150 16608 2202
rect 16788 2150 16790 2202
rect 16544 2148 16550 2150
rect 16606 2148 16630 2150
rect 16686 2148 16710 2150
rect 16766 2148 16790 2150
rect 16846 2148 16852 2150
rect 16544 2139 16852 2148
rect 20640 800 20668 2246
rect 21284 2009 21312 2382
rect 21270 2000 21326 2009
rect 21270 1935 21326 1944
rect 21560 1737 21588 2382
rect 21742 2204 22050 2213
rect 21742 2202 21748 2204
rect 21804 2202 21828 2204
rect 21884 2202 21908 2204
rect 21964 2202 21988 2204
rect 22044 2202 22050 2204
rect 21804 2150 21806 2202
rect 21986 2150 21988 2202
rect 21742 2148 21748 2150
rect 21804 2148 21828 2150
rect 21884 2148 21908 2150
rect 21964 2148 21988 2150
rect 22044 2148 22050 2150
rect 21742 2139 22050 2148
rect 21546 1728 21602 1737
rect 21546 1663 21602 1672
rect 11532 734 11744 762
rect 16026 0 16082 800
rect 20626 0 20682 800
<< via2 >>
rect 1490 20032 1546 20088
rect 1490 19660 1492 19680
rect 1492 19660 1544 19680
rect 1544 19660 1546 19680
rect 1490 19624 1546 19660
rect 1490 18808 1546 18864
rect 1490 18400 1546 18456
rect 1858 20440 1914 20496
rect 1858 19236 1914 19272
rect 1858 19216 1860 19236
rect 1860 19216 1912 19236
rect 1912 19216 1914 19236
rect 1490 18028 1492 18048
rect 1492 18028 1544 18048
rect 1544 18028 1546 18048
rect 1490 17992 1546 18028
rect 3054 21256 3110 21312
rect 2778 20848 2834 20904
rect 1490 17176 1546 17232
rect 1490 16768 1546 16824
rect 1490 16396 1492 16416
rect 1492 16396 1544 16416
rect 1544 16396 1546 16416
rect 1490 16360 1546 16396
rect 1490 15544 1546 15600
rect 1490 15136 1546 15192
rect 1490 14764 1492 14784
rect 1492 14764 1544 14784
rect 1544 14764 1546 14784
rect 1490 14728 1546 14764
rect 1858 17584 1914 17640
rect 1766 16496 1822 16552
rect 1858 15972 1914 16008
rect 1858 15952 1860 15972
rect 1860 15952 1912 15972
rect 1912 15952 1914 15972
rect 2410 16496 2466 16552
rect 2318 15952 2374 16008
rect 1490 13912 1546 13968
rect 1490 13504 1546 13560
rect 1398 13096 1454 13152
rect 1490 12280 1546 12336
rect 1490 11076 1546 11112
rect 1490 11056 1492 11076
rect 1492 11056 1544 11076
rect 1544 11056 1546 11076
rect 1398 10648 1454 10704
rect 1490 10240 1546 10296
rect 1398 9016 1454 9072
rect 1306 8200 1362 8256
rect 1674 12316 1676 12336
rect 1676 12316 1728 12336
rect 1728 12316 1730 12336
rect 1674 12280 1730 12316
rect 1858 14320 1914 14376
rect 3330 20304 3386 20360
rect 2870 19252 2872 19272
rect 2872 19252 2924 19272
rect 2924 19252 2926 19272
rect 2870 19216 2926 19252
rect 2778 18264 2834 18320
rect 2686 18128 2742 18184
rect 2226 12724 2228 12744
rect 2228 12724 2280 12744
rect 2280 12724 2282 12744
rect 2226 12688 2282 12724
rect 1858 11872 1914 11928
rect 1674 11636 1676 11656
rect 1676 11636 1728 11656
rect 1728 11636 1730 11656
rect 1674 11600 1730 11636
rect 2134 11464 2190 11520
rect 1398 7792 1454 7848
rect 1582 6704 1638 6760
rect 1674 6568 1730 6624
rect 2318 10512 2374 10568
rect 2042 10124 2098 10160
rect 2042 10104 2044 10124
rect 2044 10104 2096 10124
rect 2096 10104 2098 10124
rect 1858 9424 1914 9480
rect 2134 9832 2190 9888
rect 2226 9560 2282 9616
rect 1398 5752 1454 5808
rect 1674 5752 1730 5808
rect 1582 5616 1638 5672
rect 1398 5344 1454 5400
rect 1398 4936 1454 4992
rect 1674 4564 1676 4584
rect 1676 4564 1728 4584
rect 1728 4564 1730 4584
rect 1674 4528 1730 4564
rect 1398 3712 1454 3768
rect 1398 3304 1454 3360
rect 2226 8608 2282 8664
rect 2778 16108 2834 16144
rect 2778 16088 2780 16108
rect 2780 16088 2832 16108
rect 2832 16088 2834 16108
rect 2686 12144 2742 12200
rect 2686 10784 2742 10840
rect 3238 18944 3294 19000
rect 3330 18672 3386 18728
rect 3555 20154 3611 20156
rect 3635 20154 3691 20156
rect 3715 20154 3771 20156
rect 3795 20154 3851 20156
rect 3555 20102 3601 20154
rect 3601 20102 3611 20154
rect 3635 20102 3665 20154
rect 3665 20102 3677 20154
rect 3677 20102 3691 20154
rect 3715 20102 3729 20154
rect 3729 20102 3741 20154
rect 3741 20102 3771 20154
rect 3795 20102 3805 20154
rect 3805 20102 3851 20154
rect 3555 20100 3611 20102
rect 3635 20100 3691 20102
rect 3715 20100 3771 20102
rect 3795 20100 3851 20102
rect 3974 20032 4030 20088
rect 3790 19372 3846 19408
rect 3790 19352 3792 19372
rect 3792 19352 3844 19372
rect 3844 19352 3846 19372
rect 3555 19066 3611 19068
rect 3635 19066 3691 19068
rect 3715 19066 3771 19068
rect 3795 19066 3851 19068
rect 3555 19014 3601 19066
rect 3601 19014 3611 19066
rect 3635 19014 3665 19066
rect 3665 19014 3677 19066
rect 3677 19014 3691 19066
rect 3715 19014 3729 19066
rect 3729 19014 3741 19066
rect 3741 19014 3771 19066
rect 3795 19014 3805 19066
rect 3805 19014 3851 19066
rect 3555 19012 3611 19014
rect 3635 19012 3691 19014
rect 3715 19012 3771 19014
rect 3795 19012 3851 19014
rect 3514 18672 3570 18728
rect 4158 19116 4160 19136
rect 4160 19116 4212 19136
rect 4212 19116 4214 19136
rect 4158 19080 4214 19116
rect 2410 7248 2466 7304
rect 2226 6976 2282 7032
rect 1950 6296 2006 6352
rect 2226 6196 2228 6216
rect 2228 6196 2280 6216
rect 2280 6196 2282 6216
rect 2226 6160 2282 6196
rect 3555 17978 3611 17980
rect 3635 17978 3691 17980
rect 3715 17978 3771 17980
rect 3795 17978 3851 17980
rect 3555 17926 3601 17978
rect 3601 17926 3611 17978
rect 3635 17926 3665 17978
rect 3665 17926 3677 17978
rect 3677 17926 3691 17978
rect 3715 17926 3729 17978
rect 3729 17926 3741 17978
rect 3741 17926 3771 17978
rect 3795 17926 3805 17978
rect 3805 17926 3851 17978
rect 3555 17924 3611 17926
rect 3635 17924 3691 17926
rect 3715 17924 3771 17926
rect 3795 17924 3851 17926
rect 3555 16890 3611 16892
rect 3635 16890 3691 16892
rect 3715 16890 3771 16892
rect 3795 16890 3851 16892
rect 3555 16838 3601 16890
rect 3601 16838 3611 16890
rect 3635 16838 3665 16890
rect 3665 16838 3677 16890
rect 3677 16838 3691 16890
rect 3715 16838 3729 16890
rect 3729 16838 3741 16890
rect 3741 16838 3771 16890
rect 3795 16838 3805 16890
rect 3805 16838 3851 16890
rect 3555 16836 3611 16838
rect 3635 16836 3691 16838
rect 3715 16836 3771 16838
rect 3795 16836 3851 16838
rect 4066 18028 4068 18048
rect 4068 18028 4120 18048
rect 4120 18028 4122 18048
rect 4066 17992 4122 18028
rect 3882 16088 3938 16144
rect 3555 15802 3611 15804
rect 3635 15802 3691 15804
rect 3715 15802 3771 15804
rect 3795 15802 3851 15804
rect 3555 15750 3601 15802
rect 3601 15750 3611 15802
rect 3635 15750 3665 15802
rect 3665 15750 3677 15802
rect 3677 15750 3691 15802
rect 3715 15750 3729 15802
rect 3729 15750 3741 15802
rect 3741 15750 3771 15802
rect 3795 15750 3805 15802
rect 3805 15750 3851 15802
rect 3555 15748 3611 15750
rect 3635 15748 3691 15750
rect 3715 15748 3771 15750
rect 3795 15748 3851 15750
rect 3555 14714 3611 14716
rect 3635 14714 3691 14716
rect 3715 14714 3771 14716
rect 3795 14714 3851 14716
rect 3555 14662 3601 14714
rect 3601 14662 3611 14714
rect 3635 14662 3665 14714
rect 3665 14662 3677 14714
rect 3677 14662 3691 14714
rect 3715 14662 3729 14714
rect 3729 14662 3741 14714
rect 3741 14662 3771 14714
rect 3795 14662 3805 14714
rect 3805 14662 3851 14714
rect 3555 14660 3611 14662
rect 3635 14660 3691 14662
rect 3715 14660 3771 14662
rect 3795 14660 3851 14662
rect 3555 13626 3611 13628
rect 3635 13626 3691 13628
rect 3715 13626 3771 13628
rect 3795 13626 3851 13628
rect 3555 13574 3601 13626
rect 3601 13574 3611 13626
rect 3635 13574 3665 13626
rect 3665 13574 3677 13626
rect 3677 13574 3691 13626
rect 3715 13574 3729 13626
rect 3729 13574 3741 13626
rect 3741 13574 3771 13626
rect 3795 13574 3805 13626
rect 3805 13574 3851 13626
rect 3555 13572 3611 13574
rect 3635 13572 3691 13574
rect 3715 13572 3771 13574
rect 3795 13572 3851 13574
rect 3555 12538 3611 12540
rect 3635 12538 3691 12540
rect 3715 12538 3771 12540
rect 3795 12538 3851 12540
rect 3555 12486 3601 12538
rect 3601 12486 3611 12538
rect 3635 12486 3665 12538
rect 3665 12486 3677 12538
rect 3677 12486 3691 12538
rect 3715 12486 3729 12538
rect 3729 12486 3741 12538
rect 3741 12486 3771 12538
rect 3795 12486 3805 12538
rect 3805 12486 3851 12538
rect 3555 12484 3611 12486
rect 3635 12484 3691 12486
rect 3715 12484 3771 12486
rect 3795 12484 3851 12486
rect 3555 11450 3611 11452
rect 3635 11450 3691 11452
rect 3715 11450 3771 11452
rect 3795 11450 3851 11452
rect 3555 11398 3601 11450
rect 3601 11398 3611 11450
rect 3635 11398 3665 11450
rect 3665 11398 3677 11450
rect 3677 11398 3691 11450
rect 3715 11398 3729 11450
rect 3729 11398 3741 11450
rect 3741 11398 3771 11450
rect 3795 11398 3805 11450
rect 3805 11398 3851 11450
rect 3555 11396 3611 11398
rect 3635 11396 3691 11398
rect 3715 11396 3771 11398
rect 3795 11396 3851 11398
rect 3238 11192 3294 11248
rect 3555 10362 3611 10364
rect 3635 10362 3691 10364
rect 3715 10362 3771 10364
rect 3795 10362 3851 10364
rect 3555 10310 3601 10362
rect 3601 10310 3611 10362
rect 3635 10310 3665 10362
rect 3665 10310 3677 10362
rect 3677 10310 3691 10362
rect 3715 10310 3729 10362
rect 3729 10310 3741 10362
rect 3741 10310 3771 10362
rect 3795 10310 3805 10362
rect 3805 10310 3851 10362
rect 3555 10308 3611 10310
rect 3635 10308 3691 10310
rect 3715 10308 3771 10310
rect 3795 10308 3851 10310
rect 3514 9832 3570 9888
rect 2778 5888 2834 5944
rect 3054 6432 3110 6488
rect 1950 4120 2006 4176
rect 3555 9274 3611 9276
rect 3635 9274 3691 9276
rect 3715 9274 3771 9276
rect 3795 9274 3851 9276
rect 3555 9222 3601 9274
rect 3601 9222 3611 9274
rect 3635 9222 3665 9274
rect 3665 9222 3677 9274
rect 3677 9222 3691 9274
rect 3715 9222 3729 9274
rect 3729 9222 3741 9274
rect 3741 9222 3771 9274
rect 3795 9222 3805 9274
rect 3805 9222 3851 9274
rect 3555 9220 3611 9222
rect 3635 9220 3691 9222
rect 3715 9220 3771 9222
rect 3795 9220 3851 9222
rect 3555 8186 3611 8188
rect 3635 8186 3691 8188
rect 3715 8186 3771 8188
rect 3795 8186 3851 8188
rect 3555 8134 3601 8186
rect 3601 8134 3611 8186
rect 3635 8134 3665 8186
rect 3665 8134 3677 8186
rect 3677 8134 3691 8186
rect 3715 8134 3729 8186
rect 3729 8134 3741 8186
rect 3741 8134 3771 8186
rect 3795 8134 3805 8186
rect 3805 8134 3851 8186
rect 3555 8132 3611 8134
rect 3635 8132 3691 8134
rect 3715 8132 3771 8134
rect 3795 8132 3851 8134
rect 3422 7384 3478 7440
rect 4434 19760 4490 19816
rect 4894 20204 4896 20224
rect 4896 20204 4948 20224
rect 4948 20204 4950 20224
rect 4894 20168 4950 20204
rect 6154 20698 6210 20700
rect 6234 20698 6290 20700
rect 6314 20698 6370 20700
rect 6394 20698 6450 20700
rect 6154 20646 6200 20698
rect 6200 20646 6210 20698
rect 6234 20646 6264 20698
rect 6264 20646 6276 20698
rect 6276 20646 6290 20698
rect 6314 20646 6328 20698
rect 6328 20646 6340 20698
rect 6340 20646 6370 20698
rect 6394 20646 6404 20698
rect 6404 20646 6450 20698
rect 6154 20644 6210 20646
rect 6234 20644 6290 20646
rect 6314 20644 6370 20646
rect 6394 20644 6450 20646
rect 5354 20440 5410 20496
rect 4434 15544 4490 15600
rect 4250 11056 4306 11112
rect 4434 10784 4490 10840
rect 3974 7792 4030 7848
rect 3330 6452 3386 6488
rect 3330 6432 3332 6452
rect 3332 6432 3384 6452
rect 3384 6432 3386 6452
rect 3555 7098 3611 7100
rect 3635 7098 3691 7100
rect 3715 7098 3771 7100
rect 3795 7098 3851 7100
rect 3555 7046 3601 7098
rect 3601 7046 3611 7098
rect 3635 7046 3665 7098
rect 3665 7046 3677 7098
rect 3677 7046 3691 7098
rect 3715 7046 3729 7098
rect 3729 7046 3741 7098
rect 3741 7046 3771 7098
rect 3795 7046 3805 7098
rect 3805 7046 3851 7098
rect 3555 7044 3611 7046
rect 3635 7044 3691 7046
rect 3715 7044 3771 7046
rect 3795 7044 3851 7046
rect 4158 7148 4160 7168
rect 4160 7148 4212 7168
rect 4212 7148 4214 7168
rect 4158 7112 4214 7148
rect 3555 6010 3611 6012
rect 3635 6010 3691 6012
rect 3715 6010 3771 6012
rect 3795 6010 3851 6012
rect 3555 5958 3601 6010
rect 3601 5958 3611 6010
rect 3635 5958 3665 6010
rect 3665 5958 3677 6010
rect 3677 5958 3691 6010
rect 3715 5958 3729 6010
rect 3729 5958 3741 6010
rect 3741 5958 3771 6010
rect 3795 5958 3805 6010
rect 3805 5958 3851 6010
rect 3555 5956 3611 5958
rect 3635 5956 3691 5958
rect 3715 5956 3771 5958
rect 3795 5956 3851 5958
rect 3555 4922 3611 4924
rect 3635 4922 3691 4924
rect 3715 4922 3771 4924
rect 3795 4922 3851 4924
rect 3555 4870 3601 4922
rect 3601 4870 3611 4922
rect 3635 4870 3665 4922
rect 3665 4870 3677 4922
rect 3677 4870 3691 4922
rect 3715 4870 3729 4922
rect 3729 4870 3741 4922
rect 3741 4870 3771 4922
rect 3795 4870 3805 4922
rect 3805 4870 3851 4922
rect 3555 4868 3611 4870
rect 3635 4868 3691 4870
rect 3715 4868 3771 4870
rect 3795 4868 3851 4870
rect 3555 3834 3611 3836
rect 3635 3834 3691 3836
rect 3715 3834 3771 3836
rect 3795 3834 3851 3836
rect 3555 3782 3601 3834
rect 3601 3782 3611 3834
rect 3635 3782 3665 3834
rect 3665 3782 3677 3834
rect 3677 3782 3691 3834
rect 3715 3782 3729 3834
rect 3729 3782 3741 3834
rect 3741 3782 3771 3834
rect 3795 3782 3805 3834
rect 3805 3782 3851 3834
rect 3555 3780 3611 3782
rect 3635 3780 3691 3782
rect 3715 3780 3771 3782
rect 3795 3780 3851 3782
rect 1398 2896 1454 2952
rect 1674 2488 1730 2544
rect 2226 2080 2282 2136
rect 3555 2746 3611 2748
rect 3635 2746 3691 2748
rect 3715 2746 3771 2748
rect 3795 2746 3851 2748
rect 3555 2694 3601 2746
rect 3601 2694 3611 2746
rect 3635 2694 3665 2746
rect 3665 2694 3677 2746
rect 3677 2694 3691 2746
rect 3715 2694 3729 2746
rect 3729 2694 3741 2746
rect 3741 2694 3771 2746
rect 3795 2694 3805 2746
rect 3805 2694 3851 2746
rect 3555 2692 3611 2694
rect 3635 2692 3691 2694
rect 3715 2692 3771 2694
rect 3795 2692 3851 2694
rect 5538 19080 5594 19136
rect 5170 11056 5226 11112
rect 5170 10004 5172 10024
rect 5172 10004 5224 10024
rect 5224 10004 5226 10024
rect 5170 9968 5226 10004
rect 5354 9832 5410 9888
rect 5262 9696 5318 9752
rect 6366 19896 6422 19952
rect 6154 19610 6210 19612
rect 6234 19610 6290 19612
rect 6314 19610 6370 19612
rect 6394 19610 6450 19612
rect 6154 19558 6200 19610
rect 6200 19558 6210 19610
rect 6234 19558 6264 19610
rect 6264 19558 6276 19610
rect 6276 19558 6290 19610
rect 6314 19558 6328 19610
rect 6328 19558 6340 19610
rect 6340 19558 6370 19610
rect 6394 19558 6404 19610
rect 6404 19558 6450 19610
rect 6154 19556 6210 19558
rect 6234 19556 6290 19558
rect 6314 19556 6370 19558
rect 6394 19556 6450 19558
rect 5722 12416 5778 12472
rect 5262 6840 5318 6896
rect 7102 19488 7158 19544
rect 6550 18536 6606 18592
rect 6154 18522 6210 18524
rect 6234 18522 6290 18524
rect 6314 18522 6370 18524
rect 6394 18522 6450 18524
rect 6154 18470 6200 18522
rect 6200 18470 6210 18522
rect 6234 18470 6264 18522
rect 6264 18470 6276 18522
rect 6276 18470 6290 18522
rect 6314 18470 6328 18522
rect 6328 18470 6340 18522
rect 6340 18470 6370 18522
rect 6394 18470 6404 18522
rect 6404 18470 6450 18522
rect 6154 18468 6210 18470
rect 6234 18468 6290 18470
rect 6314 18468 6370 18470
rect 6394 18468 6450 18470
rect 6550 17992 6606 18048
rect 6154 17434 6210 17436
rect 6234 17434 6290 17436
rect 6314 17434 6370 17436
rect 6394 17434 6450 17436
rect 6154 17382 6200 17434
rect 6200 17382 6210 17434
rect 6234 17382 6264 17434
rect 6264 17382 6276 17434
rect 6276 17382 6290 17434
rect 6314 17382 6328 17434
rect 6328 17382 6340 17434
rect 6340 17382 6370 17434
rect 6394 17382 6404 17434
rect 6404 17382 6450 17434
rect 6154 17380 6210 17382
rect 6234 17380 6290 17382
rect 6314 17380 6370 17382
rect 6394 17380 6450 17382
rect 6154 16346 6210 16348
rect 6234 16346 6290 16348
rect 6314 16346 6370 16348
rect 6394 16346 6450 16348
rect 6154 16294 6200 16346
rect 6200 16294 6210 16346
rect 6234 16294 6264 16346
rect 6264 16294 6276 16346
rect 6276 16294 6290 16346
rect 6314 16294 6328 16346
rect 6328 16294 6340 16346
rect 6340 16294 6370 16346
rect 6394 16294 6404 16346
rect 6404 16294 6450 16346
rect 6154 16292 6210 16294
rect 6234 16292 6290 16294
rect 6314 16292 6370 16294
rect 6394 16292 6450 16294
rect 6550 15428 6606 15464
rect 6550 15408 6552 15428
rect 6552 15408 6604 15428
rect 6604 15408 6606 15428
rect 6154 15258 6210 15260
rect 6234 15258 6290 15260
rect 6314 15258 6370 15260
rect 6394 15258 6450 15260
rect 6154 15206 6200 15258
rect 6200 15206 6210 15258
rect 6234 15206 6264 15258
rect 6264 15206 6276 15258
rect 6276 15206 6290 15258
rect 6314 15206 6328 15258
rect 6328 15206 6340 15258
rect 6340 15206 6370 15258
rect 6394 15206 6404 15258
rect 6404 15206 6450 15258
rect 6154 15204 6210 15206
rect 6234 15204 6290 15206
rect 6314 15204 6370 15206
rect 6394 15204 6450 15206
rect 6154 14170 6210 14172
rect 6234 14170 6290 14172
rect 6314 14170 6370 14172
rect 6394 14170 6450 14172
rect 6154 14118 6200 14170
rect 6200 14118 6210 14170
rect 6234 14118 6264 14170
rect 6264 14118 6276 14170
rect 6276 14118 6290 14170
rect 6314 14118 6328 14170
rect 6328 14118 6340 14170
rect 6340 14118 6370 14170
rect 6394 14118 6404 14170
rect 6404 14118 6450 14170
rect 6154 14116 6210 14118
rect 6234 14116 6290 14118
rect 6314 14116 6370 14118
rect 6394 14116 6450 14118
rect 6154 13082 6210 13084
rect 6234 13082 6290 13084
rect 6314 13082 6370 13084
rect 6394 13082 6450 13084
rect 6154 13030 6200 13082
rect 6200 13030 6210 13082
rect 6234 13030 6264 13082
rect 6264 13030 6276 13082
rect 6276 13030 6290 13082
rect 6314 13030 6328 13082
rect 6328 13030 6340 13082
rect 6340 13030 6370 13082
rect 6394 13030 6404 13082
rect 6404 13030 6450 13082
rect 6154 13028 6210 13030
rect 6234 13028 6290 13030
rect 6314 13028 6370 13030
rect 6394 13028 6450 13030
rect 6154 11994 6210 11996
rect 6234 11994 6290 11996
rect 6314 11994 6370 11996
rect 6394 11994 6450 11996
rect 6154 11942 6200 11994
rect 6200 11942 6210 11994
rect 6234 11942 6264 11994
rect 6264 11942 6276 11994
rect 6276 11942 6290 11994
rect 6314 11942 6328 11994
rect 6328 11942 6340 11994
rect 6340 11942 6370 11994
rect 6394 11942 6404 11994
rect 6404 11942 6450 11994
rect 6154 11940 6210 11942
rect 6234 11940 6290 11942
rect 6314 11940 6370 11942
rect 6394 11940 6450 11942
rect 6154 10906 6210 10908
rect 6234 10906 6290 10908
rect 6314 10906 6370 10908
rect 6394 10906 6450 10908
rect 6154 10854 6200 10906
rect 6200 10854 6210 10906
rect 6234 10854 6264 10906
rect 6264 10854 6276 10906
rect 6276 10854 6290 10906
rect 6314 10854 6328 10906
rect 6328 10854 6340 10906
rect 6340 10854 6370 10906
rect 6394 10854 6404 10906
rect 6404 10854 6450 10906
rect 6154 10852 6210 10854
rect 6234 10852 6290 10854
rect 6314 10852 6370 10854
rect 6394 10852 6450 10854
rect 6154 9818 6210 9820
rect 6234 9818 6290 9820
rect 6314 9818 6370 9820
rect 6394 9818 6450 9820
rect 6154 9766 6200 9818
rect 6200 9766 6210 9818
rect 6234 9766 6264 9818
rect 6264 9766 6276 9818
rect 6276 9766 6290 9818
rect 6314 9766 6328 9818
rect 6328 9766 6340 9818
rect 6340 9766 6370 9818
rect 6394 9766 6404 9818
rect 6404 9766 6450 9818
rect 6154 9764 6210 9766
rect 6234 9764 6290 9766
rect 6314 9764 6370 9766
rect 6394 9764 6450 9766
rect 6154 8730 6210 8732
rect 6234 8730 6290 8732
rect 6314 8730 6370 8732
rect 6394 8730 6450 8732
rect 6154 8678 6200 8730
rect 6200 8678 6210 8730
rect 6234 8678 6264 8730
rect 6264 8678 6276 8730
rect 6276 8678 6290 8730
rect 6314 8678 6328 8730
rect 6328 8678 6340 8730
rect 6340 8678 6370 8730
rect 6394 8678 6404 8730
rect 6404 8678 6450 8730
rect 6154 8676 6210 8678
rect 6234 8676 6290 8678
rect 6314 8676 6370 8678
rect 6394 8676 6450 8678
rect 6550 7792 6606 7848
rect 6154 7642 6210 7644
rect 6234 7642 6290 7644
rect 6314 7642 6370 7644
rect 6394 7642 6450 7644
rect 6154 7590 6200 7642
rect 6200 7590 6210 7642
rect 6234 7590 6264 7642
rect 6264 7590 6276 7642
rect 6276 7590 6290 7642
rect 6314 7590 6328 7642
rect 6328 7590 6340 7642
rect 6340 7590 6370 7642
rect 6394 7590 6404 7642
rect 6404 7590 6450 7642
rect 6154 7588 6210 7590
rect 6234 7588 6290 7590
rect 6314 7588 6370 7590
rect 6394 7588 6450 7590
rect 5998 7248 6054 7304
rect 5906 7112 5962 7168
rect 6154 6554 6210 6556
rect 6234 6554 6290 6556
rect 6314 6554 6370 6556
rect 6394 6554 6450 6556
rect 6154 6502 6200 6554
rect 6200 6502 6210 6554
rect 6234 6502 6264 6554
rect 6264 6502 6276 6554
rect 6276 6502 6290 6554
rect 6314 6502 6328 6554
rect 6328 6502 6340 6554
rect 6340 6502 6370 6554
rect 6394 6502 6404 6554
rect 6404 6502 6450 6554
rect 6154 6500 6210 6502
rect 6234 6500 6290 6502
rect 6314 6500 6370 6502
rect 6394 6500 6450 6502
rect 5906 6196 5908 6216
rect 5908 6196 5960 6216
rect 5960 6196 5962 6216
rect 5906 6160 5962 6196
rect 6154 5466 6210 5468
rect 6234 5466 6290 5468
rect 6314 5466 6370 5468
rect 6394 5466 6450 5468
rect 6154 5414 6200 5466
rect 6200 5414 6210 5466
rect 6234 5414 6264 5466
rect 6264 5414 6276 5466
rect 6276 5414 6290 5466
rect 6314 5414 6328 5466
rect 6328 5414 6340 5466
rect 6340 5414 6370 5466
rect 6394 5414 6404 5466
rect 6404 5414 6450 5466
rect 6154 5412 6210 5414
rect 6234 5412 6290 5414
rect 6314 5412 6370 5414
rect 6394 5412 6450 5414
rect 6154 4378 6210 4380
rect 6234 4378 6290 4380
rect 6314 4378 6370 4380
rect 6394 4378 6450 4380
rect 6154 4326 6200 4378
rect 6200 4326 6210 4378
rect 6234 4326 6264 4378
rect 6264 4326 6276 4378
rect 6276 4326 6290 4378
rect 6314 4326 6328 4378
rect 6328 4326 6340 4378
rect 6340 4326 6370 4378
rect 6394 4326 6404 4378
rect 6404 4326 6450 4378
rect 6154 4324 6210 4326
rect 6234 4324 6290 4326
rect 6314 4324 6370 4326
rect 6394 4324 6450 4326
rect 5998 3440 6054 3496
rect 6154 3290 6210 3292
rect 6234 3290 6290 3292
rect 6314 3290 6370 3292
rect 6394 3290 6450 3292
rect 6154 3238 6200 3290
rect 6200 3238 6210 3290
rect 6234 3238 6264 3290
rect 6264 3238 6276 3290
rect 6276 3238 6290 3290
rect 6314 3238 6328 3290
rect 6328 3238 6340 3290
rect 6340 3238 6370 3290
rect 6394 3238 6404 3290
rect 6404 3238 6450 3290
rect 6154 3236 6210 3238
rect 6234 3236 6290 3238
rect 6314 3236 6370 3238
rect 6394 3236 6450 3238
rect 7286 19624 7342 19680
rect 7286 19352 7342 19408
rect 7930 19508 7986 19544
rect 7930 19488 7932 19508
rect 7932 19488 7984 19508
rect 7984 19488 7986 19508
rect 8206 20032 8262 20088
rect 8114 19488 8170 19544
rect 8298 19488 8354 19544
rect 8298 19388 8300 19408
rect 8300 19388 8352 19408
rect 8352 19388 8354 19408
rect 8298 19352 8354 19388
rect 8298 19216 8354 19272
rect 8114 19116 8116 19136
rect 8116 19116 8168 19136
rect 8168 19116 8170 19136
rect 8114 19080 8170 19116
rect 8298 17992 8354 18048
rect 8753 20154 8809 20156
rect 8833 20154 8889 20156
rect 8913 20154 8969 20156
rect 8993 20154 9049 20156
rect 8753 20102 8799 20154
rect 8799 20102 8809 20154
rect 8833 20102 8863 20154
rect 8863 20102 8875 20154
rect 8875 20102 8889 20154
rect 8913 20102 8927 20154
rect 8927 20102 8939 20154
rect 8939 20102 8969 20154
rect 8993 20102 9003 20154
rect 9003 20102 9049 20154
rect 8753 20100 8809 20102
rect 8833 20100 8889 20102
rect 8913 20100 8969 20102
rect 8993 20100 9049 20102
rect 8942 19624 8998 19680
rect 8753 19066 8809 19068
rect 8833 19066 8889 19068
rect 8913 19066 8969 19068
rect 8993 19066 9049 19068
rect 8753 19014 8799 19066
rect 8799 19014 8809 19066
rect 8833 19014 8863 19066
rect 8863 19014 8875 19066
rect 8875 19014 8889 19066
rect 8913 19014 8927 19066
rect 8927 19014 8939 19066
rect 8939 19014 8969 19066
rect 8993 19014 9003 19066
rect 9003 19014 9049 19066
rect 8753 19012 8809 19014
rect 8833 19012 8889 19014
rect 8913 19012 8969 19014
rect 8993 19012 9049 19014
rect 8753 17978 8809 17980
rect 8833 17978 8889 17980
rect 8913 17978 8969 17980
rect 8993 17978 9049 17980
rect 8753 17926 8799 17978
rect 8799 17926 8809 17978
rect 8833 17926 8863 17978
rect 8863 17926 8875 17978
rect 8875 17926 8889 17978
rect 8913 17926 8927 17978
rect 8927 17926 8939 17978
rect 8939 17926 8969 17978
rect 8993 17926 9003 17978
rect 9003 17926 9049 17978
rect 8753 17924 8809 17926
rect 8833 17924 8889 17926
rect 8913 17924 8969 17926
rect 8993 17924 9049 17926
rect 7654 12416 7710 12472
rect 8206 12824 8262 12880
rect 8753 16890 8809 16892
rect 8833 16890 8889 16892
rect 8913 16890 8969 16892
rect 8993 16890 9049 16892
rect 8753 16838 8799 16890
rect 8799 16838 8809 16890
rect 8833 16838 8863 16890
rect 8863 16838 8875 16890
rect 8875 16838 8889 16890
rect 8913 16838 8927 16890
rect 8927 16838 8939 16890
rect 8939 16838 8969 16890
rect 8993 16838 9003 16890
rect 9003 16838 9049 16890
rect 8753 16836 8809 16838
rect 8833 16836 8889 16838
rect 8913 16836 8969 16838
rect 8993 16836 9049 16838
rect 8753 15802 8809 15804
rect 8833 15802 8889 15804
rect 8913 15802 8969 15804
rect 8993 15802 9049 15804
rect 8753 15750 8799 15802
rect 8799 15750 8809 15802
rect 8833 15750 8863 15802
rect 8863 15750 8875 15802
rect 8875 15750 8889 15802
rect 8913 15750 8927 15802
rect 8927 15750 8939 15802
rect 8939 15750 8969 15802
rect 8993 15750 9003 15802
rect 9003 15750 9049 15802
rect 8753 15748 8809 15750
rect 8833 15748 8889 15750
rect 8913 15748 8969 15750
rect 8993 15748 9049 15750
rect 9218 15544 9274 15600
rect 8753 14714 8809 14716
rect 8833 14714 8889 14716
rect 8913 14714 8969 14716
rect 8993 14714 9049 14716
rect 8753 14662 8799 14714
rect 8799 14662 8809 14714
rect 8833 14662 8863 14714
rect 8863 14662 8875 14714
rect 8875 14662 8889 14714
rect 8913 14662 8927 14714
rect 8927 14662 8939 14714
rect 8939 14662 8969 14714
rect 8993 14662 9003 14714
rect 9003 14662 9049 14714
rect 8753 14660 8809 14662
rect 8833 14660 8889 14662
rect 8913 14660 8969 14662
rect 8993 14660 9049 14662
rect 8753 13626 8809 13628
rect 8833 13626 8889 13628
rect 8913 13626 8969 13628
rect 8993 13626 9049 13628
rect 8753 13574 8799 13626
rect 8799 13574 8809 13626
rect 8833 13574 8863 13626
rect 8863 13574 8875 13626
rect 8875 13574 8889 13626
rect 8913 13574 8927 13626
rect 8927 13574 8939 13626
rect 8939 13574 8969 13626
rect 8993 13574 9003 13626
rect 9003 13574 9049 13626
rect 8753 13572 8809 13574
rect 8833 13572 8889 13574
rect 8913 13572 8969 13574
rect 8993 13572 9049 13574
rect 8758 13368 8814 13424
rect 8753 12538 8809 12540
rect 8833 12538 8889 12540
rect 8913 12538 8969 12540
rect 8993 12538 9049 12540
rect 8753 12486 8799 12538
rect 8799 12486 8809 12538
rect 8833 12486 8863 12538
rect 8863 12486 8875 12538
rect 8875 12486 8889 12538
rect 8913 12486 8927 12538
rect 8927 12486 8939 12538
rect 8939 12486 8969 12538
rect 8993 12486 9003 12538
rect 9003 12486 9049 12538
rect 8753 12484 8809 12486
rect 8833 12484 8889 12486
rect 8913 12484 8969 12486
rect 8993 12484 9049 12486
rect 9678 19660 9680 19680
rect 9680 19660 9732 19680
rect 9732 19660 9734 19680
rect 9678 19624 9734 19660
rect 9402 17448 9458 17504
rect 9770 17076 9772 17096
rect 9772 17076 9824 17096
rect 9824 17076 9826 17096
rect 9770 17040 9826 17076
rect 8753 11450 8809 11452
rect 8833 11450 8889 11452
rect 8913 11450 8969 11452
rect 8993 11450 9049 11452
rect 8753 11398 8799 11450
rect 8799 11398 8809 11450
rect 8833 11398 8863 11450
rect 8863 11398 8875 11450
rect 8875 11398 8889 11450
rect 8913 11398 8927 11450
rect 8927 11398 8939 11450
rect 8939 11398 8969 11450
rect 8993 11398 9003 11450
rect 9003 11398 9049 11450
rect 8753 11396 8809 11398
rect 8833 11396 8889 11398
rect 8913 11396 8969 11398
rect 8993 11396 9049 11398
rect 8666 11192 8722 11248
rect 8206 9696 8262 9752
rect 8114 8880 8170 8936
rect 8753 10362 8809 10364
rect 8833 10362 8889 10364
rect 8913 10362 8969 10364
rect 8993 10362 9049 10364
rect 8753 10310 8799 10362
rect 8799 10310 8809 10362
rect 8833 10310 8863 10362
rect 8863 10310 8875 10362
rect 8875 10310 8889 10362
rect 8913 10310 8927 10362
rect 8927 10310 8939 10362
rect 8939 10310 8969 10362
rect 8993 10310 9003 10362
rect 9003 10310 9049 10362
rect 8753 10308 8809 10310
rect 8833 10308 8889 10310
rect 8913 10308 8969 10310
rect 8993 10308 9049 10310
rect 8753 9274 8809 9276
rect 8833 9274 8889 9276
rect 8913 9274 8969 9276
rect 8993 9274 9049 9276
rect 8753 9222 8799 9274
rect 8799 9222 8809 9274
rect 8833 9222 8863 9274
rect 8863 9222 8875 9274
rect 8875 9222 8889 9274
rect 8913 9222 8927 9274
rect 8927 9222 8939 9274
rect 8939 9222 8969 9274
rect 8993 9222 9003 9274
rect 9003 9222 9049 9274
rect 8753 9220 8809 9222
rect 8833 9220 8889 9222
rect 8913 9220 8969 9222
rect 8993 9220 9049 9222
rect 7102 6840 7158 6896
rect 8753 8186 8809 8188
rect 8833 8186 8889 8188
rect 8913 8186 8969 8188
rect 8993 8186 9049 8188
rect 8753 8134 8799 8186
rect 8799 8134 8809 8186
rect 8833 8134 8863 8186
rect 8863 8134 8875 8186
rect 8875 8134 8889 8186
rect 8913 8134 8927 8186
rect 8927 8134 8939 8186
rect 8939 8134 8969 8186
rect 8993 8134 9003 8186
rect 9003 8134 9049 8186
rect 8753 8132 8809 8134
rect 8833 8132 8889 8134
rect 8913 8132 8969 8134
rect 8993 8132 9049 8134
rect 11352 20698 11408 20700
rect 11432 20698 11488 20700
rect 11512 20698 11568 20700
rect 11592 20698 11648 20700
rect 11352 20646 11398 20698
rect 11398 20646 11408 20698
rect 11432 20646 11462 20698
rect 11462 20646 11474 20698
rect 11474 20646 11488 20698
rect 11512 20646 11526 20698
rect 11526 20646 11538 20698
rect 11538 20646 11568 20698
rect 11592 20646 11602 20698
rect 11602 20646 11648 20698
rect 11352 20644 11408 20646
rect 11432 20644 11488 20646
rect 11512 20644 11568 20646
rect 11592 20644 11648 20646
rect 10046 18808 10102 18864
rect 10046 18536 10102 18592
rect 10138 17720 10194 17776
rect 10782 18944 10838 19000
rect 9862 10104 9918 10160
rect 9954 9696 10010 9752
rect 10598 17484 10600 17504
rect 10600 17484 10652 17504
rect 10652 17484 10654 17504
rect 10598 17448 10654 17484
rect 10598 17076 10600 17096
rect 10600 17076 10652 17096
rect 10652 17076 10654 17096
rect 10598 17040 10654 17076
rect 10598 15544 10654 15600
rect 11352 19610 11408 19612
rect 11432 19610 11488 19612
rect 11512 19610 11568 19612
rect 11592 19610 11648 19612
rect 11352 19558 11398 19610
rect 11398 19558 11408 19610
rect 11432 19558 11462 19610
rect 11462 19558 11474 19610
rect 11474 19558 11488 19610
rect 11512 19558 11526 19610
rect 11526 19558 11538 19610
rect 11538 19558 11568 19610
rect 11592 19558 11602 19610
rect 11602 19558 11648 19610
rect 11352 19556 11408 19558
rect 11432 19556 11488 19558
rect 11512 19556 11568 19558
rect 11592 19556 11648 19558
rect 11334 18944 11390 19000
rect 11352 18522 11408 18524
rect 11432 18522 11488 18524
rect 11512 18522 11568 18524
rect 11592 18522 11648 18524
rect 11352 18470 11398 18522
rect 11398 18470 11408 18522
rect 11432 18470 11462 18522
rect 11462 18470 11474 18522
rect 11474 18470 11488 18522
rect 11512 18470 11526 18522
rect 11526 18470 11538 18522
rect 11538 18470 11568 18522
rect 11592 18470 11602 18522
rect 11602 18470 11648 18522
rect 11352 18468 11408 18470
rect 11432 18468 11488 18470
rect 11512 18468 11568 18470
rect 11592 18468 11648 18470
rect 11978 19372 12034 19408
rect 11978 19352 11980 19372
rect 11980 19352 12032 19372
rect 12032 19352 12034 19372
rect 11352 17434 11408 17436
rect 11432 17434 11488 17436
rect 11512 17434 11568 17436
rect 11592 17434 11648 17436
rect 11352 17382 11398 17434
rect 11398 17382 11408 17434
rect 11432 17382 11462 17434
rect 11462 17382 11474 17434
rect 11474 17382 11488 17434
rect 11512 17382 11526 17434
rect 11526 17382 11538 17434
rect 11538 17382 11568 17434
rect 11592 17382 11602 17434
rect 11602 17382 11648 17434
rect 11352 17380 11408 17382
rect 11432 17380 11488 17382
rect 11512 17380 11568 17382
rect 11592 17380 11648 17382
rect 11610 17212 11612 17232
rect 11612 17212 11664 17232
rect 11664 17212 11666 17232
rect 11610 17176 11666 17212
rect 11352 16346 11408 16348
rect 11432 16346 11488 16348
rect 11512 16346 11568 16348
rect 11592 16346 11648 16348
rect 11352 16294 11398 16346
rect 11398 16294 11408 16346
rect 11432 16294 11462 16346
rect 11462 16294 11474 16346
rect 11474 16294 11488 16346
rect 11512 16294 11526 16346
rect 11526 16294 11538 16346
rect 11538 16294 11568 16346
rect 11592 16294 11602 16346
rect 11602 16294 11648 16346
rect 11352 16292 11408 16294
rect 11432 16292 11488 16294
rect 11512 16292 11568 16294
rect 11592 16292 11648 16294
rect 11352 15258 11408 15260
rect 11432 15258 11488 15260
rect 11512 15258 11568 15260
rect 11592 15258 11648 15260
rect 11352 15206 11398 15258
rect 11398 15206 11408 15258
rect 11432 15206 11462 15258
rect 11462 15206 11474 15258
rect 11474 15206 11488 15258
rect 11512 15206 11526 15258
rect 11526 15206 11538 15258
rect 11538 15206 11568 15258
rect 11592 15206 11602 15258
rect 11602 15206 11648 15258
rect 11352 15204 11408 15206
rect 11432 15204 11488 15206
rect 11512 15204 11568 15206
rect 11592 15204 11648 15206
rect 11794 17484 11796 17504
rect 11796 17484 11848 17504
rect 11848 17484 11850 17504
rect 11794 17448 11850 17484
rect 12162 17584 12218 17640
rect 11886 16632 11942 16688
rect 11352 14170 11408 14172
rect 11432 14170 11488 14172
rect 11512 14170 11568 14172
rect 11592 14170 11648 14172
rect 11352 14118 11398 14170
rect 11398 14118 11408 14170
rect 11432 14118 11462 14170
rect 11462 14118 11474 14170
rect 11474 14118 11488 14170
rect 11512 14118 11526 14170
rect 11526 14118 11538 14170
rect 11538 14118 11568 14170
rect 11592 14118 11602 14170
rect 11602 14118 11648 14170
rect 11352 14116 11408 14118
rect 11432 14116 11488 14118
rect 11512 14116 11568 14118
rect 11592 14116 11648 14118
rect 11352 13082 11408 13084
rect 11432 13082 11488 13084
rect 11512 13082 11568 13084
rect 11592 13082 11648 13084
rect 11352 13030 11398 13082
rect 11398 13030 11408 13082
rect 11432 13030 11462 13082
rect 11462 13030 11474 13082
rect 11474 13030 11488 13082
rect 11512 13030 11526 13082
rect 11526 13030 11538 13082
rect 11538 13030 11568 13082
rect 11592 13030 11602 13082
rect 11602 13030 11648 13082
rect 11352 13028 11408 13030
rect 11432 13028 11488 13030
rect 11512 13028 11568 13030
rect 11592 13028 11648 13030
rect 10230 10648 10286 10704
rect 10966 9016 11022 9072
rect 11352 11994 11408 11996
rect 11432 11994 11488 11996
rect 11512 11994 11568 11996
rect 11592 11994 11648 11996
rect 11352 11942 11398 11994
rect 11398 11942 11408 11994
rect 11432 11942 11462 11994
rect 11462 11942 11474 11994
rect 11474 11942 11488 11994
rect 11512 11942 11526 11994
rect 11526 11942 11538 11994
rect 11538 11942 11568 11994
rect 11592 11942 11602 11994
rect 11602 11942 11648 11994
rect 11352 11940 11408 11942
rect 11432 11940 11488 11942
rect 11512 11940 11568 11942
rect 11592 11940 11648 11942
rect 11150 11736 11206 11792
rect 11352 10906 11408 10908
rect 11432 10906 11488 10908
rect 11512 10906 11568 10908
rect 11592 10906 11648 10908
rect 11352 10854 11398 10906
rect 11398 10854 11408 10906
rect 11432 10854 11462 10906
rect 11462 10854 11474 10906
rect 11474 10854 11488 10906
rect 11512 10854 11526 10906
rect 11526 10854 11538 10906
rect 11538 10854 11568 10906
rect 11592 10854 11602 10906
rect 11602 10854 11648 10906
rect 11352 10852 11408 10854
rect 11432 10852 11488 10854
rect 11512 10852 11568 10854
rect 11592 10852 11648 10854
rect 11352 9818 11408 9820
rect 11432 9818 11488 9820
rect 11512 9818 11568 9820
rect 11592 9818 11648 9820
rect 11352 9766 11398 9818
rect 11398 9766 11408 9818
rect 11432 9766 11462 9818
rect 11462 9766 11474 9818
rect 11474 9766 11488 9818
rect 11512 9766 11526 9818
rect 11526 9766 11538 9818
rect 11538 9766 11568 9818
rect 11592 9766 11602 9818
rect 11602 9766 11648 9818
rect 11352 9764 11408 9766
rect 11432 9764 11488 9766
rect 11512 9764 11568 9766
rect 11592 9764 11648 9766
rect 11352 8730 11408 8732
rect 11432 8730 11488 8732
rect 11512 8730 11568 8732
rect 11592 8730 11648 8732
rect 11352 8678 11398 8730
rect 11398 8678 11408 8730
rect 11432 8678 11462 8730
rect 11462 8678 11474 8730
rect 11474 8678 11488 8730
rect 11512 8678 11526 8730
rect 11526 8678 11538 8730
rect 11538 8678 11568 8730
rect 11592 8678 11602 8730
rect 11602 8678 11648 8730
rect 11352 8676 11408 8678
rect 11432 8676 11488 8678
rect 11512 8676 11568 8678
rect 11592 8676 11648 8678
rect 8753 7098 8809 7100
rect 8833 7098 8889 7100
rect 8913 7098 8969 7100
rect 8993 7098 9049 7100
rect 8753 7046 8799 7098
rect 8799 7046 8809 7098
rect 8833 7046 8863 7098
rect 8863 7046 8875 7098
rect 8875 7046 8889 7098
rect 8913 7046 8927 7098
rect 8927 7046 8939 7098
rect 8939 7046 8969 7098
rect 8993 7046 9003 7098
rect 9003 7046 9049 7098
rect 8753 7044 8809 7046
rect 8833 7044 8889 7046
rect 8913 7044 8969 7046
rect 8993 7044 9049 7046
rect 8753 6010 8809 6012
rect 8833 6010 8889 6012
rect 8913 6010 8969 6012
rect 8993 6010 9049 6012
rect 8753 5958 8799 6010
rect 8799 5958 8809 6010
rect 8833 5958 8863 6010
rect 8863 5958 8875 6010
rect 8875 5958 8889 6010
rect 8913 5958 8927 6010
rect 8927 5958 8939 6010
rect 8939 5958 8969 6010
rect 8993 5958 9003 6010
rect 9003 5958 9049 6010
rect 8753 5956 8809 5958
rect 8833 5956 8889 5958
rect 8913 5956 8969 5958
rect 8993 5956 9049 5958
rect 10598 7928 10654 7984
rect 9310 5752 9366 5808
rect 12070 15952 12126 16008
rect 12346 16632 12402 16688
rect 11352 7642 11408 7644
rect 11432 7642 11488 7644
rect 11512 7642 11568 7644
rect 11592 7642 11648 7644
rect 11352 7590 11398 7642
rect 11398 7590 11408 7642
rect 11432 7590 11462 7642
rect 11462 7590 11474 7642
rect 11474 7590 11488 7642
rect 11512 7590 11526 7642
rect 11526 7590 11538 7642
rect 11538 7590 11568 7642
rect 11592 7590 11602 7642
rect 11602 7590 11648 7642
rect 11352 7588 11408 7590
rect 11432 7588 11488 7590
rect 11512 7588 11568 7590
rect 11592 7588 11648 7590
rect 11352 6554 11408 6556
rect 11432 6554 11488 6556
rect 11512 6554 11568 6556
rect 11592 6554 11648 6556
rect 11352 6502 11398 6554
rect 11398 6502 11408 6554
rect 11432 6502 11462 6554
rect 11462 6502 11474 6554
rect 11474 6502 11488 6554
rect 11512 6502 11526 6554
rect 11526 6502 11538 6554
rect 11538 6502 11568 6554
rect 11592 6502 11602 6554
rect 11602 6502 11648 6554
rect 11352 6500 11408 6502
rect 11432 6500 11488 6502
rect 11512 6500 11568 6502
rect 11592 6500 11648 6502
rect 12806 14864 12862 14920
rect 12806 13776 12862 13832
rect 12806 12824 12862 12880
rect 13082 17584 13138 17640
rect 13174 17484 13176 17504
rect 13176 17484 13228 17504
rect 13228 17484 13230 17504
rect 13174 17448 13230 17484
rect 13082 16496 13138 16552
rect 12990 14864 13046 14920
rect 12254 11736 12310 11792
rect 12438 11192 12494 11248
rect 13951 20154 14007 20156
rect 14031 20154 14087 20156
rect 14111 20154 14167 20156
rect 14191 20154 14247 20156
rect 13951 20102 13997 20154
rect 13997 20102 14007 20154
rect 14031 20102 14061 20154
rect 14061 20102 14073 20154
rect 14073 20102 14087 20154
rect 14111 20102 14125 20154
rect 14125 20102 14137 20154
rect 14137 20102 14167 20154
rect 14191 20102 14201 20154
rect 14201 20102 14247 20154
rect 13951 20100 14007 20102
rect 14031 20100 14087 20102
rect 14111 20100 14167 20102
rect 14191 20100 14247 20102
rect 13951 19066 14007 19068
rect 14031 19066 14087 19068
rect 14111 19066 14167 19068
rect 14191 19066 14247 19068
rect 13951 19014 13997 19066
rect 13997 19014 14007 19066
rect 14031 19014 14061 19066
rect 14061 19014 14073 19066
rect 14073 19014 14087 19066
rect 14111 19014 14125 19066
rect 14125 19014 14137 19066
rect 14137 19014 14167 19066
rect 14191 19014 14201 19066
rect 14201 19014 14247 19066
rect 13951 19012 14007 19014
rect 14031 19012 14087 19014
rect 14111 19012 14167 19014
rect 14191 19012 14247 19014
rect 13951 17978 14007 17980
rect 14031 17978 14087 17980
rect 14111 17978 14167 17980
rect 14191 17978 14247 17980
rect 13951 17926 13997 17978
rect 13997 17926 14007 17978
rect 14031 17926 14061 17978
rect 14061 17926 14073 17978
rect 14073 17926 14087 17978
rect 14111 17926 14125 17978
rect 14125 17926 14137 17978
rect 14137 17926 14167 17978
rect 14191 17926 14201 17978
rect 14201 17926 14247 17978
rect 13951 17924 14007 17926
rect 14031 17924 14087 17926
rect 14111 17924 14167 17926
rect 14191 17924 14247 17926
rect 14370 17176 14426 17232
rect 13951 16890 14007 16892
rect 14031 16890 14087 16892
rect 14111 16890 14167 16892
rect 14191 16890 14247 16892
rect 13951 16838 13997 16890
rect 13997 16838 14007 16890
rect 14031 16838 14061 16890
rect 14061 16838 14073 16890
rect 14073 16838 14087 16890
rect 14111 16838 14125 16890
rect 14125 16838 14137 16890
rect 14137 16838 14167 16890
rect 14191 16838 14201 16890
rect 14201 16838 14247 16890
rect 13951 16836 14007 16838
rect 14031 16836 14087 16838
rect 14111 16836 14167 16838
rect 14191 16836 14247 16838
rect 13450 12688 13506 12744
rect 12898 10512 12954 10568
rect 13951 15802 14007 15804
rect 14031 15802 14087 15804
rect 14111 15802 14167 15804
rect 14191 15802 14247 15804
rect 13951 15750 13997 15802
rect 13997 15750 14007 15802
rect 14031 15750 14061 15802
rect 14061 15750 14073 15802
rect 14073 15750 14087 15802
rect 14111 15750 14125 15802
rect 14125 15750 14137 15802
rect 14137 15750 14167 15802
rect 14191 15750 14201 15802
rect 14201 15750 14247 15802
rect 13951 15748 14007 15750
rect 14031 15748 14087 15750
rect 14111 15748 14167 15750
rect 14191 15748 14247 15750
rect 13951 14714 14007 14716
rect 14031 14714 14087 14716
rect 14111 14714 14167 14716
rect 14191 14714 14247 14716
rect 13951 14662 13997 14714
rect 13997 14662 14007 14714
rect 14031 14662 14061 14714
rect 14061 14662 14073 14714
rect 14073 14662 14087 14714
rect 14111 14662 14125 14714
rect 14125 14662 14137 14714
rect 14137 14662 14167 14714
rect 14191 14662 14201 14714
rect 14201 14662 14247 14714
rect 13951 14660 14007 14662
rect 14031 14660 14087 14662
rect 14111 14660 14167 14662
rect 14191 14660 14247 14662
rect 13951 13626 14007 13628
rect 14031 13626 14087 13628
rect 14111 13626 14167 13628
rect 14191 13626 14247 13628
rect 13951 13574 13997 13626
rect 13997 13574 14007 13626
rect 14031 13574 14061 13626
rect 14061 13574 14073 13626
rect 14073 13574 14087 13626
rect 14111 13574 14125 13626
rect 14125 13574 14137 13626
rect 14137 13574 14167 13626
rect 14191 13574 14201 13626
rect 14201 13574 14247 13626
rect 13951 13572 14007 13574
rect 14031 13572 14087 13574
rect 14111 13572 14167 13574
rect 14191 13572 14247 13574
rect 13951 12538 14007 12540
rect 14031 12538 14087 12540
rect 14111 12538 14167 12540
rect 14191 12538 14247 12540
rect 13951 12486 13997 12538
rect 13997 12486 14007 12538
rect 14031 12486 14061 12538
rect 14061 12486 14073 12538
rect 14073 12486 14087 12538
rect 14111 12486 14125 12538
rect 14125 12486 14137 12538
rect 14137 12486 14167 12538
rect 14191 12486 14201 12538
rect 14201 12486 14247 12538
rect 13951 12484 14007 12486
rect 14031 12484 14087 12486
rect 14111 12484 14167 12486
rect 14191 12484 14247 12486
rect 13951 11450 14007 11452
rect 14031 11450 14087 11452
rect 14111 11450 14167 11452
rect 14191 11450 14247 11452
rect 13951 11398 13997 11450
rect 13997 11398 14007 11450
rect 14031 11398 14061 11450
rect 14061 11398 14073 11450
rect 14073 11398 14087 11450
rect 14111 11398 14125 11450
rect 14125 11398 14137 11450
rect 14137 11398 14167 11450
rect 14191 11398 14201 11450
rect 14201 11398 14247 11450
rect 13951 11396 14007 11398
rect 14031 11396 14087 11398
rect 14111 11396 14167 11398
rect 14191 11396 14247 11398
rect 15106 13368 15162 13424
rect 15842 20440 15898 20496
rect 16550 20698 16606 20700
rect 16630 20698 16686 20700
rect 16710 20698 16766 20700
rect 16790 20698 16846 20700
rect 16550 20646 16596 20698
rect 16596 20646 16606 20698
rect 16630 20646 16660 20698
rect 16660 20646 16672 20698
rect 16672 20646 16686 20698
rect 16710 20646 16724 20698
rect 16724 20646 16736 20698
rect 16736 20646 16766 20698
rect 16790 20646 16800 20698
rect 16800 20646 16846 20698
rect 16550 20644 16606 20646
rect 16630 20644 16686 20646
rect 16710 20644 16766 20646
rect 16790 20644 16846 20646
rect 16550 19610 16606 19612
rect 16630 19610 16686 19612
rect 16710 19610 16766 19612
rect 16790 19610 16846 19612
rect 16550 19558 16596 19610
rect 16596 19558 16606 19610
rect 16630 19558 16660 19610
rect 16660 19558 16672 19610
rect 16672 19558 16686 19610
rect 16710 19558 16724 19610
rect 16724 19558 16736 19610
rect 16736 19558 16766 19610
rect 16790 19558 16800 19610
rect 16800 19558 16846 19610
rect 16550 19556 16606 19558
rect 16630 19556 16686 19558
rect 16710 19556 16766 19558
rect 16790 19556 16846 19558
rect 16578 19216 16634 19272
rect 16550 18522 16606 18524
rect 16630 18522 16686 18524
rect 16710 18522 16766 18524
rect 16790 18522 16846 18524
rect 16550 18470 16596 18522
rect 16596 18470 16606 18522
rect 16630 18470 16660 18522
rect 16660 18470 16672 18522
rect 16672 18470 16686 18522
rect 16710 18470 16724 18522
rect 16724 18470 16736 18522
rect 16736 18470 16766 18522
rect 16790 18470 16800 18522
rect 16800 18470 16846 18522
rect 16550 18468 16606 18470
rect 16630 18468 16686 18470
rect 16710 18468 16766 18470
rect 16790 18468 16846 18470
rect 17222 18808 17278 18864
rect 19890 20440 19946 20496
rect 19614 20304 19670 20360
rect 19149 20154 19205 20156
rect 19229 20154 19285 20156
rect 19309 20154 19365 20156
rect 19389 20154 19445 20156
rect 19149 20102 19195 20154
rect 19195 20102 19205 20154
rect 19229 20102 19259 20154
rect 19259 20102 19271 20154
rect 19271 20102 19285 20154
rect 19309 20102 19323 20154
rect 19323 20102 19335 20154
rect 19335 20102 19365 20154
rect 19389 20102 19399 20154
rect 19399 20102 19445 20154
rect 19149 20100 19205 20102
rect 19229 20100 19285 20102
rect 19309 20100 19365 20102
rect 19389 20100 19445 20102
rect 20258 20052 20314 20088
rect 20258 20032 20260 20052
rect 20260 20032 20312 20052
rect 20312 20032 20314 20052
rect 20902 20848 20958 20904
rect 20350 19896 20406 19952
rect 18786 18672 18842 18728
rect 18694 18264 18750 18320
rect 17406 17720 17462 17776
rect 16550 17434 16606 17436
rect 16630 17434 16686 17436
rect 16710 17434 16766 17436
rect 16790 17434 16846 17436
rect 16550 17382 16596 17434
rect 16596 17382 16606 17434
rect 16630 17382 16660 17434
rect 16660 17382 16672 17434
rect 16672 17382 16686 17434
rect 16710 17382 16724 17434
rect 16724 17382 16736 17434
rect 16736 17382 16766 17434
rect 16790 17382 16800 17434
rect 16800 17382 16846 17434
rect 16550 17380 16606 17382
rect 16630 17380 16686 17382
rect 16710 17380 16766 17382
rect 16790 17380 16846 17382
rect 16550 16346 16606 16348
rect 16630 16346 16686 16348
rect 16710 16346 16766 16348
rect 16790 16346 16846 16348
rect 16550 16294 16596 16346
rect 16596 16294 16606 16346
rect 16630 16294 16660 16346
rect 16660 16294 16672 16346
rect 16672 16294 16686 16346
rect 16710 16294 16724 16346
rect 16724 16294 16736 16346
rect 16736 16294 16766 16346
rect 16790 16294 16800 16346
rect 16800 16294 16846 16346
rect 16550 16292 16606 16294
rect 16630 16292 16686 16294
rect 16710 16292 16766 16294
rect 16790 16292 16846 16294
rect 16118 15544 16174 15600
rect 15934 13368 15990 13424
rect 13951 10362 14007 10364
rect 14031 10362 14087 10364
rect 14111 10362 14167 10364
rect 14191 10362 14247 10364
rect 13951 10310 13997 10362
rect 13997 10310 14007 10362
rect 14031 10310 14061 10362
rect 14061 10310 14073 10362
rect 14073 10310 14087 10362
rect 14111 10310 14125 10362
rect 14125 10310 14137 10362
rect 14137 10310 14167 10362
rect 14191 10310 14201 10362
rect 14201 10310 14247 10362
rect 13951 10308 14007 10310
rect 14031 10308 14087 10310
rect 14111 10308 14167 10310
rect 14191 10308 14247 10310
rect 13951 9274 14007 9276
rect 14031 9274 14087 9276
rect 14111 9274 14167 9276
rect 14191 9274 14247 9276
rect 13951 9222 13997 9274
rect 13997 9222 14007 9274
rect 14031 9222 14061 9274
rect 14061 9222 14073 9274
rect 14073 9222 14087 9274
rect 14111 9222 14125 9274
rect 14125 9222 14137 9274
rect 14137 9222 14167 9274
rect 14191 9222 14201 9274
rect 14201 9222 14247 9274
rect 13951 9220 14007 9222
rect 14031 9220 14087 9222
rect 14111 9220 14167 9222
rect 14191 9220 14247 9222
rect 17314 17176 17370 17232
rect 18050 17040 18106 17096
rect 16550 15258 16606 15260
rect 16630 15258 16686 15260
rect 16710 15258 16766 15260
rect 16790 15258 16846 15260
rect 16550 15206 16596 15258
rect 16596 15206 16606 15258
rect 16630 15206 16660 15258
rect 16660 15206 16672 15258
rect 16672 15206 16686 15258
rect 16710 15206 16724 15258
rect 16724 15206 16736 15258
rect 16736 15206 16766 15258
rect 16790 15206 16800 15258
rect 16800 15206 16846 15258
rect 16550 15204 16606 15206
rect 16630 15204 16686 15206
rect 16710 15204 16766 15206
rect 16790 15204 16846 15206
rect 16550 14170 16606 14172
rect 16630 14170 16686 14172
rect 16710 14170 16766 14172
rect 16790 14170 16846 14172
rect 16550 14118 16596 14170
rect 16596 14118 16606 14170
rect 16630 14118 16660 14170
rect 16660 14118 16672 14170
rect 16672 14118 16686 14170
rect 16710 14118 16724 14170
rect 16724 14118 16736 14170
rect 16736 14118 16766 14170
rect 16790 14118 16800 14170
rect 16800 14118 16846 14170
rect 16550 14116 16606 14118
rect 16630 14116 16686 14118
rect 16710 14116 16766 14118
rect 16790 14116 16846 14118
rect 16550 13082 16606 13084
rect 16630 13082 16686 13084
rect 16710 13082 16766 13084
rect 16790 13082 16846 13084
rect 16550 13030 16596 13082
rect 16596 13030 16606 13082
rect 16630 13030 16660 13082
rect 16660 13030 16672 13082
rect 16672 13030 16686 13082
rect 16710 13030 16724 13082
rect 16724 13030 16736 13082
rect 16736 13030 16766 13082
rect 16790 13030 16800 13082
rect 16800 13030 16846 13082
rect 16550 13028 16606 13030
rect 16630 13028 16686 13030
rect 16710 13028 16766 13030
rect 16790 13028 16846 13030
rect 16550 11994 16606 11996
rect 16630 11994 16686 11996
rect 16710 11994 16766 11996
rect 16790 11994 16846 11996
rect 16550 11942 16596 11994
rect 16596 11942 16606 11994
rect 16630 11942 16660 11994
rect 16660 11942 16672 11994
rect 16672 11942 16686 11994
rect 16710 11942 16724 11994
rect 16724 11942 16736 11994
rect 16736 11942 16766 11994
rect 16790 11942 16800 11994
rect 16800 11942 16846 11994
rect 16550 11940 16606 11942
rect 16630 11940 16686 11942
rect 16710 11940 16766 11942
rect 16790 11940 16846 11942
rect 17130 13812 17132 13832
rect 17132 13812 17184 13832
rect 17184 13812 17186 13832
rect 17130 13776 17186 13812
rect 17038 11736 17094 11792
rect 15750 11192 15806 11248
rect 14554 9580 14610 9616
rect 14554 9560 14556 9580
rect 14556 9560 14608 9580
rect 14608 9560 14610 9580
rect 15290 9560 15346 9616
rect 16550 10906 16606 10908
rect 16630 10906 16686 10908
rect 16710 10906 16766 10908
rect 16790 10906 16846 10908
rect 16550 10854 16596 10906
rect 16596 10854 16606 10906
rect 16630 10854 16660 10906
rect 16660 10854 16672 10906
rect 16672 10854 16686 10906
rect 16710 10854 16724 10906
rect 16724 10854 16736 10906
rect 16736 10854 16766 10906
rect 16790 10854 16800 10906
rect 16800 10854 16846 10906
rect 16550 10852 16606 10854
rect 16630 10852 16686 10854
rect 16710 10852 16766 10854
rect 16790 10852 16846 10854
rect 16578 10124 16634 10160
rect 16578 10104 16580 10124
rect 16580 10104 16632 10124
rect 16632 10104 16634 10124
rect 17958 16088 18014 16144
rect 16550 9818 16606 9820
rect 16630 9818 16686 9820
rect 16710 9818 16766 9820
rect 16790 9818 16846 9820
rect 16550 9766 16596 9818
rect 16596 9766 16606 9818
rect 16630 9766 16660 9818
rect 16660 9766 16672 9818
rect 16672 9766 16686 9818
rect 16710 9766 16724 9818
rect 16724 9766 16736 9818
rect 16736 9766 16766 9818
rect 16790 9766 16800 9818
rect 16800 9766 16846 9818
rect 16550 9764 16606 9766
rect 16630 9764 16686 9766
rect 16710 9764 16766 9766
rect 16790 9764 16846 9766
rect 16394 9560 16450 9616
rect 16550 8730 16606 8732
rect 16630 8730 16686 8732
rect 16710 8730 16766 8732
rect 16790 8730 16846 8732
rect 16550 8678 16596 8730
rect 16596 8678 16606 8730
rect 16630 8678 16660 8730
rect 16660 8678 16672 8730
rect 16672 8678 16686 8730
rect 16710 8678 16724 8730
rect 16724 8678 16736 8730
rect 16736 8678 16766 8730
rect 16790 8678 16800 8730
rect 16800 8678 16846 8730
rect 16550 8676 16606 8678
rect 16630 8676 16686 8678
rect 16710 8676 16766 8678
rect 16790 8676 16846 8678
rect 13951 8186 14007 8188
rect 14031 8186 14087 8188
rect 14111 8186 14167 8188
rect 14191 8186 14247 8188
rect 13951 8134 13997 8186
rect 13997 8134 14007 8186
rect 14031 8134 14061 8186
rect 14061 8134 14073 8186
rect 14073 8134 14087 8186
rect 14111 8134 14125 8186
rect 14125 8134 14137 8186
rect 14137 8134 14167 8186
rect 14191 8134 14201 8186
rect 14201 8134 14247 8186
rect 13951 8132 14007 8134
rect 14031 8132 14087 8134
rect 14111 8132 14167 8134
rect 14191 8132 14247 8134
rect 17130 8608 17186 8664
rect 16550 7642 16606 7644
rect 16630 7642 16686 7644
rect 16710 7642 16766 7644
rect 16790 7642 16846 7644
rect 16550 7590 16596 7642
rect 16596 7590 16606 7642
rect 16630 7590 16660 7642
rect 16660 7590 16672 7642
rect 16672 7590 16686 7642
rect 16710 7590 16724 7642
rect 16724 7590 16736 7642
rect 16736 7590 16766 7642
rect 16790 7590 16800 7642
rect 16800 7590 16846 7642
rect 16550 7588 16606 7590
rect 16630 7588 16686 7590
rect 16710 7588 16766 7590
rect 16790 7588 16846 7590
rect 17498 8900 17554 8936
rect 17498 8880 17500 8900
rect 17500 8880 17552 8900
rect 17552 8880 17554 8900
rect 17774 11736 17830 11792
rect 17590 8780 17592 8800
rect 17592 8780 17644 8800
rect 17644 8780 17646 8800
rect 17590 8744 17646 8780
rect 17222 7928 17278 7984
rect 17866 10648 17922 10704
rect 17958 9424 18014 9480
rect 18142 16532 18144 16552
rect 18144 16532 18196 16552
rect 18196 16532 18198 16552
rect 18142 16496 18198 16532
rect 18418 15408 18474 15464
rect 18326 12144 18382 12200
rect 18234 10648 18290 10704
rect 18142 9596 18144 9616
rect 18144 9596 18196 9616
rect 18196 9596 18198 9616
rect 18142 9560 18198 9596
rect 13951 7098 14007 7100
rect 14031 7098 14087 7100
rect 14111 7098 14167 7100
rect 14191 7098 14247 7100
rect 13951 7046 13997 7098
rect 13997 7046 14007 7098
rect 14031 7046 14061 7098
rect 14061 7046 14073 7098
rect 14073 7046 14087 7098
rect 14111 7046 14125 7098
rect 14125 7046 14137 7098
rect 14137 7046 14167 7098
rect 14191 7046 14201 7098
rect 14201 7046 14247 7098
rect 13951 7044 14007 7046
rect 14031 7044 14087 7046
rect 14111 7044 14167 7046
rect 14191 7044 14247 7046
rect 14094 6296 14150 6352
rect 13951 6010 14007 6012
rect 14031 6010 14087 6012
rect 14111 6010 14167 6012
rect 14191 6010 14247 6012
rect 13951 5958 13997 6010
rect 13997 5958 14007 6010
rect 14031 5958 14061 6010
rect 14061 5958 14073 6010
rect 14073 5958 14087 6010
rect 14111 5958 14125 6010
rect 14125 5958 14137 6010
rect 14137 5958 14167 6010
rect 14191 5958 14201 6010
rect 14201 5958 14247 6010
rect 13951 5956 14007 5958
rect 14031 5956 14087 5958
rect 14111 5956 14167 5958
rect 14191 5956 14247 5958
rect 16550 6554 16606 6556
rect 16630 6554 16686 6556
rect 16710 6554 16766 6556
rect 16790 6554 16846 6556
rect 16550 6502 16596 6554
rect 16596 6502 16606 6554
rect 16630 6502 16660 6554
rect 16660 6502 16672 6554
rect 16672 6502 16686 6554
rect 16710 6502 16724 6554
rect 16724 6502 16736 6554
rect 16736 6502 16766 6554
rect 16790 6502 16800 6554
rect 16800 6502 16846 6554
rect 16550 6500 16606 6502
rect 16630 6500 16686 6502
rect 16710 6500 16766 6502
rect 16790 6500 16846 6502
rect 13082 5616 13138 5672
rect 11352 5466 11408 5468
rect 11432 5466 11488 5468
rect 11512 5466 11568 5468
rect 11592 5466 11648 5468
rect 11352 5414 11398 5466
rect 11398 5414 11408 5466
rect 11432 5414 11462 5466
rect 11462 5414 11474 5466
rect 11474 5414 11488 5466
rect 11512 5414 11526 5466
rect 11526 5414 11538 5466
rect 11538 5414 11568 5466
rect 11592 5414 11602 5466
rect 11602 5414 11648 5466
rect 11352 5412 11408 5414
rect 11432 5412 11488 5414
rect 11512 5412 11568 5414
rect 11592 5412 11648 5414
rect 16550 5466 16606 5468
rect 16630 5466 16686 5468
rect 16710 5466 16766 5468
rect 16790 5466 16846 5468
rect 16550 5414 16596 5466
rect 16596 5414 16606 5466
rect 16630 5414 16660 5466
rect 16660 5414 16672 5466
rect 16672 5414 16686 5466
rect 16710 5414 16724 5466
rect 16724 5414 16736 5466
rect 16736 5414 16766 5466
rect 16790 5414 16800 5466
rect 16800 5414 16846 5466
rect 16550 5412 16606 5414
rect 16630 5412 16686 5414
rect 16710 5412 16766 5414
rect 16790 5412 16846 5414
rect 8753 4922 8809 4924
rect 8833 4922 8889 4924
rect 8913 4922 8969 4924
rect 8993 4922 9049 4924
rect 8753 4870 8799 4922
rect 8799 4870 8809 4922
rect 8833 4870 8863 4922
rect 8863 4870 8875 4922
rect 8875 4870 8889 4922
rect 8913 4870 8927 4922
rect 8927 4870 8939 4922
rect 8939 4870 8969 4922
rect 8993 4870 9003 4922
rect 9003 4870 9049 4922
rect 8753 4868 8809 4870
rect 8833 4868 8889 4870
rect 8913 4868 8969 4870
rect 8993 4868 9049 4870
rect 13951 4922 14007 4924
rect 14031 4922 14087 4924
rect 14111 4922 14167 4924
rect 14191 4922 14247 4924
rect 13951 4870 13997 4922
rect 13997 4870 14007 4922
rect 14031 4870 14061 4922
rect 14061 4870 14073 4922
rect 14073 4870 14087 4922
rect 14111 4870 14125 4922
rect 14125 4870 14137 4922
rect 14137 4870 14167 4922
rect 14191 4870 14201 4922
rect 14201 4870 14247 4922
rect 13951 4868 14007 4870
rect 14031 4868 14087 4870
rect 14111 4868 14167 4870
rect 14191 4868 14247 4870
rect 11352 4378 11408 4380
rect 11432 4378 11488 4380
rect 11512 4378 11568 4380
rect 11592 4378 11648 4380
rect 11352 4326 11398 4378
rect 11398 4326 11408 4378
rect 11432 4326 11462 4378
rect 11462 4326 11474 4378
rect 11474 4326 11488 4378
rect 11512 4326 11526 4378
rect 11526 4326 11538 4378
rect 11538 4326 11568 4378
rect 11592 4326 11602 4378
rect 11602 4326 11648 4378
rect 11352 4324 11408 4326
rect 11432 4324 11488 4326
rect 11512 4324 11568 4326
rect 11592 4324 11648 4326
rect 16550 4378 16606 4380
rect 16630 4378 16686 4380
rect 16710 4378 16766 4380
rect 16790 4378 16846 4380
rect 16550 4326 16596 4378
rect 16596 4326 16606 4378
rect 16630 4326 16660 4378
rect 16660 4326 16672 4378
rect 16672 4326 16686 4378
rect 16710 4326 16724 4378
rect 16724 4326 16736 4378
rect 16736 4326 16766 4378
rect 16790 4326 16800 4378
rect 16800 4326 16846 4378
rect 16550 4324 16606 4326
rect 16630 4324 16686 4326
rect 16710 4324 16766 4326
rect 16790 4324 16846 4326
rect 18602 11600 18658 11656
rect 19149 19066 19205 19068
rect 19229 19066 19285 19068
rect 19309 19066 19365 19068
rect 19389 19066 19445 19068
rect 19149 19014 19195 19066
rect 19195 19014 19205 19066
rect 19229 19014 19259 19066
rect 19259 19014 19271 19066
rect 19271 19014 19285 19066
rect 19309 19014 19323 19066
rect 19323 19014 19335 19066
rect 19335 19014 19365 19066
rect 19389 19014 19399 19066
rect 19399 19014 19445 19066
rect 19149 19012 19205 19014
rect 19229 19012 19285 19014
rect 19309 19012 19365 19014
rect 19389 19012 19445 19014
rect 19149 17978 19205 17980
rect 19229 17978 19285 17980
rect 19309 17978 19365 17980
rect 19389 17978 19445 17980
rect 19149 17926 19195 17978
rect 19195 17926 19205 17978
rect 19229 17926 19259 17978
rect 19259 17926 19271 17978
rect 19271 17926 19285 17978
rect 19309 17926 19323 17978
rect 19323 17926 19335 17978
rect 19335 17926 19365 17978
rect 19389 17926 19399 17978
rect 19399 17926 19445 17978
rect 19149 17924 19205 17926
rect 19229 17924 19285 17926
rect 19309 17924 19365 17926
rect 19389 17924 19445 17926
rect 19149 16890 19205 16892
rect 19229 16890 19285 16892
rect 19309 16890 19365 16892
rect 19389 16890 19445 16892
rect 19149 16838 19195 16890
rect 19195 16838 19205 16890
rect 19229 16838 19259 16890
rect 19259 16838 19271 16890
rect 19271 16838 19285 16890
rect 19309 16838 19323 16890
rect 19323 16838 19335 16890
rect 19335 16838 19365 16890
rect 19389 16838 19399 16890
rect 19399 16838 19445 16890
rect 19149 16836 19205 16838
rect 19229 16836 19285 16838
rect 19309 16836 19365 16838
rect 19389 16836 19445 16838
rect 19149 15802 19205 15804
rect 19229 15802 19285 15804
rect 19309 15802 19365 15804
rect 19389 15802 19445 15804
rect 19149 15750 19195 15802
rect 19195 15750 19205 15802
rect 19229 15750 19259 15802
rect 19259 15750 19271 15802
rect 19271 15750 19285 15802
rect 19309 15750 19323 15802
rect 19323 15750 19335 15802
rect 19335 15750 19365 15802
rect 19389 15750 19399 15802
rect 19399 15750 19445 15802
rect 19149 15748 19205 15750
rect 19229 15748 19285 15750
rect 19309 15748 19365 15750
rect 19389 15748 19445 15750
rect 19149 14714 19205 14716
rect 19229 14714 19285 14716
rect 19309 14714 19365 14716
rect 19389 14714 19445 14716
rect 19149 14662 19195 14714
rect 19195 14662 19205 14714
rect 19229 14662 19259 14714
rect 19259 14662 19271 14714
rect 19271 14662 19285 14714
rect 19309 14662 19323 14714
rect 19323 14662 19335 14714
rect 19335 14662 19365 14714
rect 19389 14662 19399 14714
rect 19399 14662 19445 14714
rect 19149 14660 19205 14662
rect 19229 14660 19285 14662
rect 19309 14660 19365 14662
rect 19389 14660 19445 14662
rect 19149 13626 19205 13628
rect 19229 13626 19285 13628
rect 19309 13626 19365 13628
rect 19389 13626 19445 13628
rect 19149 13574 19195 13626
rect 19195 13574 19205 13626
rect 19229 13574 19259 13626
rect 19259 13574 19271 13626
rect 19271 13574 19285 13626
rect 19309 13574 19323 13626
rect 19323 13574 19335 13626
rect 19335 13574 19365 13626
rect 19389 13574 19399 13626
rect 19399 13574 19445 13626
rect 19149 13572 19205 13574
rect 19229 13572 19285 13574
rect 19309 13572 19365 13574
rect 19389 13572 19445 13574
rect 18970 13232 19026 13288
rect 18602 11192 18658 11248
rect 19149 12538 19205 12540
rect 19229 12538 19285 12540
rect 19309 12538 19365 12540
rect 19389 12538 19445 12540
rect 19149 12486 19195 12538
rect 19195 12486 19205 12538
rect 19229 12486 19259 12538
rect 19259 12486 19271 12538
rect 19271 12486 19285 12538
rect 19309 12486 19323 12538
rect 19323 12486 19335 12538
rect 19335 12486 19365 12538
rect 19389 12486 19399 12538
rect 19399 12486 19445 12538
rect 19149 12484 19205 12486
rect 19229 12484 19285 12486
rect 19309 12484 19365 12486
rect 19389 12484 19445 12486
rect 19149 11450 19205 11452
rect 19229 11450 19285 11452
rect 19309 11450 19365 11452
rect 19389 11450 19445 11452
rect 19149 11398 19195 11450
rect 19195 11398 19205 11450
rect 19229 11398 19259 11450
rect 19259 11398 19271 11450
rect 19271 11398 19285 11450
rect 19309 11398 19323 11450
rect 19323 11398 19335 11450
rect 19335 11398 19365 11450
rect 19389 11398 19399 11450
rect 19399 11398 19445 11450
rect 19149 11396 19205 11398
rect 19229 11396 19285 11398
rect 19309 11396 19365 11398
rect 19389 11396 19445 11398
rect 19246 11192 19302 11248
rect 19149 10362 19205 10364
rect 19229 10362 19285 10364
rect 19309 10362 19365 10364
rect 19389 10362 19445 10364
rect 19149 10310 19195 10362
rect 19195 10310 19205 10362
rect 19229 10310 19259 10362
rect 19259 10310 19271 10362
rect 19271 10310 19285 10362
rect 19309 10310 19323 10362
rect 19323 10310 19335 10362
rect 19335 10310 19365 10362
rect 19389 10310 19399 10362
rect 19399 10310 19445 10362
rect 19149 10308 19205 10310
rect 19229 10308 19285 10310
rect 19309 10308 19365 10310
rect 19389 10308 19445 10310
rect 19982 19760 20038 19816
rect 20626 18708 20628 18728
rect 20628 18708 20680 18728
rect 20680 18708 20682 18728
rect 20626 18672 20682 18708
rect 20166 15544 20222 15600
rect 19149 9274 19205 9276
rect 19229 9274 19285 9276
rect 19309 9274 19365 9276
rect 19389 9274 19445 9276
rect 19149 9222 19195 9274
rect 19195 9222 19205 9274
rect 19229 9222 19259 9274
rect 19259 9222 19271 9274
rect 19271 9222 19285 9274
rect 19309 9222 19323 9274
rect 19323 9222 19335 9274
rect 19335 9222 19365 9274
rect 19389 9222 19399 9274
rect 19399 9222 19445 9274
rect 19149 9220 19205 9222
rect 19229 9220 19285 9222
rect 19309 9220 19365 9222
rect 19389 9220 19445 9222
rect 19246 8608 19302 8664
rect 19246 8336 19302 8392
rect 19149 8186 19205 8188
rect 19229 8186 19285 8188
rect 19309 8186 19365 8188
rect 19389 8186 19445 8188
rect 19149 8134 19195 8186
rect 19195 8134 19205 8186
rect 19229 8134 19259 8186
rect 19259 8134 19271 8186
rect 19271 8134 19285 8186
rect 19309 8134 19323 8186
rect 19323 8134 19335 8186
rect 19335 8134 19365 8186
rect 19389 8134 19399 8186
rect 19399 8134 19445 8186
rect 19149 8132 19205 8134
rect 19229 8132 19285 8134
rect 19309 8132 19365 8134
rect 19389 8132 19445 8134
rect 19149 7098 19205 7100
rect 19229 7098 19285 7100
rect 19309 7098 19365 7100
rect 19389 7098 19445 7100
rect 19149 7046 19195 7098
rect 19195 7046 19205 7098
rect 19229 7046 19259 7098
rect 19259 7046 19271 7098
rect 19271 7046 19285 7098
rect 19309 7046 19323 7098
rect 19323 7046 19335 7098
rect 19335 7046 19365 7098
rect 19389 7046 19399 7098
rect 19399 7046 19445 7098
rect 19149 7044 19205 7046
rect 19229 7044 19285 7046
rect 19309 7044 19365 7046
rect 19389 7044 19445 7046
rect 18878 6704 18934 6760
rect 21546 21256 21602 21312
rect 20534 12164 20590 12200
rect 20534 12144 20536 12164
rect 20536 12144 20588 12164
rect 20588 12144 20590 12164
rect 21086 19216 21142 19272
rect 21086 17584 21142 17640
rect 21454 19760 21510 19816
rect 21748 20698 21804 20700
rect 21828 20698 21884 20700
rect 21908 20698 21964 20700
rect 21988 20698 22044 20700
rect 21748 20646 21794 20698
rect 21794 20646 21804 20698
rect 21828 20646 21858 20698
rect 21858 20646 21870 20698
rect 21870 20646 21884 20698
rect 21908 20646 21922 20698
rect 21922 20646 21934 20698
rect 21934 20646 21964 20698
rect 21988 20646 21998 20698
rect 21998 20646 22044 20698
rect 21748 20644 21804 20646
rect 21828 20644 21884 20646
rect 21908 20644 21964 20646
rect 21988 20644 22044 20646
rect 21748 19610 21804 19612
rect 21828 19610 21884 19612
rect 21908 19610 21964 19612
rect 21988 19610 22044 19612
rect 21748 19558 21794 19610
rect 21794 19558 21804 19610
rect 21828 19558 21858 19610
rect 21858 19558 21870 19610
rect 21870 19558 21884 19610
rect 21908 19558 21922 19610
rect 21922 19558 21934 19610
rect 21934 19558 21964 19610
rect 21988 19558 21998 19610
rect 21998 19558 22044 19610
rect 21748 19556 21804 19558
rect 21828 19556 21884 19558
rect 21908 19556 21964 19558
rect 21988 19556 22044 19558
rect 21454 18808 21510 18864
rect 21748 18522 21804 18524
rect 21828 18522 21884 18524
rect 21908 18522 21964 18524
rect 21988 18522 22044 18524
rect 21748 18470 21794 18522
rect 21794 18470 21804 18522
rect 21828 18470 21858 18522
rect 21858 18470 21870 18522
rect 21870 18470 21884 18522
rect 21908 18470 21922 18522
rect 21922 18470 21934 18522
rect 21934 18470 21964 18522
rect 21988 18470 21998 18522
rect 21998 18470 22044 18522
rect 21748 18468 21804 18470
rect 21828 18468 21884 18470
rect 21908 18468 21964 18470
rect 21988 18468 22044 18470
rect 21454 18264 21510 18320
rect 21362 18128 21418 18184
rect 21454 18028 21456 18048
rect 21456 18028 21508 18048
rect 21508 18028 21510 18048
rect 21454 17992 21510 18028
rect 21086 15972 21142 16008
rect 21086 15952 21088 15972
rect 21088 15952 21140 15972
rect 21140 15952 21142 15972
rect 21748 17434 21804 17436
rect 21828 17434 21884 17436
rect 21908 17434 21964 17436
rect 21988 17434 22044 17436
rect 21748 17382 21794 17434
rect 21794 17382 21804 17434
rect 21828 17382 21858 17434
rect 21858 17382 21870 17434
rect 21870 17382 21884 17434
rect 21908 17382 21922 17434
rect 21922 17382 21934 17434
rect 21934 17382 21964 17434
rect 21988 17382 21998 17434
rect 21998 17382 22044 17434
rect 21748 17380 21804 17382
rect 21828 17380 21884 17382
rect 21908 17380 21964 17382
rect 21988 17380 22044 17382
rect 21454 17176 21510 17232
rect 21454 16768 21510 16824
rect 21454 16496 21510 16552
rect 21748 16346 21804 16348
rect 21828 16346 21884 16348
rect 21908 16346 21964 16348
rect 21988 16346 22044 16348
rect 21748 16294 21794 16346
rect 21794 16294 21804 16346
rect 21828 16294 21858 16346
rect 21858 16294 21870 16346
rect 21870 16294 21884 16346
rect 21908 16294 21922 16346
rect 21922 16294 21934 16346
rect 21934 16294 21964 16346
rect 21988 16294 21998 16346
rect 21998 16294 22044 16346
rect 21748 16292 21804 16294
rect 21828 16292 21884 16294
rect 21908 16292 21964 16294
rect 21988 16292 22044 16294
rect 20718 12708 20774 12744
rect 20718 12688 20720 12708
rect 20720 12688 20772 12708
rect 20772 12688 20774 12708
rect 20534 10104 20590 10160
rect 20718 9968 20774 10024
rect 20074 8880 20130 8936
rect 19982 8744 20038 8800
rect 19149 6010 19205 6012
rect 19229 6010 19285 6012
rect 19309 6010 19365 6012
rect 19389 6010 19445 6012
rect 19149 5958 19195 6010
rect 19195 5958 19205 6010
rect 19229 5958 19259 6010
rect 19259 5958 19271 6010
rect 19271 5958 19285 6010
rect 19309 5958 19323 6010
rect 19323 5958 19335 6010
rect 19335 5958 19365 6010
rect 19389 5958 19399 6010
rect 19399 5958 19445 6010
rect 19149 5956 19205 5958
rect 19229 5956 19285 5958
rect 19309 5956 19365 5958
rect 19389 5956 19445 5958
rect 19149 4922 19205 4924
rect 19229 4922 19285 4924
rect 19309 4922 19365 4924
rect 19389 4922 19445 4924
rect 19149 4870 19195 4922
rect 19195 4870 19205 4922
rect 19229 4870 19259 4922
rect 19259 4870 19271 4922
rect 19271 4870 19285 4922
rect 19309 4870 19323 4922
rect 19323 4870 19335 4922
rect 19335 4870 19365 4922
rect 19389 4870 19399 4922
rect 19399 4870 19445 4922
rect 19149 4868 19205 4870
rect 19229 4868 19285 4870
rect 19309 4868 19365 4870
rect 19389 4868 19445 4870
rect 8753 3834 8809 3836
rect 8833 3834 8889 3836
rect 8913 3834 8969 3836
rect 8993 3834 9049 3836
rect 8753 3782 8799 3834
rect 8799 3782 8809 3834
rect 8833 3782 8863 3834
rect 8863 3782 8875 3834
rect 8875 3782 8889 3834
rect 8913 3782 8927 3834
rect 8927 3782 8939 3834
rect 8939 3782 8969 3834
rect 8993 3782 9003 3834
rect 9003 3782 9049 3834
rect 8753 3780 8809 3782
rect 8833 3780 8889 3782
rect 8913 3780 8969 3782
rect 8993 3780 9049 3782
rect 13951 3834 14007 3836
rect 14031 3834 14087 3836
rect 14111 3834 14167 3836
rect 14191 3834 14247 3836
rect 13951 3782 13997 3834
rect 13997 3782 14007 3834
rect 14031 3782 14061 3834
rect 14061 3782 14073 3834
rect 14073 3782 14087 3834
rect 14111 3782 14125 3834
rect 14125 3782 14137 3834
rect 14137 3782 14167 3834
rect 14191 3782 14201 3834
rect 14201 3782 14247 3834
rect 13951 3780 14007 3782
rect 14031 3780 14087 3782
rect 14111 3780 14167 3782
rect 14191 3780 14247 3782
rect 19149 3834 19205 3836
rect 19229 3834 19285 3836
rect 19309 3834 19365 3836
rect 19389 3834 19445 3836
rect 19149 3782 19195 3834
rect 19195 3782 19205 3834
rect 19229 3782 19259 3834
rect 19259 3782 19271 3834
rect 19271 3782 19285 3834
rect 19309 3782 19323 3834
rect 19323 3782 19335 3834
rect 19335 3782 19365 3834
rect 19389 3782 19399 3834
rect 19399 3782 19445 3834
rect 19149 3780 19205 3782
rect 19229 3780 19285 3782
rect 19309 3780 19365 3782
rect 19389 3780 19445 3782
rect 11352 3290 11408 3292
rect 11432 3290 11488 3292
rect 11512 3290 11568 3292
rect 11592 3290 11648 3292
rect 11352 3238 11398 3290
rect 11398 3238 11408 3290
rect 11432 3238 11462 3290
rect 11462 3238 11474 3290
rect 11474 3238 11488 3290
rect 11512 3238 11526 3290
rect 11526 3238 11538 3290
rect 11538 3238 11568 3290
rect 11592 3238 11602 3290
rect 11602 3238 11648 3290
rect 11352 3236 11408 3238
rect 11432 3236 11488 3238
rect 11512 3236 11568 3238
rect 11592 3236 11648 3238
rect 16550 3290 16606 3292
rect 16630 3290 16686 3292
rect 16710 3290 16766 3292
rect 16790 3290 16846 3292
rect 16550 3238 16596 3290
rect 16596 3238 16606 3290
rect 16630 3238 16660 3290
rect 16660 3238 16672 3290
rect 16672 3238 16686 3290
rect 16710 3238 16724 3290
rect 16724 3238 16736 3290
rect 16736 3238 16766 3290
rect 16790 3238 16800 3290
rect 16800 3238 16846 3290
rect 16550 3236 16606 3238
rect 16630 3236 16686 3238
rect 16710 3236 16766 3238
rect 16790 3236 16846 3238
rect 8753 2746 8809 2748
rect 8833 2746 8889 2748
rect 8913 2746 8969 2748
rect 8993 2746 9049 2748
rect 8753 2694 8799 2746
rect 8799 2694 8809 2746
rect 8833 2694 8863 2746
rect 8863 2694 8875 2746
rect 8875 2694 8889 2746
rect 8913 2694 8927 2746
rect 8927 2694 8939 2746
rect 8939 2694 8969 2746
rect 8993 2694 9003 2746
rect 9003 2694 9049 2746
rect 8753 2692 8809 2694
rect 8833 2692 8889 2694
rect 8913 2692 8969 2694
rect 8993 2692 9049 2694
rect 13951 2746 14007 2748
rect 14031 2746 14087 2748
rect 14111 2746 14167 2748
rect 14191 2746 14247 2748
rect 13951 2694 13997 2746
rect 13997 2694 14007 2746
rect 14031 2694 14061 2746
rect 14061 2694 14073 2746
rect 14073 2694 14087 2746
rect 14111 2694 14125 2746
rect 14125 2694 14137 2746
rect 14137 2694 14167 2746
rect 14191 2694 14201 2746
rect 14201 2694 14247 2746
rect 13951 2692 14007 2694
rect 14031 2692 14087 2694
rect 14111 2692 14167 2694
rect 14191 2692 14247 2694
rect 16854 2916 16910 2952
rect 16854 2896 16856 2916
rect 16856 2896 16908 2916
rect 16908 2896 16910 2916
rect 20258 7928 20314 7984
rect 20626 8472 20682 8528
rect 21086 14320 21142 14376
rect 20994 13368 21050 13424
rect 21086 12280 21142 12336
rect 20994 11092 20996 11112
rect 20996 11092 21048 11112
rect 21048 11092 21050 11112
rect 20994 11056 21050 11092
rect 21086 10648 21142 10704
rect 20994 9036 21050 9072
rect 20994 9016 20996 9036
rect 20996 9016 21048 9036
rect 21048 9016 21050 9036
rect 20626 7384 20682 7440
rect 20718 6976 20774 7032
rect 20810 6740 20812 6760
rect 20812 6740 20864 6760
rect 20864 6740 20866 6760
rect 20810 6704 20866 6740
rect 20718 6196 20720 6216
rect 20720 6196 20772 6216
rect 20772 6196 20774 6216
rect 20718 6160 20774 6196
rect 21454 15544 21510 15600
rect 21546 15000 21602 15056
rect 21454 14764 21456 14784
rect 21456 14764 21508 14784
rect 21508 14764 21510 14784
rect 21454 14728 21510 14764
rect 21454 13912 21510 13968
rect 21454 13504 21510 13560
rect 21546 13268 21548 13288
rect 21548 13268 21600 13288
rect 21600 13268 21602 13288
rect 21546 13232 21602 13268
rect 21748 15258 21804 15260
rect 21828 15258 21884 15260
rect 21908 15258 21964 15260
rect 21988 15258 22044 15260
rect 21748 15206 21794 15258
rect 21794 15206 21804 15258
rect 21828 15206 21858 15258
rect 21858 15206 21870 15258
rect 21870 15206 21884 15258
rect 21908 15206 21922 15258
rect 21922 15206 21934 15258
rect 21934 15206 21964 15258
rect 21988 15206 21998 15258
rect 21998 15206 22044 15258
rect 21748 15204 21804 15206
rect 21828 15204 21884 15206
rect 21908 15204 21964 15206
rect 21988 15204 22044 15206
rect 21748 14170 21804 14172
rect 21828 14170 21884 14172
rect 21908 14170 21964 14172
rect 21988 14170 22044 14172
rect 21748 14118 21794 14170
rect 21794 14118 21804 14170
rect 21828 14118 21858 14170
rect 21858 14118 21870 14170
rect 21870 14118 21884 14170
rect 21908 14118 21922 14170
rect 21922 14118 21934 14170
rect 21934 14118 21964 14170
rect 21988 14118 21998 14170
rect 21998 14118 22044 14170
rect 21748 14116 21804 14118
rect 21828 14116 21884 14118
rect 21908 14116 21964 14118
rect 21988 14116 22044 14118
rect 21748 13082 21804 13084
rect 21828 13082 21884 13084
rect 21908 13082 21964 13084
rect 21988 13082 22044 13084
rect 21748 13030 21794 13082
rect 21794 13030 21804 13082
rect 21828 13030 21858 13082
rect 21858 13030 21870 13082
rect 21870 13030 21884 13082
rect 21908 13030 21922 13082
rect 21922 13030 21934 13082
rect 21934 13030 21964 13082
rect 21988 13030 21998 13082
rect 21998 13030 22044 13082
rect 21748 13028 21804 13030
rect 21828 13028 21884 13030
rect 21908 13028 21964 13030
rect 21988 13028 22044 13030
rect 21454 12688 21510 12744
rect 21454 11736 21510 11792
rect 21546 11464 21602 11520
rect 21454 11092 21456 11112
rect 21456 11092 21508 11112
rect 21508 11092 21510 11112
rect 21454 11056 21510 11092
rect 21362 10512 21418 10568
rect 21454 10240 21510 10296
rect 21748 11994 21804 11996
rect 21828 11994 21884 11996
rect 21908 11994 21964 11996
rect 21988 11994 22044 11996
rect 21748 11942 21794 11994
rect 21794 11942 21804 11994
rect 21828 11942 21858 11994
rect 21858 11942 21870 11994
rect 21870 11942 21884 11994
rect 21908 11942 21922 11994
rect 21922 11942 21934 11994
rect 21934 11942 21964 11994
rect 21988 11942 21998 11994
rect 21998 11942 22044 11994
rect 21748 11940 21804 11942
rect 21828 11940 21884 11942
rect 21908 11940 21964 11942
rect 21988 11940 22044 11942
rect 21748 10906 21804 10908
rect 21828 10906 21884 10908
rect 21908 10906 21964 10908
rect 21988 10906 22044 10908
rect 21748 10854 21794 10906
rect 21794 10854 21804 10906
rect 21828 10854 21858 10906
rect 21858 10854 21870 10906
rect 21870 10854 21884 10906
rect 21908 10854 21922 10906
rect 21922 10854 21934 10906
rect 21934 10854 21964 10906
rect 21988 10854 21998 10906
rect 21998 10854 22044 10906
rect 21748 10852 21804 10854
rect 21828 10852 21884 10854
rect 21908 10852 21964 10854
rect 21988 10852 22044 10854
rect 21748 9818 21804 9820
rect 21828 9818 21884 9820
rect 21908 9818 21964 9820
rect 21988 9818 22044 9820
rect 21748 9766 21794 9818
rect 21794 9766 21804 9818
rect 21828 9766 21858 9818
rect 21858 9766 21870 9818
rect 21870 9766 21884 9818
rect 21908 9766 21922 9818
rect 21922 9766 21934 9818
rect 21934 9766 21964 9818
rect 21988 9766 21998 9818
rect 21998 9766 22044 9818
rect 21748 9764 21804 9766
rect 21828 9764 21884 9766
rect 21908 9764 21964 9766
rect 21988 9764 22044 9766
rect 21454 9424 21510 9480
rect 21546 9016 21602 9072
rect 21748 8730 21804 8732
rect 21828 8730 21884 8732
rect 21908 8730 21964 8732
rect 21988 8730 22044 8732
rect 21748 8678 21794 8730
rect 21794 8678 21804 8730
rect 21828 8678 21858 8730
rect 21858 8678 21870 8730
rect 21870 8678 21884 8730
rect 21908 8678 21922 8730
rect 21922 8678 21934 8730
rect 21934 8678 21964 8730
rect 21988 8678 21998 8730
rect 21998 8678 22044 8730
rect 21748 8676 21804 8678
rect 21828 8676 21884 8678
rect 21908 8676 21964 8678
rect 21988 8676 22044 8678
rect 21454 7792 21510 7848
rect 21748 7642 21804 7644
rect 21828 7642 21884 7644
rect 21908 7642 21964 7644
rect 21988 7642 22044 7644
rect 21748 7590 21794 7642
rect 21794 7590 21804 7642
rect 21828 7590 21858 7642
rect 21858 7590 21870 7642
rect 21870 7590 21884 7642
rect 21908 7590 21922 7642
rect 21922 7590 21934 7642
rect 21934 7590 21964 7642
rect 21988 7590 21998 7642
rect 21998 7590 22044 7642
rect 21748 7588 21804 7590
rect 21828 7588 21884 7590
rect 21908 7588 21964 7590
rect 21988 7588 22044 7590
rect 21748 6554 21804 6556
rect 21828 6554 21884 6556
rect 21908 6554 21964 6556
rect 21988 6554 22044 6556
rect 21748 6502 21794 6554
rect 21794 6502 21804 6554
rect 21828 6502 21858 6554
rect 21858 6502 21870 6554
rect 21870 6502 21884 6554
rect 21908 6502 21922 6554
rect 21922 6502 21934 6554
rect 21934 6502 21964 6554
rect 21988 6502 21998 6554
rect 21998 6502 22044 6554
rect 21748 6500 21804 6502
rect 21828 6500 21884 6502
rect 21908 6500 21964 6502
rect 21988 6500 22044 6502
rect 21178 6296 21234 6352
rect 21546 5752 21602 5808
rect 21748 5466 21804 5468
rect 21828 5466 21884 5468
rect 21908 5466 21964 5468
rect 21988 5466 22044 5468
rect 21748 5414 21794 5466
rect 21794 5414 21804 5466
rect 21828 5414 21858 5466
rect 21858 5414 21870 5466
rect 21870 5414 21884 5466
rect 21908 5414 21922 5466
rect 21922 5414 21934 5466
rect 21934 5414 21964 5466
rect 21988 5414 21998 5466
rect 21998 5414 22044 5466
rect 21748 5412 21804 5414
rect 21828 5412 21884 5414
rect 21908 5412 21964 5414
rect 21988 5412 22044 5414
rect 21270 5208 21326 5264
rect 21546 4936 21602 4992
rect 21546 4528 21602 4584
rect 20718 4120 20774 4176
rect 21748 4378 21804 4380
rect 21828 4378 21884 4380
rect 21908 4378 21964 4380
rect 21988 4378 22044 4380
rect 21748 4326 21794 4378
rect 21794 4326 21804 4378
rect 21828 4326 21858 4378
rect 21858 4326 21870 4378
rect 21870 4326 21884 4378
rect 21908 4326 21922 4378
rect 21922 4326 21934 4378
rect 21934 4326 21964 4378
rect 21988 4326 21998 4378
rect 21998 4326 22044 4378
rect 21748 4324 21804 4326
rect 21828 4324 21884 4326
rect 21908 4324 21964 4326
rect 21988 4324 22044 4326
rect 21270 3712 21326 3768
rect 21546 3476 21548 3496
rect 21548 3476 21600 3496
rect 21600 3476 21602 3496
rect 21546 3440 21602 3476
rect 21748 3290 21804 3292
rect 21828 3290 21884 3292
rect 21908 3290 21964 3292
rect 21988 3290 22044 3292
rect 21748 3238 21794 3290
rect 21794 3238 21804 3290
rect 21828 3238 21858 3290
rect 21858 3238 21870 3290
rect 21870 3238 21884 3290
rect 21908 3238 21922 3290
rect 21922 3238 21934 3290
rect 21934 3238 21964 3290
rect 21988 3238 21998 3290
rect 21998 3238 22044 3290
rect 21748 3236 21804 3238
rect 21828 3236 21884 3238
rect 21908 3236 21964 3238
rect 21988 3236 22044 3238
rect 19149 2746 19205 2748
rect 19229 2746 19285 2748
rect 19309 2746 19365 2748
rect 19389 2746 19445 2748
rect 19149 2694 19195 2746
rect 19195 2694 19205 2746
rect 19229 2694 19259 2746
rect 19259 2694 19271 2746
rect 19271 2694 19285 2746
rect 19309 2694 19323 2746
rect 19323 2694 19335 2746
rect 19335 2694 19365 2746
rect 19389 2694 19399 2746
rect 19399 2694 19445 2746
rect 19149 2692 19205 2694
rect 19229 2692 19285 2694
rect 19309 2692 19365 2694
rect 19389 2692 19445 2694
rect 21546 2896 21602 2952
rect 21270 2488 21326 2544
rect 6154 2202 6210 2204
rect 6234 2202 6290 2204
rect 6314 2202 6370 2204
rect 6394 2202 6450 2204
rect 6154 2150 6200 2202
rect 6200 2150 6210 2202
rect 6234 2150 6264 2202
rect 6264 2150 6276 2202
rect 6276 2150 6290 2202
rect 6314 2150 6328 2202
rect 6328 2150 6340 2202
rect 6340 2150 6370 2202
rect 6394 2150 6404 2202
rect 6404 2150 6450 2202
rect 6154 2148 6210 2150
rect 6234 2148 6290 2150
rect 6314 2148 6370 2150
rect 6394 2148 6450 2150
rect 2778 1672 2834 1728
rect 11352 2202 11408 2204
rect 11432 2202 11488 2204
rect 11512 2202 11568 2204
rect 11592 2202 11648 2204
rect 11352 2150 11398 2202
rect 11398 2150 11408 2202
rect 11432 2150 11462 2202
rect 11462 2150 11474 2202
rect 11474 2150 11488 2202
rect 11512 2150 11526 2202
rect 11526 2150 11538 2202
rect 11538 2150 11568 2202
rect 11592 2150 11602 2202
rect 11602 2150 11648 2202
rect 11352 2148 11408 2150
rect 11432 2148 11488 2150
rect 11512 2148 11568 2150
rect 11592 2148 11648 2150
rect 16550 2202 16606 2204
rect 16630 2202 16686 2204
rect 16710 2202 16766 2204
rect 16790 2202 16846 2204
rect 16550 2150 16596 2202
rect 16596 2150 16606 2202
rect 16630 2150 16660 2202
rect 16660 2150 16672 2202
rect 16672 2150 16686 2202
rect 16710 2150 16724 2202
rect 16724 2150 16736 2202
rect 16736 2150 16766 2202
rect 16790 2150 16800 2202
rect 16800 2150 16846 2202
rect 16550 2148 16606 2150
rect 16630 2148 16686 2150
rect 16710 2148 16766 2150
rect 16790 2148 16846 2150
rect 21270 1944 21326 2000
rect 21748 2202 21804 2204
rect 21828 2202 21884 2204
rect 21908 2202 21964 2204
rect 21988 2202 22044 2204
rect 21748 2150 21794 2202
rect 21794 2150 21804 2202
rect 21828 2150 21858 2202
rect 21858 2150 21870 2202
rect 21870 2150 21884 2202
rect 21908 2150 21922 2202
rect 21922 2150 21934 2202
rect 21934 2150 21964 2202
rect 21988 2150 21998 2202
rect 21998 2150 22044 2202
rect 21748 2148 21804 2150
rect 21828 2148 21884 2150
rect 21908 2148 21964 2150
rect 21988 2148 22044 2150
rect 21546 1672 21602 1728
<< metal3 >>
rect 0 21314 800 21344
rect 3049 21314 3115 21317
rect 0 21312 3115 21314
rect 0 21256 3054 21312
rect 3110 21256 3115 21312
rect 0 21254 3115 21256
rect 0 21224 800 21254
rect 3049 21251 3115 21254
rect 21541 21314 21607 21317
rect 22200 21314 23000 21344
rect 21541 21312 23000 21314
rect 21541 21256 21546 21312
rect 21602 21256 23000 21312
rect 21541 21254 23000 21256
rect 21541 21251 21607 21254
rect 22200 21224 23000 21254
rect 0 20906 800 20936
rect 2773 20906 2839 20909
rect 0 20904 2839 20906
rect 0 20848 2778 20904
rect 2834 20848 2839 20904
rect 0 20846 2839 20848
rect 0 20816 800 20846
rect 2773 20843 2839 20846
rect 20897 20906 20963 20909
rect 22200 20906 23000 20936
rect 20897 20904 23000 20906
rect 20897 20848 20902 20904
rect 20958 20848 23000 20904
rect 20897 20846 23000 20848
rect 20897 20843 20963 20846
rect 22200 20816 23000 20846
rect 6144 20704 6460 20705
rect 6144 20640 6150 20704
rect 6214 20640 6230 20704
rect 6294 20640 6310 20704
rect 6374 20640 6390 20704
rect 6454 20640 6460 20704
rect 6144 20639 6460 20640
rect 11342 20704 11658 20705
rect 11342 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11658 20704
rect 11342 20639 11658 20640
rect 16540 20704 16856 20705
rect 16540 20640 16546 20704
rect 16610 20640 16626 20704
rect 16690 20640 16706 20704
rect 16770 20640 16786 20704
rect 16850 20640 16856 20704
rect 16540 20639 16856 20640
rect 21738 20704 22054 20705
rect 21738 20640 21744 20704
rect 21808 20640 21824 20704
rect 21888 20640 21904 20704
rect 21968 20640 21984 20704
rect 22048 20640 22054 20704
rect 21738 20639 22054 20640
rect 0 20498 800 20528
rect 1853 20498 1919 20501
rect 0 20496 1919 20498
rect 0 20440 1858 20496
rect 1914 20440 1919 20496
rect 0 20438 1919 20440
rect 0 20408 800 20438
rect 1853 20435 1919 20438
rect 5349 20498 5415 20501
rect 15837 20498 15903 20501
rect 5349 20496 15903 20498
rect 5349 20440 5354 20496
rect 5410 20440 15842 20496
rect 15898 20440 15903 20496
rect 5349 20438 15903 20440
rect 5349 20435 5415 20438
rect 15837 20435 15903 20438
rect 19885 20498 19951 20501
rect 22200 20498 23000 20528
rect 19885 20496 23000 20498
rect 19885 20440 19890 20496
rect 19946 20440 23000 20496
rect 19885 20438 23000 20440
rect 19885 20435 19951 20438
rect 22200 20408 23000 20438
rect 3325 20362 3391 20365
rect 19609 20362 19675 20365
rect 3325 20360 19675 20362
rect 3325 20304 3330 20360
rect 3386 20304 19614 20360
rect 19670 20304 19675 20360
rect 3325 20302 19675 20304
rect 3325 20299 3391 20302
rect 19609 20299 19675 20302
rect 4889 20226 4955 20229
rect 5022 20226 5028 20228
rect 4889 20224 5028 20226
rect 4889 20168 4894 20224
rect 4950 20168 5028 20224
rect 4889 20166 5028 20168
rect 4889 20163 4955 20166
rect 5022 20164 5028 20166
rect 5092 20164 5098 20228
rect 3545 20160 3861 20161
rect 0 20090 800 20120
rect 3545 20096 3551 20160
rect 3615 20096 3631 20160
rect 3695 20096 3711 20160
rect 3775 20096 3791 20160
rect 3855 20096 3861 20160
rect 3545 20095 3861 20096
rect 8743 20160 9059 20161
rect 8743 20096 8749 20160
rect 8813 20096 8829 20160
rect 8893 20096 8909 20160
rect 8973 20096 8989 20160
rect 9053 20096 9059 20160
rect 8743 20095 9059 20096
rect 13941 20160 14257 20161
rect 13941 20096 13947 20160
rect 14011 20096 14027 20160
rect 14091 20096 14107 20160
rect 14171 20096 14187 20160
rect 14251 20096 14257 20160
rect 13941 20095 14257 20096
rect 19139 20160 19455 20161
rect 19139 20096 19145 20160
rect 19209 20096 19225 20160
rect 19289 20096 19305 20160
rect 19369 20096 19385 20160
rect 19449 20096 19455 20160
rect 19139 20095 19455 20096
rect 1485 20090 1551 20093
rect 0 20088 1551 20090
rect 0 20032 1490 20088
rect 1546 20032 1551 20088
rect 0 20030 1551 20032
rect 0 20000 800 20030
rect 1485 20027 1551 20030
rect 3969 20090 4035 20093
rect 8201 20092 8267 20093
rect 8150 20090 8156 20092
rect 3969 20088 6562 20090
rect 3969 20032 3974 20088
rect 4030 20032 6562 20088
rect 3969 20030 6562 20032
rect 8110 20030 8156 20090
rect 8220 20088 8267 20092
rect 8262 20032 8267 20088
rect 3969 20027 4035 20030
rect 5942 19892 5948 19956
rect 6012 19954 6018 19956
rect 6361 19954 6427 19957
rect 6012 19952 6427 19954
rect 6012 19896 6366 19952
rect 6422 19896 6427 19952
rect 6012 19894 6427 19896
rect 6502 19954 6562 20030
rect 8150 20028 8156 20030
rect 8220 20028 8267 20032
rect 8201 20027 8267 20028
rect 20253 20090 20319 20093
rect 22200 20090 23000 20120
rect 20253 20088 23000 20090
rect 20253 20032 20258 20088
rect 20314 20032 23000 20088
rect 20253 20030 23000 20032
rect 20253 20027 20319 20030
rect 22200 20000 23000 20030
rect 20345 19954 20411 19957
rect 6502 19952 20411 19954
rect 6502 19896 20350 19952
rect 20406 19896 20411 19952
rect 6502 19894 20411 19896
rect 6012 19892 6018 19894
rect 6361 19891 6427 19894
rect 20345 19891 20411 19894
rect 4429 19818 4495 19821
rect 19977 19818 20043 19821
rect 4429 19816 20043 19818
rect 4429 19760 4434 19816
rect 4490 19760 19982 19816
rect 20038 19760 20043 19816
rect 4429 19758 20043 19760
rect 4429 19755 4495 19758
rect 19977 19755 20043 19758
rect 21449 19818 21515 19821
rect 21449 19816 22202 19818
rect 21449 19760 21454 19816
rect 21510 19760 22202 19816
rect 21449 19758 22202 19760
rect 21449 19755 21515 19758
rect 22142 19712 22202 19758
rect 0 19682 800 19712
rect 1485 19682 1551 19685
rect 0 19680 1551 19682
rect 0 19624 1490 19680
rect 1546 19624 1551 19680
rect 0 19622 1551 19624
rect 0 19592 800 19622
rect 1485 19619 1551 19622
rect 7281 19682 7347 19685
rect 8937 19682 9003 19685
rect 9673 19682 9739 19685
rect 7281 19680 9003 19682
rect 7281 19624 7286 19680
rect 7342 19624 8942 19680
rect 8998 19624 9003 19680
rect 7281 19622 9003 19624
rect 7281 19619 7347 19622
rect 8937 19619 9003 19622
rect 9630 19680 9739 19682
rect 9630 19624 9678 19680
rect 9734 19624 9739 19680
rect 9630 19619 9739 19624
rect 22142 19622 23000 19712
rect 6144 19616 6460 19617
rect 6144 19552 6150 19616
rect 6214 19552 6230 19616
rect 6294 19552 6310 19616
rect 6374 19552 6390 19616
rect 6454 19552 6460 19616
rect 6144 19551 6460 19552
rect 7097 19546 7163 19549
rect 7925 19546 7991 19549
rect 8109 19546 8175 19549
rect 7097 19544 7666 19546
rect 7097 19488 7102 19544
rect 7158 19488 7666 19544
rect 7097 19486 7666 19488
rect 7097 19483 7163 19486
rect 3785 19410 3851 19413
rect 3918 19410 3924 19412
rect 3785 19408 3924 19410
rect 3785 19352 3790 19408
rect 3846 19352 3924 19408
rect 3785 19350 3924 19352
rect 3785 19347 3851 19350
rect 3918 19348 3924 19350
rect 3988 19348 3994 19412
rect 7281 19410 7347 19413
rect 4110 19408 7347 19410
rect 4110 19352 7286 19408
rect 7342 19352 7347 19408
rect 4110 19350 7347 19352
rect 7606 19410 7666 19486
rect 7925 19544 8175 19546
rect 7925 19488 7930 19544
rect 7986 19488 8114 19544
rect 8170 19488 8175 19544
rect 7925 19486 8175 19488
rect 7925 19483 7991 19486
rect 8109 19483 8175 19486
rect 8293 19548 8359 19549
rect 8293 19544 8340 19548
rect 8404 19546 8410 19548
rect 8293 19488 8298 19544
rect 8293 19484 8340 19488
rect 8404 19486 8450 19546
rect 8404 19484 8410 19486
rect 8293 19483 8359 19484
rect 8293 19410 8359 19413
rect 7606 19408 8359 19410
rect 7606 19352 8298 19408
rect 8354 19352 8359 19408
rect 7606 19350 8359 19352
rect 0 19274 800 19304
rect 1853 19274 1919 19277
rect 0 19272 1919 19274
rect 0 19216 1858 19272
rect 1914 19216 1919 19272
rect 0 19214 1919 19216
rect 0 19184 800 19214
rect 1853 19211 1919 19214
rect 2865 19274 2931 19277
rect 4110 19274 4170 19350
rect 7281 19347 7347 19350
rect 8293 19347 8359 19350
rect 2865 19272 4170 19274
rect 2865 19216 2870 19272
rect 2926 19216 4170 19272
rect 2865 19214 4170 19216
rect 8293 19274 8359 19277
rect 9630 19274 9690 19619
rect 11342 19616 11658 19617
rect 11342 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11658 19616
rect 11342 19551 11658 19552
rect 16540 19616 16856 19617
rect 16540 19552 16546 19616
rect 16610 19552 16626 19616
rect 16690 19552 16706 19616
rect 16770 19552 16786 19616
rect 16850 19552 16856 19616
rect 16540 19551 16856 19552
rect 21738 19616 22054 19617
rect 21738 19552 21744 19616
rect 21808 19552 21824 19616
rect 21888 19552 21904 19616
rect 21968 19552 21984 19616
rect 22048 19552 22054 19616
rect 22200 19592 23000 19622
rect 21738 19551 22054 19552
rect 11830 19348 11836 19412
rect 11900 19410 11906 19412
rect 11973 19410 12039 19413
rect 11900 19408 12039 19410
rect 11900 19352 11978 19408
rect 12034 19352 12039 19408
rect 11900 19350 12039 19352
rect 11900 19348 11906 19350
rect 11973 19347 12039 19350
rect 16573 19274 16639 19277
rect 8293 19272 9690 19274
rect 8293 19216 8298 19272
rect 8354 19216 9690 19272
rect 8293 19214 9690 19216
rect 9814 19272 16639 19274
rect 9814 19216 16578 19272
rect 16634 19216 16639 19272
rect 9814 19214 16639 19216
rect 2865 19211 2931 19214
rect 8293 19211 8359 19214
rect 4153 19140 4219 19141
rect 4102 19076 4108 19140
rect 4172 19138 4219 19140
rect 5533 19138 5599 19141
rect 4172 19136 5599 19138
rect 4214 19080 5538 19136
rect 5594 19080 5599 19136
rect 4172 19078 5599 19080
rect 4172 19076 4219 19078
rect 4153 19075 4219 19076
rect 5533 19075 5599 19078
rect 7966 19076 7972 19140
rect 8036 19138 8042 19140
rect 8109 19138 8175 19141
rect 8036 19136 8175 19138
rect 8036 19080 8114 19136
rect 8170 19080 8175 19136
rect 8036 19078 8175 19080
rect 8036 19076 8042 19078
rect 8109 19075 8175 19078
rect 3545 19072 3861 19073
rect 3545 19008 3551 19072
rect 3615 19008 3631 19072
rect 3695 19008 3711 19072
rect 3775 19008 3791 19072
rect 3855 19008 3861 19072
rect 3545 19007 3861 19008
rect 8743 19072 9059 19073
rect 8743 19008 8749 19072
rect 8813 19008 8829 19072
rect 8893 19008 8909 19072
rect 8973 19008 8989 19072
rect 9053 19008 9059 19072
rect 8743 19007 9059 19008
rect 3233 19002 3299 19005
rect 3190 19000 3299 19002
rect 3190 18944 3238 19000
rect 3294 18944 3299 19000
rect 3190 18939 3299 18944
rect 0 18866 800 18896
rect 1485 18866 1551 18869
rect 0 18864 1551 18866
rect 0 18808 1490 18864
rect 1546 18808 1551 18864
rect 0 18806 1551 18808
rect 0 18776 800 18806
rect 1485 18803 1551 18806
rect 3190 18730 3250 18939
rect 5022 18804 5028 18868
rect 5092 18866 5098 18868
rect 9814 18866 9874 19214
rect 16573 19211 16639 19214
rect 21081 19274 21147 19277
rect 22200 19274 23000 19304
rect 21081 19272 23000 19274
rect 21081 19216 21086 19272
rect 21142 19216 23000 19272
rect 21081 19214 23000 19216
rect 21081 19211 21147 19214
rect 22200 19184 23000 19214
rect 13941 19072 14257 19073
rect 13941 19008 13947 19072
rect 14011 19008 14027 19072
rect 14091 19008 14107 19072
rect 14171 19008 14187 19072
rect 14251 19008 14257 19072
rect 13941 19007 14257 19008
rect 19139 19072 19455 19073
rect 19139 19008 19145 19072
rect 19209 19008 19225 19072
rect 19289 19008 19305 19072
rect 19369 19008 19385 19072
rect 19449 19008 19455 19072
rect 19139 19007 19455 19008
rect 10777 19002 10843 19005
rect 11329 19002 11395 19005
rect 10777 19000 11395 19002
rect 10777 18944 10782 19000
rect 10838 18944 11334 19000
rect 11390 18944 11395 19000
rect 10777 18942 11395 18944
rect 10777 18939 10843 18942
rect 11329 18939 11395 18942
rect 5092 18806 9874 18866
rect 10041 18866 10107 18869
rect 17217 18866 17283 18869
rect 10041 18864 17283 18866
rect 10041 18808 10046 18864
rect 10102 18808 17222 18864
rect 17278 18808 17283 18864
rect 10041 18806 17283 18808
rect 5092 18804 5098 18806
rect 10041 18803 10107 18806
rect 17217 18803 17283 18806
rect 21449 18866 21515 18869
rect 22200 18866 23000 18896
rect 21449 18864 23000 18866
rect 21449 18808 21454 18864
rect 21510 18808 23000 18864
rect 21449 18806 23000 18808
rect 21449 18803 21515 18806
rect 22200 18776 23000 18806
rect 3325 18730 3391 18733
rect 3190 18728 3391 18730
rect 3190 18672 3330 18728
rect 3386 18672 3391 18728
rect 3190 18670 3391 18672
rect 3325 18667 3391 18670
rect 3509 18730 3575 18733
rect 18781 18730 18847 18733
rect 3509 18728 18847 18730
rect 3509 18672 3514 18728
rect 3570 18672 18786 18728
rect 18842 18672 18847 18728
rect 3509 18670 18847 18672
rect 3509 18667 3575 18670
rect 18781 18667 18847 18670
rect 20478 18668 20484 18732
rect 20548 18730 20554 18732
rect 20621 18730 20687 18733
rect 20548 18728 20687 18730
rect 20548 18672 20626 18728
rect 20682 18672 20687 18728
rect 20548 18670 20687 18672
rect 20548 18668 20554 18670
rect 20621 18667 20687 18670
rect 6545 18594 6611 18597
rect 10041 18594 10107 18597
rect 6545 18592 10107 18594
rect 6545 18536 6550 18592
rect 6606 18536 10046 18592
rect 10102 18536 10107 18592
rect 6545 18534 10107 18536
rect 6545 18531 6611 18534
rect 10041 18531 10107 18534
rect 6144 18528 6460 18529
rect 0 18458 800 18488
rect 6144 18464 6150 18528
rect 6214 18464 6230 18528
rect 6294 18464 6310 18528
rect 6374 18464 6390 18528
rect 6454 18464 6460 18528
rect 6144 18463 6460 18464
rect 11342 18528 11658 18529
rect 11342 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11658 18528
rect 11342 18463 11658 18464
rect 16540 18528 16856 18529
rect 16540 18464 16546 18528
rect 16610 18464 16626 18528
rect 16690 18464 16706 18528
rect 16770 18464 16786 18528
rect 16850 18464 16856 18528
rect 16540 18463 16856 18464
rect 21738 18528 22054 18529
rect 21738 18464 21744 18528
rect 21808 18464 21824 18528
rect 21888 18464 21904 18528
rect 21968 18464 21984 18528
rect 22048 18464 22054 18528
rect 21738 18463 22054 18464
rect 1485 18458 1551 18461
rect 22200 18458 23000 18488
rect 0 18456 1551 18458
rect 0 18400 1490 18456
rect 1546 18400 1551 18456
rect 0 18398 1551 18400
rect 0 18368 800 18398
rect 1485 18395 1551 18398
rect 22142 18368 23000 18458
rect 2773 18322 2839 18325
rect 18689 18322 18755 18325
rect 2773 18320 18755 18322
rect 2773 18264 2778 18320
rect 2834 18264 18694 18320
rect 18750 18264 18755 18320
rect 2773 18262 18755 18264
rect 2773 18259 2839 18262
rect 18689 18259 18755 18262
rect 21449 18322 21515 18325
rect 22142 18322 22202 18368
rect 21449 18320 22202 18322
rect 21449 18264 21454 18320
rect 21510 18264 22202 18320
rect 21449 18262 22202 18264
rect 21449 18259 21515 18262
rect 2681 18186 2747 18189
rect 21357 18186 21423 18189
rect 2681 18184 21423 18186
rect 2681 18128 2686 18184
rect 2742 18128 21362 18184
rect 21418 18128 21423 18184
rect 2681 18126 21423 18128
rect 2681 18123 2747 18126
rect 21357 18123 21423 18126
rect 0 18050 800 18080
rect 1485 18050 1551 18053
rect 0 18048 1551 18050
rect 0 17992 1490 18048
rect 1546 17992 1551 18048
rect 0 17990 1551 17992
rect 0 17960 800 17990
rect 1485 17987 1551 17990
rect 4061 18050 4127 18053
rect 6545 18050 6611 18053
rect 4061 18048 6611 18050
rect 4061 17992 4066 18048
rect 4122 17992 6550 18048
rect 6606 17992 6611 18048
rect 4061 17990 6611 17992
rect 4061 17987 4127 17990
rect 6545 17987 6611 17990
rect 8293 18050 8359 18053
rect 8518 18050 8524 18052
rect 8293 18048 8524 18050
rect 8293 17992 8298 18048
rect 8354 17992 8524 18048
rect 8293 17990 8524 17992
rect 8293 17987 8359 17990
rect 8518 17988 8524 17990
rect 8588 17988 8594 18052
rect 21449 18050 21515 18053
rect 22200 18050 23000 18080
rect 21449 18048 23000 18050
rect 21449 17992 21454 18048
rect 21510 17992 23000 18048
rect 21449 17990 23000 17992
rect 21449 17987 21515 17990
rect 3545 17984 3861 17985
rect 3545 17920 3551 17984
rect 3615 17920 3631 17984
rect 3695 17920 3711 17984
rect 3775 17920 3791 17984
rect 3855 17920 3861 17984
rect 3545 17919 3861 17920
rect 8743 17984 9059 17985
rect 8743 17920 8749 17984
rect 8813 17920 8829 17984
rect 8893 17920 8909 17984
rect 8973 17920 8989 17984
rect 9053 17920 9059 17984
rect 8743 17919 9059 17920
rect 13941 17984 14257 17985
rect 13941 17920 13947 17984
rect 14011 17920 14027 17984
rect 14091 17920 14107 17984
rect 14171 17920 14187 17984
rect 14251 17920 14257 17984
rect 13941 17919 14257 17920
rect 19139 17984 19455 17985
rect 19139 17920 19145 17984
rect 19209 17920 19225 17984
rect 19289 17920 19305 17984
rect 19369 17920 19385 17984
rect 19449 17920 19455 17984
rect 22200 17960 23000 17990
rect 19139 17919 19455 17920
rect 10133 17778 10199 17781
rect 17401 17778 17467 17781
rect 10133 17776 17467 17778
rect 10133 17720 10138 17776
rect 10194 17720 17406 17776
rect 17462 17720 17467 17776
rect 10133 17718 17467 17720
rect 10133 17715 10199 17718
rect 17401 17715 17467 17718
rect 0 17642 800 17672
rect 1853 17642 1919 17645
rect 0 17640 1919 17642
rect 0 17584 1858 17640
rect 1914 17584 1919 17640
rect 0 17582 1919 17584
rect 0 17552 800 17582
rect 1853 17579 1919 17582
rect 12157 17642 12223 17645
rect 13077 17642 13143 17645
rect 12157 17640 13143 17642
rect 12157 17584 12162 17640
rect 12218 17584 13082 17640
rect 13138 17584 13143 17640
rect 12157 17582 13143 17584
rect 12157 17579 12223 17582
rect 13077 17579 13143 17582
rect 21081 17642 21147 17645
rect 22200 17642 23000 17672
rect 21081 17640 23000 17642
rect 21081 17584 21086 17640
rect 21142 17584 23000 17640
rect 21081 17582 23000 17584
rect 21081 17579 21147 17582
rect 22200 17552 23000 17582
rect 9397 17506 9463 17509
rect 10593 17506 10659 17509
rect 9397 17504 10659 17506
rect 9397 17448 9402 17504
rect 9458 17448 10598 17504
rect 10654 17448 10659 17504
rect 9397 17446 10659 17448
rect 9397 17443 9463 17446
rect 10593 17443 10659 17446
rect 11789 17506 11855 17509
rect 13169 17506 13235 17509
rect 11789 17504 13235 17506
rect 11789 17448 11794 17504
rect 11850 17448 13174 17504
rect 13230 17448 13235 17504
rect 11789 17446 13235 17448
rect 11789 17443 11855 17446
rect 13169 17443 13235 17446
rect 6144 17440 6460 17441
rect 6144 17376 6150 17440
rect 6214 17376 6230 17440
rect 6294 17376 6310 17440
rect 6374 17376 6390 17440
rect 6454 17376 6460 17440
rect 6144 17375 6460 17376
rect 11342 17440 11658 17441
rect 11342 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11658 17440
rect 11342 17375 11658 17376
rect 16540 17440 16856 17441
rect 16540 17376 16546 17440
rect 16610 17376 16626 17440
rect 16690 17376 16706 17440
rect 16770 17376 16786 17440
rect 16850 17376 16856 17440
rect 16540 17375 16856 17376
rect 21738 17440 22054 17441
rect 21738 17376 21744 17440
rect 21808 17376 21824 17440
rect 21888 17376 21904 17440
rect 21968 17376 21984 17440
rect 22048 17376 22054 17440
rect 21738 17375 22054 17376
rect 0 17234 800 17264
rect 1485 17234 1551 17237
rect 0 17232 1551 17234
rect 0 17176 1490 17232
rect 1546 17176 1551 17232
rect 0 17174 1551 17176
rect 0 17144 800 17174
rect 1485 17171 1551 17174
rect 11605 17234 11671 17237
rect 14365 17234 14431 17237
rect 17309 17234 17375 17237
rect 11605 17232 17375 17234
rect 11605 17176 11610 17232
rect 11666 17176 14370 17232
rect 14426 17176 17314 17232
rect 17370 17176 17375 17232
rect 11605 17174 17375 17176
rect 11605 17171 11671 17174
rect 14365 17171 14431 17174
rect 17309 17171 17375 17174
rect 21449 17234 21515 17237
rect 22200 17234 23000 17264
rect 21449 17232 23000 17234
rect 21449 17176 21454 17232
rect 21510 17176 23000 17232
rect 21449 17174 23000 17176
rect 21449 17171 21515 17174
rect 22200 17144 23000 17174
rect 9765 17098 9831 17101
rect 10593 17098 10659 17101
rect 18045 17098 18111 17101
rect 9765 17096 18111 17098
rect 9765 17040 9770 17096
rect 9826 17040 10598 17096
rect 10654 17040 18050 17096
rect 18106 17040 18111 17096
rect 9765 17038 18111 17040
rect 9765 17035 9831 17038
rect 10593 17035 10659 17038
rect 18045 17035 18111 17038
rect 3545 16896 3861 16897
rect 0 16826 800 16856
rect 3545 16832 3551 16896
rect 3615 16832 3631 16896
rect 3695 16832 3711 16896
rect 3775 16832 3791 16896
rect 3855 16832 3861 16896
rect 3545 16831 3861 16832
rect 8743 16896 9059 16897
rect 8743 16832 8749 16896
rect 8813 16832 8829 16896
rect 8893 16832 8909 16896
rect 8973 16832 8989 16896
rect 9053 16832 9059 16896
rect 8743 16831 9059 16832
rect 13941 16896 14257 16897
rect 13941 16832 13947 16896
rect 14011 16832 14027 16896
rect 14091 16832 14107 16896
rect 14171 16832 14187 16896
rect 14251 16832 14257 16896
rect 13941 16831 14257 16832
rect 19139 16896 19455 16897
rect 19139 16832 19145 16896
rect 19209 16832 19225 16896
rect 19289 16832 19305 16896
rect 19369 16832 19385 16896
rect 19449 16832 19455 16896
rect 19139 16831 19455 16832
rect 1485 16826 1551 16829
rect 0 16824 1551 16826
rect 0 16768 1490 16824
rect 1546 16768 1551 16824
rect 0 16766 1551 16768
rect 0 16736 800 16766
rect 1485 16763 1551 16766
rect 21449 16826 21515 16829
rect 22200 16826 23000 16856
rect 21449 16824 23000 16826
rect 21449 16768 21454 16824
rect 21510 16768 23000 16824
rect 21449 16766 23000 16768
rect 21449 16763 21515 16766
rect 22200 16736 23000 16766
rect 11881 16690 11947 16693
rect 12341 16690 12407 16693
rect 11881 16688 12407 16690
rect 11881 16632 11886 16688
rect 11942 16632 12346 16688
rect 12402 16632 12407 16688
rect 11881 16630 12407 16632
rect 11881 16627 11947 16630
rect 12341 16627 12407 16630
rect 1761 16554 1827 16557
rect 2405 16554 2471 16557
rect 1761 16552 2471 16554
rect 1761 16496 1766 16552
rect 1822 16496 2410 16552
rect 2466 16496 2471 16552
rect 1761 16494 2471 16496
rect 1761 16491 1827 16494
rect 2405 16491 2471 16494
rect 13077 16554 13143 16557
rect 18137 16554 18203 16557
rect 13077 16552 18203 16554
rect 13077 16496 13082 16552
rect 13138 16496 18142 16552
rect 18198 16496 18203 16552
rect 13077 16494 18203 16496
rect 13077 16491 13143 16494
rect 18137 16491 18203 16494
rect 21449 16554 21515 16557
rect 21449 16552 22202 16554
rect 21449 16496 21454 16552
rect 21510 16496 22202 16552
rect 21449 16494 22202 16496
rect 21449 16491 21515 16494
rect 22142 16448 22202 16494
rect 0 16418 800 16448
rect 1485 16418 1551 16421
rect 0 16416 1551 16418
rect 0 16360 1490 16416
rect 1546 16360 1551 16416
rect 0 16358 1551 16360
rect 22142 16358 23000 16448
rect 0 16328 800 16358
rect 1485 16355 1551 16358
rect 6144 16352 6460 16353
rect 6144 16288 6150 16352
rect 6214 16288 6230 16352
rect 6294 16288 6310 16352
rect 6374 16288 6390 16352
rect 6454 16288 6460 16352
rect 6144 16287 6460 16288
rect 11342 16352 11658 16353
rect 11342 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11658 16352
rect 11342 16287 11658 16288
rect 16540 16352 16856 16353
rect 16540 16288 16546 16352
rect 16610 16288 16626 16352
rect 16690 16288 16706 16352
rect 16770 16288 16786 16352
rect 16850 16288 16856 16352
rect 16540 16287 16856 16288
rect 21738 16352 22054 16353
rect 21738 16288 21744 16352
rect 21808 16288 21824 16352
rect 21888 16288 21904 16352
rect 21968 16288 21984 16352
rect 22048 16288 22054 16352
rect 22200 16328 23000 16358
rect 21738 16287 22054 16288
rect 2773 16146 2839 16149
rect 3877 16146 3943 16149
rect 17953 16146 18019 16149
rect 2773 16144 18019 16146
rect 2773 16088 2778 16144
rect 2834 16088 3882 16144
rect 3938 16088 17958 16144
rect 18014 16088 18019 16144
rect 2773 16086 18019 16088
rect 2773 16083 2839 16086
rect 3877 16083 3943 16086
rect 17953 16083 18019 16086
rect 0 16010 800 16040
rect 1853 16010 1919 16013
rect 0 16008 1919 16010
rect 0 15952 1858 16008
rect 1914 15952 1919 16008
rect 0 15950 1919 15952
rect 0 15920 800 15950
rect 1853 15947 1919 15950
rect 2313 16010 2379 16013
rect 12065 16010 12131 16013
rect 2313 16008 12131 16010
rect 2313 15952 2318 16008
rect 2374 15952 12070 16008
rect 12126 15952 12131 16008
rect 2313 15950 12131 15952
rect 2313 15947 2379 15950
rect 12065 15947 12131 15950
rect 21081 16010 21147 16013
rect 22200 16010 23000 16040
rect 21081 16008 23000 16010
rect 21081 15952 21086 16008
rect 21142 15952 23000 16008
rect 21081 15950 23000 15952
rect 21081 15947 21147 15950
rect 22200 15920 23000 15950
rect 3545 15808 3861 15809
rect 3545 15744 3551 15808
rect 3615 15744 3631 15808
rect 3695 15744 3711 15808
rect 3775 15744 3791 15808
rect 3855 15744 3861 15808
rect 3545 15743 3861 15744
rect 8743 15808 9059 15809
rect 8743 15744 8749 15808
rect 8813 15744 8829 15808
rect 8893 15744 8909 15808
rect 8973 15744 8989 15808
rect 9053 15744 9059 15808
rect 8743 15743 9059 15744
rect 13941 15808 14257 15809
rect 13941 15744 13947 15808
rect 14011 15744 14027 15808
rect 14091 15744 14107 15808
rect 14171 15744 14187 15808
rect 14251 15744 14257 15808
rect 13941 15743 14257 15744
rect 19139 15808 19455 15809
rect 19139 15744 19145 15808
rect 19209 15744 19225 15808
rect 19289 15744 19305 15808
rect 19369 15744 19385 15808
rect 19449 15744 19455 15808
rect 19139 15743 19455 15744
rect 0 15602 800 15632
rect 1485 15602 1551 15605
rect 0 15600 1551 15602
rect 0 15544 1490 15600
rect 1546 15544 1551 15600
rect 0 15542 1551 15544
rect 0 15512 800 15542
rect 1485 15539 1551 15542
rect 4429 15602 4495 15605
rect 9213 15602 9279 15605
rect 4429 15600 9279 15602
rect 4429 15544 4434 15600
rect 4490 15544 9218 15600
rect 9274 15544 9279 15600
rect 4429 15542 9279 15544
rect 4429 15539 4495 15542
rect 9213 15539 9279 15542
rect 10593 15602 10659 15605
rect 16113 15602 16179 15605
rect 20161 15602 20227 15605
rect 10593 15600 20227 15602
rect 10593 15544 10598 15600
rect 10654 15544 16118 15600
rect 16174 15544 20166 15600
rect 20222 15544 20227 15600
rect 10593 15542 20227 15544
rect 10593 15539 10659 15542
rect 16113 15539 16179 15542
rect 20161 15539 20227 15542
rect 21449 15602 21515 15605
rect 22200 15602 23000 15632
rect 21449 15600 23000 15602
rect 21449 15544 21454 15600
rect 21510 15544 23000 15600
rect 21449 15542 23000 15544
rect 21449 15539 21515 15542
rect 22200 15512 23000 15542
rect 6545 15466 6611 15469
rect 18413 15466 18479 15469
rect 6545 15464 18479 15466
rect 6545 15408 6550 15464
rect 6606 15408 18418 15464
rect 18474 15408 18479 15464
rect 6545 15406 18479 15408
rect 6545 15403 6611 15406
rect 18413 15403 18479 15406
rect 6144 15264 6460 15265
rect 0 15194 800 15224
rect 6144 15200 6150 15264
rect 6214 15200 6230 15264
rect 6294 15200 6310 15264
rect 6374 15200 6390 15264
rect 6454 15200 6460 15264
rect 6144 15199 6460 15200
rect 11342 15264 11658 15265
rect 11342 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11658 15264
rect 11342 15199 11658 15200
rect 16540 15264 16856 15265
rect 16540 15200 16546 15264
rect 16610 15200 16626 15264
rect 16690 15200 16706 15264
rect 16770 15200 16786 15264
rect 16850 15200 16856 15264
rect 16540 15199 16856 15200
rect 21738 15264 22054 15265
rect 21738 15200 21744 15264
rect 21808 15200 21824 15264
rect 21888 15200 21904 15264
rect 21968 15200 21984 15264
rect 22048 15200 22054 15264
rect 21738 15199 22054 15200
rect 1485 15194 1551 15197
rect 22200 15194 23000 15224
rect 0 15192 1551 15194
rect 0 15136 1490 15192
rect 1546 15136 1551 15192
rect 0 15134 1551 15136
rect 0 15104 800 15134
rect 1485 15131 1551 15134
rect 22142 15104 23000 15194
rect 21541 15058 21607 15061
rect 22142 15058 22202 15104
rect 21541 15056 22202 15058
rect 21541 15000 21546 15056
rect 21602 15000 22202 15056
rect 21541 14998 22202 15000
rect 21541 14995 21607 14998
rect 12801 14922 12867 14925
rect 12985 14922 13051 14925
rect 12801 14920 13051 14922
rect 12801 14864 12806 14920
rect 12862 14864 12990 14920
rect 13046 14864 13051 14920
rect 12801 14862 13051 14864
rect 12801 14859 12867 14862
rect 12985 14859 13051 14862
rect 0 14786 800 14816
rect 1485 14786 1551 14789
rect 0 14784 1551 14786
rect 0 14728 1490 14784
rect 1546 14728 1551 14784
rect 0 14726 1551 14728
rect 0 14696 800 14726
rect 1485 14723 1551 14726
rect 21449 14786 21515 14789
rect 22200 14786 23000 14816
rect 21449 14784 23000 14786
rect 21449 14728 21454 14784
rect 21510 14728 23000 14784
rect 21449 14726 23000 14728
rect 21449 14723 21515 14726
rect 3545 14720 3861 14721
rect 3545 14656 3551 14720
rect 3615 14656 3631 14720
rect 3695 14656 3711 14720
rect 3775 14656 3791 14720
rect 3855 14656 3861 14720
rect 3545 14655 3861 14656
rect 8743 14720 9059 14721
rect 8743 14656 8749 14720
rect 8813 14656 8829 14720
rect 8893 14656 8909 14720
rect 8973 14656 8989 14720
rect 9053 14656 9059 14720
rect 8743 14655 9059 14656
rect 13941 14720 14257 14721
rect 13941 14656 13947 14720
rect 14011 14656 14027 14720
rect 14091 14656 14107 14720
rect 14171 14656 14187 14720
rect 14251 14656 14257 14720
rect 13941 14655 14257 14656
rect 19139 14720 19455 14721
rect 19139 14656 19145 14720
rect 19209 14656 19225 14720
rect 19289 14656 19305 14720
rect 19369 14656 19385 14720
rect 19449 14656 19455 14720
rect 22200 14696 23000 14726
rect 19139 14655 19455 14656
rect 0 14378 800 14408
rect 1853 14378 1919 14381
rect 0 14376 1919 14378
rect 0 14320 1858 14376
rect 1914 14320 1919 14376
rect 0 14318 1919 14320
rect 0 14288 800 14318
rect 1853 14315 1919 14318
rect 21081 14378 21147 14381
rect 22200 14378 23000 14408
rect 21081 14376 23000 14378
rect 21081 14320 21086 14376
rect 21142 14320 23000 14376
rect 21081 14318 23000 14320
rect 21081 14315 21147 14318
rect 22200 14288 23000 14318
rect 6144 14176 6460 14177
rect 6144 14112 6150 14176
rect 6214 14112 6230 14176
rect 6294 14112 6310 14176
rect 6374 14112 6390 14176
rect 6454 14112 6460 14176
rect 6144 14111 6460 14112
rect 11342 14176 11658 14177
rect 11342 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11658 14176
rect 11342 14111 11658 14112
rect 16540 14176 16856 14177
rect 16540 14112 16546 14176
rect 16610 14112 16626 14176
rect 16690 14112 16706 14176
rect 16770 14112 16786 14176
rect 16850 14112 16856 14176
rect 16540 14111 16856 14112
rect 21738 14176 22054 14177
rect 21738 14112 21744 14176
rect 21808 14112 21824 14176
rect 21888 14112 21904 14176
rect 21968 14112 21984 14176
rect 22048 14112 22054 14176
rect 21738 14111 22054 14112
rect 0 13970 800 14000
rect 1485 13970 1551 13973
rect 0 13968 1551 13970
rect 0 13912 1490 13968
rect 1546 13912 1551 13968
rect 0 13910 1551 13912
rect 0 13880 800 13910
rect 1485 13907 1551 13910
rect 21449 13970 21515 13973
rect 22200 13970 23000 14000
rect 21449 13968 23000 13970
rect 21449 13912 21454 13968
rect 21510 13912 23000 13968
rect 21449 13910 23000 13912
rect 21449 13907 21515 13910
rect 22200 13880 23000 13910
rect 12801 13834 12867 13837
rect 17125 13834 17191 13837
rect 12801 13832 17191 13834
rect 12801 13776 12806 13832
rect 12862 13776 17130 13832
rect 17186 13776 17191 13832
rect 12801 13774 17191 13776
rect 12801 13771 12867 13774
rect 17125 13771 17191 13774
rect 3545 13632 3861 13633
rect 0 13562 800 13592
rect 3545 13568 3551 13632
rect 3615 13568 3631 13632
rect 3695 13568 3711 13632
rect 3775 13568 3791 13632
rect 3855 13568 3861 13632
rect 3545 13567 3861 13568
rect 8743 13632 9059 13633
rect 8743 13568 8749 13632
rect 8813 13568 8829 13632
rect 8893 13568 8909 13632
rect 8973 13568 8989 13632
rect 9053 13568 9059 13632
rect 8743 13567 9059 13568
rect 13941 13632 14257 13633
rect 13941 13568 13947 13632
rect 14011 13568 14027 13632
rect 14091 13568 14107 13632
rect 14171 13568 14187 13632
rect 14251 13568 14257 13632
rect 13941 13567 14257 13568
rect 19139 13632 19455 13633
rect 19139 13568 19145 13632
rect 19209 13568 19225 13632
rect 19289 13568 19305 13632
rect 19369 13568 19385 13632
rect 19449 13568 19455 13632
rect 19139 13567 19455 13568
rect 1485 13562 1551 13565
rect 0 13560 1551 13562
rect 0 13504 1490 13560
rect 1546 13504 1551 13560
rect 0 13502 1551 13504
rect 0 13472 800 13502
rect 1485 13499 1551 13502
rect 21449 13562 21515 13565
rect 22200 13562 23000 13592
rect 21449 13560 23000 13562
rect 21449 13504 21454 13560
rect 21510 13504 23000 13560
rect 21449 13502 23000 13504
rect 21449 13499 21515 13502
rect 22200 13472 23000 13502
rect 8753 13426 8819 13429
rect 15101 13426 15167 13429
rect 8753 13424 15167 13426
rect 8753 13368 8758 13424
rect 8814 13368 15106 13424
rect 15162 13368 15167 13424
rect 8753 13366 15167 13368
rect 8753 13363 8819 13366
rect 15101 13363 15167 13366
rect 15929 13426 15995 13429
rect 20989 13426 21055 13429
rect 15929 13424 21055 13426
rect 15929 13368 15934 13424
rect 15990 13368 20994 13424
rect 21050 13368 21055 13424
rect 15929 13366 21055 13368
rect 15929 13363 15995 13366
rect 20989 13363 21055 13366
rect 8518 13228 8524 13292
rect 8588 13290 8594 13292
rect 18965 13290 19031 13293
rect 8588 13288 19031 13290
rect 8588 13232 18970 13288
rect 19026 13232 19031 13288
rect 8588 13230 19031 13232
rect 8588 13228 8594 13230
rect 18965 13227 19031 13230
rect 21541 13290 21607 13293
rect 21541 13288 22202 13290
rect 21541 13232 21546 13288
rect 21602 13232 22202 13288
rect 21541 13230 22202 13232
rect 21541 13227 21607 13230
rect 22142 13184 22202 13230
rect 0 13154 800 13184
rect 1393 13154 1459 13157
rect 0 13152 1459 13154
rect 0 13096 1398 13152
rect 1454 13096 1459 13152
rect 0 13094 1459 13096
rect 22142 13094 23000 13184
rect 0 13064 800 13094
rect 1393 13091 1459 13094
rect 6144 13088 6460 13089
rect 6144 13024 6150 13088
rect 6214 13024 6230 13088
rect 6294 13024 6310 13088
rect 6374 13024 6390 13088
rect 6454 13024 6460 13088
rect 6144 13023 6460 13024
rect 11342 13088 11658 13089
rect 11342 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11658 13088
rect 11342 13023 11658 13024
rect 16540 13088 16856 13089
rect 16540 13024 16546 13088
rect 16610 13024 16626 13088
rect 16690 13024 16706 13088
rect 16770 13024 16786 13088
rect 16850 13024 16856 13088
rect 16540 13023 16856 13024
rect 21738 13088 22054 13089
rect 21738 13024 21744 13088
rect 21808 13024 21824 13088
rect 21888 13024 21904 13088
rect 21968 13024 21984 13088
rect 22048 13024 22054 13088
rect 22200 13064 23000 13094
rect 21738 13023 22054 13024
rect 8201 12882 8267 12885
rect 12801 12882 12867 12885
rect 8201 12880 12867 12882
rect 8201 12824 8206 12880
rect 8262 12824 12806 12880
rect 12862 12824 12867 12880
rect 8201 12822 12867 12824
rect 8201 12819 8267 12822
rect 12801 12819 12867 12822
rect 0 12746 800 12776
rect 2221 12746 2287 12749
rect 0 12744 2287 12746
rect 0 12688 2226 12744
rect 2282 12688 2287 12744
rect 0 12686 2287 12688
rect 0 12656 800 12686
rect 2221 12683 2287 12686
rect 13445 12746 13511 12749
rect 20713 12746 20779 12749
rect 13445 12744 20779 12746
rect 13445 12688 13450 12744
rect 13506 12688 20718 12744
rect 20774 12688 20779 12744
rect 13445 12686 20779 12688
rect 13445 12683 13511 12686
rect 20713 12683 20779 12686
rect 21449 12746 21515 12749
rect 22200 12746 23000 12776
rect 21449 12744 23000 12746
rect 21449 12688 21454 12744
rect 21510 12688 23000 12744
rect 21449 12686 23000 12688
rect 21449 12683 21515 12686
rect 22200 12656 23000 12686
rect 3545 12544 3861 12545
rect 3545 12480 3551 12544
rect 3615 12480 3631 12544
rect 3695 12480 3711 12544
rect 3775 12480 3791 12544
rect 3855 12480 3861 12544
rect 3545 12479 3861 12480
rect 8743 12544 9059 12545
rect 8743 12480 8749 12544
rect 8813 12480 8829 12544
rect 8893 12480 8909 12544
rect 8973 12480 8989 12544
rect 9053 12480 9059 12544
rect 8743 12479 9059 12480
rect 13941 12544 14257 12545
rect 13941 12480 13947 12544
rect 14011 12480 14027 12544
rect 14091 12480 14107 12544
rect 14171 12480 14187 12544
rect 14251 12480 14257 12544
rect 13941 12479 14257 12480
rect 19139 12544 19455 12545
rect 19139 12480 19145 12544
rect 19209 12480 19225 12544
rect 19289 12480 19305 12544
rect 19369 12480 19385 12544
rect 19449 12480 19455 12544
rect 19139 12479 19455 12480
rect 5717 12474 5783 12477
rect 7649 12474 7715 12477
rect 5717 12472 7715 12474
rect 5717 12416 5722 12472
rect 5778 12416 7654 12472
rect 7710 12416 7715 12472
rect 5717 12414 7715 12416
rect 5717 12411 5783 12414
rect 7649 12411 7715 12414
rect 0 12338 800 12368
rect 1485 12338 1551 12341
rect 0 12336 1551 12338
rect 0 12280 1490 12336
rect 1546 12280 1551 12336
rect 0 12278 1551 12280
rect 0 12248 800 12278
rect 1485 12275 1551 12278
rect 1669 12338 1735 12341
rect 8518 12338 8524 12340
rect 1669 12336 8524 12338
rect 1669 12280 1674 12336
rect 1730 12280 8524 12336
rect 1669 12278 8524 12280
rect 1669 12275 1735 12278
rect 8518 12276 8524 12278
rect 8588 12276 8594 12340
rect 21081 12338 21147 12341
rect 22200 12338 23000 12368
rect 21081 12336 23000 12338
rect 21081 12280 21086 12336
rect 21142 12280 23000 12336
rect 21081 12278 23000 12280
rect 21081 12275 21147 12278
rect 22200 12248 23000 12278
rect 2681 12202 2747 12205
rect 18321 12202 18387 12205
rect 20529 12202 20595 12205
rect 2681 12200 20595 12202
rect 2681 12144 2686 12200
rect 2742 12144 18326 12200
rect 18382 12144 20534 12200
rect 20590 12144 20595 12200
rect 2681 12142 20595 12144
rect 2681 12139 2747 12142
rect 18321 12139 18387 12142
rect 20529 12139 20595 12142
rect 6144 12000 6460 12001
rect 0 11930 800 11960
rect 6144 11936 6150 12000
rect 6214 11936 6230 12000
rect 6294 11936 6310 12000
rect 6374 11936 6390 12000
rect 6454 11936 6460 12000
rect 6144 11935 6460 11936
rect 11342 12000 11658 12001
rect 11342 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11658 12000
rect 11342 11935 11658 11936
rect 16540 12000 16856 12001
rect 16540 11936 16546 12000
rect 16610 11936 16626 12000
rect 16690 11936 16706 12000
rect 16770 11936 16786 12000
rect 16850 11936 16856 12000
rect 16540 11935 16856 11936
rect 21738 12000 22054 12001
rect 21738 11936 21744 12000
rect 21808 11936 21824 12000
rect 21888 11936 21904 12000
rect 21968 11936 21984 12000
rect 22048 11936 22054 12000
rect 21738 11935 22054 11936
rect 1853 11930 1919 11933
rect 22200 11930 23000 11960
rect 0 11928 1919 11930
rect 0 11872 1858 11928
rect 1914 11872 1919 11928
rect 0 11870 1919 11872
rect 0 11840 800 11870
rect 1853 11867 1919 11870
rect 22142 11840 23000 11930
rect 5022 11732 5028 11796
rect 5092 11794 5098 11796
rect 11145 11794 11211 11797
rect 12249 11794 12315 11797
rect 5092 11792 12315 11794
rect 5092 11736 11150 11792
rect 11206 11736 12254 11792
rect 12310 11736 12315 11792
rect 5092 11734 12315 11736
rect 5092 11732 5098 11734
rect 11145 11731 11211 11734
rect 12249 11731 12315 11734
rect 17033 11794 17099 11797
rect 17769 11794 17835 11797
rect 17033 11792 17835 11794
rect 17033 11736 17038 11792
rect 17094 11736 17774 11792
rect 17830 11736 17835 11792
rect 17033 11734 17835 11736
rect 17033 11731 17099 11734
rect 17769 11731 17835 11734
rect 21449 11794 21515 11797
rect 22142 11794 22202 11840
rect 21449 11792 22202 11794
rect 21449 11736 21454 11792
rect 21510 11736 22202 11792
rect 21449 11734 22202 11736
rect 21449 11731 21515 11734
rect 1669 11658 1735 11661
rect 18597 11658 18663 11661
rect 1669 11656 18663 11658
rect 1669 11600 1674 11656
rect 1730 11600 18602 11656
rect 18658 11600 18663 11656
rect 1669 11598 18663 11600
rect 1669 11595 1735 11598
rect 18597 11595 18663 11598
rect 0 11522 800 11552
rect 2129 11522 2195 11525
rect 0 11520 2195 11522
rect 0 11464 2134 11520
rect 2190 11464 2195 11520
rect 0 11462 2195 11464
rect 0 11432 800 11462
rect 2129 11459 2195 11462
rect 21541 11522 21607 11525
rect 22200 11522 23000 11552
rect 21541 11520 23000 11522
rect 21541 11464 21546 11520
rect 21602 11464 23000 11520
rect 21541 11462 23000 11464
rect 21541 11459 21607 11462
rect 3545 11456 3861 11457
rect 3545 11392 3551 11456
rect 3615 11392 3631 11456
rect 3695 11392 3711 11456
rect 3775 11392 3791 11456
rect 3855 11392 3861 11456
rect 3545 11391 3861 11392
rect 8743 11456 9059 11457
rect 8743 11392 8749 11456
rect 8813 11392 8829 11456
rect 8893 11392 8909 11456
rect 8973 11392 8989 11456
rect 9053 11392 9059 11456
rect 8743 11391 9059 11392
rect 13941 11456 14257 11457
rect 13941 11392 13947 11456
rect 14011 11392 14027 11456
rect 14091 11392 14107 11456
rect 14171 11392 14187 11456
rect 14251 11392 14257 11456
rect 13941 11391 14257 11392
rect 19139 11456 19455 11457
rect 19139 11392 19145 11456
rect 19209 11392 19225 11456
rect 19289 11392 19305 11456
rect 19369 11392 19385 11456
rect 19449 11392 19455 11456
rect 22200 11432 23000 11462
rect 19139 11391 19455 11392
rect 3233 11250 3299 11253
rect 8661 11250 8727 11253
rect 12433 11250 12499 11253
rect 15745 11250 15811 11253
rect 3233 11248 3434 11250
rect 3233 11192 3238 11248
rect 3294 11192 3434 11248
rect 3233 11190 3434 11192
rect 3233 11187 3299 11190
rect 0 11114 800 11144
rect 1485 11114 1551 11117
rect 0 11112 1551 11114
rect 0 11056 1490 11112
rect 1546 11056 1551 11112
rect 0 11054 1551 11056
rect 3374 11114 3434 11190
rect 8661 11248 15811 11250
rect 8661 11192 8666 11248
rect 8722 11192 12438 11248
rect 12494 11192 15750 11248
rect 15806 11192 15811 11248
rect 8661 11190 15811 11192
rect 8661 11187 8727 11190
rect 12433 11187 12499 11190
rect 15745 11187 15811 11190
rect 18597 11250 18663 11253
rect 19241 11250 19307 11253
rect 18597 11248 19307 11250
rect 18597 11192 18602 11248
rect 18658 11192 19246 11248
rect 19302 11192 19307 11248
rect 18597 11190 19307 11192
rect 18597 11187 18663 11190
rect 19241 11187 19307 11190
rect 4245 11114 4311 11117
rect 5165 11114 5231 11117
rect 20989 11114 21055 11117
rect 3374 11112 21055 11114
rect 3374 11056 4250 11112
rect 4306 11056 5170 11112
rect 5226 11056 20994 11112
rect 21050 11056 21055 11112
rect 3374 11054 21055 11056
rect 0 11024 800 11054
rect 1485 11051 1551 11054
rect 4245 11051 4311 11054
rect 5165 11051 5231 11054
rect 20989 11051 21055 11054
rect 21449 11114 21515 11117
rect 22200 11114 23000 11144
rect 21449 11112 23000 11114
rect 21449 11056 21454 11112
rect 21510 11056 23000 11112
rect 21449 11054 23000 11056
rect 21449 11051 21515 11054
rect 22200 11024 23000 11054
rect 6144 10912 6460 10913
rect 6144 10848 6150 10912
rect 6214 10848 6230 10912
rect 6294 10848 6310 10912
rect 6374 10848 6390 10912
rect 6454 10848 6460 10912
rect 6144 10847 6460 10848
rect 11342 10912 11658 10913
rect 11342 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11658 10912
rect 11342 10847 11658 10848
rect 16540 10912 16856 10913
rect 16540 10848 16546 10912
rect 16610 10848 16626 10912
rect 16690 10848 16706 10912
rect 16770 10848 16786 10912
rect 16850 10848 16856 10912
rect 16540 10847 16856 10848
rect 21738 10912 22054 10913
rect 21738 10848 21744 10912
rect 21808 10848 21824 10912
rect 21888 10848 21904 10912
rect 21968 10848 21984 10912
rect 22048 10848 22054 10912
rect 21738 10847 22054 10848
rect 2681 10842 2747 10845
rect 4429 10842 4495 10845
rect 2681 10840 4495 10842
rect 2681 10784 2686 10840
rect 2742 10784 4434 10840
rect 4490 10784 4495 10840
rect 2681 10782 4495 10784
rect 2681 10779 2747 10782
rect 4429 10779 4495 10782
rect 0 10706 800 10736
rect 1393 10706 1459 10709
rect 0 10704 1459 10706
rect 0 10648 1398 10704
rect 1454 10648 1459 10704
rect 0 10646 1459 10648
rect 0 10616 800 10646
rect 1393 10643 1459 10646
rect 10225 10706 10291 10709
rect 17861 10706 17927 10709
rect 18229 10706 18295 10709
rect 10225 10704 18295 10706
rect 10225 10648 10230 10704
rect 10286 10648 17866 10704
rect 17922 10648 18234 10704
rect 18290 10648 18295 10704
rect 10225 10646 18295 10648
rect 10225 10643 10291 10646
rect 17861 10643 17927 10646
rect 18229 10643 18295 10646
rect 21081 10706 21147 10709
rect 22200 10706 23000 10736
rect 21081 10704 23000 10706
rect 21081 10648 21086 10704
rect 21142 10648 23000 10704
rect 21081 10646 23000 10648
rect 21081 10643 21147 10646
rect 22200 10616 23000 10646
rect 2313 10570 2379 10573
rect 3918 10570 3924 10572
rect 2313 10568 3924 10570
rect 2313 10512 2318 10568
rect 2374 10512 3924 10568
rect 2313 10510 3924 10512
rect 2313 10507 2379 10510
rect 3918 10508 3924 10510
rect 3988 10508 3994 10572
rect 12893 10570 12959 10573
rect 21357 10570 21423 10573
rect 12893 10568 21423 10570
rect 12893 10512 12898 10568
rect 12954 10512 21362 10568
rect 21418 10512 21423 10568
rect 12893 10510 21423 10512
rect 12893 10507 12959 10510
rect 21357 10507 21423 10510
rect 3545 10368 3861 10369
rect 0 10298 800 10328
rect 3545 10304 3551 10368
rect 3615 10304 3631 10368
rect 3695 10304 3711 10368
rect 3775 10304 3791 10368
rect 3855 10304 3861 10368
rect 3545 10303 3861 10304
rect 8743 10368 9059 10369
rect 8743 10304 8749 10368
rect 8813 10304 8829 10368
rect 8893 10304 8909 10368
rect 8973 10304 8989 10368
rect 9053 10304 9059 10368
rect 8743 10303 9059 10304
rect 13941 10368 14257 10369
rect 13941 10304 13947 10368
rect 14011 10304 14027 10368
rect 14091 10304 14107 10368
rect 14171 10304 14187 10368
rect 14251 10304 14257 10368
rect 13941 10303 14257 10304
rect 19139 10368 19455 10369
rect 19139 10304 19145 10368
rect 19209 10304 19225 10368
rect 19289 10304 19305 10368
rect 19369 10304 19385 10368
rect 19449 10304 19455 10368
rect 19139 10303 19455 10304
rect 1485 10298 1551 10301
rect 0 10296 1551 10298
rect 0 10240 1490 10296
rect 1546 10240 1551 10296
rect 0 10238 1551 10240
rect 0 10208 800 10238
rect 1485 10235 1551 10238
rect 21449 10298 21515 10301
rect 22200 10298 23000 10328
rect 21449 10296 23000 10298
rect 21449 10240 21454 10296
rect 21510 10240 23000 10296
rect 21449 10238 23000 10240
rect 21449 10235 21515 10238
rect 22200 10208 23000 10238
rect 2037 10162 2103 10165
rect 9857 10162 9923 10165
rect 2037 10160 9923 10162
rect 2037 10104 2042 10160
rect 2098 10104 9862 10160
rect 9918 10104 9923 10160
rect 2037 10102 9923 10104
rect 2037 10099 2103 10102
rect 9857 10099 9923 10102
rect 11830 10100 11836 10164
rect 11900 10162 11906 10164
rect 16573 10162 16639 10165
rect 11900 10160 16639 10162
rect 11900 10104 16578 10160
rect 16634 10104 16639 10160
rect 11900 10102 16639 10104
rect 11900 10100 11906 10102
rect 16573 10099 16639 10102
rect 20529 10162 20595 10165
rect 20529 10160 20914 10162
rect 20529 10104 20534 10160
rect 20590 10104 20914 10160
rect 20529 10102 20914 10104
rect 20529 10099 20595 10102
rect 5165 10026 5231 10029
rect 20713 10026 20779 10029
rect 5165 10024 20779 10026
rect 5165 9968 5170 10024
rect 5226 9968 20718 10024
rect 20774 9968 20779 10024
rect 5165 9966 20779 9968
rect 20854 10026 20914 10102
rect 20854 9966 22202 10026
rect 5165 9963 5231 9966
rect 20713 9963 20779 9966
rect 22142 9920 22202 9966
rect 0 9890 800 9920
rect 2129 9890 2195 9893
rect 0 9888 2195 9890
rect 0 9832 2134 9888
rect 2190 9832 2195 9888
rect 0 9830 2195 9832
rect 0 9800 800 9830
rect 2129 9827 2195 9830
rect 3509 9890 3575 9893
rect 5349 9890 5415 9893
rect 3509 9888 5415 9890
rect 3509 9832 3514 9888
rect 3570 9832 5354 9888
rect 5410 9832 5415 9888
rect 3509 9830 5415 9832
rect 22142 9830 23000 9920
rect 3509 9827 3575 9830
rect 5349 9827 5415 9830
rect 6144 9824 6460 9825
rect 6144 9760 6150 9824
rect 6214 9760 6230 9824
rect 6294 9760 6310 9824
rect 6374 9760 6390 9824
rect 6454 9760 6460 9824
rect 6144 9759 6460 9760
rect 11342 9824 11658 9825
rect 11342 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11658 9824
rect 11342 9759 11658 9760
rect 16540 9824 16856 9825
rect 16540 9760 16546 9824
rect 16610 9760 16626 9824
rect 16690 9760 16706 9824
rect 16770 9760 16786 9824
rect 16850 9760 16856 9824
rect 16540 9759 16856 9760
rect 21738 9824 22054 9825
rect 21738 9760 21744 9824
rect 21808 9760 21824 9824
rect 21888 9760 21904 9824
rect 21968 9760 21984 9824
rect 22048 9760 22054 9824
rect 22200 9800 23000 9830
rect 21738 9759 22054 9760
rect 5257 9754 5323 9757
rect 5214 9752 5323 9754
rect 5214 9696 5262 9752
rect 5318 9696 5323 9752
rect 5214 9691 5323 9696
rect 8201 9754 8267 9757
rect 8334 9754 8340 9756
rect 8201 9752 8340 9754
rect 8201 9696 8206 9752
rect 8262 9696 8340 9752
rect 8201 9694 8340 9696
rect 8201 9691 8267 9694
rect 8334 9692 8340 9694
rect 8404 9754 8410 9756
rect 9949 9754 10015 9757
rect 8404 9752 10015 9754
rect 8404 9696 9954 9752
rect 10010 9696 10015 9752
rect 8404 9694 10015 9696
rect 8404 9692 8410 9694
rect 9949 9691 10015 9694
rect 2221 9618 2287 9621
rect 2221 9616 2790 9618
rect 2221 9560 2226 9616
rect 2282 9560 2790 9616
rect 2221 9558 2790 9560
rect 2221 9555 2287 9558
rect 0 9482 800 9512
rect 1853 9482 1919 9485
rect 0 9480 1919 9482
rect 0 9424 1858 9480
rect 1914 9424 1919 9480
rect 0 9422 1919 9424
rect 2730 9482 2790 9558
rect 5214 9482 5274 9691
rect 14549 9618 14615 9621
rect 15285 9618 15351 9621
rect 14549 9616 15351 9618
rect 14549 9560 14554 9616
rect 14610 9560 15290 9616
rect 15346 9560 15351 9616
rect 14549 9558 15351 9560
rect 14549 9555 14615 9558
rect 15285 9555 15351 9558
rect 16389 9618 16455 9621
rect 18137 9618 18203 9621
rect 16389 9616 18203 9618
rect 16389 9560 16394 9616
rect 16450 9560 18142 9616
rect 18198 9560 18203 9616
rect 16389 9558 18203 9560
rect 16389 9555 16455 9558
rect 18137 9555 18203 9558
rect 17953 9482 18019 9485
rect 20478 9482 20484 9484
rect 2730 9480 20484 9482
rect 2730 9424 17958 9480
rect 18014 9424 20484 9480
rect 2730 9422 20484 9424
rect 0 9392 800 9422
rect 1853 9419 1919 9422
rect 17953 9419 18019 9422
rect 20478 9420 20484 9422
rect 20548 9420 20554 9484
rect 21449 9482 21515 9485
rect 22200 9482 23000 9512
rect 21449 9480 23000 9482
rect 21449 9424 21454 9480
rect 21510 9424 23000 9480
rect 21449 9422 23000 9424
rect 21449 9419 21515 9422
rect 22200 9392 23000 9422
rect 3545 9280 3861 9281
rect 3545 9216 3551 9280
rect 3615 9216 3631 9280
rect 3695 9216 3711 9280
rect 3775 9216 3791 9280
rect 3855 9216 3861 9280
rect 3545 9215 3861 9216
rect 8743 9280 9059 9281
rect 8743 9216 8749 9280
rect 8813 9216 8829 9280
rect 8893 9216 8909 9280
rect 8973 9216 8989 9280
rect 9053 9216 9059 9280
rect 8743 9215 9059 9216
rect 13941 9280 14257 9281
rect 13941 9216 13947 9280
rect 14011 9216 14027 9280
rect 14091 9216 14107 9280
rect 14171 9216 14187 9280
rect 14251 9216 14257 9280
rect 13941 9215 14257 9216
rect 19139 9280 19455 9281
rect 19139 9216 19145 9280
rect 19209 9216 19225 9280
rect 19289 9216 19305 9280
rect 19369 9216 19385 9280
rect 19449 9216 19455 9280
rect 19139 9215 19455 9216
rect 0 9074 800 9104
rect 1393 9074 1459 9077
rect 0 9072 1459 9074
rect 0 9016 1398 9072
rect 1454 9016 1459 9072
rect 0 9014 1459 9016
rect 0 8984 800 9014
rect 1393 9011 1459 9014
rect 10961 9074 11027 9077
rect 20989 9074 21055 9077
rect 10961 9072 21055 9074
rect 10961 9016 10966 9072
rect 11022 9016 20994 9072
rect 21050 9016 21055 9072
rect 10961 9014 21055 9016
rect 10961 9011 11027 9014
rect 20989 9011 21055 9014
rect 21541 9074 21607 9077
rect 22200 9074 23000 9104
rect 21541 9072 23000 9074
rect 21541 9016 21546 9072
rect 21602 9016 23000 9072
rect 21541 9014 23000 9016
rect 21541 9011 21607 9014
rect 22200 8984 23000 9014
rect 7966 8876 7972 8940
rect 8036 8938 8042 8940
rect 8109 8938 8175 8941
rect 8036 8936 8175 8938
rect 8036 8880 8114 8936
rect 8170 8880 8175 8936
rect 8036 8878 8175 8880
rect 8036 8876 8042 8878
rect 8109 8875 8175 8878
rect 17493 8938 17559 8941
rect 20069 8938 20135 8941
rect 17493 8936 20135 8938
rect 17493 8880 17498 8936
rect 17554 8880 20074 8936
rect 20130 8880 20135 8936
rect 17493 8878 20135 8880
rect 17493 8875 17559 8878
rect 20069 8875 20135 8878
rect 17585 8802 17651 8805
rect 19977 8802 20043 8805
rect 17585 8800 20043 8802
rect 17585 8744 17590 8800
rect 17646 8744 19982 8800
rect 20038 8744 20043 8800
rect 17585 8742 20043 8744
rect 17585 8739 17651 8742
rect 19977 8739 20043 8742
rect 6144 8736 6460 8737
rect 0 8666 800 8696
rect 6144 8672 6150 8736
rect 6214 8672 6230 8736
rect 6294 8672 6310 8736
rect 6374 8672 6390 8736
rect 6454 8672 6460 8736
rect 6144 8671 6460 8672
rect 11342 8736 11658 8737
rect 11342 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11658 8736
rect 11342 8671 11658 8672
rect 16540 8736 16856 8737
rect 16540 8672 16546 8736
rect 16610 8672 16626 8736
rect 16690 8672 16706 8736
rect 16770 8672 16786 8736
rect 16850 8672 16856 8736
rect 16540 8671 16856 8672
rect 21738 8736 22054 8737
rect 21738 8672 21744 8736
rect 21808 8672 21824 8736
rect 21888 8672 21904 8736
rect 21968 8672 21984 8736
rect 22048 8672 22054 8736
rect 21738 8671 22054 8672
rect 2221 8666 2287 8669
rect 0 8664 2287 8666
rect 0 8608 2226 8664
rect 2282 8608 2287 8664
rect 0 8606 2287 8608
rect 0 8576 800 8606
rect 2221 8603 2287 8606
rect 17125 8666 17191 8669
rect 19241 8666 19307 8669
rect 22200 8666 23000 8696
rect 17125 8664 19307 8666
rect 17125 8608 17130 8664
rect 17186 8608 19246 8664
rect 19302 8608 19307 8664
rect 17125 8606 19307 8608
rect 17125 8603 17191 8606
rect 19241 8603 19307 8606
rect 22142 8576 23000 8666
rect 20621 8530 20687 8533
rect 22142 8530 22202 8576
rect 20621 8528 22202 8530
rect 20621 8472 20626 8528
rect 20682 8472 22202 8528
rect 20621 8470 22202 8472
rect 20621 8467 20687 8470
rect 19241 8394 19307 8397
rect 19241 8392 19626 8394
rect 19241 8336 19246 8392
rect 19302 8336 19626 8392
rect 19241 8334 19626 8336
rect 19241 8331 19307 8334
rect 0 8258 800 8288
rect 1301 8258 1367 8261
rect 0 8256 1367 8258
rect 0 8200 1306 8256
rect 1362 8200 1367 8256
rect 0 8198 1367 8200
rect 19566 8258 19626 8334
rect 22200 8258 23000 8288
rect 19566 8198 23000 8258
rect 0 8168 800 8198
rect 1301 8195 1367 8198
rect 3545 8192 3861 8193
rect 3545 8128 3551 8192
rect 3615 8128 3631 8192
rect 3695 8128 3711 8192
rect 3775 8128 3791 8192
rect 3855 8128 3861 8192
rect 3545 8127 3861 8128
rect 8743 8192 9059 8193
rect 8743 8128 8749 8192
rect 8813 8128 8829 8192
rect 8893 8128 8909 8192
rect 8973 8128 8989 8192
rect 9053 8128 9059 8192
rect 8743 8127 9059 8128
rect 13941 8192 14257 8193
rect 13941 8128 13947 8192
rect 14011 8128 14027 8192
rect 14091 8128 14107 8192
rect 14171 8128 14187 8192
rect 14251 8128 14257 8192
rect 13941 8127 14257 8128
rect 19139 8192 19455 8193
rect 19139 8128 19145 8192
rect 19209 8128 19225 8192
rect 19289 8128 19305 8192
rect 19369 8128 19385 8192
rect 19449 8128 19455 8192
rect 22200 8168 23000 8198
rect 19139 8127 19455 8128
rect 8150 7924 8156 7988
rect 8220 7986 8226 7988
rect 10593 7986 10659 7989
rect 8220 7984 10659 7986
rect 8220 7928 10598 7984
rect 10654 7928 10659 7984
rect 8220 7926 10659 7928
rect 8220 7924 8226 7926
rect 10593 7923 10659 7926
rect 17217 7986 17283 7989
rect 20253 7986 20319 7989
rect 17217 7984 20319 7986
rect 17217 7928 17222 7984
rect 17278 7928 20258 7984
rect 20314 7928 20319 7984
rect 17217 7926 20319 7928
rect 17217 7923 17283 7926
rect 20253 7923 20319 7926
rect 0 7850 800 7880
rect 1393 7850 1459 7853
rect 3969 7850 4035 7853
rect 0 7848 4035 7850
rect 0 7792 1398 7848
rect 1454 7792 3974 7848
rect 4030 7792 4035 7848
rect 0 7790 4035 7792
rect 0 7760 800 7790
rect 1393 7787 1459 7790
rect 3969 7787 4035 7790
rect 6545 7850 6611 7853
rect 11830 7850 11836 7852
rect 6545 7848 11836 7850
rect 6545 7792 6550 7848
rect 6606 7792 11836 7848
rect 6545 7790 11836 7792
rect 6545 7787 6611 7790
rect 11830 7788 11836 7790
rect 11900 7788 11906 7852
rect 21449 7850 21515 7853
rect 22200 7850 23000 7880
rect 21449 7848 23000 7850
rect 21449 7792 21454 7848
rect 21510 7792 23000 7848
rect 21449 7790 23000 7792
rect 21449 7787 21515 7790
rect 22200 7760 23000 7790
rect 6144 7648 6460 7649
rect 6144 7584 6150 7648
rect 6214 7584 6230 7648
rect 6294 7584 6310 7648
rect 6374 7584 6390 7648
rect 6454 7584 6460 7648
rect 6144 7583 6460 7584
rect 11342 7648 11658 7649
rect 11342 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11658 7648
rect 11342 7583 11658 7584
rect 16540 7648 16856 7649
rect 16540 7584 16546 7648
rect 16610 7584 16626 7648
rect 16690 7584 16706 7648
rect 16770 7584 16786 7648
rect 16850 7584 16856 7648
rect 16540 7583 16856 7584
rect 21738 7648 22054 7649
rect 21738 7584 21744 7648
rect 21808 7584 21824 7648
rect 21888 7584 21904 7648
rect 21968 7584 21984 7648
rect 22048 7584 22054 7648
rect 21738 7583 22054 7584
rect 0 7442 800 7472
rect 3417 7442 3483 7445
rect 0 7440 3483 7442
rect 0 7384 3422 7440
rect 3478 7384 3483 7440
rect 0 7382 3483 7384
rect 0 7352 800 7382
rect 3417 7379 3483 7382
rect 20621 7442 20687 7445
rect 22200 7442 23000 7472
rect 20621 7440 23000 7442
rect 20621 7384 20626 7440
rect 20682 7384 23000 7440
rect 20621 7382 23000 7384
rect 20621 7379 20687 7382
rect 22200 7352 23000 7382
rect 2405 7306 2471 7309
rect 5993 7306 6059 7309
rect 2405 7304 6059 7306
rect 2405 7248 2410 7304
rect 2466 7248 5998 7304
rect 6054 7248 6059 7304
rect 2405 7246 6059 7248
rect 2405 7243 2471 7246
rect 5993 7243 6059 7246
rect 4153 7170 4219 7173
rect 5901 7170 5967 7173
rect 4153 7168 5967 7170
rect 4153 7112 4158 7168
rect 4214 7112 5906 7168
rect 5962 7112 5967 7168
rect 4153 7110 5967 7112
rect 4153 7107 4219 7110
rect 5901 7107 5967 7110
rect 3545 7104 3861 7105
rect 0 7034 800 7064
rect 3545 7040 3551 7104
rect 3615 7040 3631 7104
rect 3695 7040 3711 7104
rect 3775 7040 3791 7104
rect 3855 7040 3861 7104
rect 3545 7039 3861 7040
rect 8743 7104 9059 7105
rect 8743 7040 8749 7104
rect 8813 7040 8829 7104
rect 8893 7040 8909 7104
rect 8973 7040 8989 7104
rect 9053 7040 9059 7104
rect 8743 7039 9059 7040
rect 13941 7104 14257 7105
rect 13941 7040 13947 7104
rect 14011 7040 14027 7104
rect 14091 7040 14107 7104
rect 14171 7040 14187 7104
rect 14251 7040 14257 7104
rect 13941 7039 14257 7040
rect 19139 7104 19455 7105
rect 19139 7040 19145 7104
rect 19209 7040 19225 7104
rect 19289 7040 19305 7104
rect 19369 7040 19385 7104
rect 19449 7040 19455 7104
rect 19139 7039 19455 7040
rect 2221 7034 2287 7037
rect 0 7032 2287 7034
rect 0 6976 2226 7032
rect 2282 6976 2287 7032
rect 0 6974 2287 6976
rect 0 6944 800 6974
rect 2221 6971 2287 6974
rect 20713 7034 20779 7037
rect 22200 7034 23000 7064
rect 20713 7032 23000 7034
rect 20713 6976 20718 7032
rect 20774 6976 23000 7032
rect 20713 6974 23000 6976
rect 20713 6971 20779 6974
rect 22200 6944 23000 6974
rect 5257 6898 5323 6901
rect 7097 6898 7163 6901
rect 5257 6896 7163 6898
rect 5257 6840 5262 6896
rect 5318 6840 7102 6896
rect 7158 6840 7163 6896
rect 5257 6838 7163 6840
rect 5257 6835 5323 6838
rect 7097 6835 7163 6838
rect 1577 6762 1643 6765
rect 18873 6762 18939 6765
rect 1577 6760 18939 6762
rect 1577 6704 1582 6760
rect 1638 6704 18878 6760
rect 18934 6704 18939 6760
rect 1577 6702 18939 6704
rect 1577 6699 1643 6702
rect 18873 6699 18939 6702
rect 20805 6762 20871 6765
rect 20805 6760 22202 6762
rect 20805 6704 20810 6760
rect 20866 6704 22202 6760
rect 20805 6702 22202 6704
rect 20805 6699 20871 6702
rect 22142 6656 22202 6702
rect 0 6626 800 6656
rect 1669 6626 1735 6629
rect 0 6624 1735 6626
rect 0 6568 1674 6624
rect 1730 6568 1735 6624
rect 0 6566 1735 6568
rect 22142 6566 23000 6656
rect 0 6536 800 6566
rect 1669 6563 1735 6566
rect 6144 6560 6460 6561
rect 6144 6496 6150 6560
rect 6214 6496 6230 6560
rect 6294 6496 6310 6560
rect 6374 6496 6390 6560
rect 6454 6496 6460 6560
rect 6144 6495 6460 6496
rect 11342 6560 11658 6561
rect 11342 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11658 6560
rect 11342 6495 11658 6496
rect 16540 6560 16856 6561
rect 16540 6496 16546 6560
rect 16610 6496 16626 6560
rect 16690 6496 16706 6560
rect 16770 6496 16786 6560
rect 16850 6496 16856 6560
rect 16540 6495 16856 6496
rect 21738 6560 22054 6561
rect 21738 6496 21744 6560
rect 21808 6496 21824 6560
rect 21888 6496 21904 6560
rect 21968 6496 21984 6560
rect 22048 6496 22054 6560
rect 22200 6536 23000 6566
rect 21738 6495 22054 6496
rect 3049 6490 3115 6493
rect 3325 6490 3391 6493
rect 3049 6488 3391 6490
rect 3049 6432 3054 6488
rect 3110 6432 3330 6488
rect 3386 6432 3391 6488
rect 3049 6430 3391 6432
rect 3049 6427 3115 6430
rect 3325 6427 3391 6430
rect 1945 6354 2011 6357
rect 14089 6354 14155 6357
rect 21173 6354 21239 6357
rect 1945 6352 14155 6354
rect 1945 6296 1950 6352
rect 2006 6296 14094 6352
rect 14150 6296 14155 6352
rect 1945 6294 14155 6296
rect 1945 6291 2011 6294
rect 14089 6291 14155 6294
rect 16622 6352 21239 6354
rect 16622 6296 21178 6352
rect 21234 6296 21239 6352
rect 16622 6294 21239 6296
rect 0 6218 800 6248
rect 2221 6218 2287 6221
rect 0 6216 2287 6218
rect 0 6160 2226 6216
rect 2282 6160 2287 6216
rect 0 6158 2287 6160
rect 0 6128 800 6158
rect 2221 6155 2287 6158
rect 5901 6218 5967 6221
rect 16622 6218 16682 6294
rect 21173 6291 21239 6294
rect 5901 6216 16682 6218
rect 5901 6160 5906 6216
rect 5962 6160 16682 6216
rect 5901 6158 16682 6160
rect 20713 6218 20779 6221
rect 22200 6218 23000 6248
rect 20713 6216 23000 6218
rect 20713 6160 20718 6216
rect 20774 6160 23000 6216
rect 20713 6158 23000 6160
rect 5901 6155 5967 6158
rect 20713 6155 20779 6158
rect 22200 6128 23000 6158
rect 3545 6016 3861 6017
rect 3545 5952 3551 6016
rect 3615 5952 3631 6016
rect 3695 5952 3711 6016
rect 3775 5952 3791 6016
rect 3855 5952 3861 6016
rect 3545 5951 3861 5952
rect 8743 6016 9059 6017
rect 8743 5952 8749 6016
rect 8813 5952 8829 6016
rect 8893 5952 8909 6016
rect 8973 5952 8989 6016
rect 9053 5952 9059 6016
rect 8743 5951 9059 5952
rect 13941 6016 14257 6017
rect 13941 5952 13947 6016
rect 14011 5952 14027 6016
rect 14091 5952 14107 6016
rect 14171 5952 14187 6016
rect 14251 5952 14257 6016
rect 13941 5951 14257 5952
rect 19139 6016 19455 6017
rect 19139 5952 19145 6016
rect 19209 5952 19225 6016
rect 19289 5952 19305 6016
rect 19369 5952 19385 6016
rect 19449 5952 19455 6016
rect 19139 5951 19455 5952
rect 2773 5946 2839 5949
rect 1534 5944 2839 5946
rect 1534 5888 2778 5944
rect 2834 5888 2839 5944
rect 1534 5886 2839 5888
rect 0 5810 800 5840
rect 1393 5810 1459 5813
rect 1534 5810 1594 5886
rect 2773 5883 2839 5886
rect 0 5808 1594 5810
rect 0 5752 1398 5808
rect 1454 5752 1594 5808
rect 0 5750 1594 5752
rect 1669 5810 1735 5813
rect 9305 5810 9371 5813
rect 1669 5808 9371 5810
rect 1669 5752 1674 5808
rect 1730 5752 9310 5808
rect 9366 5752 9371 5808
rect 1669 5750 9371 5752
rect 0 5720 800 5750
rect 1393 5747 1459 5750
rect 1669 5747 1735 5750
rect 9305 5747 9371 5750
rect 21541 5810 21607 5813
rect 22200 5810 23000 5840
rect 21541 5808 23000 5810
rect 21541 5752 21546 5808
rect 21602 5752 23000 5808
rect 21541 5750 23000 5752
rect 21541 5747 21607 5750
rect 22200 5720 23000 5750
rect 1577 5674 1643 5677
rect 13077 5674 13143 5677
rect 1577 5672 13143 5674
rect 1577 5616 1582 5672
rect 1638 5616 13082 5672
rect 13138 5616 13143 5672
rect 1577 5614 13143 5616
rect 1577 5611 1643 5614
rect 13077 5611 13143 5614
rect 6144 5472 6460 5473
rect 0 5402 800 5432
rect 6144 5408 6150 5472
rect 6214 5408 6230 5472
rect 6294 5408 6310 5472
rect 6374 5408 6390 5472
rect 6454 5408 6460 5472
rect 6144 5407 6460 5408
rect 11342 5472 11658 5473
rect 11342 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11658 5472
rect 11342 5407 11658 5408
rect 16540 5472 16856 5473
rect 16540 5408 16546 5472
rect 16610 5408 16626 5472
rect 16690 5408 16706 5472
rect 16770 5408 16786 5472
rect 16850 5408 16856 5472
rect 16540 5407 16856 5408
rect 21738 5472 22054 5473
rect 21738 5408 21744 5472
rect 21808 5408 21824 5472
rect 21888 5408 21904 5472
rect 21968 5408 21984 5472
rect 22048 5408 22054 5472
rect 21738 5407 22054 5408
rect 1393 5402 1459 5405
rect 22200 5402 23000 5432
rect 0 5400 1459 5402
rect 0 5344 1398 5400
rect 1454 5344 1459 5400
rect 0 5342 1459 5344
rect 0 5312 800 5342
rect 1393 5339 1459 5342
rect 22142 5312 23000 5402
rect 21265 5266 21331 5269
rect 22142 5266 22202 5312
rect 21265 5264 22202 5266
rect 21265 5208 21270 5264
rect 21326 5208 22202 5264
rect 21265 5206 22202 5208
rect 21265 5203 21331 5206
rect 0 4994 800 5024
rect 1393 4994 1459 4997
rect 0 4992 1459 4994
rect 0 4936 1398 4992
rect 1454 4936 1459 4992
rect 0 4934 1459 4936
rect 0 4904 800 4934
rect 1393 4931 1459 4934
rect 21541 4994 21607 4997
rect 22200 4994 23000 5024
rect 21541 4992 23000 4994
rect 21541 4936 21546 4992
rect 21602 4936 23000 4992
rect 21541 4934 23000 4936
rect 21541 4931 21607 4934
rect 3545 4928 3861 4929
rect 3545 4864 3551 4928
rect 3615 4864 3631 4928
rect 3695 4864 3711 4928
rect 3775 4864 3791 4928
rect 3855 4864 3861 4928
rect 3545 4863 3861 4864
rect 8743 4928 9059 4929
rect 8743 4864 8749 4928
rect 8813 4864 8829 4928
rect 8893 4864 8909 4928
rect 8973 4864 8989 4928
rect 9053 4864 9059 4928
rect 8743 4863 9059 4864
rect 13941 4928 14257 4929
rect 13941 4864 13947 4928
rect 14011 4864 14027 4928
rect 14091 4864 14107 4928
rect 14171 4864 14187 4928
rect 14251 4864 14257 4928
rect 13941 4863 14257 4864
rect 19139 4928 19455 4929
rect 19139 4864 19145 4928
rect 19209 4864 19225 4928
rect 19289 4864 19305 4928
rect 19369 4864 19385 4928
rect 19449 4864 19455 4928
rect 22200 4904 23000 4934
rect 19139 4863 19455 4864
rect 0 4586 800 4616
rect 1669 4586 1735 4589
rect 0 4584 1735 4586
rect 0 4528 1674 4584
rect 1730 4528 1735 4584
rect 0 4526 1735 4528
rect 0 4496 800 4526
rect 1669 4523 1735 4526
rect 21541 4586 21607 4589
rect 22200 4586 23000 4616
rect 21541 4584 23000 4586
rect 21541 4528 21546 4584
rect 21602 4528 23000 4584
rect 21541 4526 23000 4528
rect 21541 4523 21607 4526
rect 22200 4496 23000 4526
rect 6144 4384 6460 4385
rect 6144 4320 6150 4384
rect 6214 4320 6230 4384
rect 6294 4320 6310 4384
rect 6374 4320 6390 4384
rect 6454 4320 6460 4384
rect 6144 4319 6460 4320
rect 11342 4384 11658 4385
rect 11342 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11658 4384
rect 11342 4319 11658 4320
rect 16540 4384 16856 4385
rect 16540 4320 16546 4384
rect 16610 4320 16626 4384
rect 16690 4320 16706 4384
rect 16770 4320 16786 4384
rect 16850 4320 16856 4384
rect 16540 4319 16856 4320
rect 21738 4384 22054 4385
rect 21738 4320 21744 4384
rect 21808 4320 21824 4384
rect 21888 4320 21904 4384
rect 21968 4320 21984 4384
rect 22048 4320 22054 4384
rect 21738 4319 22054 4320
rect 0 4178 800 4208
rect 1945 4178 2011 4181
rect 0 4176 2011 4178
rect 0 4120 1950 4176
rect 2006 4120 2011 4176
rect 0 4118 2011 4120
rect 0 4088 800 4118
rect 1945 4115 2011 4118
rect 20713 4178 20779 4181
rect 22200 4178 23000 4208
rect 20713 4176 23000 4178
rect 20713 4120 20718 4176
rect 20774 4120 23000 4176
rect 20713 4118 23000 4120
rect 20713 4115 20779 4118
rect 22200 4088 23000 4118
rect 3545 3840 3861 3841
rect 0 3770 800 3800
rect 3545 3776 3551 3840
rect 3615 3776 3631 3840
rect 3695 3776 3711 3840
rect 3775 3776 3791 3840
rect 3855 3776 3861 3840
rect 3545 3775 3861 3776
rect 8743 3840 9059 3841
rect 8743 3776 8749 3840
rect 8813 3776 8829 3840
rect 8893 3776 8909 3840
rect 8973 3776 8989 3840
rect 9053 3776 9059 3840
rect 8743 3775 9059 3776
rect 13941 3840 14257 3841
rect 13941 3776 13947 3840
rect 14011 3776 14027 3840
rect 14091 3776 14107 3840
rect 14171 3776 14187 3840
rect 14251 3776 14257 3840
rect 13941 3775 14257 3776
rect 19139 3840 19455 3841
rect 19139 3776 19145 3840
rect 19209 3776 19225 3840
rect 19289 3776 19305 3840
rect 19369 3776 19385 3840
rect 19449 3776 19455 3840
rect 19139 3775 19455 3776
rect 1393 3770 1459 3773
rect 0 3768 1459 3770
rect 0 3712 1398 3768
rect 1454 3712 1459 3768
rect 0 3710 1459 3712
rect 0 3680 800 3710
rect 1393 3707 1459 3710
rect 21265 3770 21331 3773
rect 22200 3770 23000 3800
rect 21265 3768 23000 3770
rect 21265 3712 21270 3768
rect 21326 3712 23000 3768
rect 21265 3710 23000 3712
rect 21265 3707 21331 3710
rect 22200 3680 23000 3710
rect 5993 3500 6059 3501
rect 5942 3436 5948 3500
rect 6012 3498 6059 3500
rect 21541 3498 21607 3501
rect 6012 3496 6104 3498
rect 6054 3440 6104 3496
rect 6012 3438 6104 3440
rect 21541 3496 22202 3498
rect 21541 3440 21546 3496
rect 21602 3440 22202 3496
rect 21541 3438 22202 3440
rect 6012 3436 6059 3438
rect 5993 3435 6059 3436
rect 21541 3435 21607 3438
rect 22142 3392 22202 3438
rect 0 3362 800 3392
rect 1393 3362 1459 3365
rect 0 3360 1459 3362
rect 0 3304 1398 3360
rect 1454 3304 1459 3360
rect 0 3302 1459 3304
rect 22142 3302 23000 3392
rect 0 3272 800 3302
rect 1393 3299 1459 3302
rect 6144 3296 6460 3297
rect 6144 3232 6150 3296
rect 6214 3232 6230 3296
rect 6294 3232 6310 3296
rect 6374 3232 6390 3296
rect 6454 3232 6460 3296
rect 6144 3231 6460 3232
rect 11342 3296 11658 3297
rect 11342 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11658 3296
rect 11342 3231 11658 3232
rect 16540 3296 16856 3297
rect 16540 3232 16546 3296
rect 16610 3232 16626 3296
rect 16690 3232 16706 3296
rect 16770 3232 16786 3296
rect 16850 3232 16856 3296
rect 16540 3231 16856 3232
rect 21738 3296 22054 3297
rect 21738 3232 21744 3296
rect 21808 3232 21824 3296
rect 21888 3232 21904 3296
rect 21968 3232 21984 3296
rect 22048 3232 22054 3296
rect 22200 3272 23000 3302
rect 21738 3231 22054 3232
rect 0 2954 800 2984
rect 1393 2954 1459 2957
rect 0 2952 1459 2954
rect 0 2896 1398 2952
rect 1454 2896 1459 2952
rect 0 2894 1459 2896
rect 0 2864 800 2894
rect 1393 2891 1459 2894
rect 4102 2892 4108 2956
rect 4172 2954 4178 2956
rect 16849 2954 16915 2957
rect 4172 2952 16915 2954
rect 4172 2896 16854 2952
rect 16910 2896 16915 2952
rect 4172 2894 16915 2896
rect 4172 2892 4178 2894
rect 16849 2891 16915 2894
rect 21541 2954 21607 2957
rect 22200 2954 23000 2984
rect 21541 2952 23000 2954
rect 21541 2896 21546 2952
rect 21602 2896 23000 2952
rect 21541 2894 23000 2896
rect 21541 2891 21607 2894
rect 22200 2864 23000 2894
rect 3545 2752 3861 2753
rect 3545 2688 3551 2752
rect 3615 2688 3631 2752
rect 3695 2688 3711 2752
rect 3775 2688 3791 2752
rect 3855 2688 3861 2752
rect 3545 2687 3861 2688
rect 8743 2752 9059 2753
rect 8743 2688 8749 2752
rect 8813 2688 8829 2752
rect 8893 2688 8909 2752
rect 8973 2688 8989 2752
rect 9053 2688 9059 2752
rect 8743 2687 9059 2688
rect 13941 2752 14257 2753
rect 13941 2688 13947 2752
rect 14011 2688 14027 2752
rect 14091 2688 14107 2752
rect 14171 2688 14187 2752
rect 14251 2688 14257 2752
rect 13941 2687 14257 2688
rect 19139 2752 19455 2753
rect 19139 2688 19145 2752
rect 19209 2688 19225 2752
rect 19289 2688 19305 2752
rect 19369 2688 19385 2752
rect 19449 2688 19455 2752
rect 19139 2687 19455 2688
rect 0 2546 800 2576
rect 1669 2546 1735 2549
rect 0 2544 1735 2546
rect 0 2488 1674 2544
rect 1730 2488 1735 2544
rect 0 2486 1735 2488
rect 0 2456 800 2486
rect 1669 2483 1735 2486
rect 21265 2546 21331 2549
rect 22200 2546 23000 2576
rect 21265 2544 23000 2546
rect 21265 2488 21270 2544
rect 21326 2488 23000 2544
rect 21265 2486 23000 2488
rect 21265 2483 21331 2486
rect 22200 2456 23000 2486
rect 6144 2208 6460 2209
rect 0 2138 800 2168
rect 6144 2144 6150 2208
rect 6214 2144 6230 2208
rect 6294 2144 6310 2208
rect 6374 2144 6390 2208
rect 6454 2144 6460 2208
rect 6144 2143 6460 2144
rect 11342 2208 11658 2209
rect 11342 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11658 2208
rect 11342 2143 11658 2144
rect 16540 2208 16856 2209
rect 16540 2144 16546 2208
rect 16610 2144 16626 2208
rect 16690 2144 16706 2208
rect 16770 2144 16786 2208
rect 16850 2144 16856 2208
rect 16540 2143 16856 2144
rect 21738 2208 22054 2209
rect 21738 2144 21744 2208
rect 21808 2144 21824 2208
rect 21888 2144 21904 2208
rect 21968 2144 21984 2208
rect 22048 2144 22054 2208
rect 21738 2143 22054 2144
rect 2221 2138 2287 2141
rect 22200 2138 23000 2168
rect 0 2136 2287 2138
rect 0 2080 2226 2136
rect 2282 2080 2287 2136
rect 0 2078 2287 2080
rect 0 2048 800 2078
rect 2221 2075 2287 2078
rect 22142 2048 23000 2138
rect 21265 2002 21331 2005
rect 22142 2002 22202 2048
rect 21265 2000 22202 2002
rect 21265 1944 21270 2000
rect 21326 1944 22202 2000
rect 21265 1942 22202 1944
rect 21265 1939 21331 1942
rect 0 1730 800 1760
rect 2773 1730 2839 1733
rect 0 1728 2839 1730
rect 0 1672 2778 1728
rect 2834 1672 2839 1728
rect 0 1670 2839 1672
rect 0 1640 800 1670
rect 2773 1667 2839 1670
rect 21541 1730 21607 1733
rect 22200 1730 23000 1760
rect 21541 1728 23000 1730
rect 21541 1672 21546 1728
rect 21602 1672 23000 1728
rect 21541 1670 23000 1672
rect 21541 1667 21607 1670
rect 22200 1640 23000 1670
<< via3 >>
rect 6150 20700 6214 20704
rect 6150 20644 6154 20700
rect 6154 20644 6210 20700
rect 6210 20644 6214 20700
rect 6150 20640 6214 20644
rect 6230 20700 6294 20704
rect 6230 20644 6234 20700
rect 6234 20644 6290 20700
rect 6290 20644 6294 20700
rect 6230 20640 6294 20644
rect 6310 20700 6374 20704
rect 6310 20644 6314 20700
rect 6314 20644 6370 20700
rect 6370 20644 6374 20700
rect 6310 20640 6374 20644
rect 6390 20700 6454 20704
rect 6390 20644 6394 20700
rect 6394 20644 6450 20700
rect 6450 20644 6454 20700
rect 6390 20640 6454 20644
rect 11348 20700 11412 20704
rect 11348 20644 11352 20700
rect 11352 20644 11408 20700
rect 11408 20644 11412 20700
rect 11348 20640 11412 20644
rect 11428 20700 11492 20704
rect 11428 20644 11432 20700
rect 11432 20644 11488 20700
rect 11488 20644 11492 20700
rect 11428 20640 11492 20644
rect 11508 20700 11572 20704
rect 11508 20644 11512 20700
rect 11512 20644 11568 20700
rect 11568 20644 11572 20700
rect 11508 20640 11572 20644
rect 11588 20700 11652 20704
rect 11588 20644 11592 20700
rect 11592 20644 11648 20700
rect 11648 20644 11652 20700
rect 11588 20640 11652 20644
rect 16546 20700 16610 20704
rect 16546 20644 16550 20700
rect 16550 20644 16606 20700
rect 16606 20644 16610 20700
rect 16546 20640 16610 20644
rect 16626 20700 16690 20704
rect 16626 20644 16630 20700
rect 16630 20644 16686 20700
rect 16686 20644 16690 20700
rect 16626 20640 16690 20644
rect 16706 20700 16770 20704
rect 16706 20644 16710 20700
rect 16710 20644 16766 20700
rect 16766 20644 16770 20700
rect 16706 20640 16770 20644
rect 16786 20700 16850 20704
rect 16786 20644 16790 20700
rect 16790 20644 16846 20700
rect 16846 20644 16850 20700
rect 16786 20640 16850 20644
rect 21744 20700 21808 20704
rect 21744 20644 21748 20700
rect 21748 20644 21804 20700
rect 21804 20644 21808 20700
rect 21744 20640 21808 20644
rect 21824 20700 21888 20704
rect 21824 20644 21828 20700
rect 21828 20644 21884 20700
rect 21884 20644 21888 20700
rect 21824 20640 21888 20644
rect 21904 20700 21968 20704
rect 21904 20644 21908 20700
rect 21908 20644 21964 20700
rect 21964 20644 21968 20700
rect 21904 20640 21968 20644
rect 21984 20700 22048 20704
rect 21984 20644 21988 20700
rect 21988 20644 22044 20700
rect 22044 20644 22048 20700
rect 21984 20640 22048 20644
rect 5028 20164 5092 20228
rect 3551 20156 3615 20160
rect 3551 20100 3555 20156
rect 3555 20100 3611 20156
rect 3611 20100 3615 20156
rect 3551 20096 3615 20100
rect 3631 20156 3695 20160
rect 3631 20100 3635 20156
rect 3635 20100 3691 20156
rect 3691 20100 3695 20156
rect 3631 20096 3695 20100
rect 3711 20156 3775 20160
rect 3711 20100 3715 20156
rect 3715 20100 3771 20156
rect 3771 20100 3775 20156
rect 3711 20096 3775 20100
rect 3791 20156 3855 20160
rect 3791 20100 3795 20156
rect 3795 20100 3851 20156
rect 3851 20100 3855 20156
rect 3791 20096 3855 20100
rect 8749 20156 8813 20160
rect 8749 20100 8753 20156
rect 8753 20100 8809 20156
rect 8809 20100 8813 20156
rect 8749 20096 8813 20100
rect 8829 20156 8893 20160
rect 8829 20100 8833 20156
rect 8833 20100 8889 20156
rect 8889 20100 8893 20156
rect 8829 20096 8893 20100
rect 8909 20156 8973 20160
rect 8909 20100 8913 20156
rect 8913 20100 8969 20156
rect 8969 20100 8973 20156
rect 8909 20096 8973 20100
rect 8989 20156 9053 20160
rect 8989 20100 8993 20156
rect 8993 20100 9049 20156
rect 9049 20100 9053 20156
rect 8989 20096 9053 20100
rect 13947 20156 14011 20160
rect 13947 20100 13951 20156
rect 13951 20100 14007 20156
rect 14007 20100 14011 20156
rect 13947 20096 14011 20100
rect 14027 20156 14091 20160
rect 14027 20100 14031 20156
rect 14031 20100 14087 20156
rect 14087 20100 14091 20156
rect 14027 20096 14091 20100
rect 14107 20156 14171 20160
rect 14107 20100 14111 20156
rect 14111 20100 14167 20156
rect 14167 20100 14171 20156
rect 14107 20096 14171 20100
rect 14187 20156 14251 20160
rect 14187 20100 14191 20156
rect 14191 20100 14247 20156
rect 14247 20100 14251 20156
rect 14187 20096 14251 20100
rect 19145 20156 19209 20160
rect 19145 20100 19149 20156
rect 19149 20100 19205 20156
rect 19205 20100 19209 20156
rect 19145 20096 19209 20100
rect 19225 20156 19289 20160
rect 19225 20100 19229 20156
rect 19229 20100 19285 20156
rect 19285 20100 19289 20156
rect 19225 20096 19289 20100
rect 19305 20156 19369 20160
rect 19305 20100 19309 20156
rect 19309 20100 19365 20156
rect 19365 20100 19369 20156
rect 19305 20096 19369 20100
rect 19385 20156 19449 20160
rect 19385 20100 19389 20156
rect 19389 20100 19445 20156
rect 19445 20100 19449 20156
rect 19385 20096 19449 20100
rect 8156 20088 8220 20092
rect 8156 20032 8206 20088
rect 8206 20032 8220 20088
rect 5948 19892 6012 19956
rect 8156 20028 8220 20032
rect 6150 19612 6214 19616
rect 6150 19556 6154 19612
rect 6154 19556 6210 19612
rect 6210 19556 6214 19612
rect 6150 19552 6214 19556
rect 6230 19612 6294 19616
rect 6230 19556 6234 19612
rect 6234 19556 6290 19612
rect 6290 19556 6294 19612
rect 6230 19552 6294 19556
rect 6310 19612 6374 19616
rect 6310 19556 6314 19612
rect 6314 19556 6370 19612
rect 6370 19556 6374 19612
rect 6310 19552 6374 19556
rect 6390 19612 6454 19616
rect 6390 19556 6394 19612
rect 6394 19556 6450 19612
rect 6450 19556 6454 19612
rect 6390 19552 6454 19556
rect 3924 19348 3988 19412
rect 8340 19544 8404 19548
rect 8340 19488 8354 19544
rect 8354 19488 8404 19544
rect 8340 19484 8404 19488
rect 11348 19612 11412 19616
rect 11348 19556 11352 19612
rect 11352 19556 11408 19612
rect 11408 19556 11412 19612
rect 11348 19552 11412 19556
rect 11428 19612 11492 19616
rect 11428 19556 11432 19612
rect 11432 19556 11488 19612
rect 11488 19556 11492 19612
rect 11428 19552 11492 19556
rect 11508 19612 11572 19616
rect 11508 19556 11512 19612
rect 11512 19556 11568 19612
rect 11568 19556 11572 19612
rect 11508 19552 11572 19556
rect 11588 19612 11652 19616
rect 11588 19556 11592 19612
rect 11592 19556 11648 19612
rect 11648 19556 11652 19612
rect 11588 19552 11652 19556
rect 16546 19612 16610 19616
rect 16546 19556 16550 19612
rect 16550 19556 16606 19612
rect 16606 19556 16610 19612
rect 16546 19552 16610 19556
rect 16626 19612 16690 19616
rect 16626 19556 16630 19612
rect 16630 19556 16686 19612
rect 16686 19556 16690 19612
rect 16626 19552 16690 19556
rect 16706 19612 16770 19616
rect 16706 19556 16710 19612
rect 16710 19556 16766 19612
rect 16766 19556 16770 19612
rect 16706 19552 16770 19556
rect 16786 19612 16850 19616
rect 16786 19556 16790 19612
rect 16790 19556 16846 19612
rect 16846 19556 16850 19612
rect 16786 19552 16850 19556
rect 21744 19612 21808 19616
rect 21744 19556 21748 19612
rect 21748 19556 21804 19612
rect 21804 19556 21808 19612
rect 21744 19552 21808 19556
rect 21824 19612 21888 19616
rect 21824 19556 21828 19612
rect 21828 19556 21884 19612
rect 21884 19556 21888 19612
rect 21824 19552 21888 19556
rect 21904 19612 21968 19616
rect 21904 19556 21908 19612
rect 21908 19556 21964 19612
rect 21964 19556 21968 19612
rect 21904 19552 21968 19556
rect 21984 19612 22048 19616
rect 21984 19556 21988 19612
rect 21988 19556 22044 19612
rect 22044 19556 22048 19612
rect 21984 19552 22048 19556
rect 11836 19348 11900 19412
rect 4108 19136 4172 19140
rect 4108 19080 4158 19136
rect 4158 19080 4172 19136
rect 4108 19076 4172 19080
rect 7972 19076 8036 19140
rect 3551 19068 3615 19072
rect 3551 19012 3555 19068
rect 3555 19012 3611 19068
rect 3611 19012 3615 19068
rect 3551 19008 3615 19012
rect 3631 19068 3695 19072
rect 3631 19012 3635 19068
rect 3635 19012 3691 19068
rect 3691 19012 3695 19068
rect 3631 19008 3695 19012
rect 3711 19068 3775 19072
rect 3711 19012 3715 19068
rect 3715 19012 3771 19068
rect 3771 19012 3775 19068
rect 3711 19008 3775 19012
rect 3791 19068 3855 19072
rect 3791 19012 3795 19068
rect 3795 19012 3851 19068
rect 3851 19012 3855 19068
rect 3791 19008 3855 19012
rect 8749 19068 8813 19072
rect 8749 19012 8753 19068
rect 8753 19012 8809 19068
rect 8809 19012 8813 19068
rect 8749 19008 8813 19012
rect 8829 19068 8893 19072
rect 8829 19012 8833 19068
rect 8833 19012 8889 19068
rect 8889 19012 8893 19068
rect 8829 19008 8893 19012
rect 8909 19068 8973 19072
rect 8909 19012 8913 19068
rect 8913 19012 8969 19068
rect 8969 19012 8973 19068
rect 8909 19008 8973 19012
rect 8989 19068 9053 19072
rect 8989 19012 8993 19068
rect 8993 19012 9049 19068
rect 9049 19012 9053 19068
rect 8989 19008 9053 19012
rect 5028 18804 5092 18868
rect 13947 19068 14011 19072
rect 13947 19012 13951 19068
rect 13951 19012 14007 19068
rect 14007 19012 14011 19068
rect 13947 19008 14011 19012
rect 14027 19068 14091 19072
rect 14027 19012 14031 19068
rect 14031 19012 14087 19068
rect 14087 19012 14091 19068
rect 14027 19008 14091 19012
rect 14107 19068 14171 19072
rect 14107 19012 14111 19068
rect 14111 19012 14167 19068
rect 14167 19012 14171 19068
rect 14107 19008 14171 19012
rect 14187 19068 14251 19072
rect 14187 19012 14191 19068
rect 14191 19012 14247 19068
rect 14247 19012 14251 19068
rect 14187 19008 14251 19012
rect 19145 19068 19209 19072
rect 19145 19012 19149 19068
rect 19149 19012 19205 19068
rect 19205 19012 19209 19068
rect 19145 19008 19209 19012
rect 19225 19068 19289 19072
rect 19225 19012 19229 19068
rect 19229 19012 19285 19068
rect 19285 19012 19289 19068
rect 19225 19008 19289 19012
rect 19305 19068 19369 19072
rect 19305 19012 19309 19068
rect 19309 19012 19365 19068
rect 19365 19012 19369 19068
rect 19305 19008 19369 19012
rect 19385 19068 19449 19072
rect 19385 19012 19389 19068
rect 19389 19012 19445 19068
rect 19445 19012 19449 19068
rect 19385 19008 19449 19012
rect 20484 18668 20548 18732
rect 6150 18524 6214 18528
rect 6150 18468 6154 18524
rect 6154 18468 6210 18524
rect 6210 18468 6214 18524
rect 6150 18464 6214 18468
rect 6230 18524 6294 18528
rect 6230 18468 6234 18524
rect 6234 18468 6290 18524
rect 6290 18468 6294 18524
rect 6230 18464 6294 18468
rect 6310 18524 6374 18528
rect 6310 18468 6314 18524
rect 6314 18468 6370 18524
rect 6370 18468 6374 18524
rect 6310 18464 6374 18468
rect 6390 18524 6454 18528
rect 6390 18468 6394 18524
rect 6394 18468 6450 18524
rect 6450 18468 6454 18524
rect 6390 18464 6454 18468
rect 11348 18524 11412 18528
rect 11348 18468 11352 18524
rect 11352 18468 11408 18524
rect 11408 18468 11412 18524
rect 11348 18464 11412 18468
rect 11428 18524 11492 18528
rect 11428 18468 11432 18524
rect 11432 18468 11488 18524
rect 11488 18468 11492 18524
rect 11428 18464 11492 18468
rect 11508 18524 11572 18528
rect 11508 18468 11512 18524
rect 11512 18468 11568 18524
rect 11568 18468 11572 18524
rect 11508 18464 11572 18468
rect 11588 18524 11652 18528
rect 11588 18468 11592 18524
rect 11592 18468 11648 18524
rect 11648 18468 11652 18524
rect 11588 18464 11652 18468
rect 16546 18524 16610 18528
rect 16546 18468 16550 18524
rect 16550 18468 16606 18524
rect 16606 18468 16610 18524
rect 16546 18464 16610 18468
rect 16626 18524 16690 18528
rect 16626 18468 16630 18524
rect 16630 18468 16686 18524
rect 16686 18468 16690 18524
rect 16626 18464 16690 18468
rect 16706 18524 16770 18528
rect 16706 18468 16710 18524
rect 16710 18468 16766 18524
rect 16766 18468 16770 18524
rect 16706 18464 16770 18468
rect 16786 18524 16850 18528
rect 16786 18468 16790 18524
rect 16790 18468 16846 18524
rect 16846 18468 16850 18524
rect 16786 18464 16850 18468
rect 21744 18524 21808 18528
rect 21744 18468 21748 18524
rect 21748 18468 21804 18524
rect 21804 18468 21808 18524
rect 21744 18464 21808 18468
rect 21824 18524 21888 18528
rect 21824 18468 21828 18524
rect 21828 18468 21884 18524
rect 21884 18468 21888 18524
rect 21824 18464 21888 18468
rect 21904 18524 21968 18528
rect 21904 18468 21908 18524
rect 21908 18468 21964 18524
rect 21964 18468 21968 18524
rect 21904 18464 21968 18468
rect 21984 18524 22048 18528
rect 21984 18468 21988 18524
rect 21988 18468 22044 18524
rect 22044 18468 22048 18524
rect 21984 18464 22048 18468
rect 8524 17988 8588 18052
rect 3551 17980 3615 17984
rect 3551 17924 3555 17980
rect 3555 17924 3611 17980
rect 3611 17924 3615 17980
rect 3551 17920 3615 17924
rect 3631 17980 3695 17984
rect 3631 17924 3635 17980
rect 3635 17924 3691 17980
rect 3691 17924 3695 17980
rect 3631 17920 3695 17924
rect 3711 17980 3775 17984
rect 3711 17924 3715 17980
rect 3715 17924 3771 17980
rect 3771 17924 3775 17980
rect 3711 17920 3775 17924
rect 3791 17980 3855 17984
rect 3791 17924 3795 17980
rect 3795 17924 3851 17980
rect 3851 17924 3855 17980
rect 3791 17920 3855 17924
rect 8749 17980 8813 17984
rect 8749 17924 8753 17980
rect 8753 17924 8809 17980
rect 8809 17924 8813 17980
rect 8749 17920 8813 17924
rect 8829 17980 8893 17984
rect 8829 17924 8833 17980
rect 8833 17924 8889 17980
rect 8889 17924 8893 17980
rect 8829 17920 8893 17924
rect 8909 17980 8973 17984
rect 8909 17924 8913 17980
rect 8913 17924 8969 17980
rect 8969 17924 8973 17980
rect 8909 17920 8973 17924
rect 8989 17980 9053 17984
rect 8989 17924 8993 17980
rect 8993 17924 9049 17980
rect 9049 17924 9053 17980
rect 8989 17920 9053 17924
rect 13947 17980 14011 17984
rect 13947 17924 13951 17980
rect 13951 17924 14007 17980
rect 14007 17924 14011 17980
rect 13947 17920 14011 17924
rect 14027 17980 14091 17984
rect 14027 17924 14031 17980
rect 14031 17924 14087 17980
rect 14087 17924 14091 17980
rect 14027 17920 14091 17924
rect 14107 17980 14171 17984
rect 14107 17924 14111 17980
rect 14111 17924 14167 17980
rect 14167 17924 14171 17980
rect 14107 17920 14171 17924
rect 14187 17980 14251 17984
rect 14187 17924 14191 17980
rect 14191 17924 14247 17980
rect 14247 17924 14251 17980
rect 14187 17920 14251 17924
rect 19145 17980 19209 17984
rect 19145 17924 19149 17980
rect 19149 17924 19205 17980
rect 19205 17924 19209 17980
rect 19145 17920 19209 17924
rect 19225 17980 19289 17984
rect 19225 17924 19229 17980
rect 19229 17924 19285 17980
rect 19285 17924 19289 17980
rect 19225 17920 19289 17924
rect 19305 17980 19369 17984
rect 19305 17924 19309 17980
rect 19309 17924 19365 17980
rect 19365 17924 19369 17980
rect 19305 17920 19369 17924
rect 19385 17980 19449 17984
rect 19385 17924 19389 17980
rect 19389 17924 19445 17980
rect 19445 17924 19449 17980
rect 19385 17920 19449 17924
rect 6150 17436 6214 17440
rect 6150 17380 6154 17436
rect 6154 17380 6210 17436
rect 6210 17380 6214 17436
rect 6150 17376 6214 17380
rect 6230 17436 6294 17440
rect 6230 17380 6234 17436
rect 6234 17380 6290 17436
rect 6290 17380 6294 17436
rect 6230 17376 6294 17380
rect 6310 17436 6374 17440
rect 6310 17380 6314 17436
rect 6314 17380 6370 17436
rect 6370 17380 6374 17436
rect 6310 17376 6374 17380
rect 6390 17436 6454 17440
rect 6390 17380 6394 17436
rect 6394 17380 6450 17436
rect 6450 17380 6454 17436
rect 6390 17376 6454 17380
rect 11348 17436 11412 17440
rect 11348 17380 11352 17436
rect 11352 17380 11408 17436
rect 11408 17380 11412 17436
rect 11348 17376 11412 17380
rect 11428 17436 11492 17440
rect 11428 17380 11432 17436
rect 11432 17380 11488 17436
rect 11488 17380 11492 17436
rect 11428 17376 11492 17380
rect 11508 17436 11572 17440
rect 11508 17380 11512 17436
rect 11512 17380 11568 17436
rect 11568 17380 11572 17436
rect 11508 17376 11572 17380
rect 11588 17436 11652 17440
rect 11588 17380 11592 17436
rect 11592 17380 11648 17436
rect 11648 17380 11652 17436
rect 11588 17376 11652 17380
rect 16546 17436 16610 17440
rect 16546 17380 16550 17436
rect 16550 17380 16606 17436
rect 16606 17380 16610 17436
rect 16546 17376 16610 17380
rect 16626 17436 16690 17440
rect 16626 17380 16630 17436
rect 16630 17380 16686 17436
rect 16686 17380 16690 17436
rect 16626 17376 16690 17380
rect 16706 17436 16770 17440
rect 16706 17380 16710 17436
rect 16710 17380 16766 17436
rect 16766 17380 16770 17436
rect 16706 17376 16770 17380
rect 16786 17436 16850 17440
rect 16786 17380 16790 17436
rect 16790 17380 16846 17436
rect 16846 17380 16850 17436
rect 16786 17376 16850 17380
rect 21744 17436 21808 17440
rect 21744 17380 21748 17436
rect 21748 17380 21804 17436
rect 21804 17380 21808 17436
rect 21744 17376 21808 17380
rect 21824 17436 21888 17440
rect 21824 17380 21828 17436
rect 21828 17380 21884 17436
rect 21884 17380 21888 17436
rect 21824 17376 21888 17380
rect 21904 17436 21968 17440
rect 21904 17380 21908 17436
rect 21908 17380 21964 17436
rect 21964 17380 21968 17436
rect 21904 17376 21968 17380
rect 21984 17436 22048 17440
rect 21984 17380 21988 17436
rect 21988 17380 22044 17436
rect 22044 17380 22048 17436
rect 21984 17376 22048 17380
rect 3551 16892 3615 16896
rect 3551 16836 3555 16892
rect 3555 16836 3611 16892
rect 3611 16836 3615 16892
rect 3551 16832 3615 16836
rect 3631 16892 3695 16896
rect 3631 16836 3635 16892
rect 3635 16836 3691 16892
rect 3691 16836 3695 16892
rect 3631 16832 3695 16836
rect 3711 16892 3775 16896
rect 3711 16836 3715 16892
rect 3715 16836 3771 16892
rect 3771 16836 3775 16892
rect 3711 16832 3775 16836
rect 3791 16892 3855 16896
rect 3791 16836 3795 16892
rect 3795 16836 3851 16892
rect 3851 16836 3855 16892
rect 3791 16832 3855 16836
rect 8749 16892 8813 16896
rect 8749 16836 8753 16892
rect 8753 16836 8809 16892
rect 8809 16836 8813 16892
rect 8749 16832 8813 16836
rect 8829 16892 8893 16896
rect 8829 16836 8833 16892
rect 8833 16836 8889 16892
rect 8889 16836 8893 16892
rect 8829 16832 8893 16836
rect 8909 16892 8973 16896
rect 8909 16836 8913 16892
rect 8913 16836 8969 16892
rect 8969 16836 8973 16892
rect 8909 16832 8973 16836
rect 8989 16892 9053 16896
rect 8989 16836 8993 16892
rect 8993 16836 9049 16892
rect 9049 16836 9053 16892
rect 8989 16832 9053 16836
rect 13947 16892 14011 16896
rect 13947 16836 13951 16892
rect 13951 16836 14007 16892
rect 14007 16836 14011 16892
rect 13947 16832 14011 16836
rect 14027 16892 14091 16896
rect 14027 16836 14031 16892
rect 14031 16836 14087 16892
rect 14087 16836 14091 16892
rect 14027 16832 14091 16836
rect 14107 16892 14171 16896
rect 14107 16836 14111 16892
rect 14111 16836 14167 16892
rect 14167 16836 14171 16892
rect 14107 16832 14171 16836
rect 14187 16892 14251 16896
rect 14187 16836 14191 16892
rect 14191 16836 14247 16892
rect 14247 16836 14251 16892
rect 14187 16832 14251 16836
rect 19145 16892 19209 16896
rect 19145 16836 19149 16892
rect 19149 16836 19205 16892
rect 19205 16836 19209 16892
rect 19145 16832 19209 16836
rect 19225 16892 19289 16896
rect 19225 16836 19229 16892
rect 19229 16836 19285 16892
rect 19285 16836 19289 16892
rect 19225 16832 19289 16836
rect 19305 16892 19369 16896
rect 19305 16836 19309 16892
rect 19309 16836 19365 16892
rect 19365 16836 19369 16892
rect 19305 16832 19369 16836
rect 19385 16892 19449 16896
rect 19385 16836 19389 16892
rect 19389 16836 19445 16892
rect 19445 16836 19449 16892
rect 19385 16832 19449 16836
rect 6150 16348 6214 16352
rect 6150 16292 6154 16348
rect 6154 16292 6210 16348
rect 6210 16292 6214 16348
rect 6150 16288 6214 16292
rect 6230 16348 6294 16352
rect 6230 16292 6234 16348
rect 6234 16292 6290 16348
rect 6290 16292 6294 16348
rect 6230 16288 6294 16292
rect 6310 16348 6374 16352
rect 6310 16292 6314 16348
rect 6314 16292 6370 16348
rect 6370 16292 6374 16348
rect 6310 16288 6374 16292
rect 6390 16348 6454 16352
rect 6390 16292 6394 16348
rect 6394 16292 6450 16348
rect 6450 16292 6454 16348
rect 6390 16288 6454 16292
rect 11348 16348 11412 16352
rect 11348 16292 11352 16348
rect 11352 16292 11408 16348
rect 11408 16292 11412 16348
rect 11348 16288 11412 16292
rect 11428 16348 11492 16352
rect 11428 16292 11432 16348
rect 11432 16292 11488 16348
rect 11488 16292 11492 16348
rect 11428 16288 11492 16292
rect 11508 16348 11572 16352
rect 11508 16292 11512 16348
rect 11512 16292 11568 16348
rect 11568 16292 11572 16348
rect 11508 16288 11572 16292
rect 11588 16348 11652 16352
rect 11588 16292 11592 16348
rect 11592 16292 11648 16348
rect 11648 16292 11652 16348
rect 11588 16288 11652 16292
rect 16546 16348 16610 16352
rect 16546 16292 16550 16348
rect 16550 16292 16606 16348
rect 16606 16292 16610 16348
rect 16546 16288 16610 16292
rect 16626 16348 16690 16352
rect 16626 16292 16630 16348
rect 16630 16292 16686 16348
rect 16686 16292 16690 16348
rect 16626 16288 16690 16292
rect 16706 16348 16770 16352
rect 16706 16292 16710 16348
rect 16710 16292 16766 16348
rect 16766 16292 16770 16348
rect 16706 16288 16770 16292
rect 16786 16348 16850 16352
rect 16786 16292 16790 16348
rect 16790 16292 16846 16348
rect 16846 16292 16850 16348
rect 16786 16288 16850 16292
rect 21744 16348 21808 16352
rect 21744 16292 21748 16348
rect 21748 16292 21804 16348
rect 21804 16292 21808 16348
rect 21744 16288 21808 16292
rect 21824 16348 21888 16352
rect 21824 16292 21828 16348
rect 21828 16292 21884 16348
rect 21884 16292 21888 16348
rect 21824 16288 21888 16292
rect 21904 16348 21968 16352
rect 21904 16292 21908 16348
rect 21908 16292 21964 16348
rect 21964 16292 21968 16348
rect 21904 16288 21968 16292
rect 21984 16348 22048 16352
rect 21984 16292 21988 16348
rect 21988 16292 22044 16348
rect 22044 16292 22048 16348
rect 21984 16288 22048 16292
rect 3551 15804 3615 15808
rect 3551 15748 3555 15804
rect 3555 15748 3611 15804
rect 3611 15748 3615 15804
rect 3551 15744 3615 15748
rect 3631 15804 3695 15808
rect 3631 15748 3635 15804
rect 3635 15748 3691 15804
rect 3691 15748 3695 15804
rect 3631 15744 3695 15748
rect 3711 15804 3775 15808
rect 3711 15748 3715 15804
rect 3715 15748 3771 15804
rect 3771 15748 3775 15804
rect 3711 15744 3775 15748
rect 3791 15804 3855 15808
rect 3791 15748 3795 15804
rect 3795 15748 3851 15804
rect 3851 15748 3855 15804
rect 3791 15744 3855 15748
rect 8749 15804 8813 15808
rect 8749 15748 8753 15804
rect 8753 15748 8809 15804
rect 8809 15748 8813 15804
rect 8749 15744 8813 15748
rect 8829 15804 8893 15808
rect 8829 15748 8833 15804
rect 8833 15748 8889 15804
rect 8889 15748 8893 15804
rect 8829 15744 8893 15748
rect 8909 15804 8973 15808
rect 8909 15748 8913 15804
rect 8913 15748 8969 15804
rect 8969 15748 8973 15804
rect 8909 15744 8973 15748
rect 8989 15804 9053 15808
rect 8989 15748 8993 15804
rect 8993 15748 9049 15804
rect 9049 15748 9053 15804
rect 8989 15744 9053 15748
rect 13947 15804 14011 15808
rect 13947 15748 13951 15804
rect 13951 15748 14007 15804
rect 14007 15748 14011 15804
rect 13947 15744 14011 15748
rect 14027 15804 14091 15808
rect 14027 15748 14031 15804
rect 14031 15748 14087 15804
rect 14087 15748 14091 15804
rect 14027 15744 14091 15748
rect 14107 15804 14171 15808
rect 14107 15748 14111 15804
rect 14111 15748 14167 15804
rect 14167 15748 14171 15804
rect 14107 15744 14171 15748
rect 14187 15804 14251 15808
rect 14187 15748 14191 15804
rect 14191 15748 14247 15804
rect 14247 15748 14251 15804
rect 14187 15744 14251 15748
rect 19145 15804 19209 15808
rect 19145 15748 19149 15804
rect 19149 15748 19205 15804
rect 19205 15748 19209 15804
rect 19145 15744 19209 15748
rect 19225 15804 19289 15808
rect 19225 15748 19229 15804
rect 19229 15748 19285 15804
rect 19285 15748 19289 15804
rect 19225 15744 19289 15748
rect 19305 15804 19369 15808
rect 19305 15748 19309 15804
rect 19309 15748 19365 15804
rect 19365 15748 19369 15804
rect 19305 15744 19369 15748
rect 19385 15804 19449 15808
rect 19385 15748 19389 15804
rect 19389 15748 19445 15804
rect 19445 15748 19449 15804
rect 19385 15744 19449 15748
rect 6150 15260 6214 15264
rect 6150 15204 6154 15260
rect 6154 15204 6210 15260
rect 6210 15204 6214 15260
rect 6150 15200 6214 15204
rect 6230 15260 6294 15264
rect 6230 15204 6234 15260
rect 6234 15204 6290 15260
rect 6290 15204 6294 15260
rect 6230 15200 6294 15204
rect 6310 15260 6374 15264
rect 6310 15204 6314 15260
rect 6314 15204 6370 15260
rect 6370 15204 6374 15260
rect 6310 15200 6374 15204
rect 6390 15260 6454 15264
rect 6390 15204 6394 15260
rect 6394 15204 6450 15260
rect 6450 15204 6454 15260
rect 6390 15200 6454 15204
rect 11348 15260 11412 15264
rect 11348 15204 11352 15260
rect 11352 15204 11408 15260
rect 11408 15204 11412 15260
rect 11348 15200 11412 15204
rect 11428 15260 11492 15264
rect 11428 15204 11432 15260
rect 11432 15204 11488 15260
rect 11488 15204 11492 15260
rect 11428 15200 11492 15204
rect 11508 15260 11572 15264
rect 11508 15204 11512 15260
rect 11512 15204 11568 15260
rect 11568 15204 11572 15260
rect 11508 15200 11572 15204
rect 11588 15260 11652 15264
rect 11588 15204 11592 15260
rect 11592 15204 11648 15260
rect 11648 15204 11652 15260
rect 11588 15200 11652 15204
rect 16546 15260 16610 15264
rect 16546 15204 16550 15260
rect 16550 15204 16606 15260
rect 16606 15204 16610 15260
rect 16546 15200 16610 15204
rect 16626 15260 16690 15264
rect 16626 15204 16630 15260
rect 16630 15204 16686 15260
rect 16686 15204 16690 15260
rect 16626 15200 16690 15204
rect 16706 15260 16770 15264
rect 16706 15204 16710 15260
rect 16710 15204 16766 15260
rect 16766 15204 16770 15260
rect 16706 15200 16770 15204
rect 16786 15260 16850 15264
rect 16786 15204 16790 15260
rect 16790 15204 16846 15260
rect 16846 15204 16850 15260
rect 16786 15200 16850 15204
rect 21744 15260 21808 15264
rect 21744 15204 21748 15260
rect 21748 15204 21804 15260
rect 21804 15204 21808 15260
rect 21744 15200 21808 15204
rect 21824 15260 21888 15264
rect 21824 15204 21828 15260
rect 21828 15204 21884 15260
rect 21884 15204 21888 15260
rect 21824 15200 21888 15204
rect 21904 15260 21968 15264
rect 21904 15204 21908 15260
rect 21908 15204 21964 15260
rect 21964 15204 21968 15260
rect 21904 15200 21968 15204
rect 21984 15260 22048 15264
rect 21984 15204 21988 15260
rect 21988 15204 22044 15260
rect 22044 15204 22048 15260
rect 21984 15200 22048 15204
rect 3551 14716 3615 14720
rect 3551 14660 3555 14716
rect 3555 14660 3611 14716
rect 3611 14660 3615 14716
rect 3551 14656 3615 14660
rect 3631 14716 3695 14720
rect 3631 14660 3635 14716
rect 3635 14660 3691 14716
rect 3691 14660 3695 14716
rect 3631 14656 3695 14660
rect 3711 14716 3775 14720
rect 3711 14660 3715 14716
rect 3715 14660 3771 14716
rect 3771 14660 3775 14716
rect 3711 14656 3775 14660
rect 3791 14716 3855 14720
rect 3791 14660 3795 14716
rect 3795 14660 3851 14716
rect 3851 14660 3855 14716
rect 3791 14656 3855 14660
rect 8749 14716 8813 14720
rect 8749 14660 8753 14716
rect 8753 14660 8809 14716
rect 8809 14660 8813 14716
rect 8749 14656 8813 14660
rect 8829 14716 8893 14720
rect 8829 14660 8833 14716
rect 8833 14660 8889 14716
rect 8889 14660 8893 14716
rect 8829 14656 8893 14660
rect 8909 14716 8973 14720
rect 8909 14660 8913 14716
rect 8913 14660 8969 14716
rect 8969 14660 8973 14716
rect 8909 14656 8973 14660
rect 8989 14716 9053 14720
rect 8989 14660 8993 14716
rect 8993 14660 9049 14716
rect 9049 14660 9053 14716
rect 8989 14656 9053 14660
rect 13947 14716 14011 14720
rect 13947 14660 13951 14716
rect 13951 14660 14007 14716
rect 14007 14660 14011 14716
rect 13947 14656 14011 14660
rect 14027 14716 14091 14720
rect 14027 14660 14031 14716
rect 14031 14660 14087 14716
rect 14087 14660 14091 14716
rect 14027 14656 14091 14660
rect 14107 14716 14171 14720
rect 14107 14660 14111 14716
rect 14111 14660 14167 14716
rect 14167 14660 14171 14716
rect 14107 14656 14171 14660
rect 14187 14716 14251 14720
rect 14187 14660 14191 14716
rect 14191 14660 14247 14716
rect 14247 14660 14251 14716
rect 14187 14656 14251 14660
rect 19145 14716 19209 14720
rect 19145 14660 19149 14716
rect 19149 14660 19205 14716
rect 19205 14660 19209 14716
rect 19145 14656 19209 14660
rect 19225 14716 19289 14720
rect 19225 14660 19229 14716
rect 19229 14660 19285 14716
rect 19285 14660 19289 14716
rect 19225 14656 19289 14660
rect 19305 14716 19369 14720
rect 19305 14660 19309 14716
rect 19309 14660 19365 14716
rect 19365 14660 19369 14716
rect 19305 14656 19369 14660
rect 19385 14716 19449 14720
rect 19385 14660 19389 14716
rect 19389 14660 19445 14716
rect 19445 14660 19449 14716
rect 19385 14656 19449 14660
rect 6150 14172 6214 14176
rect 6150 14116 6154 14172
rect 6154 14116 6210 14172
rect 6210 14116 6214 14172
rect 6150 14112 6214 14116
rect 6230 14172 6294 14176
rect 6230 14116 6234 14172
rect 6234 14116 6290 14172
rect 6290 14116 6294 14172
rect 6230 14112 6294 14116
rect 6310 14172 6374 14176
rect 6310 14116 6314 14172
rect 6314 14116 6370 14172
rect 6370 14116 6374 14172
rect 6310 14112 6374 14116
rect 6390 14172 6454 14176
rect 6390 14116 6394 14172
rect 6394 14116 6450 14172
rect 6450 14116 6454 14172
rect 6390 14112 6454 14116
rect 11348 14172 11412 14176
rect 11348 14116 11352 14172
rect 11352 14116 11408 14172
rect 11408 14116 11412 14172
rect 11348 14112 11412 14116
rect 11428 14172 11492 14176
rect 11428 14116 11432 14172
rect 11432 14116 11488 14172
rect 11488 14116 11492 14172
rect 11428 14112 11492 14116
rect 11508 14172 11572 14176
rect 11508 14116 11512 14172
rect 11512 14116 11568 14172
rect 11568 14116 11572 14172
rect 11508 14112 11572 14116
rect 11588 14172 11652 14176
rect 11588 14116 11592 14172
rect 11592 14116 11648 14172
rect 11648 14116 11652 14172
rect 11588 14112 11652 14116
rect 16546 14172 16610 14176
rect 16546 14116 16550 14172
rect 16550 14116 16606 14172
rect 16606 14116 16610 14172
rect 16546 14112 16610 14116
rect 16626 14172 16690 14176
rect 16626 14116 16630 14172
rect 16630 14116 16686 14172
rect 16686 14116 16690 14172
rect 16626 14112 16690 14116
rect 16706 14172 16770 14176
rect 16706 14116 16710 14172
rect 16710 14116 16766 14172
rect 16766 14116 16770 14172
rect 16706 14112 16770 14116
rect 16786 14172 16850 14176
rect 16786 14116 16790 14172
rect 16790 14116 16846 14172
rect 16846 14116 16850 14172
rect 16786 14112 16850 14116
rect 21744 14172 21808 14176
rect 21744 14116 21748 14172
rect 21748 14116 21804 14172
rect 21804 14116 21808 14172
rect 21744 14112 21808 14116
rect 21824 14172 21888 14176
rect 21824 14116 21828 14172
rect 21828 14116 21884 14172
rect 21884 14116 21888 14172
rect 21824 14112 21888 14116
rect 21904 14172 21968 14176
rect 21904 14116 21908 14172
rect 21908 14116 21964 14172
rect 21964 14116 21968 14172
rect 21904 14112 21968 14116
rect 21984 14172 22048 14176
rect 21984 14116 21988 14172
rect 21988 14116 22044 14172
rect 22044 14116 22048 14172
rect 21984 14112 22048 14116
rect 3551 13628 3615 13632
rect 3551 13572 3555 13628
rect 3555 13572 3611 13628
rect 3611 13572 3615 13628
rect 3551 13568 3615 13572
rect 3631 13628 3695 13632
rect 3631 13572 3635 13628
rect 3635 13572 3691 13628
rect 3691 13572 3695 13628
rect 3631 13568 3695 13572
rect 3711 13628 3775 13632
rect 3711 13572 3715 13628
rect 3715 13572 3771 13628
rect 3771 13572 3775 13628
rect 3711 13568 3775 13572
rect 3791 13628 3855 13632
rect 3791 13572 3795 13628
rect 3795 13572 3851 13628
rect 3851 13572 3855 13628
rect 3791 13568 3855 13572
rect 8749 13628 8813 13632
rect 8749 13572 8753 13628
rect 8753 13572 8809 13628
rect 8809 13572 8813 13628
rect 8749 13568 8813 13572
rect 8829 13628 8893 13632
rect 8829 13572 8833 13628
rect 8833 13572 8889 13628
rect 8889 13572 8893 13628
rect 8829 13568 8893 13572
rect 8909 13628 8973 13632
rect 8909 13572 8913 13628
rect 8913 13572 8969 13628
rect 8969 13572 8973 13628
rect 8909 13568 8973 13572
rect 8989 13628 9053 13632
rect 8989 13572 8993 13628
rect 8993 13572 9049 13628
rect 9049 13572 9053 13628
rect 8989 13568 9053 13572
rect 13947 13628 14011 13632
rect 13947 13572 13951 13628
rect 13951 13572 14007 13628
rect 14007 13572 14011 13628
rect 13947 13568 14011 13572
rect 14027 13628 14091 13632
rect 14027 13572 14031 13628
rect 14031 13572 14087 13628
rect 14087 13572 14091 13628
rect 14027 13568 14091 13572
rect 14107 13628 14171 13632
rect 14107 13572 14111 13628
rect 14111 13572 14167 13628
rect 14167 13572 14171 13628
rect 14107 13568 14171 13572
rect 14187 13628 14251 13632
rect 14187 13572 14191 13628
rect 14191 13572 14247 13628
rect 14247 13572 14251 13628
rect 14187 13568 14251 13572
rect 19145 13628 19209 13632
rect 19145 13572 19149 13628
rect 19149 13572 19205 13628
rect 19205 13572 19209 13628
rect 19145 13568 19209 13572
rect 19225 13628 19289 13632
rect 19225 13572 19229 13628
rect 19229 13572 19285 13628
rect 19285 13572 19289 13628
rect 19225 13568 19289 13572
rect 19305 13628 19369 13632
rect 19305 13572 19309 13628
rect 19309 13572 19365 13628
rect 19365 13572 19369 13628
rect 19305 13568 19369 13572
rect 19385 13628 19449 13632
rect 19385 13572 19389 13628
rect 19389 13572 19445 13628
rect 19445 13572 19449 13628
rect 19385 13568 19449 13572
rect 8524 13228 8588 13292
rect 6150 13084 6214 13088
rect 6150 13028 6154 13084
rect 6154 13028 6210 13084
rect 6210 13028 6214 13084
rect 6150 13024 6214 13028
rect 6230 13084 6294 13088
rect 6230 13028 6234 13084
rect 6234 13028 6290 13084
rect 6290 13028 6294 13084
rect 6230 13024 6294 13028
rect 6310 13084 6374 13088
rect 6310 13028 6314 13084
rect 6314 13028 6370 13084
rect 6370 13028 6374 13084
rect 6310 13024 6374 13028
rect 6390 13084 6454 13088
rect 6390 13028 6394 13084
rect 6394 13028 6450 13084
rect 6450 13028 6454 13084
rect 6390 13024 6454 13028
rect 11348 13084 11412 13088
rect 11348 13028 11352 13084
rect 11352 13028 11408 13084
rect 11408 13028 11412 13084
rect 11348 13024 11412 13028
rect 11428 13084 11492 13088
rect 11428 13028 11432 13084
rect 11432 13028 11488 13084
rect 11488 13028 11492 13084
rect 11428 13024 11492 13028
rect 11508 13084 11572 13088
rect 11508 13028 11512 13084
rect 11512 13028 11568 13084
rect 11568 13028 11572 13084
rect 11508 13024 11572 13028
rect 11588 13084 11652 13088
rect 11588 13028 11592 13084
rect 11592 13028 11648 13084
rect 11648 13028 11652 13084
rect 11588 13024 11652 13028
rect 16546 13084 16610 13088
rect 16546 13028 16550 13084
rect 16550 13028 16606 13084
rect 16606 13028 16610 13084
rect 16546 13024 16610 13028
rect 16626 13084 16690 13088
rect 16626 13028 16630 13084
rect 16630 13028 16686 13084
rect 16686 13028 16690 13084
rect 16626 13024 16690 13028
rect 16706 13084 16770 13088
rect 16706 13028 16710 13084
rect 16710 13028 16766 13084
rect 16766 13028 16770 13084
rect 16706 13024 16770 13028
rect 16786 13084 16850 13088
rect 16786 13028 16790 13084
rect 16790 13028 16846 13084
rect 16846 13028 16850 13084
rect 16786 13024 16850 13028
rect 21744 13084 21808 13088
rect 21744 13028 21748 13084
rect 21748 13028 21804 13084
rect 21804 13028 21808 13084
rect 21744 13024 21808 13028
rect 21824 13084 21888 13088
rect 21824 13028 21828 13084
rect 21828 13028 21884 13084
rect 21884 13028 21888 13084
rect 21824 13024 21888 13028
rect 21904 13084 21968 13088
rect 21904 13028 21908 13084
rect 21908 13028 21964 13084
rect 21964 13028 21968 13084
rect 21904 13024 21968 13028
rect 21984 13084 22048 13088
rect 21984 13028 21988 13084
rect 21988 13028 22044 13084
rect 22044 13028 22048 13084
rect 21984 13024 22048 13028
rect 3551 12540 3615 12544
rect 3551 12484 3555 12540
rect 3555 12484 3611 12540
rect 3611 12484 3615 12540
rect 3551 12480 3615 12484
rect 3631 12540 3695 12544
rect 3631 12484 3635 12540
rect 3635 12484 3691 12540
rect 3691 12484 3695 12540
rect 3631 12480 3695 12484
rect 3711 12540 3775 12544
rect 3711 12484 3715 12540
rect 3715 12484 3771 12540
rect 3771 12484 3775 12540
rect 3711 12480 3775 12484
rect 3791 12540 3855 12544
rect 3791 12484 3795 12540
rect 3795 12484 3851 12540
rect 3851 12484 3855 12540
rect 3791 12480 3855 12484
rect 8749 12540 8813 12544
rect 8749 12484 8753 12540
rect 8753 12484 8809 12540
rect 8809 12484 8813 12540
rect 8749 12480 8813 12484
rect 8829 12540 8893 12544
rect 8829 12484 8833 12540
rect 8833 12484 8889 12540
rect 8889 12484 8893 12540
rect 8829 12480 8893 12484
rect 8909 12540 8973 12544
rect 8909 12484 8913 12540
rect 8913 12484 8969 12540
rect 8969 12484 8973 12540
rect 8909 12480 8973 12484
rect 8989 12540 9053 12544
rect 8989 12484 8993 12540
rect 8993 12484 9049 12540
rect 9049 12484 9053 12540
rect 8989 12480 9053 12484
rect 13947 12540 14011 12544
rect 13947 12484 13951 12540
rect 13951 12484 14007 12540
rect 14007 12484 14011 12540
rect 13947 12480 14011 12484
rect 14027 12540 14091 12544
rect 14027 12484 14031 12540
rect 14031 12484 14087 12540
rect 14087 12484 14091 12540
rect 14027 12480 14091 12484
rect 14107 12540 14171 12544
rect 14107 12484 14111 12540
rect 14111 12484 14167 12540
rect 14167 12484 14171 12540
rect 14107 12480 14171 12484
rect 14187 12540 14251 12544
rect 14187 12484 14191 12540
rect 14191 12484 14247 12540
rect 14247 12484 14251 12540
rect 14187 12480 14251 12484
rect 19145 12540 19209 12544
rect 19145 12484 19149 12540
rect 19149 12484 19205 12540
rect 19205 12484 19209 12540
rect 19145 12480 19209 12484
rect 19225 12540 19289 12544
rect 19225 12484 19229 12540
rect 19229 12484 19285 12540
rect 19285 12484 19289 12540
rect 19225 12480 19289 12484
rect 19305 12540 19369 12544
rect 19305 12484 19309 12540
rect 19309 12484 19365 12540
rect 19365 12484 19369 12540
rect 19305 12480 19369 12484
rect 19385 12540 19449 12544
rect 19385 12484 19389 12540
rect 19389 12484 19445 12540
rect 19445 12484 19449 12540
rect 19385 12480 19449 12484
rect 8524 12276 8588 12340
rect 6150 11996 6214 12000
rect 6150 11940 6154 11996
rect 6154 11940 6210 11996
rect 6210 11940 6214 11996
rect 6150 11936 6214 11940
rect 6230 11996 6294 12000
rect 6230 11940 6234 11996
rect 6234 11940 6290 11996
rect 6290 11940 6294 11996
rect 6230 11936 6294 11940
rect 6310 11996 6374 12000
rect 6310 11940 6314 11996
rect 6314 11940 6370 11996
rect 6370 11940 6374 11996
rect 6310 11936 6374 11940
rect 6390 11996 6454 12000
rect 6390 11940 6394 11996
rect 6394 11940 6450 11996
rect 6450 11940 6454 11996
rect 6390 11936 6454 11940
rect 11348 11996 11412 12000
rect 11348 11940 11352 11996
rect 11352 11940 11408 11996
rect 11408 11940 11412 11996
rect 11348 11936 11412 11940
rect 11428 11996 11492 12000
rect 11428 11940 11432 11996
rect 11432 11940 11488 11996
rect 11488 11940 11492 11996
rect 11428 11936 11492 11940
rect 11508 11996 11572 12000
rect 11508 11940 11512 11996
rect 11512 11940 11568 11996
rect 11568 11940 11572 11996
rect 11508 11936 11572 11940
rect 11588 11996 11652 12000
rect 11588 11940 11592 11996
rect 11592 11940 11648 11996
rect 11648 11940 11652 11996
rect 11588 11936 11652 11940
rect 16546 11996 16610 12000
rect 16546 11940 16550 11996
rect 16550 11940 16606 11996
rect 16606 11940 16610 11996
rect 16546 11936 16610 11940
rect 16626 11996 16690 12000
rect 16626 11940 16630 11996
rect 16630 11940 16686 11996
rect 16686 11940 16690 11996
rect 16626 11936 16690 11940
rect 16706 11996 16770 12000
rect 16706 11940 16710 11996
rect 16710 11940 16766 11996
rect 16766 11940 16770 11996
rect 16706 11936 16770 11940
rect 16786 11996 16850 12000
rect 16786 11940 16790 11996
rect 16790 11940 16846 11996
rect 16846 11940 16850 11996
rect 16786 11936 16850 11940
rect 21744 11996 21808 12000
rect 21744 11940 21748 11996
rect 21748 11940 21804 11996
rect 21804 11940 21808 11996
rect 21744 11936 21808 11940
rect 21824 11996 21888 12000
rect 21824 11940 21828 11996
rect 21828 11940 21884 11996
rect 21884 11940 21888 11996
rect 21824 11936 21888 11940
rect 21904 11996 21968 12000
rect 21904 11940 21908 11996
rect 21908 11940 21964 11996
rect 21964 11940 21968 11996
rect 21904 11936 21968 11940
rect 21984 11996 22048 12000
rect 21984 11940 21988 11996
rect 21988 11940 22044 11996
rect 22044 11940 22048 11996
rect 21984 11936 22048 11940
rect 5028 11732 5092 11796
rect 3551 11452 3615 11456
rect 3551 11396 3555 11452
rect 3555 11396 3611 11452
rect 3611 11396 3615 11452
rect 3551 11392 3615 11396
rect 3631 11452 3695 11456
rect 3631 11396 3635 11452
rect 3635 11396 3691 11452
rect 3691 11396 3695 11452
rect 3631 11392 3695 11396
rect 3711 11452 3775 11456
rect 3711 11396 3715 11452
rect 3715 11396 3771 11452
rect 3771 11396 3775 11452
rect 3711 11392 3775 11396
rect 3791 11452 3855 11456
rect 3791 11396 3795 11452
rect 3795 11396 3851 11452
rect 3851 11396 3855 11452
rect 3791 11392 3855 11396
rect 8749 11452 8813 11456
rect 8749 11396 8753 11452
rect 8753 11396 8809 11452
rect 8809 11396 8813 11452
rect 8749 11392 8813 11396
rect 8829 11452 8893 11456
rect 8829 11396 8833 11452
rect 8833 11396 8889 11452
rect 8889 11396 8893 11452
rect 8829 11392 8893 11396
rect 8909 11452 8973 11456
rect 8909 11396 8913 11452
rect 8913 11396 8969 11452
rect 8969 11396 8973 11452
rect 8909 11392 8973 11396
rect 8989 11452 9053 11456
rect 8989 11396 8993 11452
rect 8993 11396 9049 11452
rect 9049 11396 9053 11452
rect 8989 11392 9053 11396
rect 13947 11452 14011 11456
rect 13947 11396 13951 11452
rect 13951 11396 14007 11452
rect 14007 11396 14011 11452
rect 13947 11392 14011 11396
rect 14027 11452 14091 11456
rect 14027 11396 14031 11452
rect 14031 11396 14087 11452
rect 14087 11396 14091 11452
rect 14027 11392 14091 11396
rect 14107 11452 14171 11456
rect 14107 11396 14111 11452
rect 14111 11396 14167 11452
rect 14167 11396 14171 11452
rect 14107 11392 14171 11396
rect 14187 11452 14251 11456
rect 14187 11396 14191 11452
rect 14191 11396 14247 11452
rect 14247 11396 14251 11452
rect 14187 11392 14251 11396
rect 19145 11452 19209 11456
rect 19145 11396 19149 11452
rect 19149 11396 19205 11452
rect 19205 11396 19209 11452
rect 19145 11392 19209 11396
rect 19225 11452 19289 11456
rect 19225 11396 19229 11452
rect 19229 11396 19285 11452
rect 19285 11396 19289 11452
rect 19225 11392 19289 11396
rect 19305 11452 19369 11456
rect 19305 11396 19309 11452
rect 19309 11396 19365 11452
rect 19365 11396 19369 11452
rect 19305 11392 19369 11396
rect 19385 11452 19449 11456
rect 19385 11396 19389 11452
rect 19389 11396 19445 11452
rect 19445 11396 19449 11452
rect 19385 11392 19449 11396
rect 6150 10908 6214 10912
rect 6150 10852 6154 10908
rect 6154 10852 6210 10908
rect 6210 10852 6214 10908
rect 6150 10848 6214 10852
rect 6230 10908 6294 10912
rect 6230 10852 6234 10908
rect 6234 10852 6290 10908
rect 6290 10852 6294 10908
rect 6230 10848 6294 10852
rect 6310 10908 6374 10912
rect 6310 10852 6314 10908
rect 6314 10852 6370 10908
rect 6370 10852 6374 10908
rect 6310 10848 6374 10852
rect 6390 10908 6454 10912
rect 6390 10852 6394 10908
rect 6394 10852 6450 10908
rect 6450 10852 6454 10908
rect 6390 10848 6454 10852
rect 11348 10908 11412 10912
rect 11348 10852 11352 10908
rect 11352 10852 11408 10908
rect 11408 10852 11412 10908
rect 11348 10848 11412 10852
rect 11428 10908 11492 10912
rect 11428 10852 11432 10908
rect 11432 10852 11488 10908
rect 11488 10852 11492 10908
rect 11428 10848 11492 10852
rect 11508 10908 11572 10912
rect 11508 10852 11512 10908
rect 11512 10852 11568 10908
rect 11568 10852 11572 10908
rect 11508 10848 11572 10852
rect 11588 10908 11652 10912
rect 11588 10852 11592 10908
rect 11592 10852 11648 10908
rect 11648 10852 11652 10908
rect 11588 10848 11652 10852
rect 16546 10908 16610 10912
rect 16546 10852 16550 10908
rect 16550 10852 16606 10908
rect 16606 10852 16610 10908
rect 16546 10848 16610 10852
rect 16626 10908 16690 10912
rect 16626 10852 16630 10908
rect 16630 10852 16686 10908
rect 16686 10852 16690 10908
rect 16626 10848 16690 10852
rect 16706 10908 16770 10912
rect 16706 10852 16710 10908
rect 16710 10852 16766 10908
rect 16766 10852 16770 10908
rect 16706 10848 16770 10852
rect 16786 10908 16850 10912
rect 16786 10852 16790 10908
rect 16790 10852 16846 10908
rect 16846 10852 16850 10908
rect 16786 10848 16850 10852
rect 21744 10908 21808 10912
rect 21744 10852 21748 10908
rect 21748 10852 21804 10908
rect 21804 10852 21808 10908
rect 21744 10848 21808 10852
rect 21824 10908 21888 10912
rect 21824 10852 21828 10908
rect 21828 10852 21884 10908
rect 21884 10852 21888 10908
rect 21824 10848 21888 10852
rect 21904 10908 21968 10912
rect 21904 10852 21908 10908
rect 21908 10852 21964 10908
rect 21964 10852 21968 10908
rect 21904 10848 21968 10852
rect 21984 10908 22048 10912
rect 21984 10852 21988 10908
rect 21988 10852 22044 10908
rect 22044 10852 22048 10908
rect 21984 10848 22048 10852
rect 3924 10508 3988 10572
rect 3551 10364 3615 10368
rect 3551 10308 3555 10364
rect 3555 10308 3611 10364
rect 3611 10308 3615 10364
rect 3551 10304 3615 10308
rect 3631 10364 3695 10368
rect 3631 10308 3635 10364
rect 3635 10308 3691 10364
rect 3691 10308 3695 10364
rect 3631 10304 3695 10308
rect 3711 10364 3775 10368
rect 3711 10308 3715 10364
rect 3715 10308 3771 10364
rect 3771 10308 3775 10364
rect 3711 10304 3775 10308
rect 3791 10364 3855 10368
rect 3791 10308 3795 10364
rect 3795 10308 3851 10364
rect 3851 10308 3855 10364
rect 3791 10304 3855 10308
rect 8749 10364 8813 10368
rect 8749 10308 8753 10364
rect 8753 10308 8809 10364
rect 8809 10308 8813 10364
rect 8749 10304 8813 10308
rect 8829 10364 8893 10368
rect 8829 10308 8833 10364
rect 8833 10308 8889 10364
rect 8889 10308 8893 10364
rect 8829 10304 8893 10308
rect 8909 10364 8973 10368
rect 8909 10308 8913 10364
rect 8913 10308 8969 10364
rect 8969 10308 8973 10364
rect 8909 10304 8973 10308
rect 8989 10364 9053 10368
rect 8989 10308 8993 10364
rect 8993 10308 9049 10364
rect 9049 10308 9053 10364
rect 8989 10304 9053 10308
rect 13947 10364 14011 10368
rect 13947 10308 13951 10364
rect 13951 10308 14007 10364
rect 14007 10308 14011 10364
rect 13947 10304 14011 10308
rect 14027 10364 14091 10368
rect 14027 10308 14031 10364
rect 14031 10308 14087 10364
rect 14087 10308 14091 10364
rect 14027 10304 14091 10308
rect 14107 10364 14171 10368
rect 14107 10308 14111 10364
rect 14111 10308 14167 10364
rect 14167 10308 14171 10364
rect 14107 10304 14171 10308
rect 14187 10364 14251 10368
rect 14187 10308 14191 10364
rect 14191 10308 14247 10364
rect 14247 10308 14251 10364
rect 14187 10304 14251 10308
rect 19145 10364 19209 10368
rect 19145 10308 19149 10364
rect 19149 10308 19205 10364
rect 19205 10308 19209 10364
rect 19145 10304 19209 10308
rect 19225 10364 19289 10368
rect 19225 10308 19229 10364
rect 19229 10308 19285 10364
rect 19285 10308 19289 10364
rect 19225 10304 19289 10308
rect 19305 10364 19369 10368
rect 19305 10308 19309 10364
rect 19309 10308 19365 10364
rect 19365 10308 19369 10364
rect 19305 10304 19369 10308
rect 19385 10364 19449 10368
rect 19385 10308 19389 10364
rect 19389 10308 19445 10364
rect 19445 10308 19449 10364
rect 19385 10304 19449 10308
rect 11836 10100 11900 10164
rect 6150 9820 6214 9824
rect 6150 9764 6154 9820
rect 6154 9764 6210 9820
rect 6210 9764 6214 9820
rect 6150 9760 6214 9764
rect 6230 9820 6294 9824
rect 6230 9764 6234 9820
rect 6234 9764 6290 9820
rect 6290 9764 6294 9820
rect 6230 9760 6294 9764
rect 6310 9820 6374 9824
rect 6310 9764 6314 9820
rect 6314 9764 6370 9820
rect 6370 9764 6374 9820
rect 6310 9760 6374 9764
rect 6390 9820 6454 9824
rect 6390 9764 6394 9820
rect 6394 9764 6450 9820
rect 6450 9764 6454 9820
rect 6390 9760 6454 9764
rect 11348 9820 11412 9824
rect 11348 9764 11352 9820
rect 11352 9764 11408 9820
rect 11408 9764 11412 9820
rect 11348 9760 11412 9764
rect 11428 9820 11492 9824
rect 11428 9764 11432 9820
rect 11432 9764 11488 9820
rect 11488 9764 11492 9820
rect 11428 9760 11492 9764
rect 11508 9820 11572 9824
rect 11508 9764 11512 9820
rect 11512 9764 11568 9820
rect 11568 9764 11572 9820
rect 11508 9760 11572 9764
rect 11588 9820 11652 9824
rect 11588 9764 11592 9820
rect 11592 9764 11648 9820
rect 11648 9764 11652 9820
rect 11588 9760 11652 9764
rect 16546 9820 16610 9824
rect 16546 9764 16550 9820
rect 16550 9764 16606 9820
rect 16606 9764 16610 9820
rect 16546 9760 16610 9764
rect 16626 9820 16690 9824
rect 16626 9764 16630 9820
rect 16630 9764 16686 9820
rect 16686 9764 16690 9820
rect 16626 9760 16690 9764
rect 16706 9820 16770 9824
rect 16706 9764 16710 9820
rect 16710 9764 16766 9820
rect 16766 9764 16770 9820
rect 16706 9760 16770 9764
rect 16786 9820 16850 9824
rect 16786 9764 16790 9820
rect 16790 9764 16846 9820
rect 16846 9764 16850 9820
rect 16786 9760 16850 9764
rect 21744 9820 21808 9824
rect 21744 9764 21748 9820
rect 21748 9764 21804 9820
rect 21804 9764 21808 9820
rect 21744 9760 21808 9764
rect 21824 9820 21888 9824
rect 21824 9764 21828 9820
rect 21828 9764 21884 9820
rect 21884 9764 21888 9820
rect 21824 9760 21888 9764
rect 21904 9820 21968 9824
rect 21904 9764 21908 9820
rect 21908 9764 21964 9820
rect 21964 9764 21968 9820
rect 21904 9760 21968 9764
rect 21984 9820 22048 9824
rect 21984 9764 21988 9820
rect 21988 9764 22044 9820
rect 22044 9764 22048 9820
rect 21984 9760 22048 9764
rect 8340 9692 8404 9756
rect 20484 9420 20548 9484
rect 3551 9276 3615 9280
rect 3551 9220 3555 9276
rect 3555 9220 3611 9276
rect 3611 9220 3615 9276
rect 3551 9216 3615 9220
rect 3631 9276 3695 9280
rect 3631 9220 3635 9276
rect 3635 9220 3691 9276
rect 3691 9220 3695 9276
rect 3631 9216 3695 9220
rect 3711 9276 3775 9280
rect 3711 9220 3715 9276
rect 3715 9220 3771 9276
rect 3771 9220 3775 9276
rect 3711 9216 3775 9220
rect 3791 9276 3855 9280
rect 3791 9220 3795 9276
rect 3795 9220 3851 9276
rect 3851 9220 3855 9276
rect 3791 9216 3855 9220
rect 8749 9276 8813 9280
rect 8749 9220 8753 9276
rect 8753 9220 8809 9276
rect 8809 9220 8813 9276
rect 8749 9216 8813 9220
rect 8829 9276 8893 9280
rect 8829 9220 8833 9276
rect 8833 9220 8889 9276
rect 8889 9220 8893 9276
rect 8829 9216 8893 9220
rect 8909 9276 8973 9280
rect 8909 9220 8913 9276
rect 8913 9220 8969 9276
rect 8969 9220 8973 9276
rect 8909 9216 8973 9220
rect 8989 9276 9053 9280
rect 8989 9220 8993 9276
rect 8993 9220 9049 9276
rect 9049 9220 9053 9276
rect 8989 9216 9053 9220
rect 13947 9276 14011 9280
rect 13947 9220 13951 9276
rect 13951 9220 14007 9276
rect 14007 9220 14011 9276
rect 13947 9216 14011 9220
rect 14027 9276 14091 9280
rect 14027 9220 14031 9276
rect 14031 9220 14087 9276
rect 14087 9220 14091 9276
rect 14027 9216 14091 9220
rect 14107 9276 14171 9280
rect 14107 9220 14111 9276
rect 14111 9220 14167 9276
rect 14167 9220 14171 9276
rect 14107 9216 14171 9220
rect 14187 9276 14251 9280
rect 14187 9220 14191 9276
rect 14191 9220 14247 9276
rect 14247 9220 14251 9276
rect 14187 9216 14251 9220
rect 19145 9276 19209 9280
rect 19145 9220 19149 9276
rect 19149 9220 19205 9276
rect 19205 9220 19209 9276
rect 19145 9216 19209 9220
rect 19225 9276 19289 9280
rect 19225 9220 19229 9276
rect 19229 9220 19285 9276
rect 19285 9220 19289 9276
rect 19225 9216 19289 9220
rect 19305 9276 19369 9280
rect 19305 9220 19309 9276
rect 19309 9220 19365 9276
rect 19365 9220 19369 9276
rect 19305 9216 19369 9220
rect 19385 9276 19449 9280
rect 19385 9220 19389 9276
rect 19389 9220 19445 9276
rect 19445 9220 19449 9276
rect 19385 9216 19449 9220
rect 7972 8876 8036 8940
rect 6150 8732 6214 8736
rect 6150 8676 6154 8732
rect 6154 8676 6210 8732
rect 6210 8676 6214 8732
rect 6150 8672 6214 8676
rect 6230 8732 6294 8736
rect 6230 8676 6234 8732
rect 6234 8676 6290 8732
rect 6290 8676 6294 8732
rect 6230 8672 6294 8676
rect 6310 8732 6374 8736
rect 6310 8676 6314 8732
rect 6314 8676 6370 8732
rect 6370 8676 6374 8732
rect 6310 8672 6374 8676
rect 6390 8732 6454 8736
rect 6390 8676 6394 8732
rect 6394 8676 6450 8732
rect 6450 8676 6454 8732
rect 6390 8672 6454 8676
rect 11348 8732 11412 8736
rect 11348 8676 11352 8732
rect 11352 8676 11408 8732
rect 11408 8676 11412 8732
rect 11348 8672 11412 8676
rect 11428 8732 11492 8736
rect 11428 8676 11432 8732
rect 11432 8676 11488 8732
rect 11488 8676 11492 8732
rect 11428 8672 11492 8676
rect 11508 8732 11572 8736
rect 11508 8676 11512 8732
rect 11512 8676 11568 8732
rect 11568 8676 11572 8732
rect 11508 8672 11572 8676
rect 11588 8732 11652 8736
rect 11588 8676 11592 8732
rect 11592 8676 11648 8732
rect 11648 8676 11652 8732
rect 11588 8672 11652 8676
rect 16546 8732 16610 8736
rect 16546 8676 16550 8732
rect 16550 8676 16606 8732
rect 16606 8676 16610 8732
rect 16546 8672 16610 8676
rect 16626 8732 16690 8736
rect 16626 8676 16630 8732
rect 16630 8676 16686 8732
rect 16686 8676 16690 8732
rect 16626 8672 16690 8676
rect 16706 8732 16770 8736
rect 16706 8676 16710 8732
rect 16710 8676 16766 8732
rect 16766 8676 16770 8732
rect 16706 8672 16770 8676
rect 16786 8732 16850 8736
rect 16786 8676 16790 8732
rect 16790 8676 16846 8732
rect 16846 8676 16850 8732
rect 16786 8672 16850 8676
rect 21744 8732 21808 8736
rect 21744 8676 21748 8732
rect 21748 8676 21804 8732
rect 21804 8676 21808 8732
rect 21744 8672 21808 8676
rect 21824 8732 21888 8736
rect 21824 8676 21828 8732
rect 21828 8676 21884 8732
rect 21884 8676 21888 8732
rect 21824 8672 21888 8676
rect 21904 8732 21968 8736
rect 21904 8676 21908 8732
rect 21908 8676 21964 8732
rect 21964 8676 21968 8732
rect 21904 8672 21968 8676
rect 21984 8732 22048 8736
rect 21984 8676 21988 8732
rect 21988 8676 22044 8732
rect 22044 8676 22048 8732
rect 21984 8672 22048 8676
rect 3551 8188 3615 8192
rect 3551 8132 3555 8188
rect 3555 8132 3611 8188
rect 3611 8132 3615 8188
rect 3551 8128 3615 8132
rect 3631 8188 3695 8192
rect 3631 8132 3635 8188
rect 3635 8132 3691 8188
rect 3691 8132 3695 8188
rect 3631 8128 3695 8132
rect 3711 8188 3775 8192
rect 3711 8132 3715 8188
rect 3715 8132 3771 8188
rect 3771 8132 3775 8188
rect 3711 8128 3775 8132
rect 3791 8188 3855 8192
rect 3791 8132 3795 8188
rect 3795 8132 3851 8188
rect 3851 8132 3855 8188
rect 3791 8128 3855 8132
rect 8749 8188 8813 8192
rect 8749 8132 8753 8188
rect 8753 8132 8809 8188
rect 8809 8132 8813 8188
rect 8749 8128 8813 8132
rect 8829 8188 8893 8192
rect 8829 8132 8833 8188
rect 8833 8132 8889 8188
rect 8889 8132 8893 8188
rect 8829 8128 8893 8132
rect 8909 8188 8973 8192
rect 8909 8132 8913 8188
rect 8913 8132 8969 8188
rect 8969 8132 8973 8188
rect 8909 8128 8973 8132
rect 8989 8188 9053 8192
rect 8989 8132 8993 8188
rect 8993 8132 9049 8188
rect 9049 8132 9053 8188
rect 8989 8128 9053 8132
rect 13947 8188 14011 8192
rect 13947 8132 13951 8188
rect 13951 8132 14007 8188
rect 14007 8132 14011 8188
rect 13947 8128 14011 8132
rect 14027 8188 14091 8192
rect 14027 8132 14031 8188
rect 14031 8132 14087 8188
rect 14087 8132 14091 8188
rect 14027 8128 14091 8132
rect 14107 8188 14171 8192
rect 14107 8132 14111 8188
rect 14111 8132 14167 8188
rect 14167 8132 14171 8188
rect 14107 8128 14171 8132
rect 14187 8188 14251 8192
rect 14187 8132 14191 8188
rect 14191 8132 14247 8188
rect 14247 8132 14251 8188
rect 14187 8128 14251 8132
rect 19145 8188 19209 8192
rect 19145 8132 19149 8188
rect 19149 8132 19205 8188
rect 19205 8132 19209 8188
rect 19145 8128 19209 8132
rect 19225 8188 19289 8192
rect 19225 8132 19229 8188
rect 19229 8132 19285 8188
rect 19285 8132 19289 8188
rect 19225 8128 19289 8132
rect 19305 8188 19369 8192
rect 19305 8132 19309 8188
rect 19309 8132 19365 8188
rect 19365 8132 19369 8188
rect 19305 8128 19369 8132
rect 19385 8188 19449 8192
rect 19385 8132 19389 8188
rect 19389 8132 19445 8188
rect 19445 8132 19449 8188
rect 19385 8128 19449 8132
rect 8156 7924 8220 7988
rect 11836 7788 11900 7852
rect 6150 7644 6214 7648
rect 6150 7588 6154 7644
rect 6154 7588 6210 7644
rect 6210 7588 6214 7644
rect 6150 7584 6214 7588
rect 6230 7644 6294 7648
rect 6230 7588 6234 7644
rect 6234 7588 6290 7644
rect 6290 7588 6294 7644
rect 6230 7584 6294 7588
rect 6310 7644 6374 7648
rect 6310 7588 6314 7644
rect 6314 7588 6370 7644
rect 6370 7588 6374 7644
rect 6310 7584 6374 7588
rect 6390 7644 6454 7648
rect 6390 7588 6394 7644
rect 6394 7588 6450 7644
rect 6450 7588 6454 7644
rect 6390 7584 6454 7588
rect 11348 7644 11412 7648
rect 11348 7588 11352 7644
rect 11352 7588 11408 7644
rect 11408 7588 11412 7644
rect 11348 7584 11412 7588
rect 11428 7644 11492 7648
rect 11428 7588 11432 7644
rect 11432 7588 11488 7644
rect 11488 7588 11492 7644
rect 11428 7584 11492 7588
rect 11508 7644 11572 7648
rect 11508 7588 11512 7644
rect 11512 7588 11568 7644
rect 11568 7588 11572 7644
rect 11508 7584 11572 7588
rect 11588 7644 11652 7648
rect 11588 7588 11592 7644
rect 11592 7588 11648 7644
rect 11648 7588 11652 7644
rect 11588 7584 11652 7588
rect 16546 7644 16610 7648
rect 16546 7588 16550 7644
rect 16550 7588 16606 7644
rect 16606 7588 16610 7644
rect 16546 7584 16610 7588
rect 16626 7644 16690 7648
rect 16626 7588 16630 7644
rect 16630 7588 16686 7644
rect 16686 7588 16690 7644
rect 16626 7584 16690 7588
rect 16706 7644 16770 7648
rect 16706 7588 16710 7644
rect 16710 7588 16766 7644
rect 16766 7588 16770 7644
rect 16706 7584 16770 7588
rect 16786 7644 16850 7648
rect 16786 7588 16790 7644
rect 16790 7588 16846 7644
rect 16846 7588 16850 7644
rect 16786 7584 16850 7588
rect 21744 7644 21808 7648
rect 21744 7588 21748 7644
rect 21748 7588 21804 7644
rect 21804 7588 21808 7644
rect 21744 7584 21808 7588
rect 21824 7644 21888 7648
rect 21824 7588 21828 7644
rect 21828 7588 21884 7644
rect 21884 7588 21888 7644
rect 21824 7584 21888 7588
rect 21904 7644 21968 7648
rect 21904 7588 21908 7644
rect 21908 7588 21964 7644
rect 21964 7588 21968 7644
rect 21904 7584 21968 7588
rect 21984 7644 22048 7648
rect 21984 7588 21988 7644
rect 21988 7588 22044 7644
rect 22044 7588 22048 7644
rect 21984 7584 22048 7588
rect 3551 7100 3615 7104
rect 3551 7044 3555 7100
rect 3555 7044 3611 7100
rect 3611 7044 3615 7100
rect 3551 7040 3615 7044
rect 3631 7100 3695 7104
rect 3631 7044 3635 7100
rect 3635 7044 3691 7100
rect 3691 7044 3695 7100
rect 3631 7040 3695 7044
rect 3711 7100 3775 7104
rect 3711 7044 3715 7100
rect 3715 7044 3771 7100
rect 3771 7044 3775 7100
rect 3711 7040 3775 7044
rect 3791 7100 3855 7104
rect 3791 7044 3795 7100
rect 3795 7044 3851 7100
rect 3851 7044 3855 7100
rect 3791 7040 3855 7044
rect 8749 7100 8813 7104
rect 8749 7044 8753 7100
rect 8753 7044 8809 7100
rect 8809 7044 8813 7100
rect 8749 7040 8813 7044
rect 8829 7100 8893 7104
rect 8829 7044 8833 7100
rect 8833 7044 8889 7100
rect 8889 7044 8893 7100
rect 8829 7040 8893 7044
rect 8909 7100 8973 7104
rect 8909 7044 8913 7100
rect 8913 7044 8969 7100
rect 8969 7044 8973 7100
rect 8909 7040 8973 7044
rect 8989 7100 9053 7104
rect 8989 7044 8993 7100
rect 8993 7044 9049 7100
rect 9049 7044 9053 7100
rect 8989 7040 9053 7044
rect 13947 7100 14011 7104
rect 13947 7044 13951 7100
rect 13951 7044 14007 7100
rect 14007 7044 14011 7100
rect 13947 7040 14011 7044
rect 14027 7100 14091 7104
rect 14027 7044 14031 7100
rect 14031 7044 14087 7100
rect 14087 7044 14091 7100
rect 14027 7040 14091 7044
rect 14107 7100 14171 7104
rect 14107 7044 14111 7100
rect 14111 7044 14167 7100
rect 14167 7044 14171 7100
rect 14107 7040 14171 7044
rect 14187 7100 14251 7104
rect 14187 7044 14191 7100
rect 14191 7044 14247 7100
rect 14247 7044 14251 7100
rect 14187 7040 14251 7044
rect 19145 7100 19209 7104
rect 19145 7044 19149 7100
rect 19149 7044 19205 7100
rect 19205 7044 19209 7100
rect 19145 7040 19209 7044
rect 19225 7100 19289 7104
rect 19225 7044 19229 7100
rect 19229 7044 19285 7100
rect 19285 7044 19289 7100
rect 19225 7040 19289 7044
rect 19305 7100 19369 7104
rect 19305 7044 19309 7100
rect 19309 7044 19365 7100
rect 19365 7044 19369 7100
rect 19305 7040 19369 7044
rect 19385 7100 19449 7104
rect 19385 7044 19389 7100
rect 19389 7044 19445 7100
rect 19445 7044 19449 7100
rect 19385 7040 19449 7044
rect 6150 6556 6214 6560
rect 6150 6500 6154 6556
rect 6154 6500 6210 6556
rect 6210 6500 6214 6556
rect 6150 6496 6214 6500
rect 6230 6556 6294 6560
rect 6230 6500 6234 6556
rect 6234 6500 6290 6556
rect 6290 6500 6294 6556
rect 6230 6496 6294 6500
rect 6310 6556 6374 6560
rect 6310 6500 6314 6556
rect 6314 6500 6370 6556
rect 6370 6500 6374 6556
rect 6310 6496 6374 6500
rect 6390 6556 6454 6560
rect 6390 6500 6394 6556
rect 6394 6500 6450 6556
rect 6450 6500 6454 6556
rect 6390 6496 6454 6500
rect 11348 6556 11412 6560
rect 11348 6500 11352 6556
rect 11352 6500 11408 6556
rect 11408 6500 11412 6556
rect 11348 6496 11412 6500
rect 11428 6556 11492 6560
rect 11428 6500 11432 6556
rect 11432 6500 11488 6556
rect 11488 6500 11492 6556
rect 11428 6496 11492 6500
rect 11508 6556 11572 6560
rect 11508 6500 11512 6556
rect 11512 6500 11568 6556
rect 11568 6500 11572 6556
rect 11508 6496 11572 6500
rect 11588 6556 11652 6560
rect 11588 6500 11592 6556
rect 11592 6500 11648 6556
rect 11648 6500 11652 6556
rect 11588 6496 11652 6500
rect 16546 6556 16610 6560
rect 16546 6500 16550 6556
rect 16550 6500 16606 6556
rect 16606 6500 16610 6556
rect 16546 6496 16610 6500
rect 16626 6556 16690 6560
rect 16626 6500 16630 6556
rect 16630 6500 16686 6556
rect 16686 6500 16690 6556
rect 16626 6496 16690 6500
rect 16706 6556 16770 6560
rect 16706 6500 16710 6556
rect 16710 6500 16766 6556
rect 16766 6500 16770 6556
rect 16706 6496 16770 6500
rect 16786 6556 16850 6560
rect 16786 6500 16790 6556
rect 16790 6500 16846 6556
rect 16846 6500 16850 6556
rect 16786 6496 16850 6500
rect 21744 6556 21808 6560
rect 21744 6500 21748 6556
rect 21748 6500 21804 6556
rect 21804 6500 21808 6556
rect 21744 6496 21808 6500
rect 21824 6556 21888 6560
rect 21824 6500 21828 6556
rect 21828 6500 21884 6556
rect 21884 6500 21888 6556
rect 21824 6496 21888 6500
rect 21904 6556 21968 6560
rect 21904 6500 21908 6556
rect 21908 6500 21964 6556
rect 21964 6500 21968 6556
rect 21904 6496 21968 6500
rect 21984 6556 22048 6560
rect 21984 6500 21988 6556
rect 21988 6500 22044 6556
rect 22044 6500 22048 6556
rect 21984 6496 22048 6500
rect 3551 6012 3615 6016
rect 3551 5956 3555 6012
rect 3555 5956 3611 6012
rect 3611 5956 3615 6012
rect 3551 5952 3615 5956
rect 3631 6012 3695 6016
rect 3631 5956 3635 6012
rect 3635 5956 3691 6012
rect 3691 5956 3695 6012
rect 3631 5952 3695 5956
rect 3711 6012 3775 6016
rect 3711 5956 3715 6012
rect 3715 5956 3771 6012
rect 3771 5956 3775 6012
rect 3711 5952 3775 5956
rect 3791 6012 3855 6016
rect 3791 5956 3795 6012
rect 3795 5956 3851 6012
rect 3851 5956 3855 6012
rect 3791 5952 3855 5956
rect 8749 6012 8813 6016
rect 8749 5956 8753 6012
rect 8753 5956 8809 6012
rect 8809 5956 8813 6012
rect 8749 5952 8813 5956
rect 8829 6012 8893 6016
rect 8829 5956 8833 6012
rect 8833 5956 8889 6012
rect 8889 5956 8893 6012
rect 8829 5952 8893 5956
rect 8909 6012 8973 6016
rect 8909 5956 8913 6012
rect 8913 5956 8969 6012
rect 8969 5956 8973 6012
rect 8909 5952 8973 5956
rect 8989 6012 9053 6016
rect 8989 5956 8993 6012
rect 8993 5956 9049 6012
rect 9049 5956 9053 6012
rect 8989 5952 9053 5956
rect 13947 6012 14011 6016
rect 13947 5956 13951 6012
rect 13951 5956 14007 6012
rect 14007 5956 14011 6012
rect 13947 5952 14011 5956
rect 14027 6012 14091 6016
rect 14027 5956 14031 6012
rect 14031 5956 14087 6012
rect 14087 5956 14091 6012
rect 14027 5952 14091 5956
rect 14107 6012 14171 6016
rect 14107 5956 14111 6012
rect 14111 5956 14167 6012
rect 14167 5956 14171 6012
rect 14107 5952 14171 5956
rect 14187 6012 14251 6016
rect 14187 5956 14191 6012
rect 14191 5956 14247 6012
rect 14247 5956 14251 6012
rect 14187 5952 14251 5956
rect 19145 6012 19209 6016
rect 19145 5956 19149 6012
rect 19149 5956 19205 6012
rect 19205 5956 19209 6012
rect 19145 5952 19209 5956
rect 19225 6012 19289 6016
rect 19225 5956 19229 6012
rect 19229 5956 19285 6012
rect 19285 5956 19289 6012
rect 19225 5952 19289 5956
rect 19305 6012 19369 6016
rect 19305 5956 19309 6012
rect 19309 5956 19365 6012
rect 19365 5956 19369 6012
rect 19305 5952 19369 5956
rect 19385 6012 19449 6016
rect 19385 5956 19389 6012
rect 19389 5956 19445 6012
rect 19445 5956 19449 6012
rect 19385 5952 19449 5956
rect 6150 5468 6214 5472
rect 6150 5412 6154 5468
rect 6154 5412 6210 5468
rect 6210 5412 6214 5468
rect 6150 5408 6214 5412
rect 6230 5468 6294 5472
rect 6230 5412 6234 5468
rect 6234 5412 6290 5468
rect 6290 5412 6294 5468
rect 6230 5408 6294 5412
rect 6310 5468 6374 5472
rect 6310 5412 6314 5468
rect 6314 5412 6370 5468
rect 6370 5412 6374 5468
rect 6310 5408 6374 5412
rect 6390 5468 6454 5472
rect 6390 5412 6394 5468
rect 6394 5412 6450 5468
rect 6450 5412 6454 5468
rect 6390 5408 6454 5412
rect 11348 5468 11412 5472
rect 11348 5412 11352 5468
rect 11352 5412 11408 5468
rect 11408 5412 11412 5468
rect 11348 5408 11412 5412
rect 11428 5468 11492 5472
rect 11428 5412 11432 5468
rect 11432 5412 11488 5468
rect 11488 5412 11492 5468
rect 11428 5408 11492 5412
rect 11508 5468 11572 5472
rect 11508 5412 11512 5468
rect 11512 5412 11568 5468
rect 11568 5412 11572 5468
rect 11508 5408 11572 5412
rect 11588 5468 11652 5472
rect 11588 5412 11592 5468
rect 11592 5412 11648 5468
rect 11648 5412 11652 5468
rect 11588 5408 11652 5412
rect 16546 5468 16610 5472
rect 16546 5412 16550 5468
rect 16550 5412 16606 5468
rect 16606 5412 16610 5468
rect 16546 5408 16610 5412
rect 16626 5468 16690 5472
rect 16626 5412 16630 5468
rect 16630 5412 16686 5468
rect 16686 5412 16690 5468
rect 16626 5408 16690 5412
rect 16706 5468 16770 5472
rect 16706 5412 16710 5468
rect 16710 5412 16766 5468
rect 16766 5412 16770 5468
rect 16706 5408 16770 5412
rect 16786 5468 16850 5472
rect 16786 5412 16790 5468
rect 16790 5412 16846 5468
rect 16846 5412 16850 5468
rect 16786 5408 16850 5412
rect 21744 5468 21808 5472
rect 21744 5412 21748 5468
rect 21748 5412 21804 5468
rect 21804 5412 21808 5468
rect 21744 5408 21808 5412
rect 21824 5468 21888 5472
rect 21824 5412 21828 5468
rect 21828 5412 21884 5468
rect 21884 5412 21888 5468
rect 21824 5408 21888 5412
rect 21904 5468 21968 5472
rect 21904 5412 21908 5468
rect 21908 5412 21964 5468
rect 21964 5412 21968 5468
rect 21904 5408 21968 5412
rect 21984 5468 22048 5472
rect 21984 5412 21988 5468
rect 21988 5412 22044 5468
rect 22044 5412 22048 5468
rect 21984 5408 22048 5412
rect 3551 4924 3615 4928
rect 3551 4868 3555 4924
rect 3555 4868 3611 4924
rect 3611 4868 3615 4924
rect 3551 4864 3615 4868
rect 3631 4924 3695 4928
rect 3631 4868 3635 4924
rect 3635 4868 3691 4924
rect 3691 4868 3695 4924
rect 3631 4864 3695 4868
rect 3711 4924 3775 4928
rect 3711 4868 3715 4924
rect 3715 4868 3771 4924
rect 3771 4868 3775 4924
rect 3711 4864 3775 4868
rect 3791 4924 3855 4928
rect 3791 4868 3795 4924
rect 3795 4868 3851 4924
rect 3851 4868 3855 4924
rect 3791 4864 3855 4868
rect 8749 4924 8813 4928
rect 8749 4868 8753 4924
rect 8753 4868 8809 4924
rect 8809 4868 8813 4924
rect 8749 4864 8813 4868
rect 8829 4924 8893 4928
rect 8829 4868 8833 4924
rect 8833 4868 8889 4924
rect 8889 4868 8893 4924
rect 8829 4864 8893 4868
rect 8909 4924 8973 4928
rect 8909 4868 8913 4924
rect 8913 4868 8969 4924
rect 8969 4868 8973 4924
rect 8909 4864 8973 4868
rect 8989 4924 9053 4928
rect 8989 4868 8993 4924
rect 8993 4868 9049 4924
rect 9049 4868 9053 4924
rect 8989 4864 9053 4868
rect 13947 4924 14011 4928
rect 13947 4868 13951 4924
rect 13951 4868 14007 4924
rect 14007 4868 14011 4924
rect 13947 4864 14011 4868
rect 14027 4924 14091 4928
rect 14027 4868 14031 4924
rect 14031 4868 14087 4924
rect 14087 4868 14091 4924
rect 14027 4864 14091 4868
rect 14107 4924 14171 4928
rect 14107 4868 14111 4924
rect 14111 4868 14167 4924
rect 14167 4868 14171 4924
rect 14107 4864 14171 4868
rect 14187 4924 14251 4928
rect 14187 4868 14191 4924
rect 14191 4868 14247 4924
rect 14247 4868 14251 4924
rect 14187 4864 14251 4868
rect 19145 4924 19209 4928
rect 19145 4868 19149 4924
rect 19149 4868 19205 4924
rect 19205 4868 19209 4924
rect 19145 4864 19209 4868
rect 19225 4924 19289 4928
rect 19225 4868 19229 4924
rect 19229 4868 19285 4924
rect 19285 4868 19289 4924
rect 19225 4864 19289 4868
rect 19305 4924 19369 4928
rect 19305 4868 19309 4924
rect 19309 4868 19365 4924
rect 19365 4868 19369 4924
rect 19305 4864 19369 4868
rect 19385 4924 19449 4928
rect 19385 4868 19389 4924
rect 19389 4868 19445 4924
rect 19445 4868 19449 4924
rect 19385 4864 19449 4868
rect 6150 4380 6214 4384
rect 6150 4324 6154 4380
rect 6154 4324 6210 4380
rect 6210 4324 6214 4380
rect 6150 4320 6214 4324
rect 6230 4380 6294 4384
rect 6230 4324 6234 4380
rect 6234 4324 6290 4380
rect 6290 4324 6294 4380
rect 6230 4320 6294 4324
rect 6310 4380 6374 4384
rect 6310 4324 6314 4380
rect 6314 4324 6370 4380
rect 6370 4324 6374 4380
rect 6310 4320 6374 4324
rect 6390 4380 6454 4384
rect 6390 4324 6394 4380
rect 6394 4324 6450 4380
rect 6450 4324 6454 4380
rect 6390 4320 6454 4324
rect 11348 4380 11412 4384
rect 11348 4324 11352 4380
rect 11352 4324 11408 4380
rect 11408 4324 11412 4380
rect 11348 4320 11412 4324
rect 11428 4380 11492 4384
rect 11428 4324 11432 4380
rect 11432 4324 11488 4380
rect 11488 4324 11492 4380
rect 11428 4320 11492 4324
rect 11508 4380 11572 4384
rect 11508 4324 11512 4380
rect 11512 4324 11568 4380
rect 11568 4324 11572 4380
rect 11508 4320 11572 4324
rect 11588 4380 11652 4384
rect 11588 4324 11592 4380
rect 11592 4324 11648 4380
rect 11648 4324 11652 4380
rect 11588 4320 11652 4324
rect 16546 4380 16610 4384
rect 16546 4324 16550 4380
rect 16550 4324 16606 4380
rect 16606 4324 16610 4380
rect 16546 4320 16610 4324
rect 16626 4380 16690 4384
rect 16626 4324 16630 4380
rect 16630 4324 16686 4380
rect 16686 4324 16690 4380
rect 16626 4320 16690 4324
rect 16706 4380 16770 4384
rect 16706 4324 16710 4380
rect 16710 4324 16766 4380
rect 16766 4324 16770 4380
rect 16706 4320 16770 4324
rect 16786 4380 16850 4384
rect 16786 4324 16790 4380
rect 16790 4324 16846 4380
rect 16846 4324 16850 4380
rect 16786 4320 16850 4324
rect 21744 4380 21808 4384
rect 21744 4324 21748 4380
rect 21748 4324 21804 4380
rect 21804 4324 21808 4380
rect 21744 4320 21808 4324
rect 21824 4380 21888 4384
rect 21824 4324 21828 4380
rect 21828 4324 21884 4380
rect 21884 4324 21888 4380
rect 21824 4320 21888 4324
rect 21904 4380 21968 4384
rect 21904 4324 21908 4380
rect 21908 4324 21964 4380
rect 21964 4324 21968 4380
rect 21904 4320 21968 4324
rect 21984 4380 22048 4384
rect 21984 4324 21988 4380
rect 21988 4324 22044 4380
rect 22044 4324 22048 4380
rect 21984 4320 22048 4324
rect 3551 3836 3615 3840
rect 3551 3780 3555 3836
rect 3555 3780 3611 3836
rect 3611 3780 3615 3836
rect 3551 3776 3615 3780
rect 3631 3836 3695 3840
rect 3631 3780 3635 3836
rect 3635 3780 3691 3836
rect 3691 3780 3695 3836
rect 3631 3776 3695 3780
rect 3711 3836 3775 3840
rect 3711 3780 3715 3836
rect 3715 3780 3771 3836
rect 3771 3780 3775 3836
rect 3711 3776 3775 3780
rect 3791 3836 3855 3840
rect 3791 3780 3795 3836
rect 3795 3780 3851 3836
rect 3851 3780 3855 3836
rect 3791 3776 3855 3780
rect 8749 3836 8813 3840
rect 8749 3780 8753 3836
rect 8753 3780 8809 3836
rect 8809 3780 8813 3836
rect 8749 3776 8813 3780
rect 8829 3836 8893 3840
rect 8829 3780 8833 3836
rect 8833 3780 8889 3836
rect 8889 3780 8893 3836
rect 8829 3776 8893 3780
rect 8909 3836 8973 3840
rect 8909 3780 8913 3836
rect 8913 3780 8969 3836
rect 8969 3780 8973 3836
rect 8909 3776 8973 3780
rect 8989 3836 9053 3840
rect 8989 3780 8993 3836
rect 8993 3780 9049 3836
rect 9049 3780 9053 3836
rect 8989 3776 9053 3780
rect 13947 3836 14011 3840
rect 13947 3780 13951 3836
rect 13951 3780 14007 3836
rect 14007 3780 14011 3836
rect 13947 3776 14011 3780
rect 14027 3836 14091 3840
rect 14027 3780 14031 3836
rect 14031 3780 14087 3836
rect 14087 3780 14091 3836
rect 14027 3776 14091 3780
rect 14107 3836 14171 3840
rect 14107 3780 14111 3836
rect 14111 3780 14167 3836
rect 14167 3780 14171 3836
rect 14107 3776 14171 3780
rect 14187 3836 14251 3840
rect 14187 3780 14191 3836
rect 14191 3780 14247 3836
rect 14247 3780 14251 3836
rect 14187 3776 14251 3780
rect 19145 3836 19209 3840
rect 19145 3780 19149 3836
rect 19149 3780 19205 3836
rect 19205 3780 19209 3836
rect 19145 3776 19209 3780
rect 19225 3836 19289 3840
rect 19225 3780 19229 3836
rect 19229 3780 19285 3836
rect 19285 3780 19289 3836
rect 19225 3776 19289 3780
rect 19305 3836 19369 3840
rect 19305 3780 19309 3836
rect 19309 3780 19365 3836
rect 19365 3780 19369 3836
rect 19305 3776 19369 3780
rect 19385 3836 19449 3840
rect 19385 3780 19389 3836
rect 19389 3780 19445 3836
rect 19445 3780 19449 3836
rect 19385 3776 19449 3780
rect 5948 3496 6012 3500
rect 5948 3440 5998 3496
rect 5998 3440 6012 3496
rect 5948 3436 6012 3440
rect 6150 3292 6214 3296
rect 6150 3236 6154 3292
rect 6154 3236 6210 3292
rect 6210 3236 6214 3292
rect 6150 3232 6214 3236
rect 6230 3292 6294 3296
rect 6230 3236 6234 3292
rect 6234 3236 6290 3292
rect 6290 3236 6294 3292
rect 6230 3232 6294 3236
rect 6310 3292 6374 3296
rect 6310 3236 6314 3292
rect 6314 3236 6370 3292
rect 6370 3236 6374 3292
rect 6310 3232 6374 3236
rect 6390 3292 6454 3296
rect 6390 3236 6394 3292
rect 6394 3236 6450 3292
rect 6450 3236 6454 3292
rect 6390 3232 6454 3236
rect 11348 3292 11412 3296
rect 11348 3236 11352 3292
rect 11352 3236 11408 3292
rect 11408 3236 11412 3292
rect 11348 3232 11412 3236
rect 11428 3292 11492 3296
rect 11428 3236 11432 3292
rect 11432 3236 11488 3292
rect 11488 3236 11492 3292
rect 11428 3232 11492 3236
rect 11508 3292 11572 3296
rect 11508 3236 11512 3292
rect 11512 3236 11568 3292
rect 11568 3236 11572 3292
rect 11508 3232 11572 3236
rect 11588 3292 11652 3296
rect 11588 3236 11592 3292
rect 11592 3236 11648 3292
rect 11648 3236 11652 3292
rect 11588 3232 11652 3236
rect 16546 3292 16610 3296
rect 16546 3236 16550 3292
rect 16550 3236 16606 3292
rect 16606 3236 16610 3292
rect 16546 3232 16610 3236
rect 16626 3292 16690 3296
rect 16626 3236 16630 3292
rect 16630 3236 16686 3292
rect 16686 3236 16690 3292
rect 16626 3232 16690 3236
rect 16706 3292 16770 3296
rect 16706 3236 16710 3292
rect 16710 3236 16766 3292
rect 16766 3236 16770 3292
rect 16706 3232 16770 3236
rect 16786 3292 16850 3296
rect 16786 3236 16790 3292
rect 16790 3236 16846 3292
rect 16846 3236 16850 3292
rect 16786 3232 16850 3236
rect 21744 3292 21808 3296
rect 21744 3236 21748 3292
rect 21748 3236 21804 3292
rect 21804 3236 21808 3292
rect 21744 3232 21808 3236
rect 21824 3292 21888 3296
rect 21824 3236 21828 3292
rect 21828 3236 21884 3292
rect 21884 3236 21888 3292
rect 21824 3232 21888 3236
rect 21904 3292 21968 3296
rect 21904 3236 21908 3292
rect 21908 3236 21964 3292
rect 21964 3236 21968 3292
rect 21904 3232 21968 3236
rect 21984 3292 22048 3296
rect 21984 3236 21988 3292
rect 21988 3236 22044 3292
rect 22044 3236 22048 3292
rect 21984 3232 22048 3236
rect 4108 2892 4172 2956
rect 3551 2748 3615 2752
rect 3551 2692 3555 2748
rect 3555 2692 3611 2748
rect 3611 2692 3615 2748
rect 3551 2688 3615 2692
rect 3631 2748 3695 2752
rect 3631 2692 3635 2748
rect 3635 2692 3691 2748
rect 3691 2692 3695 2748
rect 3631 2688 3695 2692
rect 3711 2748 3775 2752
rect 3711 2692 3715 2748
rect 3715 2692 3771 2748
rect 3771 2692 3775 2748
rect 3711 2688 3775 2692
rect 3791 2748 3855 2752
rect 3791 2692 3795 2748
rect 3795 2692 3851 2748
rect 3851 2692 3855 2748
rect 3791 2688 3855 2692
rect 8749 2748 8813 2752
rect 8749 2692 8753 2748
rect 8753 2692 8809 2748
rect 8809 2692 8813 2748
rect 8749 2688 8813 2692
rect 8829 2748 8893 2752
rect 8829 2692 8833 2748
rect 8833 2692 8889 2748
rect 8889 2692 8893 2748
rect 8829 2688 8893 2692
rect 8909 2748 8973 2752
rect 8909 2692 8913 2748
rect 8913 2692 8969 2748
rect 8969 2692 8973 2748
rect 8909 2688 8973 2692
rect 8989 2748 9053 2752
rect 8989 2692 8993 2748
rect 8993 2692 9049 2748
rect 9049 2692 9053 2748
rect 8989 2688 9053 2692
rect 13947 2748 14011 2752
rect 13947 2692 13951 2748
rect 13951 2692 14007 2748
rect 14007 2692 14011 2748
rect 13947 2688 14011 2692
rect 14027 2748 14091 2752
rect 14027 2692 14031 2748
rect 14031 2692 14087 2748
rect 14087 2692 14091 2748
rect 14027 2688 14091 2692
rect 14107 2748 14171 2752
rect 14107 2692 14111 2748
rect 14111 2692 14167 2748
rect 14167 2692 14171 2748
rect 14107 2688 14171 2692
rect 14187 2748 14251 2752
rect 14187 2692 14191 2748
rect 14191 2692 14247 2748
rect 14247 2692 14251 2748
rect 14187 2688 14251 2692
rect 19145 2748 19209 2752
rect 19145 2692 19149 2748
rect 19149 2692 19205 2748
rect 19205 2692 19209 2748
rect 19145 2688 19209 2692
rect 19225 2748 19289 2752
rect 19225 2692 19229 2748
rect 19229 2692 19285 2748
rect 19285 2692 19289 2748
rect 19225 2688 19289 2692
rect 19305 2748 19369 2752
rect 19305 2692 19309 2748
rect 19309 2692 19365 2748
rect 19365 2692 19369 2748
rect 19305 2688 19369 2692
rect 19385 2748 19449 2752
rect 19385 2692 19389 2748
rect 19389 2692 19445 2748
rect 19445 2692 19449 2748
rect 19385 2688 19449 2692
rect 6150 2204 6214 2208
rect 6150 2148 6154 2204
rect 6154 2148 6210 2204
rect 6210 2148 6214 2204
rect 6150 2144 6214 2148
rect 6230 2204 6294 2208
rect 6230 2148 6234 2204
rect 6234 2148 6290 2204
rect 6290 2148 6294 2204
rect 6230 2144 6294 2148
rect 6310 2204 6374 2208
rect 6310 2148 6314 2204
rect 6314 2148 6370 2204
rect 6370 2148 6374 2204
rect 6310 2144 6374 2148
rect 6390 2204 6454 2208
rect 6390 2148 6394 2204
rect 6394 2148 6450 2204
rect 6450 2148 6454 2204
rect 6390 2144 6454 2148
rect 11348 2204 11412 2208
rect 11348 2148 11352 2204
rect 11352 2148 11408 2204
rect 11408 2148 11412 2204
rect 11348 2144 11412 2148
rect 11428 2204 11492 2208
rect 11428 2148 11432 2204
rect 11432 2148 11488 2204
rect 11488 2148 11492 2204
rect 11428 2144 11492 2148
rect 11508 2204 11572 2208
rect 11508 2148 11512 2204
rect 11512 2148 11568 2204
rect 11568 2148 11572 2204
rect 11508 2144 11572 2148
rect 11588 2204 11652 2208
rect 11588 2148 11592 2204
rect 11592 2148 11648 2204
rect 11648 2148 11652 2204
rect 11588 2144 11652 2148
rect 16546 2204 16610 2208
rect 16546 2148 16550 2204
rect 16550 2148 16606 2204
rect 16606 2148 16610 2204
rect 16546 2144 16610 2148
rect 16626 2204 16690 2208
rect 16626 2148 16630 2204
rect 16630 2148 16686 2204
rect 16686 2148 16690 2204
rect 16626 2144 16690 2148
rect 16706 2204 16770 2208
rect 16706 2148 16710 2204
rect 16710 2148 16766 2204
rect 16766 2148 16770 2204
rect 16706 2144 16770 2148
rect 16786 2204 16850 2208
rect 16786 2148 16790 2204
rect 16790 2148 16846 2204
rect 16846 2148 16850 2204
rect 16786 2144 16850 2148
rect 21744 2204 21808 2208
rect 21744 2148 21748 2204
rect 21748 2148 21804 2204
rect 21804 2148 21808 2204
rect 21744 2144 21808 2148
rect 21824 2204 21888 2208
rect 21824 2148 21828 2204
rect 21828 2148 21884 2204
rect 21884 2148 21888 2204
rect 21824 2144 21888 2148
rect 21904 2204 21968 2208
rect 21904 2148 21908 2204
rect 21908 2148 21964 2204
rect 21964 2148 21968 2204
rect 21904 2144 21968 2148
rect 21984 2204 22048 2208
rect 21984 2148 21988 2204
rect 21988 2148 22044 2204
rect 22044 2148 22048 2204
rect 21984 2144 22048 2148
<< metal4 >>
rect 3543 20160 3863 20720
rect 6142 20704 6462 20720
rect 6142 20640 6150 20704
rect 6214 20640 6230 20704
rect 6294 20640 6310 20704
rect 6374 20640 6390 20704
rect 6454 20640 6462 20704
rect 5027 20228 5093 20229
rect 5027 20164 5028 20228
rect 5092 20164 5093 20228
rect 5027 20163 5093 20164
rect 3543 20096 3551 20160
rect 3615 20096 3631 20160
rect 3695 20096 3711 20160
rect 3775 20096 3791 20160
rect 3855 20096 3863 20160
rect 3543 19072 3863 20096
rect 3923 19412 3989 19413
rect 3923 19348 3924 19412
rect 3988 19348 3989 19412
rect 3923 19347 3989 19348
rect 3543 19008 3551 19072
rect 3615 19008 3631 19072
rect 3695 19008 3711 19072
rect 3775 19008 3791 19072
rect 3855 19008 3863 19072
rect 3543 17984 3863 19008
rect 3543 17920 3551 17984
rect 3615 17920 3631 17984
rect 3695 17920 3711 17984
rect 3775 17920 3791 17984
rect 3855 17920 3863 17984
rect 3543 16896 3863 17920
rect 3543 16832 3551 16896
rect 3615 16832 3631 16896
rect 3695 16832 3711 16896
rect 3775 16832 3791 16896
rect 3855 16832 3863 16896
rect 3543 15808 3863 16832
rect 3543 15744 3551 15808
rect 3615 15744 3631 15808
rect 3695 15744 3711 15808
rect 3775 15744 3791 15808
rect 3855 15744 3863 15808
rect 3543 14720 3863 15744
rect 3543 14656 3551 14720
rect 3615 14656 3631 14720
rect 3695 14656 3711 14720
rect 3775 14656 3791 14720
rect 3855 14656 3863 14720
rect 3543 13632 3863 14656
rect 3543 13568 3551 13632
rect 3615 13568 3631 13632
rect 3695 13568 3711 13632
rect 3775 13568 3791 13632
rect 3855 13568 3863 13632
rect 3543 12544 3863 13568
rect 3543 12480 3551 12544
rect 3615 12480 3631 12544
rect 3695 12480 3711 12544
rect 3775 12480 3791 12544
rect 3855 12480 3863 12544
rect 3543 11456 3863 12480
rect 3543 11392 3551 11456
rect 3615 11392 3631 11456
rect 3695 11392 3711 11456
rect 3775 11392 3791 11456
rect 3855 11392 3863 11456
rect 3543 10368 3863 11392
rect 3926 10573 3986 19347
rect 4107 19140 4173 19141
rect 4107 19076 4108 19140
rect 4172 19076 4173 19140
rect 4107 19075 4173 19076
rect 3923 10572 3989 10573
rect 3923 10508 3924 10572
rect 3988 10508 3989 10572
rect 3923 10507 3989 10508
rect 3543 10304 3551 10368
rect 3615 10304 3631 10368
rect 3695 10304 3711 10368
rect 3775 10304 3791 10368
rect 3855 10304 3863 10368
rect 3543 9280 3863 10304
rect 3543 9216 3551 9280
rect 3615 9216 3631 9280
rect 3695 9216 3711 9280
rect 3775 9216 3791 9280
rect 3855 9216 3863 9280
rect 3543 8192 3863 9216
rect 3543 8128 3551 8192
rect 3615 8128 3631 8192
rect 3695 8128 3711 8192
rect 3775 8128 3791 8192
rect 3855 8128 3863 8192
rect 3543 7104 3863 8128
rect 3543 7040 3551 7104
rect 3615 7040 3631 7104
rect 3695 7040 3711 7104
rect 3775 7040 3791 7104
rect 3855 7040 3863 7104
rect 3543 6016 3863 7040
rect 3543 5952 3551 6016
rect 3615 5952 3631 6016
rect 3695 5952 3711 6016
rect 3775 5952 3791 6016
rect 3855 5952 3863 6016
rect 3543 4928 3863 5952
rect 3543 4864 3551 4928
rect 3615 4864 3631 4928
rect 3695 4864 3711 4928
rect 3775 4864 3791 4928
rect 3855 4864 3863 4928
rect 3543 3840 3863 4864
rect 3543 3776 3551 3840
rect 3615 3776 3631 3840
rect 3695 3776 3711 3840
rect 3775 3776 3791 3840
rect 3855 3776 3863 3840
rect 3543 2752 3863 3776
rect 4110 2957 4170 19075
rect 5030 18869 5090 20163
rect 5947 19956 6013 19957
rect 5947 19892 5948 19956
rect 6012 19892 6013 19956
rect 5947 19891 6013 19892
rect 5027 18868 5093 18869
rect 5027 18804 5028 18868
rect 5092 18804 5093 18868
rect 5027 18803 5093 18804
rect 5030 11797 5090 18803
rect 5027 11796 5093 11797
rect 5027 11732 5028 11796
rect 5092 11732 5093 11796
rect 5027 11731 5093 11732
rect 5950 3501 6010 19891
rect 6142 19616 6462 20640
rect 8741 20160 9061 20720
rect 8741 20096 8749 20160
rect 8813 20096 8829 20160
rect 8893 20096 8909 20160
rect 8973 20096 8989 20160
rect 9053 20096 9061 20160
rect 8155 20092 8221 20093
rect 8155 20028 8156 20092
rect 8220 20028 8221 20092
rect 8155 20027 8221 20028
rect 6142 19552 6150 19616
rect 6214 19552 6230 19616
rect 6294 19552 6310 19616
rect 6374 19552 6390 19616
rect 6454 19552 6462 19616
rect 6142 18528 6462 19552
rect 7971 19140 8037 19141
rect 7971 19076 7972 19140
rect 8036 19076 8037 19140
rect 7971 19075 8037 19076
rect 6142 18464 6150 18528
rect 6214 18464 6230 18528
rect 6294 18464 6310 18528
rect 6374 18464 6390 18528
rect 6454 18464 6462 18528
rect 6142 17440 6462 18464
rect 6142 17376 6150 17440
rect 6214 17376 6230 17440
rect 6294 17376 6310 17440
rect 6374 17376 6390 17440
rect 6454 17376 6462 17440
rect 6142 16352 6462 17376
rect 6142 16288 6150 16352
rect 6214 16288 6230 16352
rect 6294 16288 6310 16352
rect 6374 16288 6390 16352
rect 6454 16288 6462 16352
rect 6142 15264 6462 16288
rect 6142 15200 6150 15264
rect 6214 15200 6230 15264
rect 6294 15200 6310 15264
rect 6374 15200 6390 15264
rect 6454 15200 6462 15264
rect 6142 14176 6462 15200
rect 6142 14112 6150 14176
rect 6214 14112 6230 14176
rect 6294 14112 6310 14176
rect 6374 14112 6390 14176
rect 6454 14112 6462 14176
rect 6142 13088 6462 14112
rect 6142 13024 6150 13088
rect 6214 13024 6230 13088
rect 6294 13024 6310 13088
rect 6374 13024 6390 13088
rect 6454 13024 6462 13088
rect 6142 12000 6462 13024
rect 6142 11936 6150 12000
rect 6214 11936 6230 12000
rect 6294 11936 6310 12000
rect 6374 11936 6390 12000
rect 6454 11936 6462 12000
rect 6142 10912 6462 11936
rect 6142 10848 6150 10912
rect 6214 10848 6230 10912
rect 6294 10848 6310 10912
rect 6374 10848 6390 10912
rect 6454 10848 6462 10912
rect 6142 9824 6462 10848
rect 6142 9760 6150 9824
rect 6214 9760 6230 9824
rect 6294 9760 6310 9824
rect 6374 9760 6390 9824
rect 6454 9760 6462 9824
rect 6142 8736 6462 9760
rect 7974 8941 8034 19075
rect 7971 8940 8037 8941
rect 7971 8876 7972 8940
rect 8036 8876 8037 8940
rect 7971 8875 8037 8876
rect 6142 8672 6150 8736
rect 6214 8672 6230 8736
rect 6294 8672 6310 8736
rect 6374 8672 6390 8736
rect 6454 8672 6462 8736
rect 6142 7648 6462 8672
rect 8158 7989 8218 20027
rect 8339 19548 8405 19549
rect 8339 19484 8340 19548
rect 8404 19484 8405 19548
rect 8339 19483 8405 19484
rect 8342 9757 8402 19483
rect 8741 19072 9061 20096
rect 8741 19008 8749 19072
rect 8813 19008 8829 19072
rect 8893 19008 8909 19072
rect 8973 19008 8989 19072
rect 9053 19008 9061 19072
rect 8523 18052 8589 18053
rect 8523 17988 8524 18052
rect 8588 17988 8589 18052
rect 8523 17987 8589 17988
rect 8526 13293 8586 17987
rect 8741 17984 9061 19008
rect 8741 17920 8749 17984
rect 8813 17920 8829 17984
rect 8893 17920 8909 17984
rect 8973 17920 8989 17984
rect 9053 17920 9061 17984
rect 8741 16896 9061 17920
rect 8741 16832 8749 16896
rect 8813 16832 8829 16896
rect 8893 16832 8909 16896
rect 8973 16832 8989 16896
rect 9053 16832 9061 16896
rect 8741 15808 9061 16832
rect 8741 15744 8749 15808
rect 8813 15744 8829 15808
rect 8893 15744 8909 15808
rect 8973 15744 8989 15808
rect 9053 15744 9061 15808
rect 8741 14720 9061 15744
rect 8741 14656 8749 14720
rect 8813 14656 8829 14720
rect 8893 14656 8909 14720
rect 8973 14656 8989 14720
rect 9053 14656 9061 14720
rect 8741 13632 9061 14656
rect 8741 13568 8749 13632
rect 8813 13568 8829 13632
rect 8893 13568 8909 13632
rect 8973 13568 8989 13632
rect 9053 13568 9061 13632
rect 8523 13292 8589 13293
rect 8523 13228 8524 13292
rect 8588 13228 8589 13292
rect 8523 13227 8589 13228
rect 8526 12341 8586 13227
rect 8741 12544 9061 13568
rect 8741 12480 8749 12544
rect 8813 12480 8829 12544
rect 8893 12480 8909 12544
rect 8973 12480 8989 12544
rect 9053 12480 9061 12544
rect 8523 12340 8589 12341
rect 8523 12276 8524 12340
rect 8588 12276 8589 12340
rect 8523 12275 8589 12276
rect 8741 11456 9061 12480
rect 8741 11392 8749 11456
rect 8813 11392 8829 11456
rect 8893 11392 8909 11456
rect 8973 11392 8989 11456
rect 9053 11392 9061 11456
rect 8741 10368 9061 11392
rect 8741 10304 8749 10368
rect 8813 10304 8829 10368
rect 8893 10304 8909 10368
rect 8973 10304 8989 10368
rect 9053 10304 9061 10368
rect 8339 9756 8405 9757
rect 8339 9692 8340 9756
rect 8404 9692 8405 9756
rect 8339 9691 8405 9692
rect 8741 9280 9061 10304
rect 8741 9216 8749 9280
rect 8813 9216 8829 9280
rect 8893 9216 8909 9280
rect 8973 9216 8989 9280
rect 9053 9216 9061 9280
rect 8741 8192 9061 9216
rect 8741 8128 8749 8192
rect 8813 8128 8829 8192
rect 8893 8128 8909 8192
rect 8973 8128 8989 8192
rect 9053 8128 9061 8192
rect 8155 7988 8221 7989
rect 8155 7924 8156 7988
rect 8220 7924 8221 7988
rect 8155 7923 8221 7924
rect 6142 7584 6150 7648
rect 6214 7584 6230 7648
rect 6294 7584 6310 7648
rect 6374 7584 6390 7648
rect 6454 7584 6462 7648
rect 6142 6560 6462 7584
rect 6142 6496 6150 6560
rect 6214 6496 6230 6560
rect 6294 6496 6310 6560
rect 6374 6496 6390 6560
rect 6454 6496 6462 6560
rect 6142 5472 6462 6496
rect 6142 5408 6150 5472
rect 6214 5408 6230 5472
rect 6294 5408 6310 5472
rect 6374 5408 6390 5472
rect 6454 5408 6462 5472
rect 6142 4384 6462 5408
rect 6142 4320 6150 4384
rect 6214 4320 6230 4384
rect 6294 4320 6310 4384
rect 6374 4320 6390 4384
rect 6454 4320 6462 4384
rect 5947 3500 6013 3501
rect 5947 3436 5948 3500
rect 6012 3436 6013 3500
rect 5947 3435 6013 3436
rect 6142 3296 6462 4320
rect 6142 3232 6150 3296
rect 6214 3232 6230 3296
rect 6294 3232 6310 3296
rect 6374 3232 6390 3296
rect 6454 3232 6462 3296
rect 4107 2956 4173 2957
rect 4107 2892 4108 2956
rect 4172 2892 4173 2956
rect 4107 2891 4173 2892
rect 3543 2688 3551 2752
rect 3615 2688 3631 2752
rect 3695 2688 3711 2752
rect 3775 2688 3791 2752
rect 3855 2688 3863 2752
rect 3543 2128 3863 2688
rect 6142 2208 6462 3232
rect 6142 2144 6150 2208
rect 6214 2144 6230 2208
rect 6294 2144 6310 2208
rect 6374 2144 6390 2208
rect 6454 2144 6462 2208
rect 6142 2128 6462 2144
rect 8741 7104 9061 8128
rect 8741 7040 8749 7104
rect 8813 7040 8829 7104
rect 8893 7040 8909 7104
rect 8973 7040 8989 7104
rect 9053 7040 9061 7104
rect 8741 6016 9061 7040
rect 8741 5952 8749 6016
rect 8813 5952 8829 6016
rect 8893 5952 8909 6016
rect 8973 5952 8989 6016
rect 9053 5952 9061 6016
rect 8741 4928 9061 5952
rect 8741 4864 8749 4928
rect 8813 4864 8829 4928
rect 8893 4864 8909 4928
rect 8973 4864 8989 4928
rect 9053 4864 9061 4928
rect 8741 3840 9061 4864
rect 8741 3776 8749 3840
rect 8813 3776 8829 3840
rect 8893 3776 8909 3840
rect 8973 3776 8989 3840
rect 9053 3776 9061 3840
rect 8741 2752 9061 3776
rect 8741 2688 8749 2752
rect 8813 2688 8829 2752
rect 8893 2688 8909 2752
rect 8973 2688 8989 2752
rect 9053 2688 9061 2752
rect 8741 2128 9061 2688
rect 11340 20704 11660 20720
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 19616 11660 20640
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 18528 11660 19552
rect 13939 20160 14259 20720
rect 13939 20096 13947 20160
rect 14011 20096 14027 20160
rect 14091 20096 14107 20160
rect 14171 20096 14187 20160
rect 14251 20096 14259 20160
rect 11835 19412 11901 19413
rect 11835 19348 11836 19412
rect 11900 19348 11901 19412
rect 11835 19347 11901 19348
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 17440 11660 18464
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 16352 11660 17376
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 15264 11660 16288
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 14176 11660 15200
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 13088 11660 14112
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 12000 11660 13024
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 10912 11660 11936
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 9824 11660 10848
rect 11838 10165 11898 19347
rect 13939 19072 14259 20096
rect 13939 19008 13947 19072
rect 14011 19008 14027 19072
rect 14091 19008 14107 19072
rect 14171 19008 14187 19072
rect 14251 19008 14259 19072
rect 13939 17984 14259 19008
rect 13939 17920 13947 17984
rect 14011 17920 14027 17984
rect 14091 17920 14107 17984
rect 14171 17920 14187 17984
rect 14251 17920 14259 17984
rect 13939 16896 14259 17920
rect 13939 16832 13947 16896
rect 14011 16832 14027 16896
rect 14091 16832 14107 16896
rect 14171 16832 14187 16896
rect 14251 16832 14259 16896
rect 13939 15808 14259 16832
rect 13939 15744 13947 15808
rect 14011 15744 14027 15808
rect 14091 15744 14107 15808
rect 14171 15744 14187 15808
rect 14251 15744 14259 15808
rect 13939 14720 14259 15744
rect 13939 14656 13947 14720
rect 14011 14656 14027 14720
rect 14091 14656 14107 14720
rect 14171 14656 14187 14720
rect 14251 14656 14259 14720
rect 13939 13632 14259 14656
rect 13939 13568 13947 13632
rect 14011 13568 14027 13632
rect 14091 13568 14107 13632
rect 14171 13568 14187 13632
rect 14251 13568 14259 13632
rect 13939 12544 14259 13568
rect 13939 12480 13947 12544
rect 14011 12480 14027 12544
rect 14091 12480 14107 12544
rect 14171 12480 14187 12544
rect 14251 12480 14259 12544
rect 13939 11456 14259 12480
rect 13939 11392 13947 11456
rect 14011 11392 14027 11456
rect 14091 11392 14107 11456
rect 14171 11392 14187 11456
rect 14251 11392 14259 11456
rect 13939 10368 14259 11392
rect 13939 10304 13947 10368
rect 14011 10304 14027 10368
rect 14091 10304 14107 10368
rect 14171 10304 14187 10368
rect 14251 10304 14259 10368
rect 11835 10164 11901 10165
rect 11835 10100 11836 10164
rect 11900 10100 11901 10164
rect 11835 10099 11901 10100
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 8736 11660 9760
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 7648 11660 8672
rect 11838 7853 11898 10099
rect 13939 9280 14259 10304
rect 13939 9216 13947 9280
rect 14011 9216 14027 9280
rect 14091 9216 14107 9280
rect 14171 9216 14187 9280
rect 14251 9216 14259 9280
rect 13939 8192 14259 9216
rect 13939 8128 13947 8192
rect 14011 8128 14027 8192
rect 14091 8128 14107 8192
rect 14171 8128 14187 8192
rect 14251 8128 14259 8192
rect 11835 7852 11901 7853
rect 11835 7788 11836 7852
rect 11900 7788 11901 7852
rect 11835 7787 11901 7788
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 6560 11660 7584
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 5472 11660 6496
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 4384 11660 5408
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 3296 11660 4320
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 2208 11660 3232
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2128 11660 2144
rect 13939 7104 14259 8128
rect 13939 7040 13947 7104
rect 14011 7040 14027 7104
rect 14091 7040 14107 7104
rect 14171 7040 14187 7104
rect 14251 7040 14259 7104
rect 13939 6016 14259 7040
rect 13939 5952 13947 6016
rect 14011 5952 14027 6016
rect 14091 5952 14107 6016
rect 14171 5952 14187 6016
rect 14251 5952 14259 6016
rect 13939 4928 14259 5952
rect 13939 4864 13947 4928
rect 14011 4864 14027 4928
rect 14091 4864 14107 4928
rect 14171 4864 14187 4928
rect 14251 4864 14259 4928
rect 13939 3840 14259 4864
rect 13939 3776 13947 3840
rect 14011 3776 14027 3840
rect 14091 3776 14107 3840
rect 14171 3776 14187 3840
rect 14251 3776 14259 3840
rect 13939 2752 14259 3776
rect 13939 2688 13947 2752
rect 14011 2688 14027 2752
rect 14091 2688 14107 2752
rect 14171 2688 14187 2752
rect 14251 2688 14259 2752
rect 13939 2128 14259 2688
rect 16538 20704 16858 20720
rect 16538 20640 16546 20704
rect 16610 20640 16626 20704
rect 16690 20640 16706 20704
rect 16770 20640 16786 20704
rect 16850 20640 16858 20704
rect 16538 19616 16858 20640
rect 16538 19552 16546 19616
rect 16610 19552 16626 19616
rect 16690 19552 16706 19616
rect 16770 19552 16786 19616
rect 16850 19552 16858 19616
rect 16538 18528 16858 19552
rect 16538 18464 16546 18528
rect 16610 18464 16626 18528
rect 16690 18464 16706 18528
rect 16770 18464 16786 18528
rect 16850 18464 16858 18528
rect 16538 17440 16858 18464
rect 16538 17376 16546 17440
rect 16610 17376 16626 17440
rect 16690 17376 16706 17440
rect 16770 17376 16786 17440
rect 16850 17376 16858 17440
rect 16538 16352 16858 17376
rect 16538 16288 16546 16352
rect 16610 16288 16626 16352
rect 16690 16288 16706 16352
rect 16770 16288 16786 16352
rect 16850 16288 16858 16352
rect 16538 15264 16858 16288
rect 16538 15200 16546 15264
rect 16610 15200 16626 15264
rect 16690 15200 16706 15264
rect 16770 15200 16786 15264
rect 16850 15200 16858 15264
rect 16538 14176 16858 15200
rect 16538 14112 16546 14176
rect 16610 14112 16626 14176
rect 16690 14112 16706 14176
rect 16770 14112 16786 14176
rect 16850 14112 16858 14176
rect 16538 13088 16858 14112
rect 16538 13024 16546 13088
rect 16610 13024 16626 13088
rect 16690 13024 16706 13088
rect 16770 13024 16786 13088
rect 16850 13024 16858 13088
rect 16538 12000 16858 13024
rect 16538 11936 16546 12000
rect 16610 11936 16626 12000
rect 16690 11936 16706 12000
rect 16770 11936 16786 12000
rect 16850 11936 16858 12000
rect 16538 10912 16858 11936
rect 16538 10848 16546 10912
rect 16610 10848 16626 10912
rect 16690 10848 16706 10912
rect 16770 10848 16786 10912
rect 16850 10848 16858 10912
rect 16538 9824 16858 10848
rect 16538 9760 16546 9824
rect 16610 9760 16626 9824
rect 16690 9760 16706 9824
rect 16770 9760 16786 9824
rect 16850 9760 16858 9824
rect 16538 8736 16858 9760
rect 16538 8672 16546 8736
rect 16610 8672 16626 8736
rect 16690 8672 16706 8736
rect 16770 8672 16786 8736
rect 16850 8672 16858 8736
rect 16538 7648 16858 8672
rect 16538 7584 16546 7648
rect 16610 7584 16626 7648
rect 16690 7584 16706 7648
rect 16770 7584 16786 7648
rect 16850 7584 16858 7648
rect 16538 6560 16858 7584
rect 16538 6496 16546 6560
rect 16610 6496 16626 6560
rect 16690 6496 16706 6560
rect 16770 6496 16786 6560
rect 16850 6496 16858 6560
rect 16538 5472 16858 6496
rect 16538 5408 16546 5472
rect 16610 5408 16626 5472
rect 16690 5408 16706 5472
rect 16770 5408 16786 5472
rect 16850 5408 16858 5472
rect 16538 4384 16858 5408
rect 16538 4320 16546 4384
rect 16610 4320 16626 4384
rect 16690 4320 16706 4384
rect 16770 4320 16786 4384
rect 16850 4320 16858 4384
rect 16538 3296 16858 4320
rect 16538 3232 16546 3296
rect 16610 3232 16626 3296
rect 16690 3232 16706 3296
rect 16770 3232 16786 3296
rect 16850 3232 16858 3296
rect 16538 2208 16858 3232
rect 16538 2144 16546 2208
rect 16610 2144 16626 2208
rect 16690 2144 16706 2208
rect 16770 2144 16786 2208
rect 16850 2144 16858 2208
rect 16538 2128 16858 2144
rect 19137 20160 19457 20720
rect 19137 20096 19145 20160
rect 19209 20096 19225 20160
rect 19289 20096 19305 20160
rect 19369 20096 19385 20160
rect 19449 20096 19457 20160
rect 19137 19072 19457 20096
rect 19137 19008 19145 19072
rect 19209 19008 19225 19072
rect 19289 19008 19305 19072
rect 19369 19008 19385 19072
rect 19449 19008 19457 19072
rect 19137 17984 19457 19008
rect 21736 20704 22056 20720
rect 21736 20640 21744 20704
rect 21808 20640 21824 20704
rect 21888 20640 21904 20704
rect 21968 20640 21984 20704
rect 22048 20640 22056 20704
rect 21736 19616 22056 20640
rect 21736 19552 21744 19616
rect 21808 19552 21824 19616
rect 21888 19552 21904 19616
rect 21968 19552 21984 19616
rect 22048 19552 22056 19616
rect 20483 18732 20549 18733
rect 20483 18668 20484 18732
rect 20548 18668 20549 18732
rect 20483 18667 20549 18668
rect 19137 17920 19145 17984
rect 19209 17920 19225 17984
rect 19289 17920 19305 17984
rect 19369 17920 19385 17984
rect 19449 17920 19457 17984
rect 19137 16896 19457 17920
rect 19137 16832 19145 16896
rect 19209 16832 19225 16896
rect 19289 16832 19305 16896
rect 19369 16832 19385 16896
rect 19449 16832 19457 16896
rect 19137 15808 19457 16832
rect 19137 15744 19145 15808
rect 19209 15744 19225 15808
rect 19289 15744 19305 15808
rect 19369 15744 19385 15808
rect 19449 15744 19457 15808
rect 19137 14720 19457 15744
rect 19137 14656 19145 14720
rect 19209 14656 19225 14720
rect 19289 14656 19305 14720
rect 19369 14656 19385 14720
rect 19449 14656 19457 14720
rect 19137 13632 19457 14656
rect 19137 13568 19145 13632
rect 19209 13568 19225 13632
rect 19289 13568 19305 13632
rect 19369 13568 19385 13632
rect 19449 13568 19457 13632
rect 19137 12544 19457 13568
rect 19137 12480 19145 12544
rect 19209 12480 19225 12544
rect 19289 12480 19305 12544
rect 19369 12480 19385 12544
rect 19449 12480 19457 12544
rect 19137 11456 19457 12480
rect 19137 11392 19145 11456
rect 19209 11392 19225 11456
rect 19289 11392 19305 11456
rect 19369 11392 19385 11456
rect 19449 11392 19457 11456
rect 19137 10368 19457 11392
rect 19137 10304 19145 10368
rect 19209 10304 19225 10368
rect 19289 10304 19305 10368
rect 19369 10304 19385 10368
rect 19449 10304 19457 10368
rect 19137 9280 19457 10304
rect 20486 9485 20546 18667
rect 21736 18528 22056 19552
rect 21736 18464 21744 18528
rect 21808 18464 21824 18528
rect 21888 18464 21904 18528
rect 21968 18464 21984 18528
rect 22048 18464 22056 18528
rect 21736 17440 22056 18464
rect 21736 17376 21744 17440
rect 21808 17376 21824 17440
rect 21888 17376 21904 17440
rect 21968 17376 21984 17440
rect 22048 17376 22056 17440
rect 21736 16352 22056 17376
rect 21736 16288 21744 16352
rect 21808 16288 21824 16352
rect 21888 16288 21904 16352
rect 21968 16288 21984 16352
rect 22048 16288 22056 16352
rect 21736 15264 22056 16288
rect 21736 15200 21744 15264
rect 21808 15200 21824 15264
rect 21888 15200 21904 15264
rect 21968 15200 21984 15264
rect 22048 15200 22056 15264
rect 21736 14176 22056 15200
rect 21736 14112 21744 14176
rect 21808 14112 21824 14176
rect 21888 14112 21904 14176
rect 21968 14112 21984 14176
rect 22048 14112 22056 14176
rect 21736 13088 22056 14112
rect 21736 13024 21744 13088
rect 21808 13024 21824 13088
rect 21888 13024 21904 13088
rect 21968 13024 21984 13088
rect 22048 13024 22056 13088
rect 21736 12000 22056 13024
rect 21736 11936 21744 12000
rect 21808 11936 21824 12000
rect 21888 11936 21904 12000
rect 21968 11936 21984 12000
rect 22048 11936 22056 12000
rect 21736 10912 22056 11936
rect 21736 10848 21744 10912
rect 21808 10848 21824 10912
rect 21888 10848 21904 10912
rect 21968 10848 21984 10912
rect 22048 10848 22056 10912
rect 21736 9824 22056 10848
rect 21736 9760 21744 9824
rect 21808 9760 21824 9824
rect 21888 9760 21904 9824
rect 21968 9760 21984 9824
rect 22048 9760 22056 9824
rect 20483 9484 20549 9485
rect 20483 9420 20484 9484
rect 20548 9420 20549 9484
rect 20483 9419 20549 9420
rect 19137 9216 19145 9280
rect 19209 9216 19225 9280
rect 19289 9216 19305 9280
rect 19369 9216 19385 9280
rect 19449 9216 19457 9280
rect 19137 8192 19457 9216
rect 19137 8128 19145 8192
rect 19209 8128 19225 8192
rect 19289 8128 19305 8192
rect 19369 8128 19385 8192
rect 19449 8128 19457 8192
rect 19137 7104 19457 8128
rect 19137 7040 19145 7104
rect 19209 7040 19225 7104
rect 19289 7040 19305 7104
rect 19369 7040 19385 7104
rect 19449 7040 19457 7104
rect 19137 6016 19457 7040
rect 19137 5952 19145 6016
rect 19209 5952 19225 6016
rect 19289 5952 19305 6016
rect 19369 5952 19385 6016
rect 19449 5952 19457 6016
rect 19137 4928 19457 5952
rect 19137 4864 19145 4928
rect 19209 4864 19225 4928
rect 19289 4864 19305 4928
rect 19369 4864 19385 4928
rect 19449 4864 19457 4928
rect 19137 3840 19457 4864
rect 19137 3776 19145 3840
rect 19209 3776 19225 3840
rect 19289 3776 19305 3840
rect 19369 3776 19385 3840
rect 19449 3776 19457 3840
rect 19137 2752 19457 3776
rect 19137 2688 19145 2752
rect 19209 2688 19225 2752
rect 19289 2688 19305 2752
rect 19369 2688 19385 2752
rect 19449 2688 19457 2752
rect 19137 2128 19457 2688
rect 21736 8736 22056 9760
rect 21736 8672 21744 8736
rect 21808 8672 21824 8736
rect 21888 8672 21904 8736
rect 21968 8672 21984 8736
rect 22048 8672 22056 8736
rect 21736 7648 22056 8672
rect 21736 7584 21744 7648
rect 21808 7584 21824 7648
rect 21888 7584 21904 7648
rect 21968 7584 21984 7648
rect 22048 7584 22056 7648
rect 21736 6560 22056 7584
rect 21736 6496 21744 6560
rect 21808 6496 21824 6560
rect 21888 6496 21904 6560
rect 21968 6496 21984 6560
rect 22048 6496 22056 6560
rect 21736 5472 22056 6496
rect 21736 5408 21744 5472
rect 21808 5408 21824 5472
rect 21888 5408 21904 5472
rect 21968 5408 21984 5472
rect 22048 5408 22056 5472
rect 21736 4384 22056 5408
rect 21736 4320 21744 4384
rect 21808 4320 21824 4384
rect 21888 4320 21904 4384
rect 21968 4320 21984 4384
rect 22048 4320 22056 4384
rect 21736 3296 22056 4320
rect 21736 3232 21744 3296
rect 21808 3232 21824 3296
rect 21888 3232 21904 3296
rect 21968 3232 21984 3296
rect 22048 3232 22056 3296
rect 21736 2208 22056 3232
rect 21736 2144 21744 2208
rect 21808 2144 21824 2208
rect 21888 2144 21904 2208
rect 21968 2144 21984 2208
rect 22048 2144 22056 2208
rect 21736 2128 22056 2144
use sky130_fd_sc_hd__diode_2  ANTENNA__060__A dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2944 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__062__A
timestamp 1649977179
transform 1 0 3772 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__063__A
timestamp 1649977179
transform -1 0 3128 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__064__A
timestamp 1649977179
transform 1 0 2668 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__066__A
timestamp 1649977179
transform 1 0 2116 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__067__A
timestamp 1649977179
transform -1 0 2944 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__068__A
timestamp 1649977179
transform -1 0 2576 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__A
timestamp 1649977179
transform 1 0 2392 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__071__A
timestamp 1649977179
transform -1 0 1932 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__072__A
timestamp 1649977179
transform 1 0 2760 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__A
timestamp 1649977179
transform 1 0 3220 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__A
timestamp 1649977179
transform 1 0 3956 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__076__A
timestamp 1649977179
transform 1 0 2944 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__080__A
timestamp 1649977179
transform 1 0 20240 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__082__A
timestamp 1649977179
transform -1 0 20792 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__083__A
timestamp 1649977179
transform -1 0 21252 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__084__A
timestamp 1649977179
transform -1 0 20240 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__A
timestamp 1649977179
transform -1 0 20792 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__087__A
timestamp 1649977179
transform -1 0 20424 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__088__A
timestamp 1649977179
transform 1 0 20148 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__A
timestamp 1649977179
transform -1 0 20148 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__A
timestamp 1649977179
transform -1 0 20332 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__A
timestamp 1649977179
transform 1 0 19320 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__094__A
timestamp 1649977179
transform 1 0 19136 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__A
timestamp 1649977179
transform -1 0 19136 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__096__A
timestamp 1649977179
transform 1 0 19504 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__110__A
timestamp 1649977179
transform -1 0 19136 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1649977179
transform -1 0 3956 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1649977179
transform -1 0 20700 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1649977179
transform -1 0 2760 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1649977179
transform -1 0 3036 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1649977179
transform -1 0 2760 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1649977179
transform -1 0 2576 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1649977179
transform -1 0 2484 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1649977179
transform -1 0 2760 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1649977179
transform -1 0 3036 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1649977179
transform -1 0 2576 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1649977179
transform -1 0 2576 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1649977179
transform -1 0 2760 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1649977179
transform -1 0 2300 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1649977179
transform -1 0 1840 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1649977179
transform -1 0 2852 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1649977179
transform -1 0 2668 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1649977179
transform -1 0 3956 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1649977179
transform -1 0 2760 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1649977179
transform -1 0 3956 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1649977179
transform -1 0 4140 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1649977179
transform -1 0 3772 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1649977179
transform -1 0 3404 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1649977179
transform -1 0 1564 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1649977179
transform -1 0 21068 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1649977179
transform -1 0 18308 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1649977179
transform -1 0 20608 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1649977179
transform -1 0 20792 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1649977179
transform -1 0 21160 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1649977179
transform -1 0 20976 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1649977179
transform -1 0 21344 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1649977179
transform -1 0 21068 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1649977179
transform -1 0 20884 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1649977179
transform -1 0 21252 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1649977179
transform -1 0 21252 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1649977179
transform -1 0 20884 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1649977179
transform -1 0 20700 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1649977179
transform -1 0 20608 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1649977179
transform -1 0 20240 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1649977179
transform -1 0 20424 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1649977179
transform -1 0 20240 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1649977179
transform -1 0 18860 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1649977179
transform -1 0 20608 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1649977179
transform -1 0 21620 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1649977179
transform -1 0 8188 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1649977179
transform -1 0 11316 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1649977179
transform -1 0 10580 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1649977179
transform -1 0 6900 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1649977179
transform -1 0 11684 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1649977179
transform -1 0 11684 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1649977179
transform -1 0 13156 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1649977179
transform -1 0 12788 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1649977179
transform -1 0 12972 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1649977179
transform -1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1649977179
transform -1 0 15732 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1649977179
transform -1 0 5612 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1649977179
transform -1 0 3680 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1649977179
transform -1 0 3956 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1649977179
transform -1 0 7820 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1649977179
transform -1 0 8004 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1649977179
transform -1 0 9292 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1649977179
transform -1 0 9108 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1649977179
transform -1 0 8648 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 1649977179
transform -1 0 9476 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 1649977179
transform -1 0 16100 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 1649977179
transform -1 0 2208 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 1649977179
transform -1 0 2392 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 1649977179
transform -1 0 1840 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input68_A
timestamp 1649977179
transform -1 0 2024 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 1649977179
transform -1 0 2392 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input70_A
timestamp 1649977179
transform -1 0 2944 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input71_A
timestamp 1649977179
transform -1 0 2024 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input72_A
timestamp 1649977179
transform -1 0 2576 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input73_A
timestamp 1649977179
transform -1 0 1840 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input74_A
timestamp 1649977179
transform -1 0 11960 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input75_A
timestamp 1649977179
transform -1 0 21068 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input76_A
timestamp 1649977179
transform -1 0 20700 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input77_A
timestamp 1649977179
transform -1 0 20884 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input78_A
timestamp 1649977179
transform -1 0 21344 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input79_A
timestamp 1649977179
transform -1 0 20332 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input80_A
timestamp 1649977179
transform -1 0 20516 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input81_A
timestamp 1649977179
transform -1 0 21068 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input82_A
timestamp 1649977179
transform -1 0 20884 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input83_A
timestamp 1649977179
transform -1 0 21344 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input84_A
timestamp 1649977179
transform -1 0 2944 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input85_A
timestamp 1649977179
transform -1 0 2760 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input86_A
timestamp 1649977179
transform -1 0 4140 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input87_A
timestamp 1649977179
transform -1 0 3588 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input88_A
timestamp 1649977179
transform -1 0 3772 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input89_A
timestamp 1649977179
transform -1 0 3956 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input90_A
timestamp 1649977179
transform -1 0 4692 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input91_A
timestamp 1649977179
transform -1 0 5060 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 14444 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 5336 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 6532 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 8004 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 7176 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 7084 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 5520 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 7820 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 5704 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 6072 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 5428 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 5244 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 6440 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 5520 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 6256 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 6440 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 6532 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 5796 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 11684 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 15916 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 15548 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13432 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11500 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 12144 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 14076 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 14260 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 8556 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 9660 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 10672 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13984 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 8280 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 13616 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13708 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11684 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13616 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 12512 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 13984 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 5980 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 7820 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 8740 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 8924 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 11684 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11132 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 9108 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 10396 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11132 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 9568 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 13340 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11316 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 15364 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 14168 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 8096 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 9200 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 7176 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 5796 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 4416 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 6348 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 8188 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 9016 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 11684 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13156 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 8188 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 10948 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 8832 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_38.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 10396 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_38.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11868 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 5152 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 4784 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 10304 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A1
timestamp 1649977179
transform -1 0 5888 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 5060 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 5428 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 4968 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 3956 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 8188 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 4600 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 7728 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 3680 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 7912 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 8648 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 17756 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 17848 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 16468 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 18768 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 17020 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_6__A0
timestamp 1649977179
transform -1 0 20332 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_6__A1
timestamp 1649977179
transform 1 0 20148 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A0
timestamp 1649977179
transform -1 0 16284 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 18860 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 20424 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 18676 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 18584 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 18032 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 16192 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 17296 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A1
timestamp 1649977179
transform -1 0 10396 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 9752 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 8188 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 11776 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 16008 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_3__A1
timestamp 1649977179
transform -1 0 14168 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 12236 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 18676 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 16744 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 10948 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 18400 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_3__A1
timestamp 1649977179
transform -1 0 16192 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 10856 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 15916 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 18860 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 17940 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 12512 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 9936 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 5336 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 5152 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 1748 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 7636 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 7452 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 18400 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 16560 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 17664 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 16008 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 8648 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 11316 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 10488 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output93_A
timestamp 1649977179
transform -1 0 4232 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output143_A
timestamp 1649977179
transform -1 0 21620 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output144_A
timestamp 1649977179
transform 1 0 18952 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output155_A
timestamp 1649977179
transform -1 0 5796 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1649977179
transform -1 0 4416 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2944 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1649977179
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6348 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67
timestamp 1649977179
transform 1 0 7268 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_79 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 8372 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1649977179
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1649977179
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118
timestamp 1649977179
transform 1 0 11960 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_130
timestamp 1649977179
transform 1 0 13064 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_153
timestamp 1649977179
transform 1 0 15180 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1649977179
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1649977179
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1649977179
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1649977179
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_197
timestamp 1649977179
transform 1 0 19228 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_205
timestamp 1649977179
transform 1 0 19964 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_216
timestamp 1649977179
transform 1 0 20976 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_16
timestamp 1649977179
transform 1 0 2576 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_28
timestamp 1649977179
transform 1 0 3680 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_40
timestamp 1649977179
transform 1 0 4784 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_52
timestamp 1649977179
transform 1 0 5888 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1649977179
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1649977179
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_81
timestamp 1649977179
transform 1 0 8556 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_88
timestamp 1649977179
transform 1 0 9200 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_100
timestamp 1649977179
transform 1 0 10304 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1649977179
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1649977179
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1649977179
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1649977179
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1649977179
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1649977179
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_175
timestamp 1649977179
transform 1 0 17204 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_187
timestamp 1649977179
transform 1 0 18308 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_199
timestamp 1649977179
transform 1 0 19412 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_211
timestamp 1649977179
transform 1 0 20516 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_10
timestamp 1649977179
transform 1 0 2024 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_22
timestamp 1649977179
transform 1 0 3128 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1649977179
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1649977179
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1649977179
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1649977179
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1649977179
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1649977179
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1649977179
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1649977179
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1649977179
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1649977179
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1649977179
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1649977179
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1649977179
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1649977179
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1649977179
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1649977179
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_209
timestamp 1649977179
transform 1 0 20332 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_217
timestamp 1649977179
transform 1 0 21068 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_12
timestamp 1649977179
transform 1 0 2208 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_24
timestamp 1649977179
transform 1 0 3312 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_36
timestamp 1649977179
transform 1 0 4416 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_48
timestamp 1649977179
transform 1 0 5520 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1649977179
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1649977179
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1649977179
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1649977179
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1649977179
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1649977179
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1649977179
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1649977179
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1649977179
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1649977179
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1649977179
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1649977179
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1649977179
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_205
timestamp 1649977179
transform 1 0 19964 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_14
timestamp 1649977179
transform 1 0 2392 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_26
timestamp 1649977179
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1649977179
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1649977179
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1649977179
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1649977179
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1649977179
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1649977179
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1649977179
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1649977179
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1649977179
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1649977179
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1649977179
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1649977179
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1649977179
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1649977179
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1649977179
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1649977179
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_209
timestamp 1649977179
transform 1 0 20332 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_21
timestamp 1649977179
transform 1 0 3036 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_33
timestamp 1649977179
transform 1 0 4140 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_45
timestamp 1649977179
transform 1 0 5244 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_53
timestamp 1649977179
transform 1 0 5980 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1649977179
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1649977179
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1649977179
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1649977179
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1649977179
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1649977179
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1649977179
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1649977179
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1649977179
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1649977179
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1649977179
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1649977179
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1649977179
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1649977179
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_217
timestamp 1649977179
transform 1 0 21068 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_6
timestamp 1649977179
transform 1 0 1656 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_25
timestamp 1649977179
transform 1 0 3404 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_29
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_37
timestamp 1649977179
transform 1 0 4508 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_47
timestamp 1649977179
transform 1 0 5428 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_59
timestamp 1649977179
transform 1 0 6532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_71
timestamp 1649977179
transform 1 0 7636 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1649977179
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1649977179
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1649977179
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1649977179
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1649977179
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1649977179
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_141
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_145
timestamp 1649977179
transform 1 0 14444 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_149
timestamp 1649977179
transform 1 0 14812 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_161
timestamp 1649977179
transform 1 0 15916 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_173
timestamp 1649977179
transform 1 0 17020 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_185
timestamp 1649977179
transform 1 0 18124 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_193
timestamp 1649977179
transform 1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1649977179
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_209
timestamp 1649977179
transform 1 0 20332 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_36
timestamp 1649977179
transform 1 0 4416 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_40
timestamp 1649977179
transform 1 0 4784 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_52
timestamp 1649977179
transform 1 0 5888 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1649977179
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1649977179
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1649977179
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1649977179
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1649977179
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_113
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_124
timestamp 1649977179
transform 1 0 12512 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_135
timestamp 1649977179
transform 1 0 13524 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_139
timestamp 1649977179
transform 1 0 13892 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_162
timestamp 1649977179
transform 1 0 16008 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1649977179
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1649977179
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1649977179
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_205
timestamp 1649977179
transform 1 0 19964 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_33
timestamp 1649977179
transform 1 0 4140 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_64
timestamp 1649977179
transform 1 0 6992 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_76
timestamp 1649977179
transform 1 0 8096 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_96
timestamp 1649977179
transform 1 0 9936 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_102
timestamp 1649977179
transform 1 0 10488 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_114
timestamp 1649977179
transform 1 0 11592 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_122
timestamp 1649977179
transform 1 0 12328 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_135
timestamp 1649977179
transform 1 0 13524 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1649977179
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1649977179
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1649977179
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1649977179
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1649977179
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1649977179
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_197
timestamp 1649977179
transform 1 0 19228 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_205
timestamp 1649977179
transform 1 0 19964 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_13
timestamp 1649977179
transform 1 0 2300 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_31
timestamp 1649977179
transform 1 0 3956 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1649977179
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_69
timestamp 1649977179
transform 1 0 7452 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1649977179
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1649977179
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1649977179
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1649977179
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1649977179
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1649977179
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_169
timestamp 1649977179
transform 1 0 16652 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_180
timestamp 1649977179
transform 1 0 17664 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_183
timestamp 1649977179
transform 1 0 17940 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_194
timestamp 1649977179
transform 1 0 18952 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_5
timestamp 1649977179
transform 1 0 1564 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_31
timestamp 1649977179
transform 1 0 3956 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_46
timestamp 1649977179
transform 1 0 5336 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_65
timestamp 1649977179
transform 1 0 7084 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_94
timestamp 1649977179
transform 1 0 9752 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_10_125
timestamp 1649977179
transform 1 0 12604 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_133
timestamp 1649977179
transform 1 0 13340 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_136
timestamp 1649977179
transform 1 0 13616 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_159
timestamp 1649977179
transform 1 0 15732 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_192
timestamp 1649977179
transform 1 0 18768 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_197
timestamp 1649977179
transform 1 0 19228 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_38
timestamp 1649977179
transform 1 0 4600 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_50
timestamp 1649977179
transform 1 0 5704 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_61
timestamp 1649977179
transform 1 0 6716 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_113
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_135
timestamp 1649977179
transform 1 0 13524 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_190
timestamp 1649977179
transform 1 0 18584 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_13
timestamp 1649977179
transform 1 0 2300 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_25
timestamp 1649977179
transform 1 0 3404 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_135
timestamp 1649977179
transform 1 0 13524 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_184
timestamp 1649977179
transform 1 0 18032 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_15
timestamp 1649977179
transform 1 0 2484 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_37
timestamp 1649977179
transform 1 0 4508 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1649977179
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_137
timestamp 1649977179
transform 1 0 13708 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_163
timestamp 1649977179
transform 1 0 16100 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1649977179
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_209
timestamp 1649977179
transform 1 0 20332 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1649977179
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_42
timestamp 1649977179
transform 1 0 4968 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_66
timestamp 1649977179
transform 1 0 7176 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_78
timestamp 1649977179
transform 1 0 8280 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_14_85
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_91
timestamp 1649977179
transform 1 0 9476 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_101
timestamp 1649977179
transform 1 0 10396 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_131
timestamp 1649977179
transform 1 0 13156 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1649977179
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_159
timestamp 1649977179
transform 1 0 15732 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_14_178
timestamp 1649977179
transform 1 0 17480 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_184
timestamp 1649977179
transform 1 0 18032 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_206
timestamp 1649977179
transform 1 0 20056 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_3
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_22
timestamp 1649977179
transform 1 0 3128 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_47
timestamp 1649977179
transform 1 0 5428 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_53
timestamp 1649977179
transform 1 0 5980 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_75
timestamp 1649977179
transform 1 0 8004 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_110
timestamp 1649977179
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_113
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_119
timestamp 1649977179
transform 1 0 12052 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_122
timestamp 1649977179
transform 1 0 12328 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_134
timestamp 1649977179
transform 1 0 13432 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_140
timestamp 1649977179
transform 1 0 13984 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_159
timestamp 1649977179
transform 1 0 15732 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1649977179
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_169
timestamp 1649977179
transform 1 0 16652 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_190
timestamp 1649977179
transform 1 0 18584 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_218
timestamp 1649977179
transform 1 0 21160 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_21
timestamp 1649977179
transform 1 0 3036 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1649977179
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_44
timestamp 1649977179
transform 1 0 5152 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_16_101
timestamp 1649977179
transform 1 0 10396 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_157
timestamp 1649977179
transform 1 0 15548 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_162
timestamp 1649977179
transform 1 0 16008 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_175
timestamp 1649977179
transform 1 0 17204 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_178
timestamp 1649977179
transform 1 0 17480 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_190
timestamp 1649977179
transform 1 0 18584 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_206
timestamp 1649977179
transform 1 0 20056 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_209
timestamp 1649977179
transform 1 0 20332 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_7
timestamp 1649977179
transform 1 0 1748 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_18
timestamp 1649977179
transform 1 0 2760 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_30
timestamp 1649977179
transform 1 0 3864 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_42
timestamp 1649977179
transform 1 0 4968 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1649977179
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_84
timestamp 1649977179
transform 1 0 8832 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_113
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_134
timestamp 1649977179
transform 1 0 13432 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_17_159
timestamp 1649977179
transform 1 0 15732 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1649977179
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_210
timestamp 1649977179
transform 1 0 20424 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1649977179
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_33
timestamp 1649977179
transform 1 0 4140 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_45
timestamp 1649977179
transform 1 0 5244 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_74
timestamp 1649977179
transform 1 0 7912 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_85
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_132
timestamp 1649977179
transform 1 0 13248 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_157
timestamp 1649977179
transform 1 0 15548 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_169
timestamp 1649977179
transform 1 0 16652 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_181
timestamp 1649977179
transform 1 0 17756 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_193
timestamp 1649977179
transform 1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_16
timestamp 1649977179
transform 1 0 2576 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_35
timestamp 1649977179
transform 1 0 4324 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_44
timestamp 1649977179
transform 1 0 5152 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_73
timestamp 1649977179
transform 1 0 7820 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_76
timestamp 1649977179
transform 1 0 8096 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_108
timestamp 1649977179
transform 1 0 11040 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_122
timestamp 1649977179
transform 1 0 12328 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_142
timestamp 1649977179
transform 1 0 14168 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_19_196
timestamp 1649977179
transform 1 0 19136 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_202
timestamp 1649977179
transform 1 0 19688 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_209
timestamp 1649977179
transform 1 0 20332 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_13
timestamp 1649977179
transform 1 0 2300 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_25
timestamp 1649977179
transform 1 0 3404 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_29
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1649977179
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_53
timestamp 1649977179
transform 1 0 5980 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_103
timestamp 1649977179
transform 1 0 10580 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_136
timestamp 1649977179
transform 1 0 13616 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_141
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_187
timestamp 1649977179
transform 1 0 18308 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_193
timestamp 1649977179
transform 1 0 18860 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_200
timestamp 1649977179
transform 1 0 19504 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_7
timestamp 1649977179
transform 1 0 1748 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_13
timestamp 1649977179
transform 1 0 2300 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_25
timestamp 1649977179
transform 1 0 3404 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_40
timestamp 1649977179
transform 1 0 4784 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_50
timestamp 1649977179
transform 1 0 5704 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_53
timestamp 1649977179
transform 1 0 5980 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_73
timestamp 1649977179
transform 1 0 7820 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_77
timestamp 1649977179
transform 1 0 8188 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_113
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_121
timestamp 1649977179
transform 1 0 12236 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_132
timestamp 1649977179
transform 1 0 13248 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_163
timestamp 1649977179
transform 1 0 16100 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1649977179
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_205
timestamp 1649977179
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_11
timestamp 1649977179
transform 1 0 2116 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_22_22
timestamp 1649977179
transform 1 0 3128 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_22_38
timestamp 1649977179
transform 1 0 4600 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_69
timestamp 1649977179
transform 1 0 7452 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_80
timestamp 1649977179
transform 1 0 8464 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_85
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_105
timestamp 1649977179
transform 1 0 10764 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_129
timestamp 1649977179
transform 1 0 12972 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_137
timestamp 1649977179
transform 1 0 13708 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_157
timestamp 1649977179
transform 1 0 15548 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_172
timestamp 1649977179
transform 1 0 16928 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_176
timestamp 1649977179
transform 1 0 17296 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_180
timestamp 1649977179
transform 1 0 17664 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_188
timestamp 1649977179
transform 1 0 18400 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_209
timestamp 1649977179
transform 1 0 20332 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_13
timestamp 1649977179
transform 1 0 2300 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_22
timestamp 1649977179
transform 1 0 3128 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_30
timestamp 1649977179
transform 1 0 3864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_49
timestamp 1649977179
transform 1 0 5612 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_53
timestamp 1649977179
transform 1 0 5980 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_86
timestamp 1649977179
transform 1 0 9016 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_23_129
timestamp 1649977179
transform 1 0 12972 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_135
timestamp 1649977179
transform 1 0 13524 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_154
timestamp 1649977179
transform 1 0 15272 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_157
timestamp 1649977179
transform 1 0 15548 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_165
timestamp 1649977179
transform 1 0 16284 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_169
timestamp 1649977179
transform 1 0 16652 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_23_183
timestamp 1649977179
transform 1 0 17940 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_189
timestamp 1649977179
transform 1 0 18492 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_199
timestamp 1649977179
transform 1 0 19412 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_7
timestamp 1649977179
transform 1 0 1748 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_22
timestamp 1649977179
transform 1 0 3128 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_24_29
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_24_38
timestamp 1649977179
transform 1 0 4600 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_46
timestamp 1649977179
transform 1 0 5336 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_74
timestamp 1649977179
transform 1 0 7912 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1649977179
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_115
timestamp 1649977179
transform 1 0 11684 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_127
timestamp 1649977179
transform 1 0 12788 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_135
timestamp 1649977179
transform 1 0 13524 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_193
timestamp 1649977179
transform 1 0 18860 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_197
timestamp 1649977179
transform 1 0 19228 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_205
timestamp 1649977179
transform 1 0 19964 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_209
timestamp 1649977179
transform 1 0 20332 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_217
timestamp 1649977179
transform 1 0 21068 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_30
timestamp 1649977179
transform 1 0 3864 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_38
timestamp 1649977179
transform 1 0 4600 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_49
timestamp 1649977179
transform 1 0 5612 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_53
timestamp 1649977179
transform 1 0 5980 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_73
timestamp 1649977179
transform 1 0 7820 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_85
timestamp 1649977179
transform 1 0 8924 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_98
timestamp 1649977179
transform 1 0 10120 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_102
timestamp 1649977179
transform 1 0 10488 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_113
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_126
timestamp 1649977179
transform 1 0 12696 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_134
timestamp 1649977179
transform 1 0 13432 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_154
timestamp 1649977179
transform 1 0 15272 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_169
timestamp 1649977179
transform 1 0 16652 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_192
timestamp 1649977179
transform 1 0 18768 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_204
timestamp 1649977179
transform 1 0 19872 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_7
timestamp 1649977179
transform 1 0 1748 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_13
timestamp 1649977179
transform 1 0 2300 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_38
timestamp 1649977179
transform 1 0 4600 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_50
timestamp 1649977179
transform 1 0 5704 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_26_78
timestamp 1649977179
transform 1 0 8280 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_26_85
timestamp 1649977179
transform 1 0 8924 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_26_109
timestamp 1649977179
transform 1 0 11132 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_136
timestamp 1649977179
transform 1 0 13616 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_157
timestamp 1649977179
transform 1 0 15548 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_161
timestamp 1649977179
transform 1 0 15916 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_176
timestamp 1649977179
transform 1 0 17296 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1649977179
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_197
timestamp 1649977179
transform 1 0 19228 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_205
timestamp 1649977179
transform 1 0 19964 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_7
timestamp 1649977179
transform 1 0 1748 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_19
timestamp 1649977179
transform 1 0 2852 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_27
timestamp 1649977179
transform 1 0 3588 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_38
timestamp 1649977179
transform 1 0 4600 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_57
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_76
timestamp 1649977179
transform 1 0 8096 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_104
timestamp 1649977179
transform 1 0 10672 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_113
timestamp 1649977179
transform 1 0 11500 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_155
timestamp 1649977179
transform 1 0 15364 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_190
timestamp 1649977179
transform 1 0 18584 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_205
timestamp 1649977179
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_217
timestamp 1649977179
transform 1 0 21068 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_20
timestamp 1649977179
transform 1 0 2944 0 1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1649977179
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_41
timestamp 1649977179
transform 1 0 4876 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_47
timestamp 1649977179
transform 1 0 5428 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_68
timestamp 1649977179
transform 1 0 7360 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_91
timestamp 1649977179
transform 1 0 9476 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_103
timestamp 1649977179
transform 1 0 10580 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_118
timestamp 1649977179
transform 1 0 11960 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1649977179
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_141
timestamp 1649977179
transform 1 0 14076 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_160
timestamp 1649977179
transform 1 0 15824 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_164
timestamp 1649977179
transform 1 0 16192 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1649977179
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_197
timestamp 1649977179
transform 1 0 19228 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_28_206
timestamp 1649977179
transform 1 0 20056 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_214
timestamp 1649977179
transform 1 0 20792 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_22
timestamp 1649977179
transform 1 0 3128 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_33
timestamp 1649977179
transform 1 0 4140 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_39
timestamp 1649977179
transform 1 0 4692 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_43
timestamp 1649977179
transform 1 0 5060 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_53
timestamp 1649977179
transform 1 0 5980 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_79
timestamp 1649977179
transform 1 0 8372 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1649977179
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_113
timestamp 1649977179
transform 1 0 11500 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_124
timestamp 1649977179
transform 1 0 12512 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_132
timestamp 1649977179
transform 1 0 13248 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_151
timestamp 1649977179
transform 1 0 14996 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_164
timestamp 1649977179
transform 1 0 16192 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_169
timestamp 1649977179
transform 1 0 16652 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_182
timestamp 1649977179
transform 1 0 17848 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_189
timestamp 1649977179
transform 1 0 18492 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_201
timestamp 1649977179
transform 1 0 19596 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_209
timestamp 1649977179
transform 1 0 20332 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_217
timestamp 1649977179
transform 1 0 21068 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1649977179
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_67
timestamp 1649977179
transform 1 0 7268 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_85
timestamp 1649977179
transform 1 0 8924 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_157
timestamp 1649977179
transform 1 0 15548 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_165
timestamp 1649977179
transform 1 0 16284 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_30_190
timestamp 1649977179
transform 1 0 18584 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_30_197
timestamp 1649977179
transform 1 0 19228 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_57
timestamp 1649977179
transform 1 0 6348 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_95
timestamp 1649977179
transform 1 0 9844 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_152
timestamp 1649977179
transform 1 0 15088 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_164
timestamp 1649977179
transform 1 0 16192 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_169
timestamp 1649977179
transform 1 0 16652 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_37
timestamp 1649977179
transform 1 0 4508 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1649977179
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_122
timestamp 1649977179
transform 1 0 12328 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_133
timestamp 1649977179
transform 1 0 13340 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_7
timestamp 1649977179
transform 1 0 1748 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_43
timestamp 1649977179
transform 1 0 5060 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1649977179
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_85
timestamp 1649977179
transform 1 0 8924 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_107
timestamp 1649977179
transform 1 0 10948 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1649977179
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_116
timestamp 1649977179
transform 1 0 11776 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1649977179
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_193
timestamp 1649977179
transform 1 0 18860 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 21896 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 21896 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 21896 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 21896 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 21896 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 21896 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 21896 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 21896 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 21896 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 21896 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 21896 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 21896 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 21896 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 21896 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 21896 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 21896 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 21896 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 21896 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 21896 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 21896 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 21896 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 21896 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 21896 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 21896 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 21896 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 21896 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 21896 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 21896 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1649977179
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1649977179
transform -1 0 21896 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1649977179
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1649977179
transform -1 0 21896 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1649977179
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1649977179
transform -1 0 21896 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1649977179
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1649977179
transform -1 0 21896 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1649977179
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1649977179
transform -1 0 21896 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1649977179
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1649977179
transform -1 0 21896 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1649977179
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1649977179
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1649977179
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1649977179
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1649977179
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1649977179
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1649977179
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1649977179
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1649977179
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1649977179
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1649977179
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1649977179
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1649977179
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1649977179
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1649977179
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1649977179
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1649977179
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1649977179
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1649977179
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1649977179
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1649977179
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1649977179
transform 1 0 3680 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1649977179
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1649977179
transform 1 0 8832 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1649977179
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1649977179
transform 1 0 13984 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1649977179
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1649977179
transform 1 0 19136 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  Test_en_N_FTB01 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 17204 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _056_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 19504 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _057_
timestamp 1649977179
transform 1 0 1840 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _058_
timestamp 1649977179
transform 1 0 1840 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _059_
timestamp 1649977179
transform 1 0 2116 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _060_
timestamp 1649977179
transform 1 0 2024 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _061_
timestamp 1649977179
transform 1 0 1748 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _062_
timestamp 1649977179
transform 1 0 3496 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _063_
timestamp 1649977179
transform 1 0 1932 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _064_
timestamp 1649977179
transform 1 0 2392 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _065_
timestamp 1649977179
transform 1 0 2208 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _066_
timestamp 1649977179
transform 1 0 1840 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _067_
timestamp 1649977179
transform 1 0 2484 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _068_
timestamp 1649977179
transform 1 0 2116 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _069_
timestamp 1649977179
transform 1 0 2116 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _070_
timestamp 1649977179
transform 1 0 2116 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _071_
timestamp 1649977179
transform 1 0 1932 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _072_
timestamp 1649977179
transform 1 0 2392 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _073_
timestamp 1649977179
transform 1 0 1932 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _074_
timestamp 1649977179
transform 1 0 2944 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _075_
timestamp 1649977179
transform 1 0 3220 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _076_
timestamp 1649977179
transform -1 0 2944 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _077_
timestamp 1649977179
transform -1 0 21252 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _078_
timestamp 1649977179
transform -1 0 21068 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _079_
timestamp 1649977179
transform -1 0 20884 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _080_
timestamp 1649977179
transform -1 0 20700 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _081_
timestamp 1649977179
transform -1 0 20792 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _082_
timestamp 1649977179
transform -1 0 21344 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _083_
timestamp 1649977179
transform -1 0 21068 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _084_
timestamp 1649977179
transform -1 0 20976 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _085_
timestamp 1649977179
transform -1 0 20608 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _086_
timestamp 1649977179
transform -1 0 21068 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _087_
timestamp 1649977179
transform -1 0 20700 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _088_
timestamp 1649977179
transform -1 0 20884 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _089_
timestamp 1649977179
transform -1 0 20792 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _090_
timestamp 1649977179
transform -1 0 20884 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _091_
timestamp 1649977179
transform -1 0 20608 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _092_
timestamp 1649977179
transform -1 0 20240 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _093_
timestamp 1649977179
transform 1 0 20792 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _094_
timestamp 1649977179
transform 1 0 20240 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _095_
timestamp 1649977179
transform -1 0 19780 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _096_
timestamp 1649977179
transform -1 0 19964 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _097_
timestamp 1649977179
transform -1 0 13708 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _098_
timestamp 1649977179
transform -1 0 11316 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _099_
timestamp 1649977179
transform -1 0 13984 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _100_
timestamp 1649977179
transform -1 0 15732 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _101_
timestamp 1649977179
transform -1 0 15088 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _102_
timestamp 1649977179
transform 1 0 16928 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _103_
timestamp 1649977179
transform -1 0 16008 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _104_
timestamp 1649977179
transform -1 0 16928 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _105_
timestamp 1649977179
transform -1 0 17480 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _106_
timestamp 1649977179
transform 1 0 17756 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _107_
timestamp 1649977179
transform 1 0 18124 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _108_
timestamp 1649977179
transform -1 0 18952 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _109_
timestamp 1649977179
transform -1 0 18676 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _110_
timestamp 1649977179
transform -1 0 18952 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _111_
timestamp 1649977179
transform -1 0 3772 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _112_
timestamp 1649977179
transform -1 0 4508 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _113_
timestamp 1649977179
transform -1 0 4048 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _114_
timestamp 1649977179
transform -1 0 2484 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _115_
timestamp 1649977179
transform -1 0 2760 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _116_
timestamp 1649977179
transform 1 0 20976 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clk_3_N_FTB01
timestamp 1649977179
transform 1 0 8924 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 11500 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1649977179
transform -1 0 3588 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1649977179
transform 1 0 20700 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1649977179
transform -1 0 2576 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1649977179
transform -1 0 1656 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 1649977179
transform 1 0 1748 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1649977179
transform -1 0 2392 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1649977179
transform 1 0 1380 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1649977179
transform -1 0 2392 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input11
timestamp 1649977179
transform 1 0 1748 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input12
timestamp 1649977179
transform 1 0 1380 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input13 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 2300 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1649977179
transform -1 0 1656 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1649977179
transform -1 0 1656 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input16
timestamp 1649977179
transform -1 0 2300 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1649977179
transform -1 0 2024 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input18
timestamp 1649977179
transform -1 0 2300 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp 1649977179
transform 1 0 3312 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input20
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1649977179
transform -1 0 1656 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input22
timestamp 1649977179
transform -1 0 2300 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input23
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1649977179
transform 1 0 21068 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input25
timestamp 1649977179
transform -1 0 21620 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1649977179
transform 1 0 20608 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input27
timestamp 1649977179
transform -1 0 21620 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input28
timestamp 1649977179
transform -1 0 21252 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input29
timestamp 1649977179
transform -1 0 21620 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1649977179
transform 1 0 21344 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input31
timestamp 1649977179
transform -1 0 21620 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input32
timestamp 1649977179
transform -1 0 21252 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input33
timestamp 1649977179
transform -1 0 21620 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1649977179
transform 1 0 21344 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1649977179
transform 1 0 21344 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input36
timestamp 1649977179
transform 1 0 20700 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1649977179
transform 1 0 20608 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input38
timestamp 1649977179
transform 1 0 20700 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input39
timestamp 1649977179
transform -1 0 21252 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input40
timestamp 1649977179
transform -1 0 21620 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1649977179
transform 1 0 18860 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input42
timestamp 1649977179
transform 1 0 20700 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input43
timestamp 1649977179
transform -1 0 21620 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1649977179
transform -1 0 8188 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1649977179
transform 1 0 9292 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1649977179
transform 1 0 9568 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1649977179
transform -1 0 10120 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1649977179
transform 1 0 11500 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input49
timestamp 1649977179
transform 1 0 11684 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input50
timestamp 1649977179
transform -1 0 12788 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input51
timestamp 1649977179
transform 1 0 12420 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input52
timestamp 1649977179
transform 1 0 12788 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1649977179
transform -1 0 13984 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input54
timestamp 1649977179
transform -1 0 14996 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1649977179
transform -1 0 5428 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1649977179
transform -1 0 7176 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1649977179
transform -1 0 7452 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1649977179
transform -1 0 7728 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1649977179
transform 1 0 7728 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1649977179
transform -1 0 8280 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1649977179
transform 1 0 8280 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1649977179
transform -1 0 8832 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1649977179
transform -1 0 9292 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1649977179
transform 1 0 16100 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1649977179
transform -1 0 1656 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1649977179
transform -1 0 2208 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input67
timestamp 1649977179
transform -1 0 1932 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input68
timestamp 1649977179
transform -1 0 1656 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input69
timestamp 1649977179
transform -1 0 2208 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input70
timestamp 1649977179
transform -1 0 2300 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input71
timestamp 1649977179
transform -1 0 1932 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input72
timestamp 1649977179
transform -1 0 1656 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input73
timestamp 1649977179
transform -1 0 1656 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input74
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input75
timestamp 1649977179
transform 1 0 21068 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input76
timestamp 1649977179
transform 1 0 20700 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input77
timestamp 1649977179
transform 1 0 21344 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input78
timestamp 1649977179
transform 1 0 21344 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input79
timestamp 1649977179
transform 1 0 21344 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input80
timestamp 1649977179
transform 1 0 21068 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input81
timestamp 1649977179
transform 1 0 21068 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input82
timestamp 1649977179
transform 1 0 21344 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input83
timestamp 1649977179
transform 1 0 21344 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input84
timestamp 1649977179
transform -1 0 2760 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input85
timestamp 1649977179
transform 1 0 2484 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input86
timestamp 1649977179
transform -1 0 3680 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input87
timestamp 1649977179
transform -1 0 3496 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input88
timestamp 1649977179
transform 1 0 3772 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input89
timestamp 1649977179
transform -1 0 4232 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input90
timestamp 1649977179
transform 1 0 4692 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input91
timestamp 1649977179
transform -1 0 4876 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 16100 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 7176 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 6348 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 8188 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 8740 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 10580 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 8832 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 8740 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 4876 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 7820 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 7820 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 6256 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 5888 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 7820 0 1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 7084 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 7820 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 7728 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 6624 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 7176 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 4784 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 6624 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 8188 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 7452 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 12052 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 15548 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 16560 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 15548 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 15088 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 11684 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 12328 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 15732 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 14444 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 15732 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 8924 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 9844 0 -1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 10856 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 15732 0 -1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 8464 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 13800 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 15364 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 11868 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 15272 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 12696 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 14168 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 7360 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 9108 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 11868 0 -1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 12604 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 9292 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 9936 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 12788 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 9752 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 12420 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 14996 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 12972 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 11500 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 15548 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 17020 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 15824 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 8188 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 10856 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 8832 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 5980 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 7912 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 8004 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 8372 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 9844 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 11868 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14076 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 14812 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 9936 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 12052 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 9200 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_38.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 10580 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_38.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 13524 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 7820 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1649977179
transform 1 0 4232 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_2_
timestamp 1649977179
transform 1 0 3956 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1649977179
transform 1 0 3772 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1649977179
transform 1 0 3404 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_2_
timestamp 1649977179
transform -1 0 2484 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_1.mux_l2_in_3__178 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3312 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_3_
timestamp 1649977179
transform 1 0 2024 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1649977179
transform 1 0 2852 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_1_
timestamp 1649977179
transform -1 0 2484 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l4_in_0_
timestamp 1649977179
transform 1 0 2392 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 2300 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1649977179
transform 1 0 10304 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1649977179
transform 1 0 9476 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1649977179
transform -1 0 5060 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_2_
timestamp 1649977179
transform -1 0 5428 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_3.mux_l2_in_3__181
timestamp 1649977179
transform 1 0 6716 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_3_
timestamp 1649977179
transform 1 0 5888 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1649977179
transform 1 0 5060 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_1_
timestamp 1649977179
transform 1 0 4876 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l4_in_0_
timestamp 1649977179
transform 1 0 4324 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 2576 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1649977179
transform 1 0 5336 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1649977179
transform 1 0 4232 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_3_
timestamp 1649977179
transform 1 0 2760 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_4_
timestamp 1649977179
transform -1 0 3588 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_5_
timestamp 1649977179
transform -1 0 3404 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_6_
timestamp 1649977179
transform 1 0 3588 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1649977179
transform 1 0 3680 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1649977179
transform 1 0 2300 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_2_
timestamp 1649977179
transform 1 0 2852 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_5.mux_l2_in_3__183
timestamp 1649977179
transform 1 0 2300 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_3_
timestamp 1649977179
transform -1 0 2484 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1649977179
transform 1 0 2024 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_1_
timestamp 1649977179
transform 1 0 1748 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l4_in_0_
timestamp 1649977179
transform -1 0 2300 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2024 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1649977179
transform -1 0 9016 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1649977179
transform 1 0 8372 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_1_
timestamp 1649977179
transform 1 0 2760 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_2_
timestamp 1649977179
transform 1 0 2484 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_9.mux_l2_in_3__184
timestamp 1649977179
transform 1 0 3220 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_3_
timestamp 1649977179
transform -1 0 3220 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_0_
timestamp 1649977179
transform -1 0 3496 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_1_
timestamp 1649977179
transform -1 0 3312 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l4_in_0_
timestamp 1649977179
transform 1 0 3496 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 2852 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1649977179
transform 1 0 5152 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_1_
timestamp 1649977179
transform 1 0 7820 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_2_
timestamp 1649977179
transform -1 0 4600 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_17.mux_l1_in_3__179
timestamp 1649977179
transform -1 0 4600 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_3_
timestamp 1649977179
transform 1 0 4784 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1649977179
transform 1 0 4876 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_1_
timestamp 1649977179
transform -1 0 4600 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l3_in_0_
timestamp 1649977179
transform 1 0 3956 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 2668 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1649977179
transform 1 0 5428 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_2_
timestamp 1649977179
transform -1 0 3680 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_25.mux_l1_in_3__180
timestamp 1649977179
transform 1 0 3404 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_3_
timestamp 1649977179
transform -1 0 3404 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1649977179
transform 1 0 4784 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_1_
timestamp 1649977179
transform -1 0 4600 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l3_in_0_
timestamp 1649977179
transform 1 0 3772 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2300 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7820 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_1_
timestamp 1649977179
transform 1 0 7084 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_2_
timestamp 1649977179
transform 1 0 5060 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1649977179
transform 1 0 5428 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_33.mux_l2_in_1__182
timestamp 1649977179
transform 1 0 4876 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_1_
timestamp 1649977179
transform 1 0 4416 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l3_in_0_
timestamp 1649977179
transform 1 0 4048 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 2392 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1649977179
transform -1 0 11132 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1649977179
transform 1 0 17020 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1649977179
transform -1 0 17112 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1649977179
transform 1 0 18124 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_2_
timestamp 1649977179
transform 1 0 17940 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_0.mux_l2_in_3__185
timestamp 1649977179
transform 1 0 18308 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_3_
timestamp 1649977179
transform 1 0 17480 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1649977179
transform 1 0 17112 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_1_
timestamp 1649977179
transform 1 0 16836 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l4_in_0_
timestamp 1649977179
transform -1 0 17480 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 20700 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1649977179
transform -1 0 10396 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1649977179
transform -1 0 17480 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1649977179
transform -1 0 17756 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1649977179
transform 1 0 18308 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_2_
timestamp 1649977179
transform 1 0 19136 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_2.mux_l2_in_3__187
timestamp 1649977179
transform 1 0 19964 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_3_
timestamp 1649977179
transform 1 0 19228 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1649977179
transform -1 0 18584 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_1_
timestamp 1649977179
transform 1 0 18308 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l4_in_0_
timestamp 1649977179
transform -1 0 18676 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 19504 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1649977179
transform -1 0 11224 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1649977179
transform -1 0 17848 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1649977179
transform 1 0 19596 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_3_
timestamp 1649977179
transform 1 0 19964 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_4_
timestamp 1649977179
transform -1 0 21436 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_5_
timestamp 1649977179
transform -1 0 19136 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_6_
timestamp 1649977179
transform 1 0 20332 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1649977179
transform -1 0 18676 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1649977179
transform 1 0 19136 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_2_
timestamp 1649977179
transform 1 0 20792 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_4.mux_l2_in_3__162
timestamp 1649977179
transform -1 0 20700 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_3_
timestamp 1649977179
transform 1 0 20148 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1649977179
transform -1 0 19504 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_1_
timestamp 1649977179
transform 1 0 19504 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l4_in_0_
timestamp 1649977179
transform -1 0 20056 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 20148 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1649977179
transform -1 0 10856 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1649977179
transform -1 0 17480 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_1_
timestamp 1649977179
transform 1 0 19228 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_2_
timestamp 1649977179
transform -1 0 19872 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_8.mux_l2_in_3__163
timestamp 1649977179
transform -1 0 20332 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_3_
timestamp 1649977179
transform 1 0 20056 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_0_
timestamp 1649977179
transform -1 0 19136 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_1_
timestamp 1649977179
transform 1 0 19228 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l4_in_0_
timestamp 1649977179
transform -1 0 19136 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 19136 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1649977179
transform -1 0 8464 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_1_
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_2_
timestamp 1649977179
transform 1 0 19228 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_16.mux_l1_in_3__186
timestamp 1649977179
transform 1 0 20056 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_3_
timestamp 1649977179
transform 1 0 19136 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1649977179
transform -1 0 16928 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_1_
timestamp 1649977179
transform 1 0 18584 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l3_in_0_
timestamp 1649977179
transform -1 0 17756 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 20332 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1649977179
transform -1 0 8832 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1649977179
transform -1 0 17296 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_2_
timestamp 1649977179
transform 1 0 18216 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_24.mux_l1_in_3__188
timestamp 1649977179
transform -1 0 18492 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_3_
timestamp 1649977179
transform 1 0 18216 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1649977179
transform 1 0 17480 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_1_
timestamp 1649977179
transform 1 0 17388 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_0_
timestamp 1649977179
transform -1 0 16560 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 20056 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1649977179
transform -1 0 10672 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_1_
timestamp 1649977179
transform -1 0 17204 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_2_
timestamp 1649977179
transform 1 0 17480 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1649977179
transform -1 0 17480 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_32.mux_l2_in_1__161
timestamp 1649977179
transform -1 0 17664 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_1_
timestamp 1649977179
transform -1 0 18308 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l3_in_0_
timestamp 1649977179
transform -1 0 18308 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 19964 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1649977179
transform -1 0 8832 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1649977179
transform -1 0 9844 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1649977179
transform -1 0 11408 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_2_
timestamp 1649977179
transform -1 0 9752 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_0.mux_l2_in_3__164
timestamp 1649977179
transform -1 0 8648 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_3_
timestamp 1649977179
transform -1 0 9476 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1649977179
transform 1 0 10672 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_1_
timestamp 1649977179
transform -1 0 9752 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l4_in_0_
timestamp 1649977179
transform -1 0 11408 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 13616 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1649977179
transform 1 0 11960 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_1_
timestamp 1649977179
transform 1 0 11592 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_2_
timestamp 1649977179
transform 1 0 14996 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_2.mux_l1_in_3__170
timestamp 1649977179
transform 1 0 14536 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_3_
timestamp 1649977179
transform 1 0 14168 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1649977179
transform -1 0 11408 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1649977179
transform 1 0 11684 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1649977179
transform 1 0 10856 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 11132 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1649977179
transform -1 0 12328 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_1_
timestamp 1649977179
transform -1 0 13248 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_2_
timestamp 1649977179
transform 1 0 16928 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_4.mux_l1_in_3__175
timestamp 1649977179
transform -1 0 16560 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_3_
timestamp 1649977179
transform 1 0 17480 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1649977179
transform 1 0 12788 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1649977179
transform 1 0 16652 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1649977179
transform -1 0 13248 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 13616 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_0_
timestamp 1649977179
transform -1 0 11960 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_1_
timestamp 1649977179
transform -1 0 12880 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_2_
timestamp 1649977179
transform 1 0 17572 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_6.mux_l1_in_3__176
timestamp 1649977179
transform 1 0 18308 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_3_
timestamp 1649977179
transform 1 0 17388 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l2_in_0_
timestamp 1649977179
transform -1 0 13708 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l2_in_1_
timestamp 1649977179
transform 1 0 16560 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l3_in_0_
timestamp 1649977179
transform -1 0 16192 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 16100 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1649977179
transform -1 0 10028 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1649977179
transform 1 0 14996 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_8.mux_l2_in_1__177
timestamp 1649977179
transform -1 0 15916 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_1_
timestamp 1649977179
transform 1 0 15824 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_0_
timestamp 1649977179
transform -1 0 14996 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 15272 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l1_in_0_
timestamp 1649977179
transform 1 0 17848 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l2_in_0_
timestamp 1649977179
transform 1 0 17020 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_10.mux_l2_in_1__165
timestamp 1649977179
transform -1 0 16468 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l2_in_1_
timestamp 1649977179
transform 1 0 16744 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l3_in_0_
timestamp 1649977179
transform 1 0 16652 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 16560 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l1_in_0_
timestamp 1649977179
transform 1 0 11684 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_12.mux_l1_in_1__166
timestamp 1649977179
transform -1 0 10028 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l1_in_1_
timestamp 1649977179
transform 1 0 10028 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l2_in_0_
timestamp 1649977179
transform -1 0 9936 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 15456 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l1_in_0_
timestamp 1649977179
transform -1 0 6256 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_14.mux_l1_in_1__167
timestamp 1649977179
transform -1 0 5612 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l1_in_1_
timestamp 1649977179
transform -1 0 6440 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l2_in_0_
timestamp 1649977179
transform -1 0 7268 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 16652 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1649977179
transform -1 0 4968 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_16.mux_l1_in_1__168
timestamp 1649977179
transform 1 0 3036 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_1_
timestamp 1649977179
transform -1 0 3036 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1649977179
transform -1 0 5428 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 16560 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l1_in_0_
timestamp 1649977179
transform -1 0 9752 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_18.mux_l1_in_1__169
timestamp 1649977179
transform 1 0 8464 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l1_in_1_
timestamp 1649977179
transform -1 0 8464 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l2_in_0_
timestamp 1649977179
transform -1 0 10948 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 17756 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l1_in_0_
timestamp 1649977179
transform -1 0 17572 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_20.mux_l1_in_1__171
timestamp 1649977179
transform -1 0 17848 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l1_in_1_
timestamp 1649977179
transform 1 0 17572 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l2_in_0_
timestamp 1649977179
transform -1 0 17572 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 18124 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l1_in_0_
timestamp 1649977179
transform 1 0 14076 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_22.mux_l1_in_1__172
timestamp 1649977179
transform 1 0 12052 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l1_in_1_
timestamp 1649977179
transform -1 0 10580 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l2_in_0_
timestamp 1649977179
transform -1 0 12512 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 18308 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1649977179
transform -1 0 9844 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_24.mux_l1_in_1__173
timestamp 1649977179
transform 1 0 10672 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_1_
timestamp 1649977179
transform 1 0 9660 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1649977179
transform -1 0 10396 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 17664 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_38.mux_l1_in_0_
timestamp 1649977179
transform 1 0 12696 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_38.mux_l2_in_0__174
timestamp 1649977179
transform 1 0 13248 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_38.mux_l2_in_0_
timestamp 1649977179
transform -1 0 13248 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_38.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 20056 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output92 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 20516 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1649977179
transform -1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1649977179
transform -1 0 7268 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1649977179
transform -1 0 1748 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1649977179
transform -1 0 2116 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1649977179
transform -1 0 1748 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1649977179
transform -1 0 1748 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1649977179
transform -1 0 1748 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp 1649977179
transform -1 0 2116 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1649977179
transform -1 0 1748 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp 1649977179
transform -1 0 1748 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp 1649977179
transform -1 0 2116 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output104
timestamp 1649977179
transform -1 0 2484 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output105
timestamp 1649977179
transform 1 0 2852 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output106
timestamp 1649977179
transform -1 0 1748 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output107
timestamp 1649977179
transform -1 0 2116 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output108
timestamp 1649977179
transform -1 0 1748 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output109
timestamp 1649977179
transform -1 0 1748 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output110
timestamp 1649977179
transform -1 0 1748 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output111
timestamp 1649977179
transform -1 0 2116 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output112
timestamp 1649977179
transform -1 0 1748 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output113
timestamp 1649977179
transform -1 0 1748 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output114
timestamp 1649977179
transform -1 0 1748 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output115
timestamp 1649977179
transform 1 0 21252 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output116
timestamp 1649977179
transform 1 0 20884 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output117
timestamp 1649977179
transform 1 0 21252 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output118
timestamp 1649977179
transform 1 0 21252 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output119
timestamp 1649977179
transform 1 0 21252 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output120
timestamp 1649977179
transform 1 0 20884 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output121
timestamp 1649977179
transform 1 0 21252 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output122
timestamp 1649977179
transform -1 0 20516 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output123
timestamp 1649977179
transform -1 0 20148 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output124
timestamp 1649977179
transform 1 0 20516 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output125
timestamp 1649977179
transform 1 0 20884 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output126
timestamp 1649977179
transform 1 0 21252 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output127
timestamp 1649977179
transform 1 0 20884 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output128
timestamp 1649977179
transform 1 0 21252 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output129
timestamp 1649977179
transform 1 0 21252 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output130
timestamp 1649977179
transform 1 0 21252 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output131
timestamp 1649977179
transform 1 0 20884 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output132
timestamp 1649977179
transform 1 0 21252 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output133
timestamp 1649977179
transform 1 0 21252 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output134
timestamp 1649977179
transform 1 0 21252 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output135
timestamp 1649977179
transform 1 0 14996 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output136
timestamp 1649977179
transform 1 0 18124 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output137
timestamp 1649977179
transform -1 0 18860 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output138
timestamp 1649977179
transform -1 0 18676 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output139
timestamp 1649977179
transform 1 0 19228 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output140
timestamp 1649977179
transform 1 0 19596 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output141
timestamp 1649977179
transform 1 0 19964 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output142
timestamp 1649977179
transform 1 0 20332 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output143
timestamp 1649977179
transform -1 0 21068 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output144
timestamp 1649977179
transform 1 0 21068 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output145
timestamp 1649977179
transform -1 0 21252 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output146
timestamp 1649977179
transform 1 0 15364 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output147
timestamp 1649977179
transform 1 0 14904 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output148
timestamp 1649977179
transform 1 0 15732 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output149
timestamp 1649977179
transform 1 0 16100 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output150
timestamp 1649977179
transform -1 0 16100 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output151
timestamp 1649977179
transform 1 0 16652 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output152
timestamp 1649977179
transform 1 0 17020 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output153
timestamp 1649977179
transform 1 0 17388 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output154
timestamp 1649977179
transform 1 0 17756 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output155
timestamp 1649977179
transform -1 0 6164 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output156
timestamp 1649977179
transform 1 0 6348 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  prog_clk_3_N_FTB01
timestamp 1649977179
transform -1 0 6256 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  repeater157
timestamp 1649977179
transform 1 0 20056 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater158
timestamp 1649977179
transform 1 0 15640 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater159
timestamp 1649977179
transform -1 0 4968 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater160
timestamp 1649977179
transform 1 0 6164 0 1 11968
box -38 -48 958 592
<< labels >>
flabel metal2 s 1674 22200 1730 23000 0 FreeSans 224 90 0 0 SC_IN_TOP
port 0 nsew signal input
flabel metal2 s 21178 22200 21234 23000 0 FreeSans 224 90 0 0 SC_OUT_TOP
port 1 nsew signal tristate
flabel metal2 s 5354 22200 5410 23000 0 FreeSans 224 90 0 0 Test_en_N_out
port 2 nsew signal tristate
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 Test_en_S_in
port 3 nsew signal input
flabel metal4 s 6142 2128 6462 20720 0 FreeSans 1920 90 0 0 VGND
port 4 nsew ground bidirectional
flabel metal4 s 11340 2128 11660 20720 0 FreeSans 1920 90 0 0 VGND
port 4 nsew ground bidirectional
flabel metal4 s 16538 2128 16858 20720 0 FreeSans 1920 90 0 0 VGND
port 4 nsew ground bidirectional
flabel metal4 s 21736 2128 22056 20720 0 FreeSans 1920 90 0 0 VGND
port 4 nsew ground bidirectional
flabel metal4 s 3543 2128 3863 20720 0 FreeSans 1920 90 0 0 VPWR
port 5 nsew power bidirectional
flabel metal4 s 8741 2128 9061 20720 0 FreeSans 1920 90 0 0 VPWR
port 5 nsew power bidirectional
flabel metal4 s 13939 2128 14259 20720 0 FreeSans 1920 90 0 0 VPWR
port 5 nsew power bidirectional
flabel metal4 s 19137 2128 19457 20720 0 FreeSans 1920 90 0 0 VPWR
port 5 nsew power bidirectional
flabel metal2 s 2226 0 2282 800 0 FreeSans 224 90 0 0 ccff_head
port 6 nsew signal input
flabel metal2 s 6826 0 6882 800 0 FreeSans 224 90 0 0 ccff_tail
port 7 nsew signal tristate
flabel metal3 s 0 5312 800 5432 0 FreeSans 480 0 0 0 chanx_left_in[0]
port 8 nsew signal input
flabel metal3 s 0 9392 800 9512 0 FreeSans 480 0 0 0 chanx_left_in[10]
port 9 nsew signal input
flabel metal3 s 0 9800 800 9920 0 FreeSans 480 0 0 0 chanx_left_in[11]
port 10 nsew signal input
flabel metal3 s 0 10208 800 10328 0 FreeSans 480 0 0 0 chanx_left_in[12]
port 11 nsew signal input
flabel metal3 s 0 10616 800 10736 0 FreeSans 480 0 0 0 chanx_left_in[13]
port 12 nsew signal input
flabel metal3 s 0 11024 800 11144 0 FreeSans 480 0 0 0 chanx_left_in[14]
port 13 nsew signal input
flabel metal3 s 0 11432 800 11552 0 FreeSans 480 0 0 0 chanx_left_in[15]
port 14 nsew signal input
flabel metal3 s 0 11840 800 11960 0 FreeSans 480 0 0 0 chanx_left_in[16]
port 15 nsew signal input
flabel metal3 s 0 12248 800 12368 0 FreeSans 480 0 0 0 chanx_left_in[17]
port 16 nsew signal input
flabel metal3 s 0 12656 800 12776 0 FreeSans 480 0 0 0 chanx_left_in[18]
port 17 nsew signal input
flabel metal3 s 0 13064 800 13184 0 FreeSans 480 0 0 0 chanx_left_in[19]
port 18 nsew signal input
flabel metal3 s 0 5720 800 5840 0 FreeSans 480 0 0 0 chanx_left_in[1]
port 19 nsew signal input
flabel metal3 s 0 6128 800 6248 0 FreeSans 480 0 0 0 chanx_left_in[2]
port 20 nsew signal input
flabel metal3 s 0 6536 800 6656 0 FreeSans 480 0 0 0 chanx_left_in[3]
port 21 nsew signal input
flabel metal3 s 0 6944 800 7064 0 FreeSans 480 0 0 0 chanx_left_in[4]
port 22 nsew signal input
flabel metal3 s 0 7352 800 7472 0 FreeSans 480 0 0 0 chanx_left_in[5]
port 23 nsew signal input
flabel metal3 s 0 7760 800 7880 0 FreeSans 480 0 0 0 chanx_left_in[6]
port 24 nsew signal input
flabel metal3 s 0 8168 800 8288 0 FreeSans 480 0 0 0 chanx_left_in[7]
port 25 nsew signal input
flabel metal3 s 0 8576 800 8696 0 FreeSans 480 0 0 0 chanx_left_in[8]
port 26 nsew signal input
flabel metal3 s 0 8984 800 9104 0 FreeSans 480 0 0 0 chanx_left_in[9]
port 27 nsew signal input
flabel metal3 s 0 13472 800 13592 0 FreeSans 480 0 0 0 chanx_left_out[0]
port 28 nsew signal tristate
flabel metal3 s 0 17552 800 17672 0 FreeSans 480 0 0 0 chanx_left_out[10]
port 29 nsew signal tristate
flabel metal3 s 0 17960 800 18080 0 FreeSans 480 0 0 0 chanx_left_out[11]
port 30 nsew signal tristate
flabel metal3 s 0 18368 800 18488 0 FreeSans 480 0 0 0 chanx_left_out[12]
port 31 nsew signal tristate
flabel metal3 s 0 18776 800 18896 0 FreeSans 480 0 0 0 chanx_left_out[13]
port 32 nsew signal tristate
flabel metal3 s 0 19184 800 19304 0 FreeSans 480 0 0 0 chanx_left_out[14]
port 33 nsew signal tristate
flabel metal3 s 0 19592 800 19712 0 FreeSans 480 0 0 0 chanx_left_out[15]
port 34 nsew signal tristate
flabel metal3 s 0 20000 800 20120 0 FreeSans 480 0 0 0 chanx_left_out[16]
port 35 nsew signal tristate
flabel metal3 s 0 20408 800 20528 0 FreeSans 480 0 0 0 chanx_left_out[17]
port 36 nsew signal tristate
flabel metal3 s 0 20816 800 20936 0 FreeSans 480 0 0 0 chanx_left_out[18]
port 37 nsew signal tristate
flabel metal3 s 0 21224 800 21344 0 FreeSans 480 0 0 0 chanx_left_out[19]
port 38 nsew signal tristate
flabel metal3 s 0 13880 800 14000 0 FreeSans 480 0 0 0 chanx_left_out[1]
port 39 nsew signal tristate
flabel metal3 s 0 14288 800 14408 0 FreeSans 480 0 0 0 chanx_left_out[2]
port 40 nsew signal tristate
flabel metal3 s 0 14696 800 14816 0 FreeSans 480 0 0 0 chanx_left_out[3]
port 41 nsew signal tristate
flabel metal3 s 0 15104 800 15224 0 FreeSans 480 0 0 0 chanx_left_out[4]
port 42 nsew signal tristate
flabel metal3 s 0 15512 800 15632 0 FreeSans 480 0 0 0 chanx_left_out[5]
port 43 nsew signal tristate
flabel metal3 s 0 15920 800 16040 0 FreeSans 480 0 0 0 chanx_left_out[6]
port 44 nsew signal tristate
flabel metal3 s 0 16328 800 16448 0 FreeSans 480 0 0 0 chanx_left_out[7]
port 45 nsew signal tristate
flabel metal3 s 0 16736 800 16856 0 FreeSans 480 0 0 0 chanx_left_out[8]
port 46 nsew signal tristate
flabel metal3 s 0 17144 800 17264 0 FreeSans 480 0 0 0 chanx_left_out[9]
port 47 nsew signal tristate
flabel metal3 s 22200 5312 23000 5432 0 FreeSans 480 0 0 0 chanx_right_in[0]
port 48 nsew signal input
flabel metal3 s 22200 9392 23000 9512 0 FreeSans 480 0 0 0 chanx_right_in[10]
port 49 nsew signal input
flabel metal3 s 22200 9800 23000 9920 0 FreeSans 480 0 0 0 chanx_right_in[11]
port 50 nsew signal input
flabel metal3 s 22200 10208 23000 10328 0 FreeSans 480 0 0 0 chanx_right_in[12]
port 51 nsew signal input
flabel metal3 s 22200 10616 23000 10736 0 FreeSans 480 0 0 0 chanx_right_in[13]
port 52 nsew signal input
flabel metal3 s 22200 11024 23000 11144 0 FreeSans 480 0 0 0 chanx_right_in[14]
port 53 nsew signal input
flabel metal3 s 22200 11432 23000 11552 0 FreeSans 480 0 0 0 chanx_right_in[15]
port 54 nsew signal input
flabel metal3 s 22200 11840 23000 11960 0 FreeSans 480 0 0 0 chanx_right_in[16]
port 55 nsew signal input
flabel metal3 s 22200 12248 23000 12368 0 FreeSans 480 0 0 0 chanx_right_in[17]
port 56 nsew signal input
flabel metal3 s 22200 12656 23000 12776 0 FreeSans 480 0 0 0 chanx_right_in[18]
port 57 nsew signal input
flabel metal3 s 22200 13064 23000 13184 0 FreeSans 480 0 0 0 chanx_right_in[19]
port 58 nsew signal input
flabel metal3 s 22200 5720 23000 5840 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 59 nsew signal input
flabel metal3 s 22200 6128 23000 6248 0 FreeSans 480 0 0 0 chanx_right_in[2]
port 60 nsew signal input
flabel metal3 s 22200 6536 23000 6656 0 FreeSans 480 0 0 0 chanx_right_in[3]
port 61 nsew signal input
flabel metal3 s 22200 6944 23000 7064 0 FreeSans 480 0 0 0 chanx_right_in[4]
port 62 nsew signal input
flabel metal3 s 22200 7352 23000 7472 0 FreeSans 480 0 0 0 chanx_right_in[5]
port 63 nsew signal input
flabel metal3 s 22200 7760 23000 7880 0 FreeSans 480 0 0 0 chanx_right_in[6]
port 64 nsew signal input
flabel metal3 s 22200 8168 23000 8288 0 FreeSans 480 0 0 0 chanx_right_in[7]
port 65 nsew signal input
flabel metal3 s 22200 8576 23000 8696 0 FreeSans 480 0 0 0 chanx_right_in[8]
port 66 nsew signal input
flabel metal3 s 22200 8984 23000 9104 0 FreeSans 480 0 0 0 chanx_right_in[9]
port 67 nsew signal input
flabel metal3 s 22200 13472 23000 13592 0 FreeSans 480 0 0 0 chanx_right_out[0]
port 68 nsew signal tristate
flabel metal3 s 22200 17552 23000 17672 0 FreeSans 480 0 0 0 chanx_right_out[10]
port 69 nsew signal tristate
flabel metal3 s 22200 17960 23000 18080 0 FreeSans 480 0 0 0 chanx_right_out[11]
port 70 nsew signal tristate
flabel metal3 s 22200 18368 23000 18488 0 FreeSans 480 0 0 0 chanx_right_out[12]
port 71 nsew signal tristate
flabel metal3 s 22200 18776 23000 18896 0 FreeSans 480 0 0 0 chanx_right_out[13]
port 72 nsew signal tristate
flabel metal3 s 22200 19184 23000 19304 0 FreeSans 480 0 0 0 chanx_right_out[14]
port 73 nsew signal tristate
flabel metal3 s 22200 19592 23000 19712 0 FreeSans 480 0 0 0 chanx_right_out[15]
port 74 nsew signal tristate
flabel metal3 s 22200 20000 23000 20120 0 FreeSans 480 0 0 0 chanx_right_out[16]
port 75 nsew signal tristate
flabel metal3 s 22200 20408 23000 20528 0 FreeSans 480 0 0 0 chanx_right_out[17]
port 76 nsew signal tristate
flabel metal3 s 22200 20816 23000 20936 0 FreeSans 480 0 0 0 chanx_right_out[18]
port 77 nsew signal tristate
flabel metal3 s 22200 21224 23000 21344 0 FreeSans 480 0 0 0 chanx_right_out[19]
port 78 nsew signal tristate
flabel metal3 s 22200 13880 23000 14000 0 FreeSans 480 0 0 0 chanx_right_out[1]
port 79 nsew signal tristate
flabel metal3 s 22200 14288 23000 14408 0 FreeSans 480 0 0 0 chanx_right_out[2]
port 80 nsew signal tristate
flabel metal3 s 22200 14696 23000 14816 0 FreeSans 480 0 0 0 chanx_right_out[3]
port 81 nsew signal tristate
flabel metal3 s 22200 15104 23000 15224 0 FreeSans 480 0 0 0 chanx_right_out[4]
port 82 nsew signal tristate
flabel metal3 s 22200 15512 23000 15632 0 FreeSans 480 0 0 0 chanx_right_out[5]
port 83 nsew signal tristate
flabel metal3 s 22200 15920 23000 16040 0 FreeSans 480 0 0 0 chanx_right_out[6]
port 84 nsew signal tristate
flabel metal3 s 22200 16328 23000 16448 0 FreeSans 480 0 0 0 chanx_right_out[7]
port 85 nsew signal tristate
flabel metal3 s 22200 16736 23000 16856 0 FreeSans 480 0 0 0 chanx_right_out[8]
port 86 nsew signal tristate
flabel metal3 s 22200 17144 23000 17264 0 FreeSans 480 0 0 0 chanx_right_out[9]
port 87 nsew signal tristate
flabel metal2 s 6458 22200 6514 23000 0 FreeSans 224 90 0 0 chany_top_in[0]
port 88 nsew signal input
flabel metal2 s 10138 22200 10194 23000 0 FreeSans 224 90 0 0 chany_top_in[10]
port 89 nsew signal input
flabel metal2 s 10506 22200 10562 23000 0 FreeSans 224 90 0 0 chany_top_in[11]
port 90 nsew signal input
flabel metal2 s 10874 22200 10930 23000 0 FreeSans 224 90 0 0 chany_top_in[12]
port 91 nsew signal input
flabel metal2 s 11242 22200 11298 23000 0 FreeSans 224 90 0 0 chany_top_in[13]
port 92 nsew signal input
flabel metal2 s 11610 22200 11666 23000 0 FreeSans 224 90 0 0 chany_top_in[14]
port 93 nsew signal input
flabel metal2 s 11978 22200 12034 23000 0 FreeSans 224 90 0 0 chany_top_in[15]
port 94 nsew signal input
flabel metal2 s 12346 22200 12402 23000 0 FreeSans 224 90 0 0 chany_top_in[16]
port 95 nsew signal input
flabel metal2 s 12714 22200 12770 23000 0 FreeSans 224 90 0 0 chany_top_in[17]
port 96 nsew signal input
flabel metal2 s 13082 22200 13138 23000 0 FreeSans 224 90 0 0 chany_top_in[18]
port 97 nsew signal input
flabel metal2 s 13450 22200 13506 23000 0 FreeSans 224 90 0 0 chany_top_in[19]
port 98 nsew signal input
flabel metal2 s 6826 22200 6882 23000 0 FreeSans 224 90 0 0 chany_top_in[1]
port 99 nsew signal input
flabel metal2 s 7194 22200 7250 23000 0 FreeSans 224 90 0 0 chany_top_in[2]
port 100 nsew signal input
flabel metal2 s 7562 22200 7618 23000 0 FreeSans 224 90 0 0 chany_top_in[3]
port 101 nsew signal input
flabel metal2 s 7930 22200 7986 23000 0 FreeSans 224 90 0 0 chany_top_in[4]
port 102 nsew signal input
flabel metal2 s 8298 22200 8354 23000 0 FreeSans 224 90 0 0 chany_top_in[5]
port 103 nsew signal input
flabel metal2 s 8666 22200 8722 23000 0 FreeSans 224 90 0 0 chany_top_in[6]
port 104 nsew signal input
flabel metal2 s 9034 22200 9090 23000 0 FreeSans 224 90 0 0 chany_top_in[7]
port 105 nsew signal input
flabel metal2 s 9402 22200 9458 23000 0 FreeSans 224 90 0 0 chany_top_in[8]
port 106 nsew signal input
flabel metal2 s 9770 22200 9826 23000 0 FreeSans 224 90 0 0 chany_top_in[9]
port 107 nsew signal input
flabel metal2 s 13818 22200 13874 23000 0 FreeSans 224 90 0 0 chany_top_out[0]
port 108 nsew signal tristate
flabel metal2 s 17498 22200 17554 23000 0 FreeSans 224 90 0 0 chany_top_out[10]
port 109 nsew signal tristate
flabel metal2 s 17866 22200 17922 23000 0 FreeSans 224 90 0 0 chany_top_out[11]
port 110 nsew signal tristate
flabel metal2 s 18234 22200 18290 23000 0 FreeSans 224 90 0 0 chany_top_out[12]
port 111 nsew signal tristate
flabel metal2 s 18602 22200 18658 23000 0 FreeSans 224 90 0 0 chany_top_out[13]
port 112 nsew signal tristate
flabel metal2 s 18970 22200 19026 23000 0 FreeSans 224 90 0 0 chany_top_out[14]
port 113 nsew signal tristate
flabel metal2 s 19338 22200 19394 23000 0 FreeSans 224 90 0 0 chany_top_out[15]
port 114 nsew signal tristate
flabel metal2 s 19706 22200 19762 23000 0 FreeSans 224 90 0 0 chany_top_out[16]
port 115 nsew signal tristate
flabel metal2 s 20074 22200 20130 23000 0 FreeSans 224 90 0 0 chany_top_out[17]
port 116 nsew signal tristate
flabel metal2 s 20442 22200 20498 23000 0 FreeSans 224 90 0 0 chany_top_out[18]
port 117 nsew signal tristate
flabel metal2 s 20810 22200 20866 23000 0 FreeSans 224 90 0 0 chany_top_out[19]
port 118 nsew signal tristate
flabel metal2 s 14186 22200 14242 23000 0 FreeSans 224 90 0 0 chany_top_out[1]
port 119 nsew signal tristate
flabel metal2 s 14554 22200 14610 23000 0 FreeSans 224 90 0 0 chany_top_out[2]
port 120 nsew signal tristate
flabel metal2 s 14922 22200 14978 23000 0 FreeSans 224 90 0 0 chany_top_out[3]
port 121 nsew signal tristate
flabel metal2 s 15290 22200 15346 23000 0 FreeSans 224 90 0 0 chany_top_out[4]
port 122 nsew signal tristate
flabel metal2 s 15658 22200 15714 23000 0 FreeSans 224 90 0 0 chany_top_out[5]
port 123 nsew signal tristate
flabel metal2 s 16026 22200 16082 23000 0 FreeSans 224 90 0 0 chany_top_out[6]
port 124 nsew signal tristate
flabel metal2 s 16394 22200 16450 23000 0 FreeSans 224 90 0 0 chany_top_out[7]
port 125 nsew signal tristate
flabel metal2 s 16762 22200 16818 23000 0 FreeSans 224 90 0 0 chany_top_out[8]
port 126 nsew signal tristate
flabel metal2 s 17130 22200 17186 23000 0 FreeSans 224 90 0 0 chany_top_out[9]
port 127 nsew signal tristate
flabel metal2 s 5722 22200 5778 23000 0 FreeSans 224 90 0 0 clk_3_N_out
port 128 nsew signal tristate
flabel metal2 s 16026 0 16082 800 0 FreeSans 224 90 0 0 clk_3_S_in
port 129 nsew signal input
flabel metal3 s 0 3680 800 3800 0 FreeSans 480 0 0 0 left_bottom_grid_pin_11_
port 130 nsew signal input
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 left_bottom_grid_pin_13_
port 131 nsew signal input
flabel metal3 s 0 4496 800 4616 0 FreeSans 480 0 0 0 left_bottom_grid_pin_15_
port 132 nsew signal input
flabel metal3 s 0 4904 800 5024 0 FreeSans 480 0 0 0 left_bottom_grid_pin_17_
port 133 nsew signal input
flabel metal3 s 0 1640 800 1760 0 FreeSans 480 0 0 0 left_bottom_grid_pin_1_
port 134 nsew signal input
flabel metal3 s 0 2048 800 2168 0 FreeSans 480 0 0 0 left_bottom_grid_pin_3_
port 135 nsew signal input
flabel metal3 s 0 2456 800 2576 0 FreeSans 480 0 0 0 left_bottom_grid_pin_5_
port 136 nsew signal input
flabel metal3 s 0 2864 800 2984 0 FreeSans 480 0 0 0 left_bottom_grid_pin_7_
port 137 nsew signal input
flabel metal3 s 0 3272 800 3392 0 FreeSans 480 0 0 0 left_bottom_grid_pin_9_
port 138 nsew signal input
flabel metal2 s 4986 22200 5042 23000 0 FreeSans 224 90 0 0 prog_clk_0_N_in
port 139 nsew signal input
flabel metal2 s 6090 22200 6146 23000 0 FreeSans 224 90 0 0 prog_clk_3_N_out
port 140 nsew signal tristate
flabel metal2 s 11426 0 11482 800 0 FreeSans 224 90 0 0 prog_clk_3_S_in
port 141 nsew signal input
flabel metal3 s 22200 3680 23000 3800 0 FreeSans 480 0 0 0 right_bottom_grid_pin_11_
port 142 nsew signal input
flabel metal3 s 22200 4088 23000 4208 0 FreeSans 480 0 0 0 right_bottom_grid_pin_13_
port 143 nsew signal input
flabel metal3 s 22200 4496 23000 4616 0 FreeSans 480 0 0 0 right_bottom_grid_pin_15_
port 144 nsew signal input
flabel metal3 s 22200 4904 23000 5024 0 FreeSans 480 0 0 0 right_bottom_grid_pin_17_
port 145 nsew signal input
flabel metal3 s 22200 1640 23000 1760 0 FreeSans 480 0 0 0 right_bottom_grid_pin_1_
port 146 nsew signal input
flabel metal3 s 22200 2048 23000 2168 0 FreeSans 480 0 0 0 right_bottom_grid_pin_3_
port 147 nsew signal input
flabel metal3 s 22200 2456 23000 2576 0 FreeSans 480 0 0 0 right_bottom_grid_pin_5_
port 148 nsew signal input
flabel metal3 s 22200 2864 23000 2984 0 FreeSans 480 0 0 0 right_bottom_grid_pin_7_
port 149 nsew signal input
flabel metal3 s 22200 3272 23000 3392 0 FreeSans 480 0 0 0 right_bottom_grid_pin_9_
port 150 nsew signal input
flabel metal2 s 2042 22200 2098 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_42_
port 151 nsew signal input
flabel metal2 s 2410 22200 2466 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_43_
port 152 nsew signal input
flabel metal2 s 2778 22200 2834 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_44_
port 153 nsew signal input
flabel metal2 s 3146 22200 3202 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_45_
port 154 nsew signal input
flabel metal2 s 3514 22200 3570 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_46_
port 155 nsew signal input
flabel metal2 s 3882 22200 3938 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_47_
port 156 nsew signal input
flabel metal2 s 4250 22200 4306 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_48_
port 157 nsew signal input
flabel metal2 s 4618 22200 4674 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_49_
port 158 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 23000 23000
<< end >>
