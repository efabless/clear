magic
tech sky130A
magscale 1 2
timestamp 1680088378
<< viali >>
rect 13829 54281 13863 54315
rect 14381 54281 14415 54315
rect 10885 54213 10919 54247
rect 15485 54213 15519 54247
rect 18429 54213 18463 54247
rect 25053 54213 25087 54247
rect 3433 54145 3467 54179
rect 6009 54145 6043 54179
rect 8585 54145 8619 54179
rect 9873 54145 9907 54179
rect 12081 54145 12115 54179
rect 14657 54145 14691 54179
rect 16129 54145 16163 54179
rect 16865 54145 16899 54179
rect 17785 54145 17819 54179
rect 19441 54145 19475 54179
rect 20361 54145 20395 54179
rect 20913 54145 20947 54179
rect 22201 54145 22235 54179
rect 23949 54145 23983 54179
rect 24777 54145 24811 54179
rect 2973 54077 3007 54111
rect 5549 54077 5583 54111
rect 8125 54077 8159 54111
rect 12541 54077 12575 54111
rect 18889 54077 18923 54111
rect 21465 54077 21499 54111
rect 23581 54077 23615 54111
rect 15669 54009 15703 54043
rect 18613 54009 18647 54043
rect 24593 54009 24627 54043
rect 14841 53941 14875 53975
rect 16313 53941 16347 53975
rect 17049 53941 17083 53975
rect 17693 53941 17727 53975
rect 19625 53941 19659 53975
rect 20269 53941 20303 53975
rect 21097 53941 21131 53975
rect 22017 53941 22051 53975
rect 15209 53737 15243 53771
rect 15485 53737 15519 53771
rect 20269 53737 20303 53771
rect 2973 53601 3007 53635
rect 6285 53601 6319 53635
rect 8309 53601 8343 53635
rect 10517 53601 10551 53635
rect 12173 53601 12207 53635
rect 23213 53601 23247 53635
rect 25053 53601 25087 53635
rect 3433 53533 3467 53567
rect 6653 53533 6687 53567
rect 7389 53533 7423 53567
rect 11069 53533 11103 53567
rect 11897 53533 11931 53567
rect 13553 53533 13587 53567
rect 14565 53533 14599 53567
rect 14841 53533 14875 53567
rect 15761 53533 15795 53567
rect 16497 53533 16531 53567
rect 17233 53533 17267 53567
rect 17969 53533 18003 53567
rect 18889 53533 18923 53567
rect 19717 53533 19751 53567
rect 19993 53533 20027 53567
rect 20545 53533 20579 53567
rect 21281 53533 21315 53567
rect 22201 53533 22235 53567
rect 24041 53533 24075 53567
rect 24777 53533 24811 53567
rect 3801 53397 3835 53431
rect 13737 53397 13771 53431
rect 14381 53397 14415 53431
rect 15945 53397 15979 53431
rect 16681 53397 16715 53431
rect 17417 53397 17451 53431
rect 18153 53397 18187 53431
rect 18705 53397 18739 53431
rect 19533 53397 19567 53431
rect 20729 53397 20763 53431
rect 21465 53397 21499 53431
rect 22017 53397 22051 53431
rect 24593 53397 24627 53431
rect 25421 53397 25455 53431
rect 2053 53193 2087 53227
rect 15945 53193 15979 53227
rect 16405 53193 16439 53227
rect 16681 53193 16715 53227
rect 17049 53193 17083 53227
rect 17877 53193 17911 53227
rect 18521 53193 18555 53227
rect 19349 53193 19383 53227
rect 20729 53193 20763 53227
rect 21097 53193 21131 53227
rect 21465 53193 21499 53227
rect 14473 53125 14507 53159
rect 14841 53125 14875 53159
rect 18245 53125 18279 53159
rect 1593 53057 1627 53091
rect 4077 53057 4111 53091
rect 5825 53057 5859 53091
rect 6837 53057 6871 53091
rect 9137 53057 9171 53091
rect 9781 53057 9815 53091
rect 11713 53057 11747 53091
rect 13829 53057 13863 53091
rect 19993 53057 20027 53091
rect 20269 53057 20303 53091
rect 21649 53057 21683 53091
rect 22017 53057 22051 53091
rect 22937 53057 22971 53091
rect 23213 53057 23247 53091
rect 25145 53057 25179 53091
rect 3709 52989 3743 53023
rect 5549 52989 5583 53023
rect 8677 52989 8711 53023
rect 10241 52989 10275 53023
rect 12173 52989 12207 53023
rect 24869 52989 24903 53023
rect 1777 52853 1811 52887
rect 6653 52853 6687 52887
rect 13645 52853 13679 52887
rect 14381 52853 14415 52887
rect 19809 52853 19843 52887
rect 22201 52853 22235 52887
rect 22753 52853 22787 52887
rect 11989 52649 12023 52683
rect 14105 52649 14139 52683
rect 21833 52649 21867 52683
rect 23949 52649 23983 52683
rect 12633 52581 12667 52615
rect 2973 52513 3007 52547
rect 3985 52513 4019 52547
rect 6101 52513 6135 52547
rect 7849 52513 7883 52547
rect 10333 52513 10367 52547
rect 25329 52513 25363 52547
rect 3433 52445 3467 52479
rect 4261 52445 4295 52479
rect 6561 52445 6595 52479
rect 8585 52445 8619 52479
rect 9873 52445 9907 52479
rect 11805 52445 11839 52479
rect 12449 52445 12483 52479
rect 13461 52445 13495 52479
rect 23121 52445 23155 52479
rect 23765 52445 23799 52479
rect 24777 52445 24811 52479
rect 25053 52445 25087 52479
rect 25421 52445 25455 52479
rect 13277 52377 13311 52411
rect 13737 52377 13771 52411
rect 23305 52309 23339 52343
rect 24593 52309 24627 52343
rect 11897 52105 11931 52139
rect 12357 52105 12391 52139
rect 23489 52105 23523 52139
rect 23949 52105 23983 52139
rect 4997 52037 5031 52071
rect 4077 51969 4111 52003
rect 6009 51969 6043 52003
rect 7021 51969 7055 52003
rect 10333 51969 10367 52003
rect 11713 51969 11747 52003
rect 23305 51969 23339 52003
rect 23765 51969 23799 52003
rect 24593 51969 24627 52003
rect 25237 51969 25271 52003
rect 3525 51901 3559 51935
rect 7389 51901 7423 51935
rect 9689 51901 9723 51935
rect 24409 51765 24443 51799
rect 25145 51765 25179 51799
rect 5917 51561 5951 51595
rect 24685 51561 24719 51595
rect 24501 51493 24535 51527
rect 2421 51425 2455 51459
rect 4169 51425 4203 51459
rect 6929 51425 6963 51459
rect 3433 51357 3467 51391
rect 5365 51357 5399 51391
rect 6101 51357 6135 51391
rect 7757 51357 7791 51391
rect 24041 51357 24075 51391
rect 25329 51357 25363 51391
rect 23857 51221 23891 51255
rect 25145 51221 25179 51255
rect 9873 51017 9907 51051
rect 10701 51017 10735 51051
rect 3065 50949 3099 50983
rect 6745 50949 6779 50983
rect 1869 50881 1903 50915
rect 4169 50881 4203 50915
rect 6929 50881 6963 50915
rect 9781 50881 9815 50915
rect 10517 50881 10551 50915
rect 24777 50881 24811 50915
rect 25329 50881 25363 50915
rect 1593 50813 1627 50847
rect 25145 50677 25179 50711
rect 1409 50405 1443 50439
rect 9413 50405 9447 50439
rect 2237 50337 2271 50371
rect 4353 50337 4387 50371
rect 3433 50269 3467 50303
rect 5365 50269 5399 50303
rect 24777 50269 24811 50303
rect 25329 50269 25363 50303
rect 9229 50201 9263 50235
rect 25145 50133 25179 50167
rect 6745 49929 6779 49963
rect 7849 49929 7883 49963
rect 25145 49929 25179 49963
rect 1961 49861 1995 49895
rect 9413 49861 9447 49895
rect 9597 49861 9631 49895
rect 3157 49793 3191 49827
rect 6561 49793 6595 49827
rect 8033 49793 8067 49827
rect 24777 49793 24811 49827
rect 25329 49793 25363 49827
rect 1777 49249 1811 49283
rect 4445 49249 4479 49283
rect 2973 49181 3007 49215
rect 6745 49181 6779 49215
rect 24777 49181 24811 49215
rect 25329 49181 25363 49215
rect 4721 49113 4755 49147
rect 6469 49113 6503 49147
rect 25145 49045 25179 49079
rect 11897 48841 11931 48875
rect 11713 48705 11747 48739
rect 24777 48705 24811 48739
rect 25329 48705 25363 48739
rect 25145 48569 25179 48603
rect 25145 48229 25179 48263
rect 25329 48093 25363 48127
rect 1685 48025 1719 48059
rect 2145 48025 2179 48059
rect 1777 47957 1811 47991
rect 23673 47957 23707 47991
rect 24501 47957 24535 47991
rect 23489 47753 23523 47787
rect 24133 47753 24167 47787
rect 24593 47685 24627 47719
rect 23305 47617 23339 47651
rect 23949 47617 23983 47651
rect 24777 47617 24811 47651
rect 25237 47481 25271 47515
rect 16957 47413 16991 47447
rect 25513 47413 25547 47447
rect 9137 47209 9171 47243
rect 11713 47209 11747 47243
rect 23857 47209 23891 47243
rect 24869 47141 24903 47175
rect 15117 47073 15151 47107
rect 17785 47073 17819 47107
rect 17877 47073 17911 47107
rect 9321 47005 9355 47039
rect 11529 47005 11563 47039
rect 16865 47005 16899 47039
rect 17693 47005 17727 47039
rect 18337 47005 18371 47039
rect 23581 47005 23615 47039
rect 24041 47005 24075 47039
rect 16589 46937 16623 46971
rect 24685 46937 24719 46971
rect 25145 46937 25179 46971
rect 17325 46869 17359 46903
rect 7113 46665 7147 46699
rect 13737 46665 13771 46699
rect 15853 46665 15887 46699
rect 17233 46665 17267 46699
rect 18521 46665 18555 46699
rect 20269 46665 20303 46699
rect 20545 46665 20579 46699
rect 15209 46597 15243 46631
rect 17325 46597 17359 46631
rect 7297 46529 7331 46563
rect 18429 46529 18463 46563
rect 19073 46529 19107 46563
rect 23489 46529 23523 46563
rect 25329 46529 25363 46563
rect 15485 46461 15519 46495
rect 17417 46461 17451 46495
rect 18613 46461 18647 46495
rect 25053 46461 25087 46495
rect 24225 46393 24259 46427
rect 16865 46325 16899 46359
rect 18061 46325 18095 46359
rect 23305 46325 23339 46359
rect 23857 46325 23891 46359
rect 15853 46121 15887 46155
rect 18153 46121 18187 46155
rect 21465 46121 21499 46155
rect 24041 46053 24075 46087
rect 17601 45985 17635 46019
rect 19625 45985 19659 46019
rect 19717 45985 19751 46019
rect 20821 45985 20855 46019
rect 21005 45985 21039 46019
rect 1593 45917 1627 45951
rect 1869 45917 1903 45951
rect 23857 45917 23891 45951
rect 24777 45917 24811 45951
rect 25053 45917 25087 45951
rect 17325 45849 17359 45883
rect 17969 45849 18003 45883
rect 19809 45849 19843 45883
rect 21097 45849 21131 45883
rect 25421 45849 25455 45883
rect 20177 45781 20211 45815
rect 24593 45781 24627 45815
rect 1409 45577 1443 45611
rect 7573 45509 7607 45543
rect 11713 45509 11747 45543
rect 14841 45509 14875 45543
rect 20177 45509 20211 45543
rect 7757 45441 7791 45475
rect 8401 45441 8435 45475
rect 9781 45441 9815 45475
rect 11161 45441 11195 45475
rect 11897 45441 11931 45475
rect 15117 45441 15151 45475
rect 20085 45441 20119 45475
rect 22661 45441 22695 45475
rect 24133 45441 24167 45475
rect 18337 45373 18371 45407
rect 18613 45373 18647 45407
rect 20361 45373 20395 45407
rect 24777 45373 24811 45407
rect 8585 45305 8619 45339
rect 9965 45305 9999 45339
rect 7205 45237 7239 45271
rect 10977 45237 11011 45271
rect 12265 45237 12299 45271
rect 13369 45237 13403 45271
rect 15393 45237 15427 45271
rect 16865 45237 16899 45271
rect 18981 45237 19015 45271
rect 19441 45237 19475 45271
rect 19717 45237 19751 45271
rect 10149 45033 10183 45067
rect 16313 45033 16347 45067
rect 7389 44965 7423 44999
rect 21833 44897 21867 44931
rect 21925 44897 21959 44931
rect 23397 44897 23431 44931
rect 7573 44829 7607 44863
rect 7941 44829 7975 44863
rect 10701 44829 10735 44863
rect 14289 44829 14323 44863
rect 21189 44829 21223 44863
rect 23213 44829 23247 44863
rect 23305 44829 23339 44863
rect 24869 44829 24903 44863
rect 25329 44829 25363 44863
rect 10057 44761 10091 44795
rect 10977 44761 11011 44795
rect 14565 44761 14599 44795
rect 20913 44761 20947 44795
rect 8401 44693 8435 44727
rect 9689 44693 9723 44727
rect 12449 44693 12483 44727
rect 12817 44693 12851 44727
rect 16037 44693 16071 44727
rect 19441 44693 19475 44727
rect 22017 44693 22051 44727
rect 22385 44693 22419 44727
rect 22845 44693 22879 44727
rect 25145 44693 25179 44727
rect 7205 44489 7239 44523
rect 8033 44489 8067 44523
rect 9045 44489 9079 44523
rect 11713 44489 11747 44523
rect 14565 44489 14599 44523
rect 17693 44489 17727 44523
rect 24133 44489 24167 44523
rect 6837 44421 6871 44455
rect 7297 44421 7331 44455
rect 8493 44421 8527 44455
rect 9689 44421 9723 44455
rect 12909 44421 12943 44455
rect 19165 44421 19199 44455
rect 7849 44353 7883 44387
rect 8677 44353 8711 44387
rect 9413 44353 9447 44387
rect 12081 44353 12115 44387
rect 13093 44353 13127 44387
rect 25053 44353 25087 44387
rect 12173 44285 12207 44319
rect 12357 44285 12391 44319
rect 14381 44285 14415 44319
rect 14473 44285 14507 44319
rect 15209 44285 15243 44319
rect 19441 44285 19475 44319
rect 21465 44285 21499 44319
rect 23489 44285 23523 44319
rect 23765 44285 23799 44319
rect 25329 44285 25363 44319
rect 14933 44217 14967 44251
rect 22017 44217 22051 44251
rect 11161 44149 11195 44183
rect 13553 44149 13587 44183
rect 19809 44149 19843 44183
rect 21281 44149 21315 44183
rect 10517 43945 10551 43979
rect 21189 43945 21223 43979
rect 22017 43945 22051 43979
rect 24133 43945 24167 43979
rect 25053 43945 25087 43979
rect 6377 43877 6411 43911
rect 8309 43877 8343 43911
rect 9689 43877 9723 43911
rect 24593 43877 24627 43911
rect 9045 43809 9079 43843
rect 15853 43809 15887 43843
rect 23765 43809 23799 43843
rect 1593 43741 1627 43775
rect 2053 43741 2087 43775
rect 8493 43741 8527 43775
rect 9413 43741 9447 43775
rect 9873 43741 9907 43775
rect 11805 43741 11839 43775
rect 19441 43741 19475 43775
rect 21465 43741 21499 43775
rect 24777 43741 24811 43775
rect 6561 43673 6595 43707
rect 10609 43673 10643 43707
rect 11069 43673 11103 43707
rect 12081 43673 12115 43707
rect 16129 43673 16163 43707
rect 17969 43673 18003 43707
rect 19717 43673 19751 43707
rect 23489 43673 23523 43707
rect 1777 43605 1811 43639
rect 7021 43605 7055 43639
rect 11253 43605 11287 43639
rect 13553 43605 13587 43639
rect 14105 43605 14139 43639
rect 17601 43605 17635 43639
rect 25513 43605 25547 43639
rect 2053 43401 2087 43435
rect 5733 43401 5767 43435
rect 8677 43401 8711 43435
rect 12265 43401 12299 43435
rect 17325 43401 17359 43435
rect 17969 43401 18003 43435
rect 23765 43401 23799 43435
rect 10793 43333 10827 43367
rect 17233 43333 17267 43367
rect 22293 43333 22327 43367
rect 24225 43333 24259 43367
rect 24317 43333 24351 43367
rect 2237 43265 2271 43299
rect 2513 43265 2547 43299
rect 5549 43265 5583 43299
rect 10425 43265 10459 43299
rect 12633 43265 12667 43299
rect 25329 43265 25363 43299
rect 10149 43197 10183 43231
rect 12725 43197 12759 43231
rect 12817 43197 12851 43231
rect 17417 43197 17451 43231
rect 22017 43197 22051 43231
rect 8217 43061 8251 43095
rect 16865 43061 16899 43095
rect 25145 43061 25179 43095
rect 14546 42857 14580 42891
rect 4169 42721 4203 42755
rect 6285 42721 6319 42755
rect 8309 42721 8343 42755
rect 9137 42721 9171 42755
rect 9505 42721 9539 42755
rect 12541 42721 12575 42755
rect 14289 42721 14323 42755
rect 18061 42721 18095 42755
rect 7021 42653 7055 42687
rect 7665 42653 7699 42687
rect 8493 42653 8527 42687
rect 9781 42653 9815 42687
rect 17969 42653 18003 42687
rect 21189 42653 21223 42687
rect 22293 42653 22327 42687
rect 24777 42653 24811 42687
rect 4353 42585 4387 42619
rect 6009 42585 6043 42619
rect 6469 42585 6503 42619
rect 20913 42585 20947 42619
rect 21741 42585 21775 42619
rect 22569 42585 22603 42619
rect 4813 42517 4847 42551
rect 7205 42517 7239 42551
rect 7849 42517 7883 42551
rect 9689 42517 9723 42551
rect 10149 42517 10183 42551
rect 11989 42517 12023 42551
rect 12357 42517 12391 42551
rect 12449 42517 12483 42551
rect 16037 42517 16071 42551
rect 16313 42517 16347 42551
rect 17509 42517 17543 42551
rect 17877 42517 17911 42551
rect 18521 42517 18555 42551
rect 19441 42517 19475 42551
rect 21557 42517 21591 42551
rect 24041 42517 24075 42551
rect 24593 42517 24627 42551
rect 25053 42517 25087 42551
rect 25513 42517 25547 42551
rect 9965 42313 9999 42347
rect 11805 42313 11839 42347
rect 22293 42313 22327 42347
rect 23305 42313 23339 42347
rect 25329 42313 25363 42347
rect 3709 42245 3743 42279
rect 12173 42245 12207 42279
rect 15669 42245 15703 42279
rect 20729 42245 20763 42279
rect 24777 42245 24811 42279
rect 3893 42177 3927 42211
rect 7849 42177 7883 42211
rect 12265 42177 12299 42211
rect 15393 42177 15427 42211
rect 17877 42177 17911 42211
rect 21465 42177 21499 42211
rect 22385 42177 22419 42211
rect 8125 42109 8159 42143
rect 12357 42109 12391 42143
rect 15117 42109 15151 42143
rect 18153 42109 18187 42143
rect 22201 42109 22235 42143
rect 25053 42109 25087 42143
rect 9597 42041 9631 42075
rect 19993 42041 20027 42075
rect 22753 42041 22787 42075
rect 4353 41973 4387 42007
rect 13645 41973 13679 42007
rect 19625 41973 19659 42007
rect 20269 41973 20303 42007
rect 4445 41769 4479 41803
rect 5365 41769 5399 41803
rect 7849 41769 7883 41803
rect 17325 41769 17359 41803
rect 16957 41701 16991 41735
rect 21465 41701 21499 41735
rect 8493 41633 8527 41667
rect 11253 41633 11287 41667
rect 11529 41633 11563 41667
rect 15209 41633 15243 41667
rect 18705 41633 18739 41667
rect 19901 41633 19935 41667
rect 19993 41633 20027 41667
rect 20821 41633 20855 41667
rect 21005 41633 21039 41667
rect 22109 41633 22143 41667
rect 25145 41633 25179 41667
rect 4537 41565 4571 41599
rect 4997 41565 5031 41599
rect 8217 41565 8251 41599
rect 17693 41565 17727 41599
rect 17969 41565 18003 41599
rect 23765 41565 23799 41599
rect 24041 41565 24075 41599
rect 24961 41565 24995 41599
rect 1685 41497 1719 41531
rect 2145 41497 2179 41531
rect 5457 41497 5491 41531
rect 15485 41497 15519 41531
rect 22293 41497 22327 41531
rect 1777 41429 1811 41463
rect 5917 41429 5951 41463
rect 8309 41429 8343 41463
rect 13001 41429 13035 41463
rect 13277 41429 13311 41463
rect 19441 41429 19475 41463
rect 19809 41429 19843 41463
rect 21097 41429 21131 41463
rect 22385 41429 22419 41463
rect 22753 41429 22787 41463
rect 24593 41429 24627 41463
rect 25053 41429 25087 41463
rect 3985 41225 4019 41259
rect 8309 41225 8343 41259
rect 12449 41225 12483 41259
rect 12817 41225 12851 41259
rect 15393 41225 15427 41259
rect 17325 41225 17359 41259
rect 22753 41225 22787 41259
rect 14841 41157 14875 41191
rect 18705 41157 18739 41191
rect 25237 41157 25271 41191
rect 4077 41089 4111 41123
rect 12081 41089 12115 41123
rect 15117 41089 15151 41123
rect 17233 41089 17267 41123
rect 18429 41089 18463 41123
rect 22385 41089 22419 41123
rect 6561 41021 6595 41055
rect 6837 41021 6871 41055
rect 9413 41021 9447 41055
rect 9689 41021 9723 41055
rect 11897 41021 11931 41055
rect 11989 41021 12023 41055
rect 17417 41021 17451 41055
rect 20545 41021 20579 41055
rect 21465 41021 21499 41055
rect 22201 41021 22235 41055
rect 22293 41021 22327 41055
rect 24685 41021 24719 41055
rect 24961 41021 24995 41055
rect 23213 40953 23247 40987
rect 4445 40885 4479 40919
rect 8585 40885 8619 40919
rect 11161 40885 11195 40919
rect 13369 40885 13403 40919
rect 16865 40885 16899 40919
rect 17877 40885 17911 40919
rect 20177 40885 20211 40919
rect 25421 40885 25455 40919
rect 14197 40681 14231 40715
rect 17417 40681 17451 40715
rect 25145 40681 25179 40715
rect 2973 40613 3007 40647
rect 20821 40613 20855 40647
rect 23949 40613 23983 40647
rect 24501 40613 24535 40647
rect 8125 40545 8159 40579
rect 12081 40545 12115 40579
rect 13093 40545 13127 40579
rect 16037 40545 16071 40579
rect 16129 40545 16163 40579
rect 17141 40545 17175 40579
rect 17969 40545 18003 40579
rect 19533 40545 19567 40579
rect 19717 40545 19751 40579
rect 20545 40545 20579 40579
rect 22937 40545 22971 40579
rect 6377 40477 6411 40511
rect 13185 40477 13219 40511
rect 13277 40477 13311 40511
rect 19809 40477 19843 40511
rect 23397 40477 23431 40511
rect 25329 40477 25363 40511
rect 2789 40409 2823 40443
rect 6653 40409 6687 40443
rect 11345 40409 11379 40443
rect 14381 40409 14415 40443
rect 17785 40409 17819 40443
rect 22661 40409 22695 40443
rect 3341 40341 3375 40375
rect 8401 40341 8435 40375
rect 12541 40341 12575 40375
rect 13645 40341 13679 40375
rect 16221 40341 16255 40375
rect 16589 40341 16623 40375
rect 17877 40341 17911 40375
rect 20177 40341 20211 40375
rect 21189 40341 21223 40375
rect 24225 40341 24259 40375
rect 24869 40341 24903 40375
rect 8125 40137 8159 40171
rect 8493 40137 8527 40171
rect 14841 40137 14875 40171
rect 15577 40137 15611 40171
rect 21005 40137 21039 40171
rect 21465 40137 21499 40171
rect 22385 40137 22419 40171
rect 22753 40137 22787 40171
rect 9045 40069 9079 40103
rect 15669 40069 15703 40103
rect 21097 40069 21131 40103
rect 7389 40001 7423 40035
rect 8033 40001 8067 40035
rect 9873 40001 9907 40035
rect 12173 40001 12207 40035
rect 7849 39933 7883 39967
rect 12449 39933 12483 39967
rect 14381 39933 14415 39967
rect 15853 39933 15887 39967
rect 20821 39933 20855 39967
rect 22201 39933 22235 39967
rect 22293 39933 22327 39967
rect 23765 39933 23799 39967
rect 24041 39933 24075 39967
rect 25053 39933 25087 39967
rect 25329 39933 25363 39967
rect 20361 39865 20395 39899
rect 10241 39797 10275 39831
rect 13921 39797 13955 39831
rect 15209 39797 15243 39831
rect 20177 39797 20211 39831
rect 8401 39593 8435 39627
rect 14289 39593 14323 39627
rect 19533 39593 19567 39627
rect 23581 39593 23615 39627
rect 15761 39525 15795 39559
rect 7757 39457 7791 39491
rect 9229 39457 9263 39491
rect 10425 39457 10459 39491
rect 11897 39457 11931 39491
rect 12173 39457 12207 39491
rect 13185 39457 13219 39491
rect 14841 39457 14875 39491
rect 16405 39457 16439 39491
rect 17601 39457 17635 39491
rect 17693 39457 17727 39491
rect 20177 39457 20211 39491
rect 20913 39457 20947 39491
rect 22477 39457 22511 39491
rect 23029 39457 23063 39491
rect 25145 39457 25179 39491
rect 8677 39389 8711 39423
rect 9505 39389 9539 39423
rect 13093 39389 13127 39423
rect 14749 39389 14783 39423
rect 24041 39389 24075 39423
rect 7941 39321 7975 39355
rect 9413 39321 9447 39355
rect 13001 39321 13035 39355
rect 16221 39321 16255 39355
rect 21097 39321 21131 39355
rect 22293 39321 22327 39355
rect 22385 39321 22419 39355
rect 24961 39321 24995 39355
rect 25053 39321 25087 39355
rect 8033 39253 8067 39287
rect 9873 39253 9907 39287
rect 12633 39253 12667 39287
rect 14657 39253 14691 39287
rect 16129 39253 16163 39287
rect 17785 39253 17819 39287
rect 18153 39253 18187 39287
rect 19901 39253 19935 39287
rect 19993 39253 20027 39287
rect 21005 39253 21039 39287
rect 21465 39253 21499 39287
rect 21925 39253 21959 39287
rect 23857 39253 23891 39287
rect 24593 39253 24627 39287
rect 6009 39049 6043 39083
rect 9781 39049 9815 39083
rect 12541 39049 12575 39083
rect 12909 39049 12943 39083
rect 14105 39049 14139 39083
rect 14473 39049 14507 39083
rect 15761 39049 15795 39083
rect 20177 39049 20211 39083
rect 21097 39049 21131 39083
rect 23489 39049 23523 39083
rect 6377 38981 6411 39015
rect 10149 38981 10183 39015
rect 20269 38981 20303 39015
rect 22477 38981 22511 39015
rect 24961 38981 24995 39015
rect 1593 38913 1627 38947
rect 2053 38913 2087 38947
rect 12173 38913 12207 38947
rect 15853 38913 15887 38947
rect 21005 38913 21039 38947
rect 22385 38913 22419 38947
rect 4261 38845 4295 38879
rect 4537 38845 4571 38879
rect 8585 38845 8619 38879
rect 10241 38845 10275 38879
rect 10425 38845 10459 38879
rect 10977 38845 11011 38879
rect 11897 38845 11931 38879
rect 12081 38845 12115 38879
rect 13921 38845 13955 38879
rect 14013 38845 14047 38879
rect 15577 38845 15611 38879
rect 19441 38845 19475 38879
rect 19993 38845 20027 38879
rect 21557 38845 21591 38879
rect 22569 38845 22603 38879
rect 25237 38845 25271 38879
rect 17693 38777 17727 38811
rect 1777 38709 1811 38743
rect 13369 38709 13403 38743
rect 15209 38709 15243 38743
rect 16221 38709 16255 38743
rect 19177 38709 19211 38743
rect 20637 38709 20671 38743
rect 22017 38709 22051 38743
rect 23029 38709 23063 38743
rect 4905 38505 4939 38539
rect 8585 38505 8619 38539
rect 9505 38505 9539 38539
rect 11437 38505 11471 38539
rect 16405 38505 16439 38539
rect 16865 38505 16899 38539
rect 20177 38505 20211 38539
rect 11989 38437 12023 38471
rect 6653 38369 6687 38403
rect 8033 38369 8067 38403
rect 9965 38369 9999 38403
rect 10149 38369 10183 38403
rect 10885 38369 10919 38403
rect 12541 38369 12575 38403
rect 15117 38369 15151 38403
rect 15853 38369 15887 38403
rect 17417 38369 17451 38403
rect 19625 38369 19659 38403
rect 23213 38369 23247 38403
rect 23305 38369 23339 38403
rect 7573 38301 7607 38335
rect 8125 38301 8159 38335
rect 8217 38301 8251 38335
rect 11069 38301 11103 38335
rect 14841 38301 14875 38335
rect 19717 38301 19751 38335
rect 22293 38301 22327 38335
rect 24869 38301 24903 38335
rect 25329 38301 25363 38335
rect 6377 38233 6411 38267
rect 14105 38233 14139 38267
rect 14933 38233 14967 38267
rect 15945 38233 15979 38267
rect 17325 38233 17359 38267
rect 21465 38233 21499 38267
rect 6929 38165 6963 38199
rect 9873 38165 9907 38199
rect 10977 38165 11011 38199
rect 12357 38165 12391 38199
rect 12449 38165 12483 38199
rect 14473 38165 14507 38199
rect 16037 38165 16071 38199
rect 17233 38165 17267 38199
rect 18889 38165 18923 38199
rect 19809 38165 19843 38199
rect 21097 38165 21131 38199
rect 22661 38165 22695 38199
rect 23397 38165 23431 38199
rect 23765 38165 23799 38199
rect 24501 38165 24535 38199
rect 24685 38165 24719 38199
rect 25145 38165 25179 38199
rect 10885 37961 10919 37995
rect 12265 37961 12299 37995
rect 13185 37961 13219 37995
rect 13645 37961 13679 37995
rect 15393 37961 15427 37995
rect 16129 37961 16163 37995
rect 22017 37961 22051 37995
rect 22385 37961 22419 37995
rect 9413 37893 9447 37927
rect 20637 37893 20671 37927
rect 22477 37893 22511 37927
rect 9689 37825 9723 37859
rect 10517 37825 10551 37859
rect 13277 37825 13311 37859
rect 14105 37825 14139 37859
rect 15301 37825 15335 37859
rect 16681 37825 16715 37859
rect 17049 37825 17083 37859
rect 20545 37825 20579 37859
rect 23213 37825 23247 37859
rect 7665 37757 7699 37791
rect 10241 37757 10275 37791
rect 10425 37757 10459 37791
rect 13001 37757 13035 37791
rect 15485 37757 15519 37791
rect 17325 37757 17359 37791
rect 18797 37757 18831 37791
rect 19441 37757 19475 37791
rect 20453 37757 20487 37791
rect 22661 37757 22695 37791
rect 21005 37689 21039 37723
rect 25421 37689 25455 37723
rect 11161 37621 11195 37655
rect 11529 37621 11563 37655
rect 14933 37621 14967 37655
rect 19073 37621 19107 37655
rect 19901 37621 19935 37655
rect 23476 37621 23510 37655
rect 24961 37621 24995 37655
rect 25329 37621 25363 37655
rect 8953 37417 8987 37451
rect 9321 37417 9355 37451
rect 12817 37417 12851 37451
rect 9413 37349 9447 37383
rect 5549 37281 5583 37315
rect 8309 37281 8343 37315
rect 10425 37281 10459 37315
rect 10885 37281 10919 37315
rect 11897 37281 11931 37315
rect 12449 37281 12483 37315
rect 15577 37281 15611 37315
rect 16681 37281 16715 37315
rect 17785 37281 17819 37315
rect 18337 37281 18371 37315
rect 18429 37281 18463 37315
rect 21465 37281 21499 37315
rect 23581 37281 23615 37315
rect 24685 37281 24719 37315
rect 5273 37213 5307 37247
rect 8125 37213 8159 37247
rect 10241 37213 10275 37247
rect 11713 37213 11747 37247
rect 16865 37213 16899 37247
rect 19533 37213 19567 37247
rect 24041 37213 24075 37247
rect 25329 37213 25363 37247
rect 7297 37145 7331 37179
rect 8217 37145 8251 37179
rect 10149 37145 10183 37179
rect 11805 37145 11839 37179
rect 15393 37145 15427 37179
rect 18521 37145 18555 37179
rect 20361 37145 20395 37179
rect 21741 37145 21775 37179
rect 24501 37145 24535 37179
rect 7757 37077 7791 37111
rect 9781 37077 9815 37111
rect 11345 37077 11379 37111
rect 15025 37077 15059 37111
rect 15485 37077 15519 37111
rect 16037 37077 16071 37111
rect 16773 37077 16807 37111
rect 17233 37077 17267 37111
rect 18889 37077 18923 37111
rect 23213 37077 23247 37111
rect 23857 37077 23891 37111
rect 25145 37077 25179 37111
rect 5181 36873 5215 36907
rect 5641 36873 5675 36907
rect 9321 36873 9355 36907
rect 9781 36873 9815 36907
rect 10977 36873 11011 36907
rect 12081 36873 12115 36907
rect 12173 36873 12207 36907
rect 13001 36873 13035 36907
rect 13461 36873 13495 36907
rect 15301 36873 15335 36907
rect 15761 36873 15795 36907
rect 18429 36873 18463 36907
rect 19717 36873 19751 36907
rect 20177 36873 20211 36907
rect 13369 36805 13403 36839
rect 16313 36805 16347 36839
rect 23029 36805 23063 36839
rect 1593 36737 1627 36771
rect 2053 36737 2087 36771
rect 5549 36737 5583 36771
rect 10149 36737 10183 36771
rect 10241 36737 10275 36771
rect 14841 36737 14875 36771
rect 15669 36737 15703 36771
rect 20085 36737 20119 36771
rect 22753 36737 22787 36771
rect 25329 36737 25363 36771
rect 5733 36669 5767 36703
rect 7573 36669 7607 36703
rect 7849 36669 7883 36703
rect 10333 36669 10367 36703
rect 12265 36669 12299 36703
rect 13553 36669 13587 36703
rect 15853 36669 15887 36703
rect 16865 36669 16899 36703
rect 18245 36669 18279 36703
rect 18337 36669 18371 36703
rect 20269 36669 20303 36703
rect 19349 36601 19383 36635
rect 25145 36601 25179 36635
rect 1777 36533 1811 36567
rect 11713 36533 11747 36567
rect 18797 36533 18831 36567
rect 19165 36533 19199 36567
rect 24501 36533 24535 36567
rect 6101 36329 6135 36363
rect 8217 36329 8251 36363
rect 15393 36329 15427 36363
rect 16681 36329 16715 36363
rect 19625 36329 19659 36363
rect 22201 36329 22235 36363
rect 15577 36261 15611 36295
rect 17141 36261 17175 36295
rect 20729 36261 20763 36295
rect 7849 36193 7883 36227
rect 9229 36193 9263 36227
rect 10517 36193 10551 36227
rect 14933 36193 14967 36227
rect 16037 36193 16071 36227
rect 17693 36193 17727 36227
rect 20177 36193 20211 36227
rect 21557 36193 21591 36227
rect 23489 36193 23523 36227
rect 23581 36193 23615 36227
rect 8769 36125 8803 36159
rect 10057 36125 10091 36159
rect 12173 36125 12207 36159
rect 12449 36125 12483 36159
rect 16221 36125 16255 36159
rect 16313 36125 16347 36159
rect 17601 36125 17635 36159
rect 20361 36125 20395 36159
rect 22477 36125 22511 36159
rect 24869 36125 24903 36159
rect 25329 36125 25363 36159
rect 7573 36057 7607 36091
rect 11345 36057 11379 36091
rect 17509 36057 17543 36091
rect 14289 35989 14323 36023
rect 14657 35989 14691 36023
rect 14749 35989 14783 36023
rect 20269 35989 20303 36023
rect 21005 35989 21039 36023
rect 21741 35989 21775 36023
rect 21833 35989 21867 36023
rect 22661 35989 22695 36023
rect 23673 35989 23707 36023
rect 24041 35989 24075 36023
rect 25145 35989 25179 36023
rect 6009 35785 6043 35819
rect 9413 35785 9447 35819
rect 14197 35785 14231 35819
rect 15577 35785 15611 35819
rect 16865 35785 16899 35819
rect 17233 35785 17267 35819
rect 6469 35717 6503 35751
rect 12173 35717 12207 35751
rect 15669 35717 15703 35751
rect 18981 35717 19015 35751
rect 17325 35649 17359 35683
rect 18705 35649 18739 35683
rect 25329 35649 25363 35683
rect 4261 35581 4295 35615
rect 4537 35581 4571 35615
rect 10885 35581 10919 35615
rect 11161 35581 11195 35615
rect 11897 35581 11931 35615
rect 13645 35581 13679 35615
rect 14749 35581 14783 35615
rect 15761 35581 15795 35615
rect 17417 35581 17451 35615
rect 23581 35581 23615 35615
rect 25053 35581 25087 35615
rect 15209 35513 15243 35547
rect 20729 35513 20763 35547
rect 11529 35445 11563 35479
rect 13921 35445 13955 35479
rect 20453 35445 20487 35479
rect 5273 35241 5307 35275
rect 7665 35241 7699 35275
rect 10333 35241 10367 35275
rect 13479 35241 13513 35275
rect 14473 35241 14507 35275
rect 15577 35241 15611 35275
rect 23489 35241 23523 35275
rect 18153 35173 18187 35207
rect 8217 35105 8251 35139
rect 9689 35105 9723 35139
rect 11989 35105 12023 35139
rect 15025 35105 15059 35139
rect 18705 35105 18739 35139
rect 20545 35105 20579 35139
rect 21741 35105 21775 35139
rect 21833 35105 21867 35139
rect 22937 35105 22971 35139
rect 7021 35037 7055 35071
rect 9965 35037 9999 35071
rect 13737 35037 13771 35071
rect 15209 35037 15243 35071
rect 18521 35037 18555 35071
rect 24869 35037 24903 35071
rect 25329 35037 25363 35071
rect 6745 34969 6779 35003
rect 14105 34969 14139 35003
rect 15117 34969 15151 35003
rect 20361 34969 20395 35003
rect 23029 34969 23063 35003
rect 7297 34901 7331 34935
rect 8033 34901 8067 34935
rect 8125 34901 8159 34935
rect 9873 34901 9907 34935
rect 18613 34901 18647 34935
rect 19993 34901 20027 34935
rect 20453 34901 20487 34935
rect 21925 34901 21959 34935
rect 22293 34901 22327 34935
rect 23121 34901 23155 34935
rect 24685 34901 24719 34935
rect 25145 34901 25179 34935
rect 1777 34697 1811 34731
rect 3525 34697 3559 34731
rect 5641 34697 5675 34731
rect 9045 34697 9079 34731
rect 9413 34697 9447 34731
rect 14105 34697 14139 34731
rect 14473 34697 14507 34731
rect 19441 34697 19475 34731
rect 22385 34697 22419 34731
rect 22477 34697 22511 34731
rect 23213 34697 23247 34731
rect 7021 34629 7055 34663
rect 13829 34629 13863 34663
rect 14565 34629 14599 34663
rect 1593 34561 1627 34595
rect 2053 34561 2087 34595
rect 9505 34561 9539 34595
rect 13461 34561 13495 34595
rect 18613 34561 18647 34595
rect 25329 34561 25363 34595
rect 5273 34493 5307 34527
rect 6745 34493 6779 34527
rect 9689 34493 9723 34527
rect 13185 34493 13219 34527
rect 14657 34493 14691 34527
rect 16865 34493 16899 34527
rect 18337 34493 18371 34527
rect 19533 34493 19567 34527
rect 19625 34493 19659 34527
rect 20269 34493 20303 34527
rect 22569 34493 22603 34527
rect 8493 34425 8527 34459
rect 25145 34425 25179 34459
rect 5009 34357 5043 34391
rect 11713 34357 11747 34391
rect 19073 34357 19107 34391
rect 22017 34357 22051 34391
rect 7021 34153 7055 34187
rect 8677 34153 8711 34187
rect 9137 34153 9171 34187
rect 12265 34153 12299 34187
rect 20177 34153 20211 34187
rect 4905 34017 4939 34051
rect 9597 34017 9631 34051
rect 9689 34017 9723 34051
rect 12817 34017 12851 34051
rect 19625 34017 19659 34051
rect 20821 34017 20855 34051
rect 6653 33949 6687 33983
rect 12725 33949 12759 33983
rect 19809 33949 19843 33983
rect 23581 33949 23615 33983
rect 24593 33949 24627 33983
rect 6377 33881 6411 33915
rect 12633 33881 12667 33915
rect 21097 33881 21131 33915
rect 22937 33881 22971 33915
rect 25421 33881 25455 33915
rect 9505 33813 9539 33847
rect 13645 33813 13679 33847
rect 18797 33813 18831 33847
rect 18981 33813 19015 33847
rect 19717 33813 19751 33847
rect 22569 33813 22603 33847
rect 23765 33813 23799 33847
rect 24777 33813 24811 33847
rect 25329 33813 25363 33847
rect 9505 33609 9539 33643
rect 9965 33609 9999 33643
rect 11897 33609 11931 33643
rect 13921 33609 13955 33643
rect 14933 33609 14967 33643
rect 18613 33609 18647 33643
rect 22385 33609 22419 33643
rect 25237 33609 25271 33643
rect 10333 33541 10367 33575
rect 12265 33473 12299 33507
rect 13829 33473 13863 33507
rect 15025 33473 15059 33507
rect 23489 33473 23523 33507
rect 7757 33405 7791 33439
rect 8033 33405 8067 33439
rect 10425 33405 10459 33439
rect 10609 33405 10643 33439
rect 11621 33405 11655 33439
rect 12357 33405 12391 33439
rect 12541 33405 12575 33439
rect 14013 33405 14047 33439
rect 14749 33405 14783 33439
rect 18705 33405 18739 33439
rect 18797 33405 18831 33439
rect 23765 33405 23799 33439
rect 18245 33337 18279 33371
rect 11253 33269 11287 33303
rect 13461 33269 13495 33303
rect 15393 33269 15427 33303
rect 7297 33065 7331 33099
rect 9873 33065 9907 33099
rect 13645 33065 13679 33099
rect 18613 33065 18647 33099
rect 19717 33065 19751 33099
rect 11713 32997 11747 33031
rect 20453 32997 20487 33031
rect 5549 32929 5583 32963
rect 9229 32929 9263 32963
rect 12173 32929 12207 32963
rect 12265 32929 12299 32963
rect 13093 32929 13127 32963
rect 16865 32929 16899 32963
rect 22201 32929 22235 32963
rect 23213 32929 23247 32963
rect 13185 32861 13219 32895
rect 19533 32861 19567 32895
rect 23029 32861 23063 32895
rect 24869 32861 24903 32895
rect 25329 32861 25363 32895
rect 5825 32793 5859 32827
rect 7665 32793 7699 32827
rect 9413 32793 9447 32827
rect 12081 32793 12115 32827
rect 17141 32793 17175 32827
rect 21925 32793 21959 32827
rect 9505 32725 9539 32759
rect 10149 32725 10183 32759
rect 13277 32725 13311 32759
rect 14289 32725 14323 32759
rect 16313 32725 16347 32759
rect 18889 32725 18923 32759
rect 22661 32725 22695 32759
rect 23121 32725 23155 32759
rect 25145 32725 25179 32759
rect 7113 32521 7147 32555
rect 8677 32521 8711 32555
rect 11253 32521 11287 32555
rect 12725 32521 12759 32555
rect 13369 32521 13403 32555
rect 18061 32521 18095 32555
rect 18429 32521 18463 32555
rect 19625 32521 19659 32555
rect 21005 32521 21039 32555
rect 21097 32521 21131 32555
rect 22661 32521 22695 32555
rect 17233 32453 17267 32487
rect 18521 32453 18555 32487
rect 1593 32385 1627 32419
rect 2053 32385 2087 32419
rect 16221 32385 16255 32419
rect 19717 32385 19751 32419
rect 22017 32385 22051 32419
rect 23029 32385 23063 32419
rect 23857 32385 23891 32419
rect 24869 32385 24903 32419
rect 25329 32385 25363 32419
rect 4997 32317 5031 32351
rect 7481 32317 7515 32351
rect 9137 32317 9171 32351
rect 9413 32317 9447 32351
rect 15945 32317 15979 32351
rect 17049 32317 17083 32351
rect 17141 32317 17175 32351
rect 18613 32317 18647 32351
rect 19809 32317 19843 32351
rect 21189 32317 21223 32351
rect 23121 32317 23155 32351
rect 23213 32317 23247 32351
rect 19257 32249 19291 32283
rect 25145 32249 25179 32283
rect 1777 32181 1811 32215
rect 10885 32181 10919 32215
rect 14473 32181 14507 32215
rect 17601 32181 17635 32215
rect 20637 32181 20671 32215
rect 22201 32181 22235 32215
rect 24041 32181 24075 32215
rect 5181 31977 5215 32011
rect 11253 31977 11287 32011
rect 12357 31977 12391 32011
rect 15209 31977 15243 32011
rect 17693 31977 17727 32011
rect 20269 31977 20303 32011
rect 25145 31977 25179 32011
rect 8217 31909 8251 31943
rect 21465 31909 21499 31943
rect 22661 31909 22695 31943
rect 23857 31909 23891 31943
rect 6653 31841 6687 31875
rect 7665 31841 7699 31875
rect 9137 31841 9171 31875
rect 12909 31841 12943 31875
rect 16957 31841 16991 31875
rect 17417 31841 17451 31875
rect 19717 31841 19751 31875
rect 19809 31841 19843 31875
rect 20821 31841 20855 31875
rect 22017 31841 22051 31875
rect 23121 31841 23155 31875
rect 6929 31773 6963 31807
rect 7757 31773 7791 31807
rect 10885 31773 10919 31807
rect 12081 31773 12115 31807
rect 12817 31773 12851 31807
rect 22201 31773 22235 31807
rect 23581 31773 23615 31807
rect 24869 31773 24903 31807
rect 25329 31773 25363 31807
rect 10609 31705 10643 31739
rect 12725 31705 12759 31739
rect 16681 31705 16715 31739
rect 17325 31705 17359 31739
rect 22293 31705 22327 31739
rect 7849 31637 7883 31671
rect 18981 31637 19015 31671
rect 19901 31637 19935 31671
rect 21005 31637 21039 31671
rect 21097 31637 21131 31671
rect 4905 31433 4939 31467
rect 5273 31433 5307 31467
rect 7757 31433 7791 31467
rect 8217 31433 8251 31467
rect 10149 31433 10183 31467
rect 17693 31433 17727 31467
rect 20453 31433 20487 31467
rect 24225 31433 24259 31467
rect 6745 31297 6779 31331
rect 7297 31297 7331 31331
rect 7389 31297 7423 31331
rect 8861 31297 8895 31331
rect 10517 31297 10551 31331
rect 12541 31297 12575 31331
rect 17601 31297 17635 31331
rect 19441 31297 19475 31331
rect 22017 31297 22051 31331
rect 23397 31297 23431 31331
rect 25329 31297 25363 31331
rect 4721 31229 4755 31263
rect 4813 31229 4847 31263
rect 7205 31229 7239 31263
rect 9873 31229 9907 31263
rect 10609 31229 10643 31263
rect 10793 31229 10827 31263
rect 17785 31229 17819 31263
rect 25053 31229 25087 31263
rect 4261 31161 4295 31195
rect 19625 31161 19659 31195
rect 22477 31161 22511 31195
rect 23581 31161 23615 31195
rect 9689 31093 9723 31127
rect 12909 31093 12943 31127
rect 17233 31093 17267 31127
rect 21557 31093 21591 31127
rect 22201 31093 22235 31127
rect 7849 30889 7883 30923
rect 13001 30889 13035 30923
rect 25237 30889 25271 30923
rect 25421 30889 25455 30923
rect 7297 30753 7331 30787
rect 10701 30753 10735 30787
rect 13553 30753 13587 30787
rect 16681 30753 16715 30787
rect 18153 30753 18187 30787
rect 18337 30753 18371 30787
rect 21005 30753 21039 30787
rect 22293 30753 22327 30787
rect 7481 30685 7515 30719
rect 14289 30685 14323 30719
rect 18061 30685 18095 30719
rect 19625 30685 19659 30719
rect 20913 30685 20947 30719
rect 24593 30685 24627 30719
rect 10977 30617 11011 30651
rect 13369 30617 13403 30651
rect 14565 30617 14599 30651
rect 16773 30617 16807 30651
rect 22569 30617 22603 30651
rect 6837 30549 6871 30583
rect 7389 30549 7423 30583
rect 12449 30549 12483 30583
rect 13461 30549 13495 30583
rect 16037 30549 16071 30583
rect 16865 30549 16899 30583
rect 17233 30549 17267 30583
rect 17693 30549 17727 30583
rect 18797 30549 18831 30583
rect 19441 30549 19475 30583
rect 20453 30549 20487 30583
rect 20821 30549 20855 30583
rect 24041 30549 24075 30583
rect 24777 30549 24811 30583
rect 7665 30345 7699 30379
rect 15301 30345 15335 30379
rect 16129 30345 16163 30379
rect 17325 30345 17359 30379
rect 17693 30345 17727 30379
rect 20085 30345 20119 30379
rect 12265 30277 12299 30311
rect 13001 30277 13035 30311
rect 18981 30277 19015 30311
rect 22293 30277 22327 30311
rect 22385 30277 22419 30311
rect 9413 30209 9447 30243
rect 9781 30209 9815 30243
rect 13093 30209 13127 30243
rect 15209 30209 15243 30243
rect 16681 30209 16715 30243
rect 17785 30209 17819 30243
rect 18889 30209 18923 30243
rect 9137 30141 9171 30175
rect 11713 30141 11747 30175
rect 13277 30141 13311 30175
rect 15393 30141 15427 30175
rect 17877 30141 17911 30175
rect 19073 30141 19107 30175
rect 19901 30141 19935 30175
rect 19993 30141 20027 30175
rect 22201 30141 22235 30175
rect 23489 30141 23523 30175
rect 24961 30141 24995 30175
rect 25237 30141 25271 30175
rect 12633 30073 12667 30107
rect 18521 30073 18555 30107
rect 14841 30005 14875 30039
rect 15945 30005 15979 30039
rect 16313 30005 16347 30039
rect 20453 30005 20487 30039
rect 22753 30005 22787 30039
rect 8493 29801 8527 29835
rect 9137 29801 9171 29835
rect 25145 29801 25179 29835
rect 11345 29733 11379 29767
rect 17877 29733 17911 29767
rect 2053 29665 2087 29699
rect 3985 29665 4019 29699
rect 9689 29665 9723 29699
rect 10701 29665 10735 29699
rect 12357 29665 12391 29699
rect 13093 29665 13127 29699
rect 13277 29665 13311 29699
rect 17325 29665 17359 29699
rect 18245 29665 18279 29699
rect 19901 29665 19935 29699
rect 19993 29665 20027 29699
rect 21373 29665 21407 29699
rect 22109 29665 22143 29699
rect 22293 29665 22327 29699
rect 23305 29665 23339 29699
rect 23489 29665 23523 29699
rect 1777 29597 1811 29631
rect 9505 29597 9539 29631
rect 10977 29597 11011 29631
rect 13369 29597 13403 29631
rect 17417 29597 17451 29631
rect 19809 29597 19843 29631
rect 21281 29597 21315 29631
rect 22385 29597 22419 29631
rect 25329 29597 25363 29631
rect 4169 29529 4203 29563
rect 5825 29529 5859 29563
rect 8769 29529 8803 29563
rect 9597 29529 9631 29563
rect 16773 29529 16807 29563
rect 17509 29529 17543 29563
rect 21189 29529 21223 29563
rect 10241 29461 10275 29495
rect 10885 29461 10919 29495
rect 11805 29461 11839 29495
rect 12173 29461 12207 29495
rect 12265 29461 12299 29495
rect 13737 29461 13771 29495
rect 19441 29461 19475 29495
rect 20821 29461 20855 29495
rect 22753 29461 22787 29495
rect 23581 29461 23615 29495
rect 23949 29461 23983 29495
rect 8217 29257 8251 29291
rect 13093 29257 13127 29291
rect 19809 29257 19843 29291
rect 25421 29257 25455 29291
rect 12265 29189 12299 29223
rect 13369 29189 13403 29223
rect 24777 29189 24811 29223
rect 10241 29121 10275 29155
rect 12173 29121 12207 29155
rect 16313 29121 16347 29155
rect 19533 29121 19567 29155
rect 23673 29121 23707 29155
rect 24133 29121 24167 29155
rect 9965 29053 9999 29087
rect 12357 29053 12391 29087
rect 13277 29053 13311 29087
rect 19257 29053 19291 29087
rect 22201 29053 22235 29087
rect 11805 28985 11839 29019
rect 12909 28985 12943 29019
rect 15025 28985 15059 29019
rect 16773 28985 16807 29019
rect 23949 28985 23983 29019
rect 24593 28985 24627 29019
rect 9707 28917 9741 28951
rect 17785 28917 17819 28951
rect 8493 28713 8527 28747
rect 9873 28713 9907 28747
rect 13461 28713 13495 28747
rect 16313 28713 16347 28747
rect 22569 28713 22603 28747
rect 25145 28713 25179 28747
rect 8401 28645 8435 28679
rect 23857 28645 23891 28679
rect 3985 28577 4019 28611
rect 8033 28577 8067 28611
rect 9321 28577 9355 28611
rect 11253 28577 11287 28611
rect 11529 28577 11563 28611
rect 13001 28577 13035 28611
rect 14565 28577 14599 28611
rect 14841 28577 14875 28611
rect 17601 28577 17635 28611
rect 19533 28577 19567 28611
rect 20821 28577 20855 28611
rect 22017 28577 22051 28611
rect 24501 28577 24535 28611
rect 8769 28509 8803 28543
rect 9413 28509 9447 28543
rect 19717 28509 19751 28543
rect 19809 28509 19843 28543
rect 22201 28509 22235 28543
rect 24041 28509 24075 28543
rect 25329 28509 25363 28543
rect 4169 28441 4203 28475
rect 5825 28441 5859 28475
rect 7757 28441 7791 28475
rect 17417 28441 17451 28475
rect 18245 28441 18279 28475
rect 21005 28441 21039 28475
rect 22109 28441 22143 28475
rect 22845 28441 22879 28475
rect 6285 28373 6319 28407
rect 9505 28373 9539 28407
rect 13369 28373 13403 28407
rect 16589 28373 16623 28407
rect 17049 28373 17083 28407
rect 17509 28373 17543 28407
rect 18705 28373 18739 28407
rect 20177 28373 20211 28407
rect 20913 28373 20947 28407
rect 21373 28373 21407 28407
rect 24685 28373 24719 28407
rect 8585 28169 8619 28203
rect 9229 28169 9263 28203
rect 11345 28169 11379 28203
rect 14657 28169 14691 28203
rect 15393 28169 15427 28203
rect 16865 28169 16899 28203
rect 17325 28169 17359 28203
rect 18061 28169 18095 28203
rect 18521 28169 18555 28203
rect 22293 28169 22327 28203
rect 22385 28169 22419 28203
rect 22753 28169 22787 28203
rect 25421 28169 25455 28203
rect 12265 28101 12299 28135
rect 17233 28101 17267 28135
rect 21465 28101 21499 28135
rect 24777 28101 24811 28135
rect 6561 28033 6595 28067
rect 10977 28033 11011 28067
rect 13737 28033 13771 28067
rect 18429 28033 18463 28067
rect 19257 28033 19291 28067
rect 20453 28033 20487 28067
rect 23489 28033 23523 28067
rect 23949 28033 23983 28067
rect 6837 27965 6871 27999
rect 8309 27965 8343 27999
rect 10701 27965 10735 27999
rect 12357 27965 12391 27999
rect 12449 27965 12483 27999
rect 13185 27965 13219 27999
rect 14013 27965 14047 27999
rect 14749 27965 14783 27999
rect 14841 27965 14875 27999
rect 17417 27965 17451 27999
rect 18705 27965 18739 27999
rect 22201 27965 22235 27999
rect 19441 27897 19475 27931
rect 23305 27897 23339 27931
rect 24593 27897 24627 27931
rect 11897 27829 11931 27863
rect 14289 27829 14323 27863
rect 24133 27829 24167 27863
rect 19441 27625 19475 27659
rect 20931 27625 20965 27659
rect 8401 27557 8435 27591
rect 24041 27557 24075 27591
rect 2053 27489 2087 27523
rect 3985 27489 4019 27523
rect 5825 27489 5859 27523
rect 8033 27489 8067 27523
rect 12909 27489 12943 27523
rect 14841 27489 14875 27523
rect 16221 27489 16255 27523
rect 17325 27489 17359 27523
rect 18153 27489 18187 27523
rect 18245 27489 18279 27523
rect 19073 27489 19107 27523
rect 21557 27489 21591 27523
rect 1777 27421 1811 27455
rect 13093 27421 13127 27455
rect 14749 27421 14783 27455
rect 17141 27421 17175 27455
rect 21189 27421 21223 27455
rect 22293 27421 22327 27455
rect 24777 27421 24811 27455
rect 4169 27353 4203 27387
rect 7757 27353 7791 27387
rect 14657 27353 14691 27387
rect 22569 27353 22603 27387
rect 24593 27353 24627 27387
rect 6285 27285 6319 27319
rect 10701 27285 10735 27319
rect 12357 27285 12391 27319
rect 13001 27285 13035 27319
rect 13461 27285 13495 27319
rect 14289 27285 14323 27319
rect 15577 27285 15611 27319
rect 15945 27285 15979 27319
rect 16037 27285 16071 27319
rect 16773 27285 16807 27319
rect 17233 27285 17267 27319
rect 18337 27285 18371 27319
rect 18705 27285 18739 27319
rect 2053 27081 2087 27115
rect 3479 27081 3513 27115
rect 10333 27081 10367 27115
rect 15761 27081 15795 27115
rect 18429 27081 18463 27115
rect 18705 27081 18739 27115
rect 25421 27081 25455 27115
rect 13829 27013 13863 27047
rect 15117 27013 15151 27047
rect 17049 27013 17083 27047
rect 17785 27013 17819 27047
rect 24777 27013 24811 27047
rect 2237 26945 2271 26979
rect 3376 26945 3410 26979
rect 7849 26945 7883 26979
rect 7941 26945 7975 26979
rect 10425 26945 10459 26979
rect 13461 26945 13495 26979
rect 15025 26945 15059 26979
rect 16405 26945 16439 26979
rect 17693 26945 17727 26979
rect 23949 26945 23983 26979
rect 7757 26877 7791 26911
rect 8769 26877 8803 26911
rect 10149 26877 10183 26911
rect 11713 26877 11747 26911
rect 13185 26877 13219 26911
rect 15209 26877 15243 26911
rect 17601 26877 17635 26911
rect 22201 26877 22235 26911
rect 23673 26877 23707 26911
rect 24593 26809 24627 26843
rect 7205 26741 7239 26775
rect 8309 26741 8343 26775
rect 10793 26741 10827 26775
rect 14657 26741 14691 26775
rect 15853 26741 15887 26775
rect 16681 26741 16715 26775
rect 18153 26741 18187 26775
rect 24225 26741 24259 26775
rect 25145 26741 25179 26775
rect 8033 26537 8067 26571
rect 8401 26537 8435 26571
rect 16313 26537 16347 26571
rect 20545 26537 20579 26571
rect 23213 26537 23247 26571
rect 10977 26469 11011 26503
rect 13553 26469 13587 26503
rect 18153 26469 18187 26503
rect 23857 26469 23891 26503
rect 25145 26469 25179 26503
rect 3985 26401 4019 26435
rect 5825 26401 5859 26435
rect 6285 26401 6319 26435
rect 6561 26401 6595 26435
rect 10425 26401 10459 26435
rect 12909 26401 12943 26435
rect 17601 26401 17635 26435
rect 19993 26401 20027 26435
rect 9137 26333 9171 26367
rect 9689 26333 9723 26367
rect 10609 26333 10643 26367
rect 13185 26333 13219 26367
rect 14565 26333 14599 26367
rect 16589 26333 16623 26367
rect 17693 26333 17727 26367
rect 21465 26333 21499 26367
rect 24041 26333 24075 26367
rect 24685 26333 24719 26367
rect 4169 26265 4203 26299
rect 9505 26265 9539 26299
rect 10517 26265 10551 26299
rect 13093 26265 13127 26299
rect 14841 26265 14875 26299
rect 17141 26265 17175 26299
rect 17785 26265 17819 26299
rect 19441 26265 19475 26299
rect 20085 26265 20119 26299
rect 20177 26265 20211 26299
rect 21741 26265 21775 26299
rect 24869 26265 24903 26299
rect 2605 25993 2639 26027
rect 3847 25993 3881 26027
rect 7849 25993 7883 26027
rect 8677 25993 8711 26027
rect 10333 25993 10367 26027
rect 13921 25993 13955 26027
rect 19717 25993 19751 26027
rect 22385 25993 22419 26027
rect 10241 25925 10275 25959
rect 19625 25925 19659 25959
rect 22477 25925 22511 25959
rect 23121 25925 23155 25959
rect 23581 25925 23615 25959
rect 24317 25925 24351 25959
rect 25053 25925 25087 25959
rect 3744 25857 3778 25891
rect 13553 25857 13587 25891
rect 21005 25857 21039 25891
rect 21465 25857 21499 25891
rect 25421 25857 25455 25891
rect 3065 25789 3099 25823
rect 3249 25789 3283 25823
rect 7573 25789 7607 25823
rect 7757 25789 7791 25823
rect 10057 25789 10091 25823
rect 13277 25789 13311 25823
rect 16957 25789 16991 25823
rect 17233 25789 17267 25823
rect 18705 25789 18739 25823
rect 19901 25789 19935 25823
rect 20453 25789 20487 25823
rect 22569 25789 22603 25823
rect 23397 25789 23431 25823
rect 8217 25721 8251 25755
rect 21281 25721 21315 25755
rect 24133 25721 24167 25755
rect 24869 25721 24903 25755
rect 7113 25653 7147 25687
rect 10701 25653 10735 25687
rect 11805 25653 11839 25687
rect 16129 25653 16163 25687
rect 19257 25653 19291 25687
rect 22017 25653 22051 25687
rect 3617 25449 3651 25483
rect 4169 25449 4203 25483
rect 18153 25449 18187 25483
rect 8401 25381 8435 25415
rect 18889 25381 18923 25415
rect 23397 25381 23431 25415
rect 2053 25313 2087 25347
rect 3985 25313 4019 25347
rect 6377 25313 6411 25347
rect 6653 25313 6687 25347
rect 15577 25313 15611 25347
rect 15669 25313 15703 25347
rect 16773 25313 16807 25347
rect 16957 25313 16991 25347
rect 20453 25313 20487 25347
rect 22753 25313 22787 25347
rect 22937 25313 22971 25347
rect 1777 25245 1811 25279
rect 4445 25245 4479 25279
rect 15485 25245 15519 25279
rect 17969 25245 18003 25279
rect 24777 25245 24811 25279
rect 16681 25177 16715 25211
rect 20729 25177 20763 25211
rect 23029 25177 23063 25211
rect 23857 25177 23891 25211
rect 25053 25177 25087 25211
rect 8125 25109 8159 25143
rect 9137 25109 9171 25143
rect 12633 25109 12667 25143
rect 15117 25109 15151 25143
rect 16313 25109 16347 25143
rect 22201 25109 22235 25143
rect 24593 25109 24627 25143
rect 12541 24905 12575 24939
rect 18337 24905 18371 24939
rect 19625 24905 19659 24939
rect 22385 24905 22419 24939
rect 12449 24837 12483 24871
rect 2237 24769 2271 24803
rect 4813 24769 4847 24803
rect 7941 24769 7975 24803
rect 9965 24769 9999 24803
rect 10701 24769 10735 24803
rect 10793 24769 10827 24803
rect 11897 24769 11931 24803
rect 16681 24769 16715 24803
rect 18429 24769 18463 24803
rect 19533 24769 19567 24803
rect 22293 24769 22327 24803
rect 25237 24769 25271 24803
rect 3065 24701 3099 24735
rect 4537 24701 4571 24735
rect 7481 24701 7515 24735
rect 8217 24701 8251 24735
rect 10517 24701 10551 24735
rect 12357 24701 12391 24735
rect 14565 24701 14599 24735
rect 14841 24701 14875 24735
rect 16313 24701 16347 24735
rect 18613 24701 18647 24735
rect 19349 24701 19383 24735
rect 22109 24701 22143 24735
rect 23213 24701 23247 24735
rect 23489 24701 23523 24735
rect 24961 24701 24995 24735
rect 2053 24633 2087 24667
rect 9689 24633 9723 24667
rect 11161 24633 11195 24667
rect 12909 24633 12943 24667
rect 5181 24565 5215 24599
rect 13277 24565 13311 24599
rect 17969 24565 18003 24599
rect 19993 24565 20027 24599
rect 22753 24565 22787 24599
rect 2881 24361 2915 24395
rect 3157 24361 3191 24395
rect 4537 24361 4571 24395
rect 7481 24361 7515 24395
rect 8585 24361 8619 24395
rect 11253 24361 11287 24395
rect 12633 24361 12667 24395
rect 15025 24293 15059 24327
rect 7941 24225 7975 24259
rect 8125 24225 8159 24259
rect 10609 24225 10643 24259
rect 12081 24225 12115 24259
rect 13185 24225 13219 24259
rect 14381 24225 14415 24259
rect 14565 24225 14599 24259
rect 15669 24225 15703 24259
rect 15761 24225 15795 24259
rect 17969 24225 18003 24259
rect 18061 24225 18095 24259
rect 19993 24225 20027 24259
rect 20177 24225 20211 24259
rect 21373 24225 21407 24259
rect 23397 24225 23431 24259
rect 3341 24157 3375 24191
rect 4052 24157 4086 24191
rect 8217 24157 8251 24191
rect 10885 24157 10919 24191
rect 11897 24157 11931 24191
rect 19901 24157 19935 24191
rect 24041 24157 24075 24191
rect 2605 24089 2639 24123
rect 11989 24089 12023 24123
rect 13277 24089 13311 24123
rect 15853 24089 15887 24123
rect 21189 24089 21223 24123
rect 24777 24089 24811 24123
rect 4123 24021 4157 24055
rect 9137 24021 9171 24055
rect 11529 24021 11563 24055
rect 13369 24021 13403 24055
rect 13737 24021 13771 24055
rect 14657 24021 14691 24055
rect 16221 24021 16255 24055
rect 17417 24021 17451 24055
rect 18153 24021 18187 24055
rect 18521 24021 18555 24055
rect 19533 24021 19567 24055
rect 20729 24021 20763 24055
rect 21097 24021 21131 24055
rect 24685 24021 24719 24055
rect 8861 23817 8895 23851
rect 9965 23817 9999 23851
rect 10425 23817 10459 23851
rect 12725 23817 12759 23851
rect 13553 23817 13587 23851
rect 15945 23817 15979 23851
rect 16037 23817 16071 23851
rect 20545 23817 20579 23851
rect 3525 23749 3559 23783
rect 8953 23749 8987 23783
rect 12633 23749 12667 23783
rect 25145 23749 25179 23783
rect 6009 23681 6043 23715
rect 10057 23681 10091 23715
rect 10885 23681 10919 23715
rect 17509 23681 17543 23715
rect 23305 23681 23339 23715
rect 24133 23681 24167 23715
rect 3801 23613 3835 23647
rect 5733 23613 5767 23647
rect 9045 23613 9079 23647
rect 9781 23613 9815 23647
rect 12449 23613 12483 23647
rect 16221 23613 16255 23647
rect 23029 23613 23063 23647
rect 6469 23545 6503 23579
rect 2053 23477 2087 23511
rect 4261 23477 4295 23511
rect 8493 23477 8527 23511
rect 11529 23477 11563 23511
rect 13093 23477 13127 23511
rect 15577 23477 15611 23511
rect 17693 23477 17727 23511
rect 4169 23273 4203 23307
rect 9045 23273 9079 23307
rect 9229 23273 9263 23307
rect 13737 23273 13771 23307
rect 18889 23273 18923 23307
rect 20177 23273 20211 23307
rect 22293 23273 22327 23307
rect 11437 23205 11471 23239
rect 7021 23137 7055 23171
rect 7297 23137 7331 23171
rect 7665 23137 7699 23171
rect 10241 23137 10275 23171
rect 11989 23137 12023 23171
rect 13277 23137 13311 23171
rect 17417 23137 17451 23171
rect 21649 23137 21683 23171
rect 23397 23137 23431 23171
rect 25237 23137 25271 23171
rect 2789 23069 2823 23103
rect 4353 23069 4387 23103
rect 11897 23069 11931 23103
rect 17141 23069 17175 23103
rect 21925 23069 21959 23103
rect 24041 23069 24075 23103
rect 24961 23069 24995 23103
rect 1777 23001 1811 23035
rect 9965 23001 9999 23035
rect 10793 23001 10827 23035
rect 11805 23001 11839 23035
rect 13093 23001 13127 23035
rect 19349 23001 19383 23035
rect 5549 22933 5583 22967
rect 8401 22933 8435 22967
rect 9597 22933 9631 22967
rect 10057 22933 10091 22967
rect 12633 22933 12667 22967
rect 13001 22933 13035 22967
rect 24593 22933 24627 22967
rect 25053 22933 25087 22967
rect 1961 22729 1995 22763
rect 2605 22729 2639 22763
rect 4031 22729 4065 22763
rect 10793 22729 10827 22763
rect 12725 22729 12759 22763
rect 15117 22729 15151 22763
rect 15761 22729 15795 22763
rect 25145 22729 25179 22763
rect 7389 22661 7423 22695
rect 8217 22661 8251 22695
rect 10149 22661 10183 22695
rect 10977 22661 11011 22695
rect 12541 22661 12575 22695
rect 12909 22661 12943 22695
rect 13645 22661 13679 22695
rect 16129 22661 16163 22695
rect 16497 22661 16531 22695
rect 17141 22661 17175 22695
rect 21373 22661 21407 22695
rect 22293 22661 22327 22695
rect 23213 22661 23247 22695
rect 2145 22593 2179 22627
rect 3065 22593 3099 22627
rect 3928 22593 3962 22627
rect 5549 22593 5583 22627
rect 5641 22593 5675 22627
rect 10425 22593 10459 22627
rect 13369 22593 13403 22627
rect 15577 22593 15611 22627
rect 17233 22593 17267 22627
rect 18061 22593 18095 22627
rect 22937 22593 22971 22627
rect 25329 22593 25363 22627
rect 3249 22525 3283 22559
rect 5733 22525 5767 22559
rect 8677 22525 8711 22559
rect 12357 22525 12391 22559
rect 17049 22525 17083 22559
rect 19073 22525 19107 22559
rect 20821 22525 20855 22559
rect 21097 22525 21131 22559
rect 5181 22389 5215 22423
rect 17601 22389 17635 22423
rect 22385 22389 22419 22423
rect 24685 22389 24719 22423
rect 6193 22185 6227 22219
rect 17417 22185 17451 22219
rect 22017 22185 22051 22219
rect 25421 22185 25455 22219
rect 24777 22117 24811 22151
rect 6837 22049 6871 22083
rect 8033 22049 8067 22083
rect 11345 22049 11379 22083
rect 12449 22049 12483 22083
rect 14841 22049 14875 22083
rect 15669 22049 15703 22083
rect 18705 22049 18739 22083
rect 19625 22049 19659 22083
rect 21465 22049 21499 22083
rect 23397 22049 23431 22083
rect 2237 21981 2271 22015
rect 2881 21981 2915 22015
rect 6561 21981 6595 22015
rect 7757 21981 7791 22015
rect 13369 21981 13403 22015
rect 14657 21981 14691 22015
rect 19717 21981 19751 22015
rect 24041 21981 24075 22015
rect 10517 21913 10551 21947
rect 12357 21913 12391 21947
rect 15945 21913 15979 21947
rect 17969 21913 18003 21947
rect 20637 21913 20671 21947
rect 21833 21913 21867 21947
rect 2053 21845 2087 21879
rect 2697 21845 2731 21879
rect 6653 21845 6687 21879
rect 7389 21845 7423 21879
rect 7849 21845 7883 21879
rect 11897 21845 11931 21879
rect 12265 21845 12299 21879
rect 13185 21845 13219 21879
rect 13829 21845 13863 21879
rect 14289 21845 14323 21879
rect 14749 21845 14783 21879
rect 15393 21845 15427 21879
rect 19809 21845 19843 21879
rect 20177 21845 20211 21879
rect 2513 21641 2547 21675
rect 6561 21641 6595 21675
rect 6929 21641 6963 21675
rect 7757 21641 7791 21675
rect 8217 21641 8251 21675
rect 10333 21641 10367 21675
rect 11069 21641 11103 21675
rect 11621 21641 11655 21675
rect 17785 21641 17819 21675
rect 18521 21641 18555 21675
rect 22017 21641 22051 21675
rect 25053 21641 25087 21675
rect 11713 21573 11747 21607
rect 13001 21573 13035 21607
rect 15025 21573 15059 21607
rect 22661 21573 22695 21607
rect 3893 21505 3927 21539
rect 4905 21505 4939 21539
rect 7021 21505 7055 21539
rect 8125 21505 8159 21539
rect 13093 21505 13127 21539
rect 14289 21505 14323 21539
rect 15485 21505 15519 21539
rect 18429 21505 18463 21539
rect 21373 21505 21407 21539
rect 2973 21437 3007 21471
rect 3157 21437 3191 21471
rect 7113 21437 7147 21471
rect 8309 21437 8343 21471
rect 9689 21437 9723 21471
rect 10425 21437 10459 21471
rect 10609 21437 10643 21471
rect 12909 21437 12943 21471
rect 14381 21437 14415 21471
rect 14473 21437 14507 21471
rect 15117 21437 15151 21471
rect 18337 21437 18371 21471
rect 21097 21437 21131 21471
rect 24409 21437 24443 21471
rect 24685 21437 24719 21471
rect 4445 21369 4479 21403
rect 9965 21369 9999 21403
rect 13921 21369 13955 21403
rect 15669 21369 15703 21403
rect 3709 21301 3743 21335
rect 4813 21301 4847 21335
rect 13461 21301 13495 21335
rect 17509 21301 17543 21335
rect 18889 21301 18923 21335
rect 19625 21301 19659 21335
rect 2881 21097 2915 21131
rect 7665 21097 7699 21131
rect 10333 21097 10367 21131
rect 11437 21097 11471 21131
rect 12633 21097 12667 21131
rect 16313 21097 16347 21131
rect 19625 21097 19659 21131
rect 22293 21029 22327 21063
rect 23489 21029 23523 21063
rect 3433 20961 3467 20995
rect 5273 20961 5307 20995
rect 8217 20961 8251 20995
rect 10793 20961 10827 20995
rect 10885 20961 10919 20995
rect 11989 20961 12023 20995
rect 14289 20961 14323 20995
rect 14565 20961 14599 20995
rect 18613 20961 18647 20995
rect 18797 20961 18831 20995
rect 20545 20961 20579 20995
rect 3249 20893 3283 20927
rect 4997 20893 5031 20927
rect 7021 20893 7055 20927
rect 13553 20893 13587 20927
rect 18521 20893 18555 20927
rect 19441 20893 19475 20927
rect 8125 20825 8159 20859
rect 10701 20825 10735 20859
rect 12173 20825 12207 20859
rect 20821 20825 20855 20859
rect 22937 20825 22971 20859
rect 23121 20825 23155 20859
rect 4353 20757 4387 20791
rect 6745 20757 6779 20791
rect 7297 20757 7331 20791
rect 8033 20757 8067 20791
rect 11529 20757 11563 20791
rect 12265 20757 12299 20791
rect 16037 20757 16071 20791
rect 16865 20757 16899 20791
rect 18153 20757 18187 20791
rect 10333 20553 10367 20587
rect 12081 20553 12115 20587
rect 14749 20553 14783 20587
rect 14841 20553 14875 20587
rect 16405 20553 16439 20587
rect 17233 20553 17267 20587
rect 20729 20553 20763 20587
rect 22385 20553 22419 20587
rect 22477 20553 22511 20587
rect 23305 20553 23339 20587
rect 25329 20553 25363 20587
rect 4169 20485 4203 20519
rect 17141 20485 17175 20519
rect 18981 20485 19015 20519
rect 1777 20417 1811 20451
rect 3893 20417 3927 20451
rect 7757 20417 7791 20451
rect 8585 20417 8619 20451
rect 12173 20417 12207 20451
rect 15761 20417 15795 20451
rect 18705 20417 18739 20451
rect 25053 20417 25087 20451
rect 2053 20349 2087 20383
rect 7573 20349 7607 20383
rect 7665 20349 7699 20383
rect 8861 20349 8895 20383
rect 11161 20349 11195 20383
rect 12265 20349 12299 20383
rect 15025 20349 15059 20383
rect 17049 20349 17083 20383
rect 20453 20349 20487 20383
rect 22661 20349 22695 20383
rect 24777 20349 24811 20383
rect 8125 20281 8159 20315
rect 22017 20281 22051 20315
rect 5641 20213 5675 20247
rect 6009 20213 6043 20247
rect 7021 20213 7055 20247
rect 11713 20213 11747 20247
rect 14381 20213 14415 20247
rect 15577 20213 15611 20247
rect 17601 20213 17635 20247
rect 5457 20009 5491 20043
rect 6947 20009 6981 20043
rect 9137 20009 9171 20043
rect 10517 20009 10551 20043
rect 12449 20009 12483 20043
rect 16129 19941 16163 19975
rect 7205 19873 7239 19907
rect 8401 19873 8435 19907
rect 9689 19873 9723 19907
rect 11805 19873 11839 19907
rect 11989 19873 12023 19907
rect 18337 19873 18371 19907
rect 18521 19873 18555 19907
rect 23397 19873 23431 19907
rect 2237 19805 2271 19839
rect 8309 19805 8343 19839
rect 9505 19805 9539 19839
rect 11713 19805 11747 19839
rect 15945 19805 15979 19839
rect 16865 19805 16899 19839
rect 17233 19805 17267 19839
rect 18245 19805 18279 19839
rect 19625 19805 19659 19839
rect 21281 19805 21315 19839
rect 24041 19805 24075 19839
rect 8217 19737 8251 19771
rect 22017 19737 22051 19771
rect 22201 19737 22235 19771
rect 2053 19669 2087 19703
rect 7481 19669 7515 19703
rect 7849 19669 7883 19703
rect 9597 19669 9631 19703
rect 11345 19669 11379 19703
rect 17325 19669 17359 19703
rect 17877 19669 17911 19703
rect 19441 19669 19475 19703
rect 21373 19669 21407 19703
rect 4905 19465 4939 19499
rect 10425 19465 10459 19499
rect 13093 19465 13127 19499
rect 18153 19465 18187 19499
rect 6929 19397 6963 19431
rect 9229 19397 9263 19431
rect 10885 19397 10919 19431
rect 16957 19397 16991 19431
rect 17325 19397 17359 19431
rect 20545 19397 20579 19431
rect 22569 19397 22603 19431
rect 5089 19329 5123 19363
rect 7205 19329 7239 19363
rect 10793 19329 10827 19363
rect 13461 19329 13495 19363
rect 17969 19329 18003 19363
rect 18797 19329 18831 19363
rect 21465 19329 21499 19363
rect 23397 19329 23431 19363
rect 24409 19329 24443 19363
rect 25237 19329 25271 19363
rect 7481 19261 7515 19295
rect 9597 19261 9631 19295
rect 10977 19261 11011 19295
rect 12817 19261 12851 19295
rect 13553 19261 13587 19295
rect 13645 19261 13679 19295
rect 14197 19193 14231 19227
rect 17417 19125 17451 19159
rect 18613 19125 18647 19159
rect 3985 18921 4019 18955
rect 10701 18921 10735 18955
rect 12449 18921 12483 18955
rect 23593 18921 23627 18955
rect 24225 18921 24259 18955
rect 9781 18853 9815 18887
rect 12725 18853 12759 18887
rect 17877 18853 17911 18887
rect 20177 18853 20211 18887
rect 21741 18853 21775 18887
rect 8309 18785 8343 18819
rect 11345 18785 11379 18819
rect 13185 18785 13219 18819
rect 13369 18785 13403 18819
rect 17325 18785 17359 18819
rect 17417 18785 17451 18819
rect 18153 18785 18187 18819
rect 19625 18785 19659 18819
rect 19717 18785 19751 18819
rect 20913 18785 20947 18819
rect 23857 18785 23891 18819
rect 2237 18717 2271 18751
rect 4169 18717 4203 18751
rect 8585 18717 8619 18751
rect 13093 18717 13127 18751
rect 16865 18717 16899 18751
rect 17509 18717 17543 18751
rect 21005 18717 21039 18751
rect 24777 18717 24811 18751
rect 11069 18649 11103 18683
rect 24593 18649 24627 18683
rect 2053 18581 2087 18615
rect 6837 18581 6871 18615
rect 9229 18581 9263 18615
rect 10333 18581 10367 18615
rect 11161 18581 11195 18615
rect 19073 18581 19107 18615
rect 19809 18581 19843 18615
rect 21097 18581 21131 18615
rect 21465 18581 21499 18615
rect 22109 18581 22143 18615
rect 11529 18377 11563 18411
rect 12449 18377 12483 18411
rect 13645 18377 13679 18411
rect 17693 18377 17727 18411
rect 19993 18377 20027 18411
rect 24409 18377 24443 18411
rect 10885 18309 10919 18343
rect 17141 18309 17175 18343
rect 18889 18309 18923 18343
rect 20361 18309 20395 18343
rect 24685 18309 24719 18343
rect 1777 18241 1811 18275
rect 7941 18241 7975 18275
rect 12817 18241 12851 18275
rect 14013 18241 14047 18275
rect 21189 18241 21223 18275
rect 22661 18241 22695 18275
rect 2053 18173 2087 18207
rect 8677 18173 8711 18207
rect 11161 18173 11195 18207
rect 12173 18173 12207 18207
rect 12909 18173 12943 18207
rect 13093 18173 13127 18207
rect 14105 18173 14139 18207
rect 14197 18173 14231 18207
rect 18061 18173 18095 18207
rect 22937 18173 22971 18207
rect 9413 18037 9447 18071
rect 17049 18037 17083 18071
rect 21649 18037 21683 18071
rect 8677 17833 8711 17867
rect 9505 17833 9539 17867
rect 13553 17833 13587 17867
rect 16037 17833 16071 17867
rect 18981 17833 19015 17867
rect 6929 17765 6963 17799
rect 6561 17697 6595 17731
rect 7665 17697 7699 17731
rect 11529 17697 11563 17731
rect 13093 17697 13127 17731
rect 14749 17697 14783 17731
rect 14933 17697 14967 17731
rect 17785 17697 17819 17731
rect 19441 17697 19475 17731
rect 23397 17697 23431 17731
rect 7849 17629 7883 17663
rect 9597 17629 9631 17663
rect 9873 17629 9907 17663
rect 11253 17629 11287 17663
rect 13001 17629 13035 17663
rect 24041 17629 24075 17663
rect 6285 17561 6319 17595
rect 7205 17561 7239 17595
rect 7941 17561 7975 17595
rect 10517 17561 10551 17595
rect 12909 17561 12943 17595
rect 17509 17561 17543 17595
rect 18337 17561 18371 17595
rect 18521 17561 18555 17595
rect 19717 17561 19751 17595
rect 21741 17561 21775 17595
rect 21925 17561 21959 17595
rect 4813 17493 4847 17527
rect 8309 17493 8343 17527
rect 9137 17493 9171 17527
rect 12541 17493 12575 17527
rect 14289 17493 14323 17527
rect 14657 17493 14691 17527
rect 15393 17493 15427 17527
rect 18797 17493 18831 17527
rect 21189 17493 21223 17527
rect 22201 17493 22235 17527
rect 5273 17289 5307 17323
rect 5641 17289 5675 17323
rect 7021 17289 7055 17323
rect 7481 17289 7515 17323
rect 10149 17289 10183 17323
rect 11713 17289 11747 17323
rect 12081 17289 12115 17323
rect 12173 17289 12207 17323
rect 13645 17289 13679 17323
rect 15853 17289 15887 17323
rect 16681 17289 16715 17323
rect 19073 17289 19107 17323
rect 19717 17289 19751 17323
rect 23765 17289 23799 17323
rect 24133 17289 24167 17323
rect 9137 17221 9171 17255
rect 10609 17221 10643 17255
rect 14749 17221 14783 17255
rect 22293 17221 22327 17255
rect 7389 17153 7423 17187
rect 9229 17153 9263 17187
rect 10517 17153 10551 17187
rect 15945 17153 15979 17187
rect 5733 17085 5767 17119
rect 5825 17085 5859 17119
rect 7573 17085 7607 17119
rect 9321 17085 9355 17119
rect 10701 17085 10735 17119
rect 12265 17085 12299 17119
rect 13001 17085 13035 17119
rect 13737 17085 13771 17119
rect 13829 17085 13863 17119
rect 15761 17085 15795 17119
rect 17325 17085 17359 17119
rect 17601 17085 17635 17119
rect 19441 17085 19475 17119
rect 21189 17085 21223 17119
rect 21465 17085 21499 17119
rect 22017 17085 22051 17119
rect 8769 17017 8803 17051
rect 13277 17017 13311 17051
rect 16313 17017 16347 17051
rect 14841 16949 14875 16983
rect 5904 16745 5938 16779
rect 7941 16745 7975 16779
rect 11437 16745 11471 16779
rect 16221 16745 16255 16779
rect 24409 16745 24443 16779
rect 2421 16609 2455 16643
rect 5641 16609 5675 16643
rect 9597 16609 9631 16643
rect 9689 16609 9723 16643
rect 10793 16609 10827 16643
rect 10885 16609 10919 16643
rect 11897 16609 11931 16643
rect 12173 16609 12207 16643
rect 14105 16609 14139 16643
rect 20085 16609 20119 16643
rect 23121 16609 23155 16643
rect 23397 16609 23431 16643
rect 2605 16541 2639 16575
rect 15761 16541 15795 16575
rect 20177 16541 20211 16575
rect 7665 16473 7699 16507
rect 9505 16473 9539 16507
rect 10701 16473 10735 16507
rect 9137 16405 9171 16439
rect 10333 16405 10367 16439
rect 13645 16405 13679 16439
rect 15945 16405 15979 16439
rect 20269 16405 20303 16439
rect 20637 16405 20671 16439
rect 21649 16405 21683 16439
rect 23857 16405 23891 16439
rect 7573 16201 7607 16235
rect 7941 16201 7975 16235
rect 10793 16201 10827 16235
rect 16221 16133 16255 16167
rect 20545 16133 20579 16167
rect 1777 16065 1811 16099
rect 9137 16065 9171 16099
rect 15209 16065 15243 16099
rect 21281 16065 21315 16099
rect 23397 16065 23431 16099
rect 23949 16065 23983 16099
rect 2053 15997 2087 16031
rect 8033 15997 8067 16031
rect 8125 15997 8159 16031
rect 9229 15997 9263 16031
rect 9321 15997 9355 16031
rect 10885 15997 10919 16031
rect 10977 15997 11011 16031
rect 15301 15997 15335 16031
rect 15485 15997 15519 16031
rect 19533 15997 19567 16031
rect 21465 15997 21499 16031
rect 23029 15997 23063 16031
rect 24777 15997 24811 16031
rect 10425 15929 10459 15963
rect 16037 15929 16071 15963
rect 17785 15929 17819 15963
rect 20729 15929 20763 15963
rect 8769 15861 8803 15895
rect 14841 15861 14875 15895
rect 16773 15861 16807 15895
rect 19993 15861 20027 15895
rect 6193 15657 6227 15691
rect 11989 15657 12023 15691
rect 12817 15657 12851 15691
rect 17693 15657 17727 15691
rect 21097 15657 21131 15691
rect 8309 15589 8343 15623
rect 10241 15521 10275 15555
rect 12449 15521 12483 15555
rect 15945 15521 15979 15555
rect 18245 15521 18279 15555
rect 18429 15521 18463 15555
rect 19625 15521 19659 15555
rect 20637 15521 20671 15555
rect 21649 15521 21683 15555
rect 23857 15521 23891 15555
rect 7941 15453 7975 15487
rect 14473 15453 14507 15487
rect 14841 15453 14875 15487
rect 19717 15453 19751 15487
rect 21741 15453 21775 15487
rect 21833 15453 21867 15487
rect 22661 15453 22695 15487
rect 7665 15385 7699 15419
rect 10517 15385 10551 15419
rect 16221 15385 16255 15419
rect 19809 15385 19843 15419
rect 14381 15317 14415 15351
rect 18521 15317 18555 15351
rect 18889 15317 18923 15351
rect 20177 15317 20211 15351
rect 22201 15317 22235 15351
rect 13093 15113 13127 15147
rect 13461 15113 13495 15147
rect 18521 15113 18555 15147
rect 19533 15113 19567 15147
rect 19901 15113 19935 15147
rect 10977 15045 11011 15079
rect 12541 15045 12575 15079
rect 16129 15045 16163 15079
rect 16681 15045 16715 15079
rect 19441 15045 19475 15079
rect 23305 15045 23339 15079
rect 13553 14977 13587 15011
rect 17417 14977 17451 15011
rect 20545 14977 20579 15011
rect 21465 14977 21499 15011
rect 22109 14977 22143 15011
rect 23949 14977 23983 15011
rect 10333 14909 10367 14943
rect 10609 14909 10643 14943
rect 13645 14909 13679 14943
rect 17141 14909 17175 14943
rect 17325 14909 17359 14943
rect 18061 14909 18095 14943
rect 19349 14909 19383 14943
rect 24685 14909 24719 14943
rect 12357 14841 12391 14875
rect 16313 14841 16347 14875
rect 17785 14841 17819 14875
rect 8861 14773 8895 14807
rect 20361 14773 20395 14807
rect 21281 14773 21315 14807
rect 9229 14569 9263 14603
rect 10517 14569 10551 14603
rect 12817 14569 12851 14603
rect 15025 14569 15059 14603
rect 18797 14569 18831 14603
rect 8309 14433 8343 14467
rect 9689 14433 9723 14467
rect 9873 14433 9907 14467
rect 11989 14433 12023 14467
rect 13277 14433 13311 14467
rect 13369 14433 13403 14467
rect 8585 14365 8619 14399
rect 12265 14365 12299 14399
rect 16773 14365 16807 14399
rect 17509 14365 17543 14399
rect 18061 14365 18095 14399
rect 23121 14365 23155 14399
rect 16497 14297 16531 14331
rect 18245 14297 18279 14331
rect 6837 14229 6871 14263
rect 9597 14229 9631 14263
rect 13185 14229 13219 14263
rect 17325 14229 17359 14263
rect 18521 14229 18555 14263
rect 18889 14229 18923 14263
rect 23305 14229 23339 14263
rect 8493 14025 8527 14059
rect 12725 14025 12759 14059
rect 13093 14025 13127 14059
rect 13185 14025 13219 14059
rect 14657 14025 14691 14059
rect 18613 14025 18647 14059
rect 21005 14025 21039 14059
rect 21465 14025 21499 14059
rect 22201 14025 22235 14059
rect 10885 13957 10919 13991
rect 11253 13957 11287 13991
rect 14289 13957 14323 13991
rect 15301 13957 15335 13991
rect 16037 13957 16071 13991
rect 19901 13957 19935 13991
rect 20361 13957 20395 13991
rect 21097 13957 21131 13991
rect 25145 13957 25179 13991
rect 2789 13889 2823 13923
rect 12357 13889 12391 13923
rect 14197 13889 14231 13923
rect 20085 13889 20119 13923
rect 22017 13889 22051 13923
rect 22661 13889 22695 13923
rect 23949 13889 23983 13923
rect 1777 13821 1811 13855
rect 8861 13821 8895 13855
rect 9137 13821 9171 13855
rect 13277 13821 13311 13855
rect 14105 13821 14139 13855
rect 15485 13821 15519 13855
rect 15853 13821 15887 13855
rect 16865 13821 16899 13855
rect 17141 13821 17175 13855
rect 19073 13821 19107 13855
rect 20821 13821 20855 13855
rect 22845 13753 22879 13787
rect 23121 13685 23155 13719
rect 8953 13481 8987 13515
rect 13829 13481 13863 13515
rect 14197 13481 14231 13515
rect 15485 13481 15519 13515
rect 18889 13481 18923 13515
rect 12817 13413 12851 13447
rect 19349 13413 19383 13447
rect 19901 13413 19935 13447
rect 7113 13345 7147 13379
rect 12265 13345 12299 13379
rect 13185 13345 13219 13379
rect 18337 13345 18371 13379
rect 18429 13345 18463 13379
rect 22569 13345 22603 13379
rect 23029 13345 23063 13379
rect 6837 13277 6871 13311
rect 14933 13277 14967 13311
rect 18521 13277 18555 13311
rect 19717 13277 19751 13311
rect 20177 13277 20211 13311
rect 23673 13277 23707 13311
rect 12449 13209 12483 13243
rect 17509 13209 17543 13243
rect 22293 13209 22327 13243
rect 8585 13141 8619 13175
rect 12357 13141 12391 13175
rect 15025 13141 15059 13175
rect 16865 13141 16899 13175
rect 17601 13141 17635 13175
rect 20821 13141 20855 13175
rect 23857 13141 23891 13175
rect 9137 12937 9171 12971
rect 11805 12937 11839 12971
rect 13185 12937 13219 12971
rect 17141 12937 17175 12971
rect 17233 12937 17267 12971
rect 12265 12869 12299 12903
rect 14473 12869 14507 12903
rect 16313 12869 16347 12903
rect 19073 12869 19107 12903
rect 21189 12869 21223 12903
rect 23305 12869 23339 12903
rect 9229 12801 9263 12835
rect 12173 12801 12207 12835
rect 13553 12801 13587 12835
rect 14197 12801 14231 12835
rect 18337 12801 18371 12835
rect 18429 12801 18463 12835
rect 22109 12801 22143 12835
rect 23949 12801 23983 12835
rect 8953 12733 8987 12767
rect 12357 12733 12391 12767
rect 15945 12733 15979 12767
rect 16957 12733 16991 12767
rect 18245 12733 18279 12767
rect 19717 12733 19751 12767
rect 21465 12733 21499 12767
rect 24777 12733 24811 12767
rect 18797 12665 18831 12699
rect 9597 12597 9631 12631
rect 13645 12597 13679 12631
rect 17601 12597 17635 12631
rect 11069 12393 11103 12427
rect 14289 12393 14323 12427
rect 17141 12393 17175 12427
rect 21005 12393 21039 12427
rect 16405 12325 16439 12359
rect 19993 12325 20027 12359
rect 9321 12257 9355 12291
rect 14933 12257 14967 12291
rect 18889 12257 18923 12291
rect 12817 12189 12851 12223
rect 14657 12189 14691 12223
rect 15577 12189 15611 12223
rect 16221 12189 16255 12223
rect 19533 12189 19567 12223
rect 20821 12189 20855 12223
rect 22661 12189 22695 12223
rect 24777 12189 24811 12223
rect 9597 12121 9631 12155
rect 13553 12121 13587 12155
rect 13737 12121 13771 12155
rect 16681 12121 16715 12155
rect 18613 12121 18647 12155
rect 23857 12121 23891 12155
rect 11345 12053 11379 12087
rect 12909 12053 12943 12087
rect 14749 12053 14783 12087
rect 15669 12053 15703 12087
rect 19625 12053 19659 12087
rect 21557 12053 21591 12087
rect 24593 12053 24627 12087
rect 14381 11849 14415 11883
rect 14933 11849 14967 11883
rect 19809 11849 19843 11883
rect 22661 11849 22695 11883
rect 15301 11781 15335 11815
rect 19625 11713 19659 11747
rect 20361 11713 20395 11747
rect 20821 11713 20855 11747
rect 22477 11713 22511 11747
rect 23213 11713 23247 11747
rect 23949 11713 23983 11747
rect 12633 11645 12667 11679
rect 12909 11645 12943 11679
rect 15393 11645 15427 11679
rect 15485 11645 15519 11679
rect 16129 11645 16163 11679
rect 24685 11645 24719 11679
rect 20545 11577 20579 11611
rect 19073 11509 19107 11543
rect 23397 11509 23431 11543
rect 13277 11305 13311 11339
rect 15485 11305 15519 11339
rect 18337 11305 18371 11339
rect 13829 11237 13863 11271
rect 15025 11237 15059 11271
rect 20177 11237 20211 11271
rect 22937 11237 22971 11271
rect 11253 11169 11287 11203
rect 11529 11169 11563 11203
rect 13001 11169 13035 11203
rect 14381 11169 14415 11203
rect 14565 11169 14599 11203
rect 16037 11169 16071 11203
rect 19533 11169 19567 11203
rect 19717 11169 19751 11203
rect 14657 11101 14691 11135
rect 15853 11101 15887 11135
rect 18153 11101 18187 11135
rect 22753 11101 22787 11135
rect 23857 11101 23891 11135
rect 24777 11101 24811 11135
rect 19809 11033 19843 11067
rect 20637 11033 20671 11067
rect 24593 11033 24627 11067
rect 15945 10965 15979 10999
rect 24041 10965 24075 10999
rect 14473 10761 14507 10795
rect 18061 10761 18095 10795
rect 19533 10693 19567 10727
rect 21097 10625 21131 10659
rect 23949 10625 23983 10659
rect 19809 10557 19843 10591
rect 24777 10557 24811 10591
rect 20177 10489 20211 10523
rect 15393 10421 15427 10455
rect 21281 10421 21315 10455
rect 23397 10081 23431 10115
rect 11621 10013 11655 10047
rect 17049 10013 17083 10047
rect 24041 10013 24075 10047
rect 24777 10013 24811 10047
rect 11805 9945 11839 9979
rect 16865 9945 16899 9979
rect 24593 9877 24627 9911
rect 6837 9605 6871 9639
rect 14381 9605 14415 9639
rect 6009 9537 6043 9571
rect 6929 9537 6963 9571
rect 22017 9537 22051 9571
rect 23949 9537 23983 9571
rect 6745 9469 6779 9503
rect 24777 9469 24811 9503
rect 7297 9401 7331 9435
rect 14565 9401 14599 9435
rect 22201 9333 22235 9367
rect 16129 8925 16163 8959
rect 18521 8925 18555 8959
rect 23121 8925 23155 8959
rect 24869 8925 24903 8959
rect 25329 8925 25363 8959
rect 16313 8857 16347 8891
rect 18705 8857 18739 8891
rect 23765 8857 23799 8891
rect 23949 8857 23983 8891
rect 23305 8789 23339 8823
rect 24685 8789 24719 8823
rect 25237 8789 25271 8823
rect 5917 8517 5951 8551
rect 25145 8517 25179 8551
rect 3893 8449 3927 8483
rect 6377 8449 6411 8483
rect 23489 8449 23523 8483
rect 24041 8449 24075 8483
rect 4169 8381 4203 8415
rect 23029 8381 23063 8415
rect 23397 7905 23431 7939
rect 18705 7837 18739 7871
rect 20361 7837 20395 7871
rect 24041 7837 24075 7871
rect 24869 7837 24903 7871
rect 18889 7769 18923 7803
rect 20545 7769 20579 7803
rect 24685 7701 24719 7735
rect 21465 7361 21499 7395
rect 22109 7361 22143 7395
rect 24133 7361 24167 7395
rect 21005 7293 21039 7327
rect 22569 7293 22603 7327
rect 24777 7293 24811 7327
rect 23397 6817 23431 6851
rect 18245 6749 18279 6783
rect 19441 6749 19475 6783
rect 20821 6749 20855 6783
rect 24041 6749 24075 6783
rect 24777 6749 24811 6783
rect 18429 6681 18463 6715
rect 22017 6681 22051 6715
rect 19625 6613 19659 6647
rect 24593 6613 24627 6647
rect 19533 6409 19567 6443
rect 21281 6341 21315 6375
rect 19441 6273 19475 6307
rect 20085 6273 20119 6307
rect 22109 6273 22143 6307
rect 23949 6273 23983 6307
rect 22569 6205 22603 6239
rect 24777 6205 24811 6239
rect 20177 5865 20211 5899
rect 21189 5729 21223 5763
rect 23029 5729 23063 5763
rect 19993 5661 20027 5695
rect 20729 5661 20763 5695
rect 22569 5661 22603 5695
rect 16221 5253 16255 5287
rect 16037 5185 16071 5219
rect 19165 5185 19199 5219
rect 19625 5185 19659 5219
rect 22017 5185 22051 5219
rect 24133 5185 24167 5219
rect 18705 5117 18739 5151
rect 20085 5117 20119 5151
rect 22477 5117 22511 5151
rect 24777 5117 24811 5151
rect 25329 4777 25363 4811
rect 19901 4641 19935 4675
rect 21741 4641 21775 4675
rect 17417 4573 17451 4607
rect 19441 4573 19475 4607
rect 21281 4573 21315 4607
rect 18337 4505 18371 4539
rect 1409 4437 1443 4471
rect 1593 4097 1627 4131
rect 8125 4097 8159 4131
rect 9321 4097 9355 4131
rect 9873 4097 9907 4131
rect 13001 4097 13035 4131
rect 16865 4097 16899 4131
rect 18705 4097 18739 4131
rect 22109 4097 22143 4131
rect 23857 4097 23891 4131
rect 13461 4029 13495 4063
rect 17325 4029 17359 4063
rect 19165 4029 19199 4063
rect 22477 4029 22511 4063
rect 24317 4029 24351 4063
rect 1777 3961 1811 3995
rect 7941 3961 7975 3995
rect 9505 3961 9539 3995
rect 2237 3893 2271 3927
rect 2881 3893 2915 3927
rect 3249 3893 3283 3927
rect 5549 3893 5583 3927
rect 8493 3893 8527 3927
rect 11253 3893 11287 3927
rect 12633 3893 12667 3927
rect 2513 3689 2547 3723
rect 3249 3689 3283 3723
rect 5089 3689 5123 3723
rect 6561 3689 6595 3723
rect 7665 3689 7699 3723
rect 8401 3689 8435 3723
rect 11529 3689 11563 3723
rect 25237 3689 25271 3723
rect 1869 3621 1903 3655
rect 5825 3621 5859 3655
rect 10333 3553 10367 3587
rect 14749 3553 14783 3587
rect 16589 3553 16623 3587
rect 19901 3553 19935 3587
rect 21741 3553 21775 3587
rect 23489 3553 23523 3587
rect 2329 3485 2363 3519
rect 3065 3485 3099 3519
rect 4905 3485 4939 3519
rect 5641 3485 5675 3519
rect 6377 3485 6411 3519
rect 6929 3485 6963 3519
rect 7481 3485 7515 3519
rect 8217 3485 8251 3519
rect 9597 3485 9631 3519
rect 10057 3485 10091 3519
rect 11345 3485 11379 3519
rect 11897 3485 11931 3519
rect 13737 3485 13771 3519
rect 14289 3485 14323 3519
rect 16129 3485 16163 3519
rect 19441 3485 19475 3519
rect 21281 3485 21315 3519
rect 23213 3485 23247 3519
rect 24409 3485 24443 3519
rect 24777 3485 24811 3519
rect 25053 3485 25087 3519
rect 1685 3417 1719 3451
rect 12541 3417 12575 3451
rect 3893 3349 3927 3383
rect 4169 3349 4203 3383
rect 4445 3349 4479 3383
rect 4629 3349 4663 3383
rect 7205 3349 7239 3383
rect 9413 3349 9447 3383
rect 2145 3145 2179 3179
rect 4445 3145 4479 3179
rect 5089 3145 5123 3179
rect 5917 3145 5951 3179
rect 23857 3145 23891 3179
rect 1961 3009 1995 3043
rect 2881 3009 2915 3043
rect 3801 3009 3835 3043
rect 4261 3009 4295 3043
rect 5273 3009 5307 3043
rect 5825 3009 5859 3043
rect 6377 3009 6411 3043
rect 7389 3009 7423 3043
rect 8861 3009 8895 3043
rect 11161 3009 11195 3043
rect 12265 3009 12299 3043
rect 14197 3009 14231 3043
rect 16221 3009 16255 3043
rect 16865 3009 16899 3043
rect 18705 3009 18739 3043
rect 25329 3009 25363 3043
rect 3065 2941 3099 2975
rect 7113 2941 7147 2975
rect 8585 2941 8619 2975
rect 10885 2941 10919 2975
rect 12541 2941 12575 2975
rect 13645 2941 13679 2975
rect 15025 2941 15059 2975
rect 17325 2941 17359 2975
rect 19165 2941 19199 2975
rect 3617 2873 3651 2907
rect 1501 2805 1535 2839
rect 1685 2805 1719 2839
rect 6837 2805 6871 2839
rect 8217 2805 8251 2839
rect 9689 2805 9723 2839
rect 9965 2805 9999 2839
rect 11897 2601 11931 2635
rect 24685 2601 24719 2635
rect 25421 2601 25455 2635
rect 2053 2533 2087 2567
rect 5825 2533 5859 2567
rect 7297 2533 7331 2567
rect 3433 2465 3467 2499
rect 4445 2465 4479 2499
rect 10701 2465 10735 2499
rect 14105 2465 14139 2499
rect 17325 2465 17359 2499
rect 19901 2465 19935 2499
rect 22477 2465 22511 2499
rect 1593 2397 1627 2431
rect 1869 2397 1903 2431
rect 3157 2397 3191 2431
rect 4169 2397 4203 2431
rect 6009 2397 6043 2431
rect 8309 2397 8343 2431
rect 8585 2397 8619 2431
rect 11069 2397 11103 2431
rect 11713 2397 11747 2431
rect 12357 2397 12391 2431
rect 15669 2397 15703 2431
rect 16865 2397 16899 2431
rect 19441 2397 19475 2431
rect 22017 2397 22051 2431
rect 24869 2397 24903 2431
rect 25145 2397 25179 2431
rect 6745 2329 6779 2363
rect 7113 2329 7147 2363
rect 13277 2329 13311 2363
rect 14657 2329 14691 2363
rect 3893 2261 3927 2295
rect 5365 2261 5399 2295
rect 6469 2261 6503 2295
rect 8953 2261 8987 2295
rect 9229 2261 9263 2295
<< metal1 >>
rect 1104 54426 25852 54448
rect 1104 54374 7950 54426
rect 8002 54374 8014 54426
rect 8066 54374 8078 54426
rect 8130 54374 8142 54426
rect 8194 54374 8206 54426
rect 8258 54374 17950 54426
rect 18002 54374 18014 54426
rect 18066 54374 18078 54426
rect 18130 54374 18142 54426
rect 18194 54374 18206 54426
rect 18258 54374 25852 54426
rect 1104 54352 25852 54374
rect 13814 54272 13820 54324
rect 13872 54272 13878 54324
rect 14369 54315 14427 54321
rect 14369 54281 14381 54315
rect 14415 54312 14427 54315
rect 14550 54312 14556 54324
rect 14415 54284 14556 54312
rect 14415 54281 14427 54284
rect 14369 54275 14427 54281
rect 14550 54272 14556 54284
rect 14608 54272 14614 54324
rect 19334 54272 19340 54324
rect 19392 54272 19398 54324
rect 8478 54244 8484 54256
rect 6886 54216 8484 54244
rect 3421 54179 3479 54185
rect 3421 54145 3433 54179
rect 3467 54176 3479 54179
rect 5902 54176 5908 54188
rect 3467 54148 5908 54176
rect 3467 54145 3479 54148
rect 3421 54139 3479 54145
rect 5902 54136 5908 54148
rect 5960 54136 5966 54188
rect 5997 54179 6055 54185
rect 5997 54145 6009 54179
rect 6043 54176 6055 54179
rect 6886 54176 6914 54216
rect 8478 54204 8484 54216
rect 8536 54204 8542 54256
rect 10870 54204 10876 54256
rect 10928 54204 10934 54256
rect 6043 54148 6914 54176
rect 8573 54179 8631 54185
rect 6043 54145 6055 54148
rect 5997 54139 6055 54145
rect 8573 54145 8585 54179
rect 8619 54176 8631 54179
rect 8619 54148 9812 54176
rect 8619 54145 8631 54148
rect 8573 54139 8631 54145
rect 2961 54111 3019 54117
rect 2961 54077 2973 54111
rect 3007 54108 3019 54111
rect 5350 54108 5356 54120
rect 3007 54080 5356 54108
rect 3007 54077 3019 54080
rect 2961 54071 3019 54077
rect 5350 54068 5356 54080
rect 5408 54068 5414 54120
rect 5537 54111 5595 54117
rect 5537 54077 5549 54111
rect 5583 54108 5595 54111
rect 7190 54108 7196 54120
rect 5583 54080 7196 54108
rect 5583 54077 5595 54080
rect 5537 54071 5595 54077
rect 7190 54068 7196 54080
rect 7248 54068 7254 54120
rect 8113 54111 8171 54117
rect 8113 54077 8125 54111
rect 8159 54108 8171 54111
rect 9398 54108 9404 54120
rect 8159 54080 9404 54108
rect 8159 54077 8171 54080
rect 8113 54071 8171 54077
rect 9398 54068 9404 54080
rect 9456 54068 9462 54120
rect 9784 54108 9812 54148
rect 9858 54136 9864 54188
rect 9916 54136 9922 54188
rect 12066 54136 12072 54188
rect 12124 54136 12130 54188
rect 14568 54176 14596 54272
rect 14918 54204 14924 54256
rect 14976 54244 14982 54256
rect 15473 54247 15531 54253
rect 15473 54244 15485 54247
rect 14976 54216 15485 54244
rect 14976 54204 14982 54216
rect 15473 54213 15485 54216
rect 15519 54213 15531 54247
rect 15473 54207 15531 54213
rect 16022 54204 16028 54256
rect 16080 54244 16086 54256
rect 16666 54244 16672 54256
rect 16080 54216 16672 54244
rect 16080 54204 16086 54216
rect 16666 54204 16672 54216
rect 16724 54244 16730 54256
rect 16724 54216 16896 54244
rect 16724 54204 16730 54216
rect 14645 54179 14703 54185
rect 14645 54176 14657 54179
rect 14568 54148 14657 54176
rect 14645 54145 14657 54148
rect 14691 54145 14703 54179
rect 14645 54139 14703 54145
rect 15286 54136 15292 54188
rect 15344 54176 15350 54188
rect 15838 54176 15844 54188
rect 15344 54148 15844 54176
rect 15344 54136 15350 54148
rect 15838 54136 15844 54148
rect 15896 54176 15902 54188
rect 16868 54185 16896 54216
rect 17494 54204 17500 54256
rect 17552 54244 17558 54256
rect 18414 54244 18420 54256
rect 17552 54216 18420 54244
rect 17552 54204 17558 54216
rect 18414 54204 18420 54216
rect 18472 54204 18478 54256
rect 19352 54244 19380 54272
rect 19352 54216 20024 54244
rect 16117 54179 16175 54185
rect 16117 54176 16129 54179
rect 15896 54148 16129 54176
rect 15896 54136 15902 54148
rect 16117 54145 16129 54148
rect 16163 54145 16175 54179
rect 16117 54139 16175 54145
rect 16853 54179 16911 54185
rect 16853 54145 16865 54179
rect 16899 54145 16911 54179
rect 16853 54139 16911 54145
rect 17126 54136 17132 54188
rect 17184 54176 17190 54188
rect 17773 54179 17831 54185
rect 17773 54176 17785 54179
rect 17184 54148 17785 54176
rect 17184 54136 17190 54148
rect 17773 54145 17785 54148
rect 17819 54145 17831 54179
rect 17773 54139 17831 54145
rect 11882 54108 11888 54120
rect 9784 54080 11888 54108
rect 11882 54068 11888 54080
rect 11940 54068 11946 54120
rect 11974 54068 11980 54120
rect 12032 54108 12038 54120
rect 12529 54111 12587 54117
rect 12529 54108 12541 54111
rect 12032 54080 12541 54108
rect 12032 54068 12038 54080
rect 12529 54077 12541 54080
rect 12575 54077 12587 54111
rect 17788 54108 17816 54139
rect 18598 54136 18604 54188
rect 18656 54176 18662 54188
rect 19334 54176 19340 54188
rect 18656 54148 19340 54176
rect 18656 54136 18662 54148
rect 19334 54136 19340 54148
rect 19392 54176 19398 54188
rect 19429 54179 19487 54185
rect 19429 54176 19441 54179
rect 19392 54148 19441 54176
rect 19392 54136 19398 54148
rect 19429 54145 19441 54148
rect 19475 54145 19487 54179
rect 19996 54176 20024 54216
rect 20070 54204 20076 54256
rect 20128 54244 20134 54256
rect 20714 54244 20720 54256
rect 20128 54216 20720 54244
rect 20128 54204 20134 54216
rect 20714 54204 20720 54216
rect 20772 54244 20778 54256
rect 20772 54216 20944 54244
rect 20772 54204 20778 54216
rect 20916 54185 20944 54216
rect 22646 54204 22652 54256
rect 22704 54244 22710 54256
rect 25041 54247 25099 54253
rect 25041 54244 25053 54247
rect 22704 54216 25053 54244
rect 22704 54204 22710 54216
rect 20349 54179 20407 54185
rect 20349 54176 20361 54179
rect 19996 54148 20361 54176
rect 19429 54139 19487 54145
rect 20349 54145 20361 54148
rect 20395 54145 20407 54179
rect 20349 54139 20407 54145
rect 20901 54179 20959 54185
rect 20901 54145 20913 54179
rect 20947 54145 20959 54179
rect 20901 54139 20959 54145
rect 18877 54111 18935 54117
rect 18877 54108 18889 54111
rect 17788 54080 18889 54108
rect 12529 54071 12587 54077
rect 18877 54077 18889 54080
rect 18923 54077 18935 54111
rect 20364 54108 20392 54139
rect 21174 54136 21180 54188
rect 21232 54176 21238 54188
rect 21818 54176 21824 54188
rect 21232 54148 21824 54176
rect 21232 54136 21238 54148
rect 21818 54136 21824 54148
rect 21876 54176 21882 54188
rect 22189 54179 22247 54185
rect 22189 54176 22201 54179
rect 21876 54148 22201 54176
rect 21876 54136 21882 54148
rect 22189 54145 22201 54148
rect 22235 54145 22247 54179
rect 22189 54139 22247 54145
rect 23934 54136 23940 54188
rect 23992 54136 23998 54188
rect 24780 54185 24808 54216
rect 25041 54213 25053 54216
rect 25087 54213 25099 54247
rect 25041 54207 25099 54213
rect 24765 54179 24823 54185
rect 24765 54145 24777 54179
rect 24811 54145 24823 54179
rect 24765 54139 24823 54145
rect 21453 54111 21511 54117
rect 21453 54108 21465 54111
rect 20364 54080 21465 54108
rect 18877 54071 18935 54077
rect 21453 54077 21465 54080
rect 21499 54077 21511 54111
rect 21453 54071 21511 54077
rect 23569 54111 23627 54117
rect 23569 54077 23581 54111
rect 23615 54108 23627 54111
rect 24118 54108 24124 54120
rect 23615 54080 24124 54108
rect 23615 54077 23627 54080
rect 23569 54071 23627 54077
rect 24118 54068 24124 54080
rect 24176 54068 24182 54120
rect 15654 54000 15660 54052
rect 15712 54000 15718 54052
rect 18598 54000 18604 54052
rect 18656 54000 18662 54052
rect 21726 54000 21732 54052
rect 21784 54040 21790 54052
rect 24581 54043 24639 54049
rect 24581 54040 24593 54043
rect 21784 54012 24593 54040
rect 21784 54000 21790 54012
rect 24581 54009 24593 54012
rect 24627 54009 24639 54043
rect 24581 54003 24639 54009
rect 14829 53975 14887 53981
rect 14829 53941 14841 53975
rect 14875 53972 14887 53975
rect 15102 53972 15108 53984
rect 14875 53944 15108 53972
rect 14875 53941 14887 53944
rect 14829 53935 14887 53941
rect 15102 53932 15108 53944
rect 15160 53932 15166 53984
rect 16301 53975 16359 53981
rect 16301 53941 16313 53975
rect 16347 53972 16359 53975
rect 16482 53972 16488 53984
rect 16347 53944 16488 53972
rect 16347 53941 16359 53944
rect 16301 53935 16359 53941
rect 16482 53932 16488 53944
rect 16540 53932 16546 53984
rect 16942 53932 16948 53984
rect 17000 53972 17006 53984
rect 17037 53975 17095 53981
rect 17037 53972 17049 53975
rect 17000 53944 17049 53972
rect 17000 53932 17006 53944
rect 17037 53941 17049 53944
rect 17083 53941 17095 53975
rect 17037 53935 17095 53941
rect 17681 53975 17739 53981
rect 17681 53941 17693 53975
rect 17727 53972 17739 53975
rect 17770 53972 17776 53984
rect 17727 53944 17776 53972
rect 17727 53941 17739 53944
rect 17681 53935 17739 53941
rect 17770 53932 17776 53944
rect 17828 53932 17834 53984
rect 19610 53932 19616 53984
rect 19668 53932 19674 53984
rect 20257 53975 20315 53981
rect 20257 53941 20269 53975
rect 20303 53972 20315 53975
rect 20530 53972 20536 53984
rect 20303 53944 20536 53972
rect 20303 53941 20315 53944
rect 20257 53935 20315 53941
rect 20530 53932 20536 53944
rect 20588 53932 20594 53984
rect 21085 53975 21143 53981
rect 21085 53941 21097 53975
rect 21131 53972 21143 53975
rect 21174 53972 21180 53984
rect 21131 53944 21180 53972
rect 21131 53941 21143 53944
rect 21085 53935 21143 53941
rect 21174 53932 21180 53944
rect 21232 53932 21238 53984
rect 22002 53932 22008 53984
rect 22060 53932 22066 53984
rect 1104 53882 25852 53904
rect 1104 53830 2950 53882
rect 3002 53830 3014 53882
rect 3066 53830 3078 53882
rect 3130 53830 3142 53882
rect 3194 53830 3206 53882
rect 3258 53830 12950 53882
rect 13002 53830 13014 53882
rect 13066 53830 13078 53882
rect 13130 53830 13142 53882
rect 13194 53830 13206 53882
rect 13258 53830 22950 53882
rect 23002 53830 23014 53882
rect 23066 53830 23078 53882
rect 23130 53830 23142 53882
rect 23194 53830 23206 53882
rect 23258 53830 25852 53882
rect 1104 53808 25852 53830
rect 14918 53728 14924 53780
rect 14976 53768 14982 53780
rect 15197 53771 15255 53777
rect 15197 53768 15209 53771
rect 14976 53740 15209 53768
rect 14976 53728 14982 53740
rect 15197 53737 15209 53740
rect 15243 53737 15255 53771
rect 15197 53731 15255 53737
rect 15473 53771 15531 53777
rect 15473 53737 15485 53771
rect 15519 53768 15531 53771
rect 15562 53768 15568 53780
rect 15519 53740 15568 53768
rect 15519 53737 15531 53740
rect 15473 53731 15531 53737
rect 15562 53728 15568 53740
rect 15620 53728 15626 53780
rect 20257 53771 20315 53777
rect 20257 53737 20269 53771
rect 20303 53768 20315 53771
rect 20438 53768 20444 53780
rect 20303 53740 20444 53768
rect 20303 53737 20315 53740
rect 20257 53731 20315 53737
rect 20438 53728 20444 53740
rect 20496 53728 20502 53780
rect 25590 53700 25596 53712
rect 23216 53672 25596 53700
rect 2961 53635 3019 53641
rect 2961 53601 2973 53635
rect 3007 53632 3019 53635
rect 4614 53632 4620 53644
rect 3007 53604 4620 53632
rect 3007 53601 3019 53604
rect 2961 53595 3019 53601
rect 4614 53592 4620 53604
rect 4672 53592 4678 53644
rect 6273 53635 6331 53641
rect 6273 53601 6285 53635
rect 6319 53632 6331 53635
rect 7558 53632 7564 53644
rect 6319 53604 7564 53632
rect 6319 53601 6331 53604
rect 6273 53595 6331 53601
rect 7558 53592 7564 53604
rect 7616 53592 7622 53644
rect 8294 53592 8300 53644
rect 8352 53592 8358 53644
rect 10502 53592 10508 53644
rect 10560 53592 10566 53644
rect 11606 53592 11612 53644
rect 11664 53632 11670 53644
rect 23216 53641 23244 53672
rect 25590 53660 25596 53672
rect 25648 53660 25654 53712
rect 12161 53635 12219 53641
rect 12161 53632 12173 53635
rect 11664 53604 12173 53632
rect 11664 53592 11670 53604
rect 12161 53601 12173 53604
rect 12207 53601 12219 53635
rect 12161 53595 12219 53601
rect 23201 53635 23259 53641
rect 23201 53601 23213 53635
rect 23247 53601 23259 53635
rect 23201 53595 23259 53601
rect 23290 53592 23296 53644
rect 23348 53632 23354 53644
rect 25041 53635 25099 53641
rect 25041 53632 25053 53635
rect 23348 53604 25053 53632
rect 23348 53592 23354 53604
rect 3421 53567 3479 53573
rect 3421 53533 3433 53567
rect 3467 53564 3479 53567
rect 6178 53564 6184 53576
rect 3467 53536 6184 53564
rect 3467 53533 3479 53536
rect 3421 53527 3479 53533
rect 6178 53524 6184 53536
rect 6236 53524 6242 53576
rect 6638 53524 6644 53576
rect 6696 53524 6702 53576
rect 7374 53524 7380 53576
rect 7432 53524 7438 53576
rect 9030 53524 9036 53576
rect 9088 53564 9094 53576
rect 9674 53564 9680 53576
rect 9088 53536 9680 53564
rect 9088 53524 9094 53536
rect 9674 53524 9680 53536
rect 9732 53524 9738 53576
rect 11054 53524 11060 53576
rect 11112 53524 11118 53576
rect 11882 53524 11888 53576
rect 11940 53524 11946 53576
rect 13541 53567 13599 53573
rect 13541 53533 13553 53567
rect 13587 53564 13599 53567
rect 13814 53564 13820 53576
rect 13587 53536 13820 53564
rect 13587 53533 13599 53536
rect 13541 53527 13599 53533
rect 13814 53524 13820 53536
rect 13872 53524 13878 53576
rect 14182 53524 14188 53576
rect 14240 53564 14246 53576
rect 14553 53567 14611 53573
rect 14553 53564 14565 53567
rect 14240 53536 14565 53564
rect 14240 53524 14246 53536
rect 14553 53533 14565 53536
rect 14599 53564 14611 53567
rect 14829 53567 14887 53573
rect 14829 53564 14841 53567
rect 14599 53536 14841 53564
rect 14599 53533 14611 53536
rect 14553 53527 14611 53533
rect 14829 53533 14841 53536
rect 14875 53533 14887 53567
rect 14829 53527 14887 53533
rect 15562 53524 15568 53576
rect 15620 53564 15626 53576
rect 15749 53567 15807 53573
rect 15749 53564 15761 53567
rect 15620 53536 15761 53564
rect 15620 53524 15626 53536
rect 15749 53533 15761 53536
rect 15795 53533 15807 53567
rect 15749 53527 15807 53533
rect 16390 53524 16396 53576
rect 16448 53564 16454 53576
rect 16485 53567 16543 53573
rect 16485 53564 16497 53567
rect 16448 53536 16497 53564
rect 16448 53524 16454 53536
rect 16485 53533 16497 53536
rect 16531 53533 16543 53567
rect 16485 53527 16543 53533
rect 16758 53524 16764 53576
rect 16816 53564 16822 53576
rect 17221 53567 17279 53573
rect 17221 53564 17233 53567
rect 16816 53536 17233 53564
rect 16816 53524 16822 53536
rect 17221 53533 17233 53536
rect 17267 53533 17279 53567
rect 17221 53527 17279 53533
rect 17862 53524 17868 53576
rect 17920 53564 17926 53576
rect 17957 53567 18015 53573
rect 17957 53564 17969 53567
rect 17920 53536 17969 53564
rect 17920 53524 17926 53536
rect 17957 53533 17969 53536
rect 18003 53533 18015 53567
rect 17957 53527 18015 53533
rect 18322 53524 18328 53576
rect 18380 53564 18386 53576
rect 18877 53567 18935 53573
rect 18877 53564 18889 53567
rect 18380 53536 18889 53564
rect 18380 53524 18386 53536
rect 18877 53533 18889 53536
rect 18923 53533 18935 53567
rect 18877 53527 18935 53533
rect 18966 53524 18972 53576
rect 19024 53564 19030 53576
rect 19705 53567 19763 53573
rect 19705 53564 19717 53567
rect 19024 53536 19717 53564
rect 19024 53524 19030 53536
rect 19705 53533 19717 53536
rect 19751 53564 19763 53567
rect 19981 53567 20039 53573
rect 19981 53564 19993 53567
rect 19751 53536 19993 53564
rect 19751 53533 19763 53536
rect 19705 53527 19763 53533
rect 19981 53533 19993 53536
rect 20027 53533 20039 53567
rect 19981 53527 20039 53533
rect 20438 53524 20444 53576
rect 20496 53564 20502 53576
rect 20533 53567 20591 53573
rect 20533 53564 20545 53567
rect 20496 53536 20545 53564
rect 20496 53524 20502 53536
rect 20533 53533 20545 53536
rect 20579 53533 20591 53567
rect 20533 53527 20591 53533
rect 20806 53524 20812 53576
rect 20864 53564 20870 53576
rect 21269 53567 21327 53573
rect 21269 53564 21281 53567
rect 20864 53536 21281 53564
rect 20864 53524 20870 53536
rect 21269 53533 21281 53536
rect 21315 53533 21327 53567
rect 21269 53527 21327 53533
rect 21542 53524 21548 53576
rect 21600 53564 21606 53576
rect 22189 53567 22247 53573
rect 22189 53564 22201 53567
rect 21600 53536 22201 53564
rect 21600 53524 21606 53536
rect 22189 53533 22201 53536
rect 22235 53533 22247 53567
rect 22189 53527 22247 53533
rect 24026 53524 24032 53576
rect 24084 53524 24090 53576
rect 24780 53573 24808 53604
rect 25041 53601 25053 53604
rect 25087 53601 25099 53635
rect 25041 53595 25099 53601
rect 24765 53567 24823 53573
rect 24765 53533 24777 53567
rect 24811 53533 24823 53567
rect 24765 53527 24823 53533
rect 3786 53388 3792 53440
rect 3844 53388 3850 53440
rect 13630 53388 13636 53440
rect 13688 53428 13694 53440
rect 13725 53431 13783 53437
rect 13725 53428 13737 53431
rect 13688 53400 13737 53428
rect 13688 53388 13694 53400
rect 13725 53397 13737 53400
rect 13771 53397 13783 53431
rect 13725 53391 13783 53397
rect 14369 53431 14427 53437
rect 14369 53397 14381 53431
rect 14415 53428 14427 53431
rect 15746 53428 15752 53440
rect 14415 53400 15752 53428
rect 14415 53397 14427 53400
rect 14369 53391 14427 53397
rect 15746 53388 15752 53400
rect 15804 53388 15810 53440
rect 15930 53388 15936 53440
rect 15988 53388 15994 53440
rect 16669 53431 16727 53437
rect 16669 53397 16681 53431
rect 16715 53428 16727 53431
rect 17034 53428 17040 53440
rect 16715 53400 17040 53428
rect 16715 53397 16727 53400
rect 16669 53391 16727 53397
rect 17034 53388 17040 53400
rect 17092 53388 17098 53440
rect 17402 53388 17408 53440
rect 17460 53388 17466 53440
rect 18141 53431 18199 53437
rect 18141 53397 18153 53431
rect 18187 53428 18199 53431
rect 18506 53428 18512 53440
rect 18187 53400 18512 53428
rect 18187 53397 18199 53400
rect 18141 53391 18199 53397
rect 18506 53388 18512 53400
rect 18564 53388 18570 53440
rect 18690 53388 18696 53440
rect 18748 53388 18754 53440
rect 19518 53388 19524 53440
rect 19576 53388 19582 53440
rect 20717 53431 20775 53437
rect 20717 53397 20729 53431
rect 20763 53428 20775 53431
rect 21266 53428 21272 53440
rect 20763 53400 21272 53428
rect 20763 53397 20775 53400
rect 20717 53391 20775 53397
rect 21266 53388 21272 53400
rect 21324 53388 21330 53440
rect 21450 53388 21456 53440
rect 21508 53388 21514 53440
rect 21542 53388 21548 53440
rect 21600 53428 21606 53440
rect 22005 53431 22063 53437
rect 22005 53428 22017 53431
rect 21600 53400 22017 53428
rect 21600 53388 21606 53400
rect 22005 53397 22017 53400
rect 22051 53397 22063 53431
rect 22005 53391 22063 53397
rect 24486 53388 24492 53440
rect 24544 53428 24550 53440
rect 24581 53431 24639 53437
rect 24581 53428 24593 53431
rect 24544 53400 24593 53428
rect 24544 53388 24550 53400
rect 24581 53397 24593 53400
rect 24627 53397 24639 53431
rect 24581 53391 24639 53397
rect 25314 53388 25320 53440
rect 25372 53428 25378 53440
rect 25409 53431 25467 53437
rect 25409 53428 25421 53431
rect 25372 53400 25421 53428
rect 25372 53388 25378 53400
rect 25409 53397 25421 53400
rect 25455 53397 25467 53431
rect 25409 53391 25467 53397
rect 1104 53338 25852 53360
rect 1104 53286 7950 53338
rect 8002 53286 8014 53338
rect 8066 53286 8078 53338
rect 8130 53286 8142 53338
rect 8194 53286 8206 53338
rect 8258 53286 17950 53338
rect 18002 53286 18014 53338
rect 18066 53286 18078 53338
rect 18130 53286 18142 53338
rect 18194 53286 18206 53338
rect 18258 53286 25852 53338
rect 1104 53264 25852 53286
rect 2041 53227 2099 53233
rect 2041 53193 2053 53227
rect 2087 53224 2099 53227
rect 2774 53224 2780 53236
rect 2087 53196 2780 53224
rect 2087 53193 2099 53196
rect 2041 53187 2099 53193
rect 1581 53091 1639 53097
rect 1581 53057 1593 53091
rect 1627 53088 1639 53091
rect 2056 53088 2084 53187
rect 2774 53184 2780 53196
rect 2832 53184 2838 53236
rect 15838 53184 15844 53236
rect 15896 53224 15902 53236
rect 15933 53227 15991 53233
rect 15933 53224 15945 53227
rect 15896 53196 15945 53224
rect 15896 53184 15902 53196
rect 15933 53193 15945 53196
rect 15979 53193 15991 53227
rect 15933 53187 15991 53193
rect 16390 53184 16396 53236
rect 16448 53184 16454 53236
rect 16666 53184 16672 53236
rect 16724 53184 16730 53236
rect 16758 53184 16764 53236
rect 16816 53224 16822 53236
rect 17037 53227 17095 53233
rect 17037 53224 17049 53227
rect 16816 53196 17049 53224
rect 16816 53184 16822 53196
rect 17037 53193 17049 53196
rect 17083 53193 17095 53227
rect 17037 53187 17095 53193
rect 17862 53184 17868 53236
rect 17920 53184 17926 53236
rect 18322 53184 18328 53236
rect 18380 53224 18386 53236
rect 18509 53227 18567 53233
rect 18509 53224 18521 53227
rect 18380 53196 18521 53224
rect 18380 53184 18386 53196
rect 18509 53193 18521 53196
rect 18555 53193 18567 53227
rect 18509 53187 18567 53193
rect 19334 53184 19340 53236
rect 19392 53184 19398 53236
rect 20714 53184 20720 53236
rect 20772 53184 20778 53236
rect 20806 53184 20812 53236
rect 20864 53224 20870 53236
rect 21085 53227 21143 53233
rect 21085 53224 21097 53227
rect 20864 53196 21097 53224
rect 20864 53184 20870 53196
rect 21085 53193 21097 53196
rect 21131 53193 21143 53227
rect 21085 53187 21143 53193
rect 21453 53227 21511 53233
rect 21453 53193 21465 53227
rect 21499 53224 21511 53227
rect 21634 53224 21640 53236
rect 21499 53196 21640 53224
rect 21499 53193 21511 53196
rect 21453 53187 21511 53193
rect 21634 53184 21640 53196
rect 21692 53184 21698 53236
rect 6362 53156 6368 53168
rect 4080 53128 6368 53156
rect 4080 53097 4108 53128
rect 6362 53116 6368 53128
rect 6420 53116 6426 53168
rect 12710 53116 12716 53168
rect 12768 53156 12774 53168
rect 14461 53159 14519 53165
rect 14461 53156 14473 53159
rect 12768 53128 14473 53156
rect 12768 53116 12774 53128
rect 14461 53125 14473 53128
rect 14507 53156 14519 53159
rect 14829 53159 14887 53165
rect 14829 53156 14841 53159
rect 14507 53128 14841 53156
rect 14507 53125 14519 53128
rect 14461 53119 14519 53125
rect 14829 53125 14841 53128
rect 14875 53125 14887 53159
rect 14829 53119 14887 53125
rect 18233 53159 18291 53165
rect 18233 53125 18245 53159
rect 18279 53156 18291 53159
rect 18414 53156 18420 53168
rect 18279 53128 18420 53156
rect 18279 53125 18291 53128
rect 18233 53119 18291 53125
rect 18414 53116 18420 53128
rect 18472 53116 18478 53168
rect 1627 53060 2084 53088
rect 4065 53091 4123 53097
rect 1627 53057 1639 53060
rect 1581 53051 1639 53057
rect 4065 53057 4077 53091
rect 4111 53057 4123 53091
rect 4065 53051 4123 53057
rect 5810 53048 5816 53100
rect 5868 53048 5874 53100
rect 6730 53048 6736 53100
rect 6788 53088 6794 53100
rect 6825 53091 6883 53097
rect 6825 53088 6837 53091
rect 6788 53060 6837 53088
rect 6788 53048 6794 53060
rect 6825 53057 6837 53060
rect 6871 53057 6883 53091
rect 6825 53051 6883 53057
rect 9122 53048 9128 53100
rect 9180 53048 9186 53100
rect 9398 53048 9404 53100
rect 9456 53088 9462 53100
rect 9769 53091 9827 53097
rect 9769 53088 9781 53091
rect 9456 53060 9781 53088
rect 9456 53048 9462 53060
rect 9769 53057 9781 53060
rect 9815 53057 9827 53091
rect 9769 53051 9827 53057
rect 10686 53048 10692 53100
rect 10744 53088 10750 53100
rect 11701 53091 11759 53097
rect 11701 53088 11713 53091
rect 10744 53060 11713 53088
rect 10744 53048 10750 53060
rect 11701 53057 11713 53060
rect 11747 53057 11759 53091
rect 11701 53051 11759 53057
rect 13446 53048 13452 53100
rect 13504 53088 13510 53100
rect 13817 53091 13875 53097
rect 13817 53088 13829 53091
rect 13504 53060 13829 53088
rect 13504 53048 13510 53060
rect 13817 53057 13829 53060
rect 13863 53057 13875 53091
rect 13817 53051 13875 53057
rect 19702 53048 19708 53100
rect 19760 53088 19766 53100
rect 19981 53091 20039 53097
rect 19981 53088 19993 53091
rect 19760 53060 19993 53088
rect 19760 53048 19766 53060
rect 19981 53057 19993 53060
rect 20027 53088 20039 53091
rect 20257 53091 20315 53097
rect 20257 53088 20269 53091
rect 20027 53060 20269 53088
rect 20027 53057 20039 53060
rect 19981 53051 20039 53057
rect 20257 53057 20269 53060
rect 20303 53057 20315 53091
rect 20257 53051 20315 53057
rect 21637 53091 21695 53097
rect 21637 53057 21649 53091
rect 21683 53088 21695 53091
rect 21910 53088 21916 53100
rect 21683 53060 21916 53088
rect 21683 53057 21695 53060
rect 21637 53051 21695 53057
rect 21910 53048 21916 53060
rect 21968 53088 21974 53100
rect 22005 53091 22063 53097
rect 22005 53088 22017 53091
rect 21968 53060 22017 53088
rect 21968 53048 21974 53060
rect 22005 53057 22017 53060
rect 22051 53057 22063 53091
rect 22005 53051 22063 53057
rect 22278 53048 22284 53100
rect 22336 53088 22342 53100
rect 22925 53091 22983 53097
rect 22925 53088 22937 53091
rect 22336 53060 22937 53088
rect 22336 53048 22342 53060
rect 22925 53057 22937 53060
rect 22971 53088 22983 53091
rect 23201 53091 23259 53097
rect 23201 53088 23213 53091
rect 22971 53060 23213 53088
rect 22971 53057 22983 53060
rect 22925 53051 22983 53057
rect 23201 53057 23213 53060
rect 23247 53057 23259 53091
rect 23201 53051 23259 53057
rect 24946 53048 24952 53100
rect 25004 53088 25010 53100
rect 25133 53091 25191 53097
rect 25133 53088 25145 53091
rect 25004 53060 25145 53088
rect 25004 53048 25010 53060
rect 25133 53057 25145 53060
rect 25179 53057 25191 53091
rect 25133 53051 25191 53057
rect 3697 53023 3755 53029
rect 3697 52989 3709 53023
rect 3743 53020 3755 53023
rect 4246 53020 4252 53032
rect 3743 52992 4252 53020
rect 3743 52989 3755 52992
rect 3697 52983 3755 52989
rect 4246 52980 4252 52992
rect 4304 52980 4310 53032
rect 5537 53023 5595 53029
rect 5537 52989 5549 53023
rect 5583 53020 5595 53023
rect 5718 53020 5724 53032
rect 5583 52992 5724 53020
rect 5583 52989 5595 52992
rect 5537 52983 5595 52989
rect 5718 52980 5724 52992
rect 5776 52980 5782 53032
rect 8662 52980 8668 53032
rect 8720 52980 8726 53032
rect 10134 52980 10140 53032
rect 10192 53020 10198 53032
rect 10229 53023 10287 53029
rect 10229 53020 10241 53023
rect 10192 52992 10241 53020
rect 10192 52980 10198 52992
rect 10229 52989 10241 52992
rect 10275 52989 10287 53023
rect 10229 52983 10287 52989
rect 11238 52980 11244 53032
rect 11296 53020 11302 53032
rect 12161 53023 12219 53029
rect 12161 53020 12173 53023
rect 11296 52992 12173 53020
rect 11296 52980 11302 52992
rect 12161 52989 12173 52992
rect 12207 52989 12219 53023
rect 12161 52983 12219 52989
rect 24854 52980 24860 53032
rect 24912 52980 24918 53032
rect 1765 52887 1823 52893
rect 1765 52853 1777 52887
rect 1811 52884 1823 52887
rect 4062 52884 4068 52896
rect 1811 52856 4068 52884
rect 1811 52853 1823 52856
rect 1765 52847 1823 52853
rect 4062 52844 4068 52856
rect 4120 52844 4126 52896
rect 5994 52844 6000 52896
rect 6052 52884 6058 52896
rect 6641 52887 6699 52893
rect 6641 52884 6653 52887
rect 6052 52856 6653 52884
rect 6052 52844 6058 52856
rect 6641 52853 6653 52856
rect 6687 52853 6699 52887
rect 6641 52847 6699 52853
rect 12802 52844 12808 52896
rect 12860 52884 12866 52896
rect 13633 52887 13691 52893
rect 13633 52884 13645 52887
rect 12860 52856 13645 52884
rect 12860 52844 12866 52856
rect 13633 52853 13645 52856
rect 13679 52853 13691 52887
rect 13633 52847 13691 52853
rect 14366 52844 14372 52896
rect 14424 52844 14430 52896
rect 19794 52844 19800 52896
rect 19852 52844 19858 52896
rect 22186 52844 22192 52896
rect 22244 52844 22250 52896
rect 22738 52844 22744 52896
rect 22796 52844 22802 52896
rect 23474 52844 23480 52896
rect 23532 52884 23538 52896
rect 25222 52884 25228 52896
rect 23532 52856 25228 52884
rect 23532 52844 23538 52856
rect 25222 52844 25228 52856
rect 25280 52844 25286 52896
rect 1104 52794 25852 52816
rect 1104 52742 2950 52794
rect 3002 52742 3014 52794
rect 3066 52742 3078 52794
rect 3130 52742 3142 52794
rect 3194 52742 3206 52794
rect 3258 52742 12950 52794
rect 13002 52742 13014 52794
rect 13066 52742 13078 52794
rect 13130 52742 13142 52794
rect 13194 52742 13206 52794
rect 13258 52742 22950 52794
rect 23002 52742 23014 52794
rect 23066 52742 23078 52794
rect 23130 52742 23142 52794
rect 23194 52742 23206 52794
rect 23258 52742 25852 52794
rect 1104 52720 25852 52742
rect 934 52640 940 52692
rect 992 52680 998 52692
rect 4338 52680 4344 52692
rect 992 52652 4344 52680
rect 992 52640 998 52652
rect 4338 52640 4344 52652
rect 4396 52640 4402 52692
rect 11977 52683 12035 52689
rect 11977 52649 11989 52683
rect 12023 52680 12035 52683
rect 12066 52680 12072 52692
rect 12023 52652 12072 52680
rect 12023 52649 12035 52652
rect 11977 52643 12035 52649
rect 12066 52640 12072 52652
rect 12124 52640 12130 52692
rect 13446 52640 13452 52692
rect 13504 52680 13510 52692
rect 14093 52683 14151 52689
rect 14093 52680 14105 52683
rect 13504 52652 14105 52680
rect 13504 52640 13510 52652
rect 14093 52649 14105 52652
rect 14139 52649 14151 52683
rect 14093 52643 14151 52649
rect 21818 52640 21824 52692
rect 21876 52640 21882 52692
rect 23934 52640 23940 52692
rect 23992 52640 23998 52692
rect 1210 52572 1216 52624
rect 1268 52612 1274 52624
rect 3786 52612 3792 52624
rect 1268 52584 3792 52612
rect 1268 52572 1274 52584
rect 3786 52572 3792 52584
rect 3844 52612 3850 52624
rect 12621 52615 12679 52621
rect 3844 52584 4016 52612
rect 3844 52572 3850 52584
rect 2961 52547 3019 52553
rect 2961 52513 2973 52547
rect 3007 52544 3019 52547
rect 3326 52544 3332 52556
rect 3007 52516 3332 52544
rect 3007 52513 3019 52516
rect 2961 52507 3019 52513
rect 3326 52504 3332 52516
rect 3384 52504 3390 52556
rect 3988 52553 4016 52584
rect 12621 52581 12633 52615
rect 12667 52612 12679 52615
rect 13354 52612 13360 52624
rect 12667 52584 13360 52612
rect 12667 52581 12679 52584
rect 12621 52575 12679 52581
rect 13354 52572 13360 52584
rect 13412 52572 13418 52624
rect 24762 52572 24768 52624
rect 24820 52612 24826 52624
rect 25958 52612 25964 52624
rect 24820 52584 25964 52612
rect 24820 52572 24826 52584
rect 25958 52572 25964 52584
rect 26016 52572 26022 52624
rect 3973 52547 4031 52553
rect 3973 52513 3985 52547
rect 4019 52513 4031 52547
rect 4430 52544 4436 52556
rect 3973 52507 4031 52513
rect 4080 52516 4436 52544
rect 3421 52479 3479 52485
rect 3421 52445 3433 52479
rect 3467 52476 3479 52479
rect 4080 52476 4108 52516
rect 4430 52504 4436 52516
rect 4488 52504 4494 52556
rect 6086 52504 6092 52556
rect 6144 52504 6150 52556
rect 6454 52504 6460 52556
rect 6512 52544 6518 52556
rect 6914 52544 6920 52556
rect 6512 52516 6920 52544
rect 6512 52504 6518 52516
rect 6914 52504 6920 52516
rect 6972 52504 6978 52556
rect 7834 52504 7840 52556
rect 7892 52504 7898 52556
rect 9766 52504 9772 52556
rect 9824 52544 9830 52556
rect 10321 52547 10379 52553
rect 10321 52544 10333 52547
rect 9824 52516 10333 52544
rect 9824 52504 9830 52516
rect 10321 52513 10333 52516
rect 10367 52513 10379 52547
rect 25317 52547 25375 52553
rect 25317 52544 25329 52547
rect 10321 52507 10379 52513
rect 25056 52516 25329 52544
rect 3467 52448 4108 52476
rect 4249 52479 4307 52485
rect 3467 52445 3479 52448
rect 3421 52439 3479 52445
rect 4249 52445 4261 52479
rect 4295 52476 4307 52479
rect 4522 52476 4528 52488
rect 4295 52448 4528 52476
rect 4295 52445 4307 52448
rect 4249 52439 4307 52445
rect 4522 52436 4528 52448
rect 4580 52436 4586 52488
rect 6546 52436 6552 52488
rect 6604 52436 6610 52488
rect 8573 52479 8631 52485
rect 8573 52445 8585 52479
rect 8619 52476 8631 52479
rect 9490 52476 9496 52488
rect 8619 52448 9496 52476
rect 8619 52445 8631 52448
rect 8573 52439 8631 52445
rect 9490 52436 9496 52448
rect 9548 52436 9554 52488
rect 9582 52436 9588 52488
rect 9640 52476 9646 52488
rect 9861 52479 9919 52485
rect 9861 52476 9873 52479
rect 9640 52448 9873 52476
rect 9640 52436 9646 52448
rect 9861 52445 9873 52448
rect 9907 52445 9919 52479
rect 9861 52439 9919 52445
rect 11790 52436 11796 52488
rect 11848 52436 11854 52488
rect 12342 52436 12348 52488
rect 12400 52476 12406 52488
rect 12437 52479 12495 52485
rect 12437 52476 12449 52479
rect 12400 52448 12449 52476
rect 12400 52436 12406 52448
rect 12437 52445 12449 52448
rect 12483 52445 12495 52479
rect 12437 52439 12495 52445
rect 13446 52436 13452 52488
rect 13504 52436 13510 52488
rect 23109 52479 23167 52485
rect 23109 52445 23121 52479
rect 23155 52476 23167 52479
rect 23474 52476 23480 52488
rect 23155 52448 23480 52476
rect 23155 52445 23167 52448
rect 23109 52439 23167 52445
rect 23474 52436 23480 52448
rect 23532 52436 23538 52488
rect 23753 52479 23811 52485
rect 23753 52445 23765 52479
rect 23799 52476 23811 52479
rect 24210 52476 24216 52488
rect 23799 52448 24216 52476
rect 23799 52445 23811 52448
rect 23753 52439 23811 52445
rect 24210 52436 24216 52448
rect 24268 52476 24274 52488
rect 25056 52485 25084 52516
rect 25317 52513 25329 52516
rect 25363 52513 25375 52547
rect 25317 52507 25375 52513
rect 24765 52479 24823 52485
rect 24765 52476 24777 52479
rect 24268 52448 24777 52476
rect 24268 52436 24274 52448
rect 24765 52445 24777 52448
rect 24811 52476 24823 52479
rect 25041 52479 25099 52485
rect 25041 52476 25053 52479
rect 24811 52448 25053 52476
rect 24811 52445 24823 52448
rect 24765 52439 24823 52445
rect 25041 52445 25053 52448
rect 25087 52445 25099 52479
rect 25041 52439 25099 52445
rect 25222 52436 25228 52488
rect 25280 52476 25286 52488
rect 25409 52479 25467 52485
rect 25409 52476 25421 52479
rect 25280 52448 25421 52476
rect 25280 52436 25286 52448
rect 25409 52445 25421 52448
rect 25455 52445 25467 52479
rect 25409 52439 25467 52445
rect 12710 52368 12716 52420
rect 12768 52408 12774 52420
rect 13265 52411 13323 52417
rect 13265 52408 13277 52411
rect 12768 52380 13277 52408
rect 12768 52368 12774 52380
rect 13265 52377 13277 52380
rect 13311 52408 13323 52411
rect 13725 52411 13783 52417
rect 13725 52408 13737 52411
rect 13311 52380 13737 52408
rect 13311 52377 13323 52380
rect 13265 52371 13323 52377
rect 13725 52377 13737 52380
rect 13771 52377 13783 52411
rect 13725 52371 13783 52377
rect 23290 52300 23296 52352
rect 23348 52300 23354 52352
rect 24578 52300 24584 52352
rect 24636 52300 24642 52352
rect 1104 52250 25852 52272
rect 1104 52198 7950 52250
rect 8002 52198 8014 52250
rect 8066 52198 8078 52250
rect 8130 52198 8142 52250
rect 8194 52198 8206 52250
rect 8258 52198 17950 52250
rect 18002 52198 18014 52250
rect 18066 52198 18078 52250
rect 18130 52198 18142 52250
rect 18194 52198 18206 52250
rect 18258 52198 25852 52250
rect 1104 52176 25852 52198
rect 11882 52096 11888 52148
rect 11940 52096 11946 52148
rect 12342 52096 12348 52148
rect 12400 52096 12406 52148
rect 23474 52096 23480 52148
rect 23532 52096 23538 52148
rect 23937 52139 23995 52145
rect 23937 52105 23949 52139
rect 23983 52136 23995 52139
rect 24578 52136 24584 52148
rect 23983 52108 24584 52136
rect 23983 52105 23995 52108
rect 23937 52099 23995 52105
rect 24578 52096 24584 52108
rect 24636 52096 24642 52148
rect 4982 52028 4988 52080
rect 5040 52028 5046 52080
rect 7190 52068 7196 52080
rect 6012 52040 7196 52068
rect 4065 52003 4123 52009
rect 4065 51969 4077 52003
rect 4111 52000 4123 52003
rect 5350 52000 5356 52012
rect 4111 51972 5356 52000
rect 4111 51969 4123 51972
rect 4065 51963 4123 51969
rect 5350 51960 5356 51972
rect 5408 51960 5414 52012
rect 6012 52009 6040 52040
rect 7190 52028 7196 52040
rect 7248 52028 7254 52080
rect 5997 52003 6055 52009
rect 5997 51969 6009 52003
rect 6043 51969 6055 52003
rect 5997 51963 6055 51969
rect 7006 51960 7012 52012
rect 7064 51960 7070 52012
rect 10134 51960 10140 52012
rect 10192 52000 10198 52012
rect 10321 52003 10379 52009
rect 10321 52000 10333 52003
rect 10192 51972 10333 52000
rect 10192 51960 10198 51972
rect 10321 51969 10333 51972
rect 10367 51969 10379 52003
rect 10321 51963 10379 51969
rect 11606 51960 11612 52012
rect 11664 52000 11670 52012
rect 11701 52003 11759 52009
rect 11701 52000 11713 52003
rect 11664 51972 11713 52000
rect 11664 51960 11670 51972
rect 11701 51969 11713 51972
rect 11747 51969 11759 52003
rect 11701 51963 11759 51969
rect 23293 52003 23351 52009
rect 23293 51969 23305 52003
rect 23339 52000 23351 52003
rect 23753 52003 23811 52009
rect 23753 52000 23765 52003
rect 23339 51972 23765 52000
rect 23339 51969 23351 51972
rect 23293 51963 23351 51969
rect 23753 51969 23765 51972
rect 23799 52000 23811 52003
rect 24394 52000 24400 52012
rect 23799 51972 24400 52000
rect 23799 51969 23811 51972
rect 23753 51963 23811 51969
rect 24394 51960 24400 51972
rect 24452 51960 24458 52012
rect 24581 52003 24639 52009
rect 24581 51969 24593 52003
rect 24627 52000 24639 52003
rect 24670 52000 24676 52012
rect 24627 51972 24676 52000
rect 24627 51969 24639 51972
rect 24581 51963 24639 51969
rect 24670 51960 24676 51972
rect 24728 51960 24734 52012
rect 25222 51960 25228 52012
rect 25280 51960 25286 52012
rect 3510 51892 3516 51944
rect 3568 51892 3574 51944
rect 7098 51892 7104 51944
rect 7156 51932 7162 51944
rect 7377 51935 7435 51941
rect 7377 51932 7389 51935
rect 7156 51904 7389 51932
rect 7156 51892 7162 51904
rect 7377 51901 7389 51904
rect 7423 51901 7435 51935
rect 7377 51895 7435 51901
rect 9674 51892 9680 51944
rect 9732 51892 9738 51944
rect 24394 51756 24400 51808
rect 24452 51756 24458 51808
rect 25133 51799 25191 51805
rect 25133 51765 25145 51799
rect 25179 51796 25191 51799
rect 25682 51796 25688 51808
rect 25179 51768 25688 51796
rect 25179 51765 25191 51768
rect 25133 51759 25191 51765
rect 25682 51756 25688 51768
rect 25740 51756 25746 51808
rect 1104 51706 25852 51728
rect 1104 51654 2950 51706
rect 3002 51654 3014 51706
rect 3066 51654 3078 51706
rect 3130 51654 3142 51706
rect 3194 51654 3206 51706
rect 3258 51654 12950 51706
rect 13002 51654 13014 51706
rect 13066 51654 13078 51706
rect 13130 51654 13142 51706
rect 13194 51654 13206 51706
rect 13258 51654 22950 51706
rect 23002 51654 23014 51706
rect 23066 51654 23078 51706
rect 23130 51654 23142 51706
rect 23194 51654 23206 51706
rect 23258 51654 25852 51706
rect 1104 51632 25852 51654
rect 5902 51552 5908 51604
rect 5960 51552 5966 51604
rect 24670 51552 24676 51604
rect 24728 51552 24734 51604
rect 24489 51527 24547 51533
rect 24489 51493 24501 51527
rect 24535 51524 24547 51527
rect 24762 51524 24768 51536
rect 24535 51496 24768 51524
rect 24535 51493 24547 51496
rect 24489 51487 24547 51493
rect 2406 51416 2412 51468
rect 2464 51416 2470 51468
rect 4154 51416 4160 51468
rect 4212 51416 4218 51468
rect 6914 51416 6920 51468
rect 6972 51416 6978 51468
rect 3421 51391 3479 51397
rect 3421 51357 3433 51391
rect 3467 51357 3479 51391
rect 3421 51351 3479 51357
rect 5353 51391 5411 51397
rect 5353 51357 5365 51391
rect 5399 51388 5411 51391
rect 5994 51388 6000 51400
rect 5399 51360 6000 51388
rect 5399 51357 5411 51360
rect 5353 51351 5411 51357
rect 3436 51320 3464 51351
rect 5994 51348 6000 51360
rect 6052 51348 6058 51400
rect 6089 51391 6147 51397
rect 6089 51357 6101 51391
rect 6135 51388 6147 51391
rect 7098 51388 7104 51400
rect 6135 51360 7104 51388
rect 6135 51357 6147 51360
rect 6089 51351 6147 51357
rect 7098 51348 7104 51360
rect 7156 51348 7162 51400
rect 7742 51348 7748 51400
rect 7800 51348 7806 51400
rect 24029 51391 24087 51397
rect 24029 51357 24041 51391
rect 24075 51388 24087 51391
rect 24504 51388 24532 51487
rect 24762 51484 24768 51496
rect 24820 51484 24826 51536
rect 24075 51360 24532 51388
rect 24075 51357 24087 51360
rect 24029 51351 24087 51357
rect 25314 51348 25320 51400
rect 25372 51348 25378 51400
rect 6730 51320 6736 51332
rect 3436 51292 6736 51320
rect 6730 51280 6736 51292
rect 6788 51280 6794 51332
rect 20990 51212 20996 51264
rect 21048 51252 21054 51264
rect 22738 51252 22744 51264
rect 21048 51224 22744 51252
rect 21048 51212 21054 51224
rect 22738 51212 22744 51224
rect 22796 51212 22802 51264
rect 23842 51212 23848 51264
rect 23900 51212 23906 51264
rect 25133 51255 25191 51261
rect 25133 51221 25145 51255
rect 25179 51252 25191 51255
rect 25590 51252 25596 51264
rect 25179 51224 25596 51252
rect 25179 51221 25191 51224
rect 25133 51215 25191 51221
rect 25590 51212 25596 51224
rect 25648 51212 25654 51264
rect 1104 51162 25852 51184
rect 1104 51110 7950 51162
rect 8002 51110 8014 51162
rect 8066 51110 8078 51162
rect 8130 51110 8142 51162
rect 8194 51110 8206 51162
rect 8258 51110 17950 51162
rect 18002 51110 18014 51162
rect 18066 51110 18078 51162
rect 18130 51110 18142 51162
rect 18194 51110 18206 51162
rect 18258 51110 25852 51162
rect 1104 51088 25852 51110
rect 9858 51008 9864 51060
rect 9916 51008 9922 51060
rect 10686 51008 10692 51060
rect 10744 51008 10750 51060
rect 2866 50940 2872 50992
rect 2924 50980 2930 50992
rect 3053 50983 3111 50989
rect 3053 50980 3065 50983
rect 2924 50952 3065 50980
rect 2924 50940 2930 50952
rect 3053 50949 3065 50952
rect 3099 50949 3111 50983
rect 3053 50943 3111 50949
rect 6730 50940 6736 50992
rect 6788 50940 6794 50992
rect 1857 50915 1915 50921
rect 1857 50881 1869 50915
rect 1903 50912 1915 50915
rect 1903 50884 2774 50912
rect 1903 50881 1915 50884
rect 1857 50875 1915 50881
rect 1118 50804 1124 50856
rect 1176 50844 1182 50856
rect 1581 50847 1639 50853
rect 1581 50844 1593 50847
rect 1176 50816 1593 50844
rect 1176 50804 1182 50816
rect 1581 50813 1593 50816
rect 1627 50813 1639 50847
rect 1581 50807 1639 50813
rect 2746 50776 2774 50884
rect 4154 50872 4160 50924
rect 4212 50872 4218 50924
rect 6917 50915 6975 50921
rect 6917 50881 6929 50915
rect 6963 50912 6975 50915
rect 8294 50912 8300 50924
rect 6963 50884 8300 50912
rect 6963 50881 6975 50884
rect 6917 50875 6975 50881
rect 8294 50872 8300 50884
rect 8352 50872 8358 50924
rect 8570 50872 8576 50924
rect 8628 50912 8634 50924
rect 9769 50915 9827 50921
rect 9769 50912 9781 50915
rect 8628 50884 9781 50912
rect 8628 50872 8634 50884
rect 9769 50881 9781 50884
rect 9815 50881 9827 50915
rect 9769 50875 9827 50881
rect 9950 50872 9956 50924
rect 10008 50912 10014 50924
rect 10505 50915 10563 50921
rect 10505 50912 10517 50915
rect 10008 50884 10517 50912
rect 10008 50872 10014 50884
rect 10505 50881 10517 50884
rect 10551 50881 10563 50915
rect 10505 50875 10563 50881
rect 24765 50915 24823 50921
rect 24765 50881 24777 50915
rect 24811 50912 24823 50915
rect 25314 50912 25320 50924
rect 24811 50884 25320 50912
rect 24811 50881 24823 50884
rect 24765 50875 24823 50881
rect 25314 50872 25320 50884
rect 25372 50872 25378 50924
rect 6914 50776 6920 50788
rect 2746 50748 6920 50776
rect 6914 50736 6920 50748
rect 6972 50736 6978 50788
rect 25130 50668 25136 50720
rect 25188 50668 25194 50720
rect 1104 50618 25852 50640
rect 1104 50566 2950 50618
rect 3002 50566 3014 50618
rect 3066 50566 3078 50618
rect 3130 50566 3142 50618
rect 3194 50566 3206 50618
rect 3258 50566 12950 50618
rect 13002 50566 13014 50618
rect 13066 50566 13078 50618
rect 13130 50566 13142 50618
rect 13194 50566 13206 50618
rect 13258 50566 22950 50618
rect 23002 50566 23014 50618
rect 23066 50566 23078 50618
rect 23130 50566 23142 50618
rect 23194 50566 23206 50618
rect 23258 50566 25852 50618
rect 1104 50544 25852 50566
rect 1118 50396 1124 50448
rect 1176 50436 1182 50448
rect 1397 50439 1455 50445
rect 1397 50436 1409 50439
rect 1176 50408 1409 50436
rect 1176 50396 1182 50408
rect 1397 50405 1409 50408
rect 1443 50405 1455 50439
rect 1397 50399 1455 50405
rect 9398 50396 9404 50448
rect 9456 50396 9462 50448
rect 2038 50328 2044 50380
rect 2096 50368 2102 50380
rect 2225 50371 2283 50377
rect 2225 50368 2237 50371
rect 2096 50340 2237 50368
rect 2096 50328 2102 50340
rect 2225 50337 2237 50340
rect 2271 50337 2283 50371
rect 2225 50331 2283 50337
rect 4338 50328 4344 50380
rect 4396 50328 4402 50380
rect 3421 50303 3479 50309
rect 3421 50269 3433 50303
rect 3467 50300 3479 50303
rect 3970 50300 3976 50312
rect 3467 50272 3976 50300
rect 3467 50269 3479 50272
rect 3421 50263 3479 50269
rect 3970 50260 3976 50272
rect 4028 50260 4034 50312
rect 5353 50303 5411 50309
rect 5353 50269 5365 50303
rect 5399 50300 5411 50303
rect 8662 50300 8668 50312
rect 5399 50272 8668 50300
rect 5399 50269 5411 50272
rect 5353 50263 5411 50269
rect 8662 50260 8668 50272
rect 8720 50260 8726 50312
rect 24765 50303 24823 50309
rect 24765 50269 24777 50303
rect 24811 50300 24823 50303
rect 25314 50300 25320 50312
rect 24811 50272 25320 50300
rect 24811 50269 24823 50272
rect 24765 50263 24823 50269
rect 25314 50260 25320 50272
rect 25372 50260 25378 50312
rect 7742 50192 7748 50244
rect 7800 50232 7806 50244
rect 9217 50235 9275 50241
rect 9217 50232 9229 50235
rect 7800 50204 9229 50232
rect 7800 50192 7806 50204
rect 9217 50201 9229 50204
rect 9263 50201 9275 50235
rect 9217 50195 9275 50201
rect 23382 50124 23388 50176
rect 23440 50164 23446 50176
rect 25133 50167 25191 50173
rect 25133 50164 25145 50167
rect 23440 50136 25145 50164
rect 23440 50124 23446 50136
rect 25133 50133 25145 50136
rect 25179 50133 25191 50167
rect 25133 50127 25191 50133
rect 1104 50074 25852 50096
rect 1104 50022 7950 50074
rect 8002 50022 8014 50074
rect 8066 50022 8078 50074
rect 8130 50022 8142 50074
rect 8194 50022 8206 50074
rect 8258 50022 17950 50074
rect 18002 50022 18014 50074
rect 18066 50022 18078 50074
rect 18130 50022 18142 50074
rect 18194 50022 18206 50074
rect 18258 50022 25852 50074
rect 1104 50000 25852 50022
rect 6733 49963 6791 49969
rect 6733 49929 6745 49963
rect 6779 49960 6791 49963
rect 7006 49960 7012 49972
rect 6779 49932 7012 49960
rect 6779 49929 6791 49932
rect 6733 49923 6791 49929
rect 7006 49920 7012 49932
rect 7064 49920 7070 49972
rect 7374 49920 7380 49972
rect 7432 49960 7438 49972
rect 7837 49963 7895 49969
rect 7837 49960 7849 49963
rect 7432 49932 7849 49960
rect 7432 49920 7438 49932
rect 7837 49929 7849 49932
rect 7883 49929 7895 49963
rect 7837 49923 7895 49929
rect 21358 49920 21364 49972
rect 21416 49960 21422 49972
rect 25133 49963 25191 49969
rect 25133 49960 25145 49963
rect 21416 49932 25145 49960
rect 21416 49920 21422 49932
rect 25133 49929 25145 49932
rect 25179 49929 25191 49963
rect 25133 49923 25191 49929
rect 1670 49852 1676 49904
rect 1728 49892 1734 49904
rect 1949 49895 2007 49901
rect 1949 49892 1961 49895
rect 1728 49864 1961 49892
rect 1728 49852 1734 49864
rect 1949 49861 1961 49864
rect 1995 49861 2007 49895
rect 1949 49855 2007 49861
rect 7650 49852 7656 49904
rect 7708 49892 7714 49904
rect 9401 49895 9459 49901
rect 9401 49892 9413 49895
rect 7708 49864 9413 49892
rect 7708 49852 7714 49864
rect 9401 49861 9413 49864
rect 9447 49861 9459 49895
rect 9401 49855 9459 49861
rect 9582 49852 9588 49904
rect 9640 49852 9646 49904
rect 3145 49827 3203 49833
rect 3145 49793 3157 49827
rect 3191 49824 3203 49827
rect 3694 49824 3700 49836
rect 3191 49796 3700 49824
rect 3191 49793 3203 49796
rect 3145 49787 3203 49793
rect 3694 49784 3700 49796
rect 3752 49784 3758 49836
rect 6546 49784 6552 49836
rect 6604 49784 6610 49836
rect 7374 49784 7380 49836
rect 7432 49824 7438 49836
rect 8021 49827 8079 49833
rect 8021 49824 8033 49827
rect 7432 49796 8033 49824
rect 7432 49784 7438 49796
rect 8021 49793 8033 49796
rect 8067 49793 8079 49827
rect 8021 49787 8079 49793
rect 24762 49784 24768 49836
rect 24820 49824 24826 49836
rect 25317 49827 25375 49833
rect 25317 49824 25329 49827
rect 24820 49796 25329 49824
rect 24820 49784 24826 49796
rect 25317 49793 25329 49796
rect 25363 49793 25375 49827
rect 25317 49787 25375 49793
rect 1104 49530 25852 49552
rect 1104 49478 2950 49530
rect 3002 49478 3014 49530
rect 3066 49478 3078 49530
rect 3130 49478 3142 49530
rect 3194 49478 3206 49530
rect 3258 49478 12950 49530
rect 13002 49478 13014 49530
rect 13066 49478 13078 49530
rect 13130 49478 13142 49530
rect 13194 49478 13206 49530
rect 13258 49478 22950 49530
rect 23002 49478 23014 49530
rect 23066 49478 23078 49530
rect 23130 49478 23142 49530
rect 23194 49478 23206 49530
rect 23258 49478 25852 49530
rect 1104 49456 25852 49478
rect 1302 49240 1308 49292
rect 1360 49280 1366 49292
rect 1765 49283 1823 49289
rect 1765 49280 1777 49283
rect 1360 49252 1777 49280
rect 1360 49240 1366 49252
rect 1765 49249 1777 49252
rect 1811 49249 1823 49283
rect 1765 49243 1823 49249
rect 4433 49283 4491 49289
rect 4433 49249 4445 49283
rect 4479 49280 4491 49283
rect 9398 49280 9404 49292
rect 4479 49252 9404 49280
rect 4479 49249 4491 49252
rect 4433 49243 4491 49249
rect 9398 49240 9404 49252
rect 9456 49240 9462 49292
rect 2961 49215 3019 49221
rect 2961 49181 2973 49215
rect 3007 49212 3019 49215
rect 3326 49212 3332 49224
rect 3007 49184 3332 49212
rect 3007 49181 3019 49184
rect 2961 49175 3019 49181
rect 3326 49172 3332 49184
rect 3384 49172 3390 49224
rect 6733 49215 6791 49221
rect 6733 49212 6745 49215
rect 5842 49184 6745 49212
rect 6733 49181 6745 49184
rect 6779 49212 6791 49215
rect 10042 49212 10048 49224
rect 6779 49184 10048 49212
rect 6779 49181 6791 49184
rect 6733 49175 6791 49181
rect 10042 49172 10048 49184
rect 10100 49172 10106 49224
rect 24765 49215 24823 49221
rect 24765 49181 24777 49215
rect 24811 49212 24823 49215
rect 25314 49212 25320 49224
rect 24811 49184 25320 49212
rect 24811 49181 24823 49184
rect 24765 49175 24823 49181
rect 25314 49172 25320 49184
rect 25372 49172 25378 49224
rect 4062 49104 4068 49156
rect 4120 49144 4126 49156
rect 4709 49147 4767 49153
rect 4709 49144 4721 49147
rect 4120 49116 4721 49144
rect 4120 49104 4126 49116
rect 4709 49113 4721 49116
rect 4755 49113 4767 49147
rect 4709 49107 4767 49113
rect 6457 49147 6515 49153
rect 6457 49113 6469 49147
rect 6503 49144 6515 49147
rect 9030 49144 9036 49156
rect 6503 49116 9036 49144
rect 6503 49113 6515 49116
rect 6457 49107 6515 49113
rect 9030 49104 9036 49116
rect 9088 49104 9094 49156
rect 22066 49116 25176 49144
rect 19886 49036 19892 49088
rect 19944 49076 19950 49088
rect 22066 49076 22094 49116
rect 25148 49085 25176 49116
rect 19944 49048 22094 49076
rect 25133 49079 25191 49085
rect 19944 49036 19950 49048
rect 25133 49045 25145 49079
rect 25179 49045 25191 49079
rect 25133 49039 25191 49045
rect 1104 48986 25852 49008
rect 1104 48934 7950 48986
rect 8002 48934 8014 48986
rect 8066 48934 8078 48986
rect 8130 48934 8142 48986
rect 8194 48934 8206 48986
rect 8258 48934 17950 48986
rect 18002 48934 18014 48986
rect 18066 48934 18078 48986
rect 18130 48934 18142 48986
rect 18194 48934 18206 48986
rect 18258 48934 25852 48986
rect 1104 48912 25852 48934
rect 11790 48832 11796 48884
rect 11848 48872 11854 48884
rect 11885 48875 11943 48881
rect 11885 48872 11897 48875
rect 11848 48844 11897 48872
rect 11848 48832 11854 48844
rect 11885 48841 11897 48844
rect 11931 48841 11943 48875
rect 11885 48835 11943 48841
rect 11698 48696 11704 48748
rect 11756 48696 11762 48748
rect 24762 48696 24768 48748
rect 24820 48736 24826 48748
rect 25317 48739 25375 48745
rect 25317 48736 25329 48739
rect 24820 48708 25329 48736
rect 24820 48696 24826 48708
rect 25317 48705 25329 48708
rect 25363 48705 25375 48739
rect 25317 48699 25375 48705
rect 25133 48603 25191 48609
rect 25133 48600 25145 48603
rect 22066 48572 25145 48600
rect 21634 48492 21640 48544
rect 21692 48532 21698 48544
rect 22066 48532 22094 48572
rect 25133 48569 25145 48572
rect 25179 48569 25191 48603
rect 25133 48563 25191 48569
rect 21692 48504 22094 48532
rect 21692 48492 21698 48504
rect 1104 48442 25852 48464
rect 1104 48390 2950 48442
rect 3002 48390 3014 48442
rect 3066 48390 3078 48442
rect 3130 48390 3142 48442
rect 3194 48390 3206 48442
rect 3258 48390 12950 48442
rect 13002 48390 13014 48442
rect 13066 48390 13078 48442
rect 13130 48390 13142 48442
rect 13194 48390 13206 48442
rect 13258 48390 22950 48442
rect 23002 48390 23014 48442
rect 23066 48390 23078 48442
rect 23130 48390 23142 48442
rect 23194 48390 23206 48442
rect 23258 48390 25852 48442
rect 1104 48368 25852 48390
rect 20714 48220 20720 48272
rect 20772 48260 20778 48272
rect 25133 48263 25191 48269
rect 25133 48260 25145 48263
rect 20772 48232 25145 48260
rect 20772 48220 20778 48232
rect 25133 48229 25145 48232
rect 25179 48229 25191 48263
rect 25133 48223 25191 48229
rect 25317 48127 25375 48133
rect 25317 48093 25329 48127
rect 25363 48124 25375 48127
rect 25498 48124 25504 48136
rect 25363 48096 25504 48124
rect 25363 48093 25375 48096
rect 25317 48087 25375 48093
rect 25498 48084 25504 48096
rect 25556 48084 25562 48136
rect 1302 48016 1308 48068
rect 1360 48056 1366 48068
rect 1673 48059 1731 48065
rect 1673 48056 1685 48059
rect 1360 48028 1685 48056
rect 1360 48016 1366 48028
rect 1673 48025 1685 48028
rect 1719 48056 1731 48059
rect 2133 48059 2191 48065
rect 2133 48056 2145 48059
rect 1719 48028 2145 48056
rect 1719 48025 1731 48028
rect 1673 48019 1731 48025
rect 2133 48025 2145 48028
rect 2179 48025 2191 48059
rect 2133 48019 2191 48025
rect 1765 47991 1823 47997
rect 1765 47957 1777 47991
rect 1811 47988 1823 47991
rect 4062 47988 4068 48000
rect 1811 47960 4068 47988
rect 1811 47957 1823 47960
rect 1765 47951 1823 47957
rect 4062 47948 4068 47960
rect 4120 47948 4126 48000
rect 23661 47991 23719 47997
rect 23661 47957 23673 47991
rect 23707 47988 23719 47991
rect 24489 47991 24547 47997
rect 24489 47988 24501 47991
rect 23707 47960 24501 47988
rect 23707 47957 23719 47960
rect 23661 47951 23719 47957
rect 24489 47957 24501 47960
rect 24535 47988 24547 47991
rect 24854 47988 24860 48000
rect 24535 47960 24860 47988
rect 24535 47957 24547 47960
rect 24489 47951 24547 47957
rect 24854 47948 24860 47960
rect 24912 47948 24918 48000
rect 1104 47898 25852 47920
rect 1104 47846 7950 47898
rect 8002 47846 8014 47898
rect 8066 47846 8078 47898
rect 8130 47846 8142 47898
rect 8194 47846 8206 47898
rect 8258 47846 17950 47898
rect 18002 47846 18014 47898
rect 18066 47846 18078 47898
rect 18130 47846 18142 47898
rect 18194 47846 18206 47898
rect 18258 47846 25852 47898
rect 1104 47824 25852 47846
rect 23477 47787 23535 47793
rect 23477 47753 23489 47787
rect 23523 47784 23535 47787
rect 23842 47784 23848 47796
rect 23523 47756 23848 47784
rect 23523 47753 23535 47756
rect 23477 47747 23535 47753
rect 23842 47744 23848 47756
rect 23900 47744 23906 47796
rect 24121 47787 24179 47793
rect 24121 47753 24133 47787
rect 24167 47784 24179 47787
rect 24394 47784 24400 47796
rect 24167 47756 24400 47784
rect 24167 47753 24179 47756
rect 24121 47747 24179 47753
rect 24394 47744 24400 47756
rect 24452 47744 24458 47796
rect 24026 47676 24032 47728
rect 24084 47716 24090 47728
rect 24581 47719 24639 47725
rect 24581 47716 24593 47719
rect 24084 47688 24593 47716
rect 24084 47676 24090 47688
rect 24581 47685 24593 47688
rect 24627 47685 24639 47719
rect 24581 47679 24639 47685
rect 23293 47651 23351 47657
rect 23293 47617 23305 47651
rect 23339 47648 23351 47651
rect 23937 47651 23995 47657
rect 23937 47648 23949 47651
rect 23339 47620 23949 47648
rect 23339 47617 23351 47620
rect 23293 47611 23351 47617
rect 23937 47617 23949 47620
rect 23983 47648 23995 47651
rect 24765 47651 24823 47657
rect 24765 47648 24777 47651
rect 23983 47620 24777 47648
rect 23983 47617 23995 47620
rect 23937 47611 23995 47617
rect 24765 47617 24777 47620
rect 24811 47648 24823 47651
rect 24854 47648 24860 47660
rect 24811 47620 24860 47648
rect 24811 47617 24823 47620
rect 24765 47611 24823 47617
rect 24854 47608 24860 47620
rect 24912 47648 24918 47660
rect 24912 47620 25268 47648
rect 24912 47608 24918 47620
rect 25240 47521 25268 47620
rect 25225 47515 25283 47521
rect 25225 47481 25237 47515
rect 25271 47512 25283 47515
rect 25866 47512 25872 47524
rect 25271 47484 25872 47512
rect 25271 47481 25283 47484
rect 25225 47475 25283 47481
rect 25866 47472 25872 47484
rect 25924 47472 25930 47524
rect 16114 47404 16120 47456
rect 16172 47444 16178 47456
rect 16945 47447 17003 47453
rect 16945 47444 16957 47447
rect 16172 47416 16957 47444
rect 16172 47404 16178 47416
rect 16945 47413 16957 47416
rect 16991 47413 17003 47447
rect 16945 47407 17003 47413
rect 25498 47404 25504 47456
rect 25556 47404 25562 47456
rect 1104 47354 25852 47376
rect 1104 47302 2950 47354
rect 3002 47302 3014 47354
rect 3066 47302 3078 47354
rect 3130 47302 3142 47354
rect 3194 47302 3206 47354
rect 3258 47302 12950 47354
rect 13002 47302 13014 47354
rect 13066 47302 13078 47354
rect 13130 47302 13142 47354
rect 13194 47302 13206 47354
rect 13258 47302 22950 47354
rect 23002 47302 23014 47354
rect 23066 47302 23078 47354
rect 23130 47302 23142 47354
rect 23194 47302 23206 47354
rect 23258 47302 25852 47354
rect 1104 47280 25852 47302
rect 6822 47200 6828 47252
rect 6880 47240 6886 47252
rect 9125 47243 9183 47249
rect 9125 47240 9137 47243
rect 6880 47212 9137 47240
rect 6880 47200 6886 47212
rect 9125 47209 9137 47212
rect 9171 47209 9183 47243
rect 9125 47203 9183 47209
rect 11606 47200 11612 47252
rect 11664 47240 11670 47252
rect 11701 47243 11759 47249
rect 11701 47240 11713 47243
rect 11664 47212 11713 47240
rect 11664 47200 11670 47212
rect 11701 47209 11713 47212
rect 11747 47209 11759 47243
rect 11701 47203 11759 47209
rect 13814 47200 13820 47252
rect 13872 47240 13878 47252
rect 14826 47240 14832 47252
rect 13872 47212 14832 47240
rect 13872 47200 13878 47212
rect 14826 47200 14832 47212
rect 14884 47240 14890 47252
rect 14884 47212 17908 47240
rect 14884 47200 14890 47212
rect 14550 47064 14556 47116
rect 14608 47104 14614 47116
rect 15105 47107 15163 47113
rect 15105 47104 15117 47107
rect 14608 47076 15117 47104
rect 14608 47064 14614 47076
rect 15105 47073 15117 47076
rect 15151 47073 15163 47107
rect 15105 47067 15163 47073
rect 16482 47064 16488 47116
rect 16540 47104 16546 47116
rect 16540 47076 17724 47104
rect 16540 47064 16546 47076
rect 9309 47039 9367 47045
rect 9309 47005 9321 47039
rect 9355 47036 9367 47039
rect 10962 47036 10968 47048
rect 9355 47008 10968 47036
rect 9355 47005 9367 47008
rect 9309 46999 9367 47005
rect 10962 46996 10968 47008
rect 11020 46996 11026 47048
rect 11514 46996 11520 47048
rect 11572 46996 11578 47048
rect 16850 46996 16856 47048
rect 16908 46996 16914 47048
rect 17696 47045 17724 47076
rect 17770 47064 17776 47116
rect 17828 47064 17834 47116
rect 17880 47113 17908 47212
rect 23290 47200 23296 47252
rect 23348 47240 23354 47252
rect 23845 47243 23903 47249
rect 23845 47240 23857 47243
rect 23348 47212 23857 47240
rect 23348 47200 23354 47212
rect 23845 47209 23857 47212
rect 23891 47209 23903 47243
rect 23845 47203 23903 47209
rect 24857 47175 24915 47181
rect 24857 47141 24869 47175
rect 24903 47172 24915 47175
rect 24946 47172 24952 47184
rect 24903 47144 24952 47172
rect 24903 47141 24915 47144
rect 24857 47135 24915 47141
rect 24946 47132 24952 47144
rect 25004 47132 25010 47184
rect 17865 47107 17923 47113
rect 17865 47073 17877 47107
rect 17911 47073 17923 47107
rect 17865 47067 17923 47073
rect 17681 47039 17739 47045
rect 17681 47005 17693 47039
rect 17727 47005 17739 47039
rect 17788 47036 17816 47064
rect 18325 47039 18383 47045
rect 18325 47036 18337 47039
rect 17788 47008 18337 47036
rect 17681 46999 17739 47005
rect 18325 47005 18337 47008
rect 18371 47036 18383 47039
rect 18966 47036 18972 47048
rect 18371 47008 18972 47036
rect 18371 47005 18383 47008
rect 18325 46999 18383 47005
rect 18966 46996 18972 47008
rect 19024 46996 19030 47048
rect 23569 47039 23627 47045
rect 23569 47005 23581 47039
rect 23615 47036 23627 47039
rect 24029 47039 24087 47045
rect 24029 47036 24041 47039
rect 23615 47008 24041 47036
rect 23615 47005 23627 47008
rect 23569 46999 23627 47005
rect 24029 47005 24041 47008
rect 24075 47036 24087 47039
rect 24075 47008 24716 47036
rect 24075 47005 24087 47008
rect 24029 46999 24087 47005
rect 16114 46928 16120 46980
rect 16172 46928 16178 46980
rect 16574 46928 16580 46980
rect 16632 46928 16638 46980
rect 24688 46977 24716 47008
rect 24673 46971 24731 46977
rect 24673 46937 24685 46971
rect 24719 46968 24731 46971
rect 24946 46968 24952 46980
rect 24719 46940 24952 46968
rect 24719 46937 24731 46940
rect 24673 46931 24731 46937
rect 24946 46928 24952 46940
rect 25004 46968 25010 46980
rect 25133 46971 25191 46977
rect 25133 46968 25145 46971
rect 25004 46940 25145 46968
rect 25004 46928 25010 46940
rect 25133 46937 25145 46940
rect 25179 46937 25191 46971
rect 25133 46931 25191 46937
rect 17310 46860 17316 46912
rect 17368 46860 17374 46912
rect 1104 46810 25852 46832
rect 1104 46758 7950 46810
rect 8002 46758 8014 46810
rect 8066 46758 8078 46810
rect 8130 46758 8142 46810
rect 8194 46758 8206 46810
rect 8258 46758 17950 46810
rect 18002 46758 18014 46810
rect 18066 46758 18078 46810
rect 18130 46758 18142 46810
rect 18194 46758 18206 46810
rect 18258 46758 25852 46810
rect 1104 46736 25852 46758
rect 7098 46656 7104 46708
rect 7156 46656 7162 46708
rect 13725 46699 13783 46705
rect 13725 46665 13737 46699
rect 13771 46696 13783 46699
rect 13814 46696 13820 46708
rect 13771 46668 13820 46696
rect 13771 46665 13783 46668
rect 13725 46659 13783 46665
rect 13814 46656 13820 46668
rect 13872 46656 13878 46708
rect 15841 46699 15899 46705
rect 15841 46696 15853 46699
rect 15120 46668 15853 46696
rect 15120 46628 15148 46668
rect 15841 46665 15853 46668
rect 15887 46696 15899 46699
rect 16114 46696 16120 46708
rect 15887 46668 16120 46696
rect 15887 46665 15899 46668
rect 15841 46659 15899 46665
rect 16114 46656 16120 46668
rect 16172 46656 16178 46708
rect 17221 46699 17279 46705
rect 17221 46665 17233 46699
rect 17267 46696 17279 46699
rect 17402 46696 17408 46708
rect 17267 46668 17408 46696
rect 17267 46665 17279 46668
rect 17221 46659 17279 46665
rect 17402 46656 17408 46668
rect 17460 46656 17466 46708
rect 18509 46699 18567 46705
rect 18509 46665 18521 46699
rect 18555 46696 18567 46699
rect 18690 46696 18696 46708
rect 18555 46668 18696 46696
rect 18555 46665 18567 46668
rect 18509 46659 18567 46665
rect 18690 46656 18696 46668
rect 18748 46656 18754 46708
rect 19610 46656 19616 46708
rect 19668 46696 19674 46708
rect 20257 46699 20315 46705
rect 20257 46696 20269 46699
rect 19668 46668 20269 46696
rect 19668 46656 19674 46668
rect 20257 46665 20269 46668
rect 20303 46665 20315 46699
rect 20257 46659 20315 46665
rect 20530 46656 20536 46708
rect 20588 46656 20594 46708
rect 14766 46600 15148 46628
rect 15197 46631 15255 46637
rect 15197 46597 15209 46631
rect 15243 46628 15255 46631
rect 16022 46628 16028 46640
rect 15243 46600 16028 46628
rect 15243 46597 15255 46600
rect 15197 46591 15255 46597
rect 16022 46588 16028 46600
rect 16080 46588 16086 46640
rect 17313 46631 17371 46637
rect 17313 46597 17325 46631
rect 17359 46628 17371 46631
rect 18598 46628 18604 46640
rect 17359 46600 18604 46628
rect 17359 46597 17371 46600
rect 17313 46591 17371 46597
rect 18598 46588 18604 46600
rect 18656 46588 18662 46640
rect 7282 46520 7288 46572
rect 7340 46520 7346 46572
rect 16574 46520 16580 46572
rect 16632 46560 16638 46572
rect 16632 46532 17448 46560
rect 16632 46520 16638 46532
rect 15470 46452 15476 46504
rect 15528 46492 15534 46504
rect 16850 46492 16856 46504
rect 15528 46464 16856 46492
rect 15528 46452 15534 46464
rect 16850 46452 16856 46464
rect 16908 46452 16914 46504
rect 17420 46501 17448 46532
rect 17770 46520 17776 46572
rect 17828 46560 17834 46572
rect 18417 46563 18475 46569
rect 18417 46560 18429 46563
rect 17828 46532 18429 46560
rect 17828 46520 17834 46532
rect 18417 46529 18429 46532
rect 18463 46560 18475 46563
rect 18506 46560 18512 46572
rect 18463 46532 18512 46560
rect 18463 46529 18475 46532
rect 18417 46523 18475 46529
rect 18506 46520 18512 46532
rect 18564 46560 18570 46572
rect 19061 46563 19119 46569
rect 19061 46560 19073 46563
rect 18564 46532 19073 46560
rect 18564 46520 18570 46532
rect 19061 46529 19073 46532
rect 19107 46529 19119 46563
rect 19061 46523 19119 46529
rect 23477 46563 23535 46569
rect 23477 46529 23489 46563
rect 23523 46560 23535 46563
rect 23842 46560 23848 46572
rect 23523 46532 23848 46560
rect 23523 46529 23535 46532
rect 23477 46523 23535 46529
rect 23842 46520 23848 46532
rect 23900 46520 23906 46572
rect 24670 46520 24676 46572
rect 24728 46560 24734 46572
rect 25317 46563 25375 46569
rect 25317 46560 25329 46563
rect 24728 46532 25329 46560
rect 24728 46520 24734 46532
rect 25317 46529 25329 46532
rect 25363 46529 25375 46563
rect 25317 46523 25375 46529
rect 17405 46495 17463 46501
rect 17405 46461 17417 46495
rect 17451 46461 17463 46495
rect 17405 46455 17463 46461
rect 18598 46452 18604 46504
rect 18656 46452 18662 46504
rect 25041 46495 25099 46501
rect 25041 46461 25053 46495
rect 25087 46492 25099 46495
rect 26050 46492 26056 46504
rect 25087 46464 26056 46492
rect 25087 46461 25099 46464
rect 25041 46455 25099 46461
rect 26050 46452 26056 46464
rect 26108 46452 26114 46504
rect 24213 46427 24271 46433
rect 24213 46393 24225 46427
rect 24259 46424 24271 46427
rect 24854 46424 24860 46436
rect 24259 46396 24860 46424
rect 24259 46393 24271 46396
rect 24213 46387 24271 46393
rect 24854 46384 24860 46396
rect 24912 46384 24918 46436
rect 16853 46359 16911 46365
rect 16853 46325 16865 46359
rect 16899 46356 16911 46359
rect 17126 46356 17132 46368
rect 16899 46328 17132 46356
rect 16899 46325 16911 46328
rect 16853 46319 16911 46325
rect 17126 46316 17132 46328
rect 17184 46316 17190 46368
rect 18049 46359 18107 46365
rect 18049 46325 18061 46359
rect 18095 46356 18107 46359
rect 18322 46356 18328 46368
rect 18095 46328 18328 46356
rect 18095 46325 18107 46328
rect 18049 46319 18107 46325
rect 18322 46316 18328 46328
rect 18380 46316 18386 46368
rect 23290 46316 23296 46368
rect 23348 46316 23354 46368
rect 23842 46316 23848 46368
rect 23900 46316 23906 46368
rect 1104 46266 25852 46288
rect 1104 46214 2950 46266
rect 3002 46214 3014 46266
rect 3066 46214 3078 46266
rect 3130 46214 3142 46266
rect 3194 46214 3206 46266
rect 3258 46214 12950 46266
rect 13002 46214 13014 46266
rect 13066 46214 13078 46266
rect 13130 46214 13142 46266
rect 13194 46214 13206 46266
rect 13258 46214 22950 46266
rect 23002 46214 23014 46266
rect 23066 46214 23078 46266
rect 23130 46214 23142 46266
rect 23194 46214 23206 46266
rect 23258 46214 25852 46266
rect 1104 46192 25852 46214
rect 15841 46155 15899 46161
rect 15841 46121 15853 46155
rect 15887 46152 15899 46155
rect 16574 46152 16580 46164
rect 15887 46124 16580 46152
rect 15887 46121 15899 46124
rect 15841 46115 15899 46121
rect 16574 46112 16580 46124
rect 16632 46112 16638 46164
rect 18141 46155 18199 46161
rect 18141 46121 18153 46155
rect 18187 46152 18199 46155
rect 18414 46152 18420 46164
rect 18187 46124 18420 46152
rect 18187 46121 18199 46124
rect 18141 46115 18199 46121
rect 18414 46112 18420 46124
rect 18472 46152 18478 46164
rect 18690 46152 18696 46164
rect 18472 46124 18696 46152
rect 18472 46112 18478 46124
rect 18690 46112 18696 46124
rect 18748 46112 18754 46164
rect 21453 46155 21511 46161
rect 21453 46121 21465 46155
rect 21499 46152 21511 46155
rect 25038 46152 25044 46164
rect 21499 46124 25044 46152
rect 21499 46121 21511 46124
rect 21453 46115 21511 46121
rect 25038 46112 25044 46124
rect 25096 46112 25102 46164
rect 22278 46084 22284 46096
rect 20824 46056 22284 46084
rect 15838 45976 15844 46028
rect 15896 46016 15902 46028
rect 16114 46016 16120 46028
rect 15896 45988 16120 46016
rect 15896 45976 15902 45988
rect 16114 45976 16120 45988
rect 16172 46016 16178 46028
rect 16172 45988 16252 46016
rect 16172 45976 16178 45988
rect 1210 45908 1216 45960
rect 1268 45948 1274 45960
rect 1581 45951 1639 45957
rect 1581 45948 1593 45951
rect 1268 45920 1593 45948
rect 1268 45908 1274 45920
rect 1581 45917 1593 45920
rect 1627 45917 1639 45951
rect 1581 45911 1639 45917
rect 1857 45951 1915 45957
rect 1857 45917 1869 45951
rect 1903 45948 1915 45951
rect 9858 45948 9864 45960
rect 1903 45920 9864 45948
rect 1903 45917 1915 45920
rect 1857 45911 1915 45917
rect 9858 45908 9864 45920
rect 9916 45908 9922 45960
rect 16224 45934 16252 45988
rect 16850 45976 16856 46028
rect 16908 46016 16914 46028
rect 17589 46019 17647 46025
rect 17589 46016 17601 46019
rect 16908 45988 17601 46016
rect 16908 45976 16914 45988
rect 17589 45985 17601 45988
rect 17635 45985 17647 46019
rect 17589 45979 17647 45985
rect 19613 46019 19671 46025
rect 19613 45985 19625 46019
rect 19659 45985 19671 46019
rect 19613 45979 19671 45985
rect 19705 46019 19763 46025
rect 19705 45985 19717 46019
rect 19751 46016 19763 46019
rect 19794 46016 19800 46028
rect 19751 45988 19800 46016
rect 19751 45985 19763 45988
rect 19705 45979 19763 45985
rect 19628 45948 19656 45979
rect 19794 45976 19800 45988
rect 19852 45976 19858 46028
rect 20824 46025 20852 46056
rect 22278 46044 22284 46056
rect 22336 46044 22342 46096
rect 24029 46087 24087 46093
rect 24029 46053 24041 46087
rect 24075 46084 24087 46087
rect 24578 46084 24584 46096
rect 24075 46056 24584 46084
rect 24075 46053 24087 46056
rect 24029 46047 24087 46053
rect 24578 46044 24584 46056
rect 24636 46044 24642 46096
rect 20809 46019 20867 46025
rect 20809 45985 20821 46019
rect 20855 45985 20867 46019
rect 20809 45979 20867 45985
rect 20993 46019 21051 46025
rect 20993 45985 21005 46019
rect 21039 46016 21051 46019
rect 21542 46016 21548 46028
rect 21039 45988 21548 46016
rect 21039 45985 21051 45988
rect 20993 45979 21051 45985
rect 21542 45976 21548 45988
rect 21600 45976 21606 46028
rect 24854 46016 24860 46028
rect 23860 45988 24860 46016
rect 20898 45948 20904 45960
rect 19628 45920 20904 45948
rect 20898 45908 20904 45920
rect 20956 45908 20962 45960
rect 23860 45957 23888 45988
rect 24854 45976 24860 45988
rect 24912 45976 24918 46028
rect 23845 45951 23903 45957
rect 23845 45917 23857 45951
rect 23891 45917 23903 45951
rect 23845 45911 23903 45917
rect 24210 45908 24216 45960
rect 24268 45948 24274 45960
rect 24765 45951 24823 45957
rect 24765 45948 24777 45951
rect 24268 45920 24777 45948
rect 24268 45908 24274 45920
rect 24765 45917 24777 45920
rect 24811 45948 24823 45951
rect 25041 45951 25099 45957
rect 25041 45948 25053 45951
rect 24811 45920 25053 45948
rect 24811 45917 24823 45920
rect 24765 45911 24823 45917
rect 25041 45917 25053 45920
rect 25087 45917 25099 45951
rect 25041 45911 25099 45917
rect 17313 45883 17371 45889
rect 17313 45849 17325 45883
rect 17359 45880 17371 45883
rect 17586 45880 17592 45892
rect 17359 45852 17592 45880
rect 17359 45849 17371 45852
rect 17313 45843 17371 45849
rect 17586 45840 17592 45852
rect 17644 45840 17650 45892
rect 17957 45883 18015 45889
rect 17957 45849 17969 45883
rect 18003 45880 18015 45883
rect 18598 45880 18604 45892
rect 18003 45852 18604 45880
rect 18003 45849 18015 45852
rect 17957 45843 18015 45849
rect 18598 45840 18604 45852
rect 18656 45840 18662 45892
rect 19610 45840 19616 45892
rect 19668 45880 19674 45892
rect 19797 45883 19855 45889
rect 19797 45880 19809 45883
rect 19668 45852 19809 45880
rect 19668 45840 19674 45852
rect 19797 45849 19809 45852
rect 19843 45880 19855 45883
rect 20254 45880 20260 45892
rect 19843 45852 20260 45880
rect 19843 45849 19855 45852
rect 19797 45843 19855 45849
rect 20254 45840 20260 45852
rect 20312 45840 20318 45892
rect 20530 45840 20536 45892
rect 20588 45880 20594 45892
rect 21085 45883 21143 45889
rect 21085 45880 21097 45883
rect 20588 45852 21097 45880
rect 20588 45840 20594 45852
rect 21085 45849 21097 45852
rect 21131 45849 21143 45883
rect 21085 45843 21143 45849
rect 24670 45840 24676 45892
rect 24728 45880 24734 45892
rect 25409 45883 25467 45889
rect 25409 45880 25421 45883
rect 24728 45852 25421 45880
rect 24728 45840 24734 45852
rect 25409 45849 25421 45852
rect 25455 45849 25467 45883
rect 25409 45843 25467 45849
rect 20070 45772 20076 45824
rect 20128 45812 20134 45824
rect 20165 45815 20223 45821
rect 20165 45812 20177 45815
rect 20128 45784 20177 45812
rect 20128 45772 20134 45784
rect 20165 45781 20177 45784
rect 20211 45781 20223 45815
rect 20165 45775 20223 45781
rect 24118 45772 24124 45824
rect 24176 45812 24182 45824
rect 24581 45815 24639 45821
rect 24581 45812 24593 45815
rect 24176 45784 24593 45812
rect 24176 45772 24182 45784
rect 24581 45781 24593 45784
rect 24627 45781 24639 45815
rect 24581 45775 24639 45781
rect 1104 45722 25852 45744
rect 1104 45670 7950 45722
rect 8002 45670 8014 45722
rect 8066 45670 8078 45722
rect 8130 45670 8142 45722
rect 8194 45670 8206 45722
rect 8258 45670 17950 45722
rect 18002 45670 18014 45722
rect 18066 45670 18078 45722
rect 18130 45670 18142 45722
rect 18194 45670 18206 45722
rect 18258 45670 25852 45722
rect 1104 45648 25852 45670
rect 1210 45568 1216 45620
rect 1268 45608 1274 45620
rect 1397 45611 1455 45617
rect 1397 45608 1409 45611
rect 1268 45580 1409 45608
rect 1268 45568 1274 45580
rect 1397 45577 1409 45580
rect 1443 45577 1455 45611
rect 1397 45571 1455 45577
rect 6638 45500 6644 45552
rect 6696 45540 6702 45552
rect 7561 45543 7619 45549
rect 7561 45540 7573 45543
rect 6696 45512 7573 45540
rect 6696 45500 6702 45512
rect 7561 45509 7573 45512
rect 7607 45509 7619 45543
rect 7561 45503 7619 45509
rect 11701 45543 11759 45549
rect 11701 45509 11713 45543
rect 11747 45540 11759 45543
rect 11974 45540 11980 45552
rect 11747 45512 11980 45540
rect 11747 45509 11759 45512
rect 11701 45503 11759 45509
rect 11974 45500 11980 45512
rect 12032 45500 12038 45552
rect 14826 45500 14832 45552
rect 14884 45500 14890 45552
rect 20165 45543 20223 45549
rect 20165 45509 20177 45543
rect 20211 45540 20223 45543
rect 22002 45540 22008 45552
rect 20211 45512 22008 45540
rect 20211 45509 20223 45512
rect 20165 45503 20223 45509
rect 22002 45500 22008 45512
rect 22060 45500 22066 45552
rect 7745 45475 7803 45481
rect 7745 45472 7757 45475
rect 7208 45444 7757 45472
rect 7098 45228 7104 45280
rect 7156 45268 7162 45280
rect 7208 45277 7236 45444
rect 7745 45441 7757 45444
rect 7791 45441 7803 45475
rect 7745 45435 7803 45441
rect 8386 45432 8392 45484
rect 8444 45432 8450 45484
rect 9766 45432 9772 45484
rect 9824 45432 9830 45484
rect 11149 45475 11207 45481
rect 11149 45441 11161 45475
rect 11195 45441 11207 45475
rect 11149 45435 11207 45441
rect 11885 45475 11943 45481
rect 11885 45441 11897 45475
rect 11931 45472 11943 45475
rect 12250 45472 12256 45484
rect 11931 45444 12256 45472
rect 11931 45441 11943 45444
rect 11885 45435 11943 45441
rect 11164 45404 11192 45435
rect 12250 45432 12256 45444
rect 12308 45432 12314 45484
rect 13722 45432 13728 45484
rect 13780 45432 13786 45484
rect 15105 45475 15163 45481
rect 15105 45441 15117 45475
rect 15151 45472 15163 45475
rect 15470 45472 15476 45484
rect 15151 45444 15476 45472
rect 15151 45441 15163 45444
rect 15105 45435 15163 45441
rect 15470 45432 15476 45444
rect 15528 45432 15534 45484
rect 17218 45432 17224 45484
rect 17276 45432 17282 45484
rect 19518 45432 19524 45484
rect 19576 45472 19582 45484
rect 20073 45475 20131 45481
rect 20073 45472 20085 45475
rect 19576 45444 20085 45472
rect 19576 45432 19582 45444
rect 20073 45441 20085 45444
rect 20119 45441 20131 45475
rect 20073 45435 20131 45441
rect 22646 45432 22652 45484
rect 22704 45432 22710 45484
rect 24118 45432 24124 45484
rect 24176 45432 24182 45484
rect 13538 45404 13544 45416
rect 11164 45376 13544 45404
rect 13538 45364 13544 45376
rect 13596 45364 13602 45416
rect 18325 45407 18383 45413
rect 18325 45373 18337 45407
rect 18371 45404 18383 45407
rect 18601 45407 18659 45413
rect 18371 45376 18552 45404
rect 18371 45373 18383 45376
rect 18325 45367 18383 45373
rect 8570 45296 8576 45348
rect 8628 45296 8634 45348
rect 9950 45296 9956 45348
rect 10008 45296 10014 45348
rect 18524 45280 18552 45376
rect 18601 45373 18613 45407
rect 18647 45404 18659 45407
rect 19426 45404 19432 45416
rect 18647 45376 19432 45404
rect 18647 45373 18659 45376
rect 18601 45367 18659 45373
rect 19426 45364 19432 45376
rect 19484 45364 19490 45416
rect 20349 45407 20407 45413
rect 20349 45373 20361 45407
rect 20395 45404 20407 45407
rect 20806 45404 20812 45416
rect 20395 45376 20812 45404
rect 20395 45373 20407 45376
rect 20349 45367 20407 45373
rect 20806 45364 20812 45376
rect 20864 45364 20870 45416
rect 24762 45364 24768 45416
rect 24820 45364 24826 45416
rect 7193 45271 7251 45277
rect 7193 45268 7205 45271
rect 7156 45240 7205 45268
rect 7156 45228 7162 45240
rect 7193 45237 7205 45240
rect 7239 45237 7251 45271
rect 7193 45231 7251 45237
rect 8294 45228 8300 45280
rect 8352 45268 8358 45280
rect 10965 45271 11023 45277
rect 10965 45268 10977 45271
rect 8352 45240 10977 45268
rect 8352 45228 8358 45240
rect 10965 45237 10977 45240
rect 11011 45237 11023 45271
rect 10965 45231 11023 45237
rect 12250 45228 12256 45280
rect 12308 45228 12314 45280
rect 12710 45228 12716 45280
rect 12768 45268 12774 45280
rect 13357 45271 13415 45277
rect 13357 45268 13369 45271
rect 12768 45240 13369 45268
rect 12768 45228 12774 45240
rect 13357 45237 13369 45240
rect 13403 45237 13415 45271
rect 13357 45231 13415 45237
rect 15286 45228 15292 45280
rect 15344 45268 15350 45280
rect 15381 45271 15439 45277
rect 15381 45268 15393 45271
rect 15344 45240 15393 45268
rect 15344 45228 15350 45240
rect 15381 45237 15393 45240
rect 15427 45268 15439 45271
rect 15838 45268 15844 45280
rect 15427 45240 15844 45268
rect 15427 45237 15439 45240
rect 15381 45231 15439 45237
rect 15838 45228 15844 45240
rect 15896 45228 15902 45280
rect 16850 45228 16856 45280
rect 16908 45228 16914 45280
rect 18506 45228 18512 45280
rect 18564 45228 18570 45280
rect 18598 45228 18604 45280
rect 18656 45268 18662 45280
rect 18969 45271 19027 45277
rect 18969 45268 18981 45271
rect 18656 45240 18981 45268
rect 18656 45228 18662 45240
rect 18969 45237 18981 45240
rect 19015 45268 19027 45271
rect 19058 45268 19064 45280
rect 19015 45240 19064 45268
rect 19015 45237 19027 45240
rect 18969 45231 19027 45237
rect 19058 45228 19064 45240
rect 19116 45228 19122 45280
rect 19429 45271 19487 45277
rect 19429 45237 19441 45271
rect 19475 45268 19487 45271
rect 19518 45268 19524 45280
rect 19475 45240 19524 45268
rect 19475 45237 19487 45240
rect 19429 45231 19487 45237
rect 19518 45228 19524 45240
rect 19576 45228 19582 45280
rect 19702 45228 19708 45280
rect 19760 45228 19766 45280
rect 1104 45178 25852 45200
rect 1104 45126 2950 45178
rect 3002 45126 3014 45178
rect 3066 45126 3078 45178
rect 3130 45126 3142 45178
rect 3194 45126 3206 45178
rect 3258 45126 12950 45178
rect 13002 45126 13014 45178
rect 13066 45126 13078 45178
rect 13130 45126 13142 45178
rect 13194 45126 13206 45178
rect 13258 45126 22950 45178
rect 23002 45126 23014 45178
rect 23066 45126 23078 45178
rect 23130 45126 23142 45178
rect 23194 45126 23206 45178
rect 23258 45126 25852 45178
rect 1104 45104 25852 45126
rect 10134 45024 10140 45076
rect 10192 45024 10198 45076
rect 15838 45024 15844 45076
rect 15896 45064 15902 45076
rect 16301 45067 16359 45073
rect 16301 45064 16313 45067
rect 15896 45036 16313 45064
rect 15896 45024 15902 45036
rect 16301 45033 16313 45036
rect 16347 45033 16359 45067
rect 16301 45027 16359 45033
rect 5810 44956 5816 45008
rect 5868 44996 5874 45008
rect 7377 44999 7435 45005
rect 7377 44996 7389 44999
rect 5868 44968 7389 44996
rect 5868 44956 5874 44968
rect 7377 44965 7389 44968
rect 7423 44965 7435 44999
rect 7377 44959 7435 44965
rect 7466 44820 7472 44872
rect 7524 44860 7530 44872
rect 7561 44863 7619 44869
rect 7561 44860 7573 44863
rect 7524 44832 7573 44860
rect 7524 44820 7530 44832
rect 7561 44829 7573 44832
rect 7607 44860 7619 44863
rect 7929 44863 7987 44869
rect 7929 44860 7941 44863
rect 7607 44832 7941 44860
rect 7607 44829 7619 44832
rect 7561 44823 7619 44829
rect 7929 44829 7941 44832
rect 7975 44829 7987 44863
rect 7929 44823 7987 44829
rect 10686 44820 10692 44872
rect 10744 44820 10750 44872
rect 14274 44820 14280 44872
rect 14332 44820 14338 44872
rect 10045 44795 10103 44801
rect 10045 44761 10057 44795
rect 10091 44761 10103 44795
rect 10045 44755 10103 44761
rect 10965 44795 11023 44801
rect 10965 44761 10977 44795
rect 11011 44792 11023 44795
rect 11238 44792 11244 44804
rect 11011 44764 11244 44792
rect 11011 44761 11023 44764
rect 10965 44755 11023 44761
rect 8389 44727 8447 44733
rect 8389 44693 8401 44727
rect 8435 44724 8447 44727
rect 8754 44724 8760 44736
rect 8435 44696 8760 44724
rect 8435 44693 8447 44696
rect 8389 44687 8447 44693
rect 8754 44684 8760 44696
rect 8812 44684 8818 44736
rect 9674 44684 9680 44736
rect 9732 44724 9738 44736
rect 10060 44724 10088 44755
rect 11238 44752 11244 44764
rect 11296 44752 11302 44804
rect 12190 44764 12848 44792
rect 9732 44696 10088 44724
rect 9732 44684 9738 44696
rect 12342 44684 12348 44736
rect 12400 44724 12406 44736
rect 12820 44733 12848 44764
rect 14090 44752 14096 44804
rect 14148 44792 14154 44804
rect 14550 44792 14556 44804
rect 14148 44764 14556 44792
rect 14148 44752 14154 44764
rect 14550 44752 14556 44764
rect 14608 44752 14614 44804
rect 15286 44752 15292 44804
rect 15344 44752 15350 44804
rect 12437 44727 12495 44733
rect 12437 44724 12449 44727
rect 12400 44696 12449 44724
rect 12400 44684 12406 44696
rect 12437 44693 12449 44696
rect 12483 44693 12495 44727
rect 12437 44687 12495 44693
rect 12805 44727 12863 44733
rect 12805 44693 12817 44727
rect 12851 44724 12863 44727
rect 13722 44724 13728 44736
rect 12851 44696 13728 44724
rect 12851 44693 12863 44696
rect 12805 44687 12863 44693
rect 13722 44684 13728 44696
rect 13780 44684 13786 44736
rect 16022 44684 16028 44736
rect 16080 44684 16086 44736
rect 16316 44724 16344 45027
rect 22738 44996 22744 45008
rect 21836 44968 22744 44996
rect 21836 44937 21864 44968
rect 22738 44956 22744 44968
rect 22796 44956 22802 45008
rect 21821 44931 21879 44937
rect 21821 44897 21833 44931
rect 21867 44897 21879 44931
rect 21821 44891 21879 44897
rect 21910 44888 21916 44940
rect 21968 44888 21974 44940
rect 23385 44931 23443 44937
rect 23385 44897 23397 44931
rect 23431 44928 23443 44931
rect 24118 44928 24124 44940
rect 23431 44900 24124 44928
rect 23431 44897 23443 44900
rect 23385 44891 23443 44897
rect 24118 44888 24124 44900
rect 24176 44888 24182 44940
rect 21174 44820 21180 44872
rect 21232 44820 21238 44872
rect 22646 44820 22652 44872
rect 22704 44860 22710 44872
rect 23201 44863 23259 44869
rect 23201 44860 23213 44863
rect 22704 44832 23213 44860
rect 22704 44820 22710 44832
rect 23201 44829 23213 44832
rect 23247 44829 23259 44863
rect 23201 44823 23259 44829
rect 23293 44863 23351 44869
rect 23293 44829 23305 44863
rect 23339 44860 23351 44863
rect 24486 44860 24492 44872
rect 23339 44832 24492 44860
rect 23339 44829 23351 44832
rect 23293 44823 23351 44829
rect 24486 44820 24492 44832
rect 24544 44820 24550 44872
rect 24857 44863 24915 44869
rect 24857 44829 24869 44863
rect 24903 44860 24915 44863
rect 25314 44860 25320 44872
rect 24903 44832 25320 44860
rect 24903 44829 24915 44832
rect 24857 44823 24915 44829
rect 25314 44820 25320 44832
rect 25372 44820 25378 44872
rect 20470 44764 20760 44792
rect 17218 44724 17224 44736
rect 16316 44696 17224 44724
rect 17218 44684 17224 44696
rect 17276 44724 17282 44736
rect 17494 44724 17500 44736
rect 17276 44696 17500 44724
rect 17276 44684 17282 44696
rect 17494 44684 17500 44696
rect 17552 44684 17558 44736
rect 19334 44684 19340 44736
rect 19392 44724 19398 44736
rect 19429 44727 19487 44733
rect 19429 44724 19441 44727
rect 19392 44696 19441 44724
rect 19392 44684 19398 44696
rect 19429 44693 19441 44696
rect 19475 44693 19487 44727
rect 20732 44724 20760 44764
rect 20898 44752 20904 44804
rect 20956 44752 20962 44804
rect 21082 44724 21088 44736
rect 20732 44696 21088 44724
rect 19429 44687 19487 44693
rect 21082 44684 21088 44696
rect 21140 44684 21146 44736
rect 21450 44684 21456 44736
rect 21508 44724 21514 44736
rect 22005 44727 22063 44733
rect 22005 44724 22017 44727
rect 21508 44696 22017 44724
rect 21508 44684 21514 44696
rect 22005 44693 22017 44696
rect 22051 44693 22063 44727
rect 22005 44687 22063 44693
rect 22373 44727 22431 44733
rect 22373 44693 22385 44727
rect 22419 44724 22431 44727
rect 22462 44724 22468 44736
rect 22419 44696 22468 44724
rect 22419 44693 22431 44696
rect 22373 44687 22431 44693
rect 22462 44684 22468 44696
rect 22520 44684 22526 44736
rect 22830 44684 22836 44736
rect 22888 44684 22894 44736
rect 23566 44684 23572 44736
rect 23624 44724 23630 44736
rect 25133 44727 25191 44733
rect 25133 44724 25145 44727
rect 23624 44696 25145 44724
rect 23624 44684 23630 44696
rect 25133 44693 25145 44696
rect 25179 44693 25191 44727
rect 25133 44687 25191 44693
rect 1104 44634 25852 44656
rect 1104 44582 7950 44634
rect 8002 44582 8014 44634
rect 8066 44582 8078 44634
rect 8130 44582 8142 44634
rect 8194 44582 8206 44634
rect 8258 44582 17950 44634
rect 18002 44582 18014 44634
rect 18066 44582 18078 44634
rect 18130 44582 18142 44634
rect 18194 44582 18206 44634
rect 18258 44582 25852 44634
rect 1104 44560 25852 44582
rect 7190 44480 7196 44532
rect 7248 44480 7254 44532
rect 7742 44480 7748 44532
rect 7800 44520 7806 44532
rect 8021 44523 8079 44529
rect 8021 44520 8033 44523
rect 7800 44492 8033 44520
rect 7800 44480 7806 44492
rect 8021 44489 8033 44492
rect 8067 44489 8079 44523
rect 8021 44483 8079 44489
rect 9030 44480 9036 44532
rect 9088 44520 9094 44532
rect 9214 44520 9220 44532
rect 9088 44492 9220 44520
rect 9088 44480 9094 44492
rect 9214 44480 9220 44492
rect 9272 44520 9278 44532
rect 9272 44492 9720 44520
rect 9272 44480 9278 44492
rect 6825 44455 6883 44461
rect 6825 44421 6837 44455
rect 6871 44452 6883 44455
rect 7285 44455 7343 44461
rect 7285 44452 7297 44455
rect 6871 44424 7297 44452
rect 6871 44421 6883 44424
rect 6825 44415 6883 44421
rect 7285 44421 7297 44424
rect 7331 44452 7343 44455
rect 7331 44424 8432 44452
rect 7331 44421 7343 44424
rect 7285 44415 7343 44421
rect 7742 44344 7748 44396
rect 7800 44384 7806 44396
rect 7837 44387 7895 44393
rect 7837 44384 7849 44387
rect 7800 44356 7849 44384
rect 7800 44344 7806 44356
rect 7837 44353 7849 44356
rect 7883 44353 7895 44387
rect 8404 44384 8432 44424
rect 8478 44412 8484 44464
rect 8536 44412 8542 44464
rect 9692 44461 9720 44492
rect 10042 44480 10048 44532
rect 10100 44480 10106 44532
rect 11698 44480 11704 44532
rect 11756 44480 11762 44532
rect 13630 44480 13636 44532
rect 13688 44520 13694 44532
rect 14553 44523 14611 44529
rect 14553 44520 14565 44523
rect 13688 44492 14565 44520
rect 13688 44480 13694 44492
rect 14553 44489 14565 44492
rect 14599 44489 14611 44523
rect 17034 44520 17040 44532
rect 14553 44483 14611 44489
rect 16546 44492 17040 44520
rect 9677 44455 9735 44461
rect 9677 44421 9689 44455
rect 9723 44421 9735 44455
rect 10060 44452 10088 44480
rect 10060 44424 10166 44452
rect 9677 44415 9735 44421
rect 11054 44412 11060 44464
rect 11112 44452 11118 44464
rect 12897 44455 12955 44461
rect 12897 44452 12909 44455
rect 11112 44424 12909 44452
rect 11112 44412 11118 44424
rect 12897 44421 12909 44424
rect 12943 44421 12955 44455
rect 12897 44415 12955 44421
rect 8665 44387 8723 44393
rect 8404 44356 8524 44384
rect 7837 44347 7895 44353
rect 6730 44276 6736 44328
rect 6788 44316 6794 44328
rect 8294 44316 8300 44328
rect 6788 44288 8300 44316
rect 6788 44276 6794 44288
rect 8294 44276 8300 44288
rect 8352 44276 8358 44328
rect 8496 44316 8524 44356
rect 8665 44353 8677 44387
rect 8711 44384 8723 44387
rect 8754 44384 8760 44396
rect 8711 44356 8760 44384
rect 8711 44353 8723 44356
rect 8665 44347 8723 44353
rect 8754 44344 8760 44356
rect 8812 44344 8818 44396
rect 9398 44344 9404 44396
rect 9456 44344 9462 44396
rect 12069 44387 12127 44393
rect 12069 44353 12081 44387
rect 12115 44384 12127 44387
rect 12618 44384 12624 44396
rect 12115 44356 12624 44384
rect 12115 44353 12127 44356
rect 12069 44347 12127 44353
rect 12618 44344 12624 44356
rect 12676 44344 12682 44396
rect 13081 44387 13139 44393
rect 13081 44353 13093 44387
rect 13127 44384 13139 44387
rect 13127 44356 13584 44384
rect 13127 44353 13139 44356
rect 13081 44347 13139 44353
rect 11330 44316 11336 44328
rect 8496 44288 11336 44316
rect 11330 44276 11336 44288
rect 11388 44276 11394 44328
rect 12158 44276 12164 44328
rect 12216 44276 12222 44328
rect 12342 44276 12348 44328
rect 12400 44276 12406 44328
rect 11149 44183 11207 44189
rect 11149 44149 11161 44183
rect 11195 44180 11207 44183
rect 11238 44180 11244 44192
rect 11195 44152 11244 44180
rect 11195 44149 11207 44152
rect 11149 44143 11207 44149
rect 11238 44140 11244 44152
rect 11296 44180 11302 44192
rect 11882 44180 11888 44192
rect 11296 44152 11888 44180
rect 11296 44140 11302 44152
rect 11882 44140 11888 44152
rect 11940 44140 11946 44192
rect 13556 44189 13584 44356
rect 14369 44319 14427 44325
rect 14369 44285 14381 44319
rect 14415 44285 14427 44319
rect 14369 44279 14427 44285
rect 14461 44319 14519 44325
rect 14461 44285 14473 44319
rect 14507 44316 14519 44319
rect 15197 44319 15255 44325
rect 15197 44316 15209 44319
rect 14507 44288 15209 44316
rect 14507 44285 14519 44288
rect 14461 44279 14519 44285
rect 15197 44285 15209 44288
rect 15243 44316 15255 44319
rect 15930 44316 15936 44328
rect 15243 44288 15936 44316
rect 15243 44285 15255 44288
rect 15197 44279 15255 44285
rect 14384 44248 14412 44279
rect 15930 44276 15936 44288
rect 15988 44316 15994 44328
rect 16546 44316 16574 44492
rect 17034 44480 17040 44492
rect 17092 44480 17098 44532
rect 17681 44523 17739 44529
rect 17681 44489 17693 44523
rect 17727 44520 17739 44523
rect 18506 44520 18512 44532
rect 17727 44492 18512 44520
rect 17727 44489 17739 44492
rect 17681 44483 17739 44489
rect 18506 44480 18512 44492
rect 18564 44480 18570 44532
rect 24121 44523 24179 44529
rect 24121 44489 24133 44523
rect 24167 44520 24179 44523
rect 24210 44520 24216 44532
rect 24167 44492 24216 44520
rect 24167 44489 24179 44492
rect 24121 44483 24179 44489
rect 24210 44480 24216 44492
rect 24268 44480 24274 44532
rect 19153 44455 19211 44461
rect 19153 44421 19165 44455
rect 19199 44452 19211 44455
rect 19610 44452 19616 44464
rect 19199 44424 19616 44452
rect 19199 44421 19211 44424
rect 19153 44415 19211 44421
rect 19610 44412 19616 44424
rect 19668 44412 19674 44464
rect 21082 44412 21088 44464
rect 21140 44452 21146 44464
rect 21140 44424 22310 44452
rect 21140 44412 21146 44424
rect 18046 44344 18052 44396
rect 18104 44344 18110 44396
rect 25041 44387 25099 44393
rect 25041 44353 25053 44387
rect 25087 44384 25099 44387
rect 25958 44384 25964 44396
rect 25087 44356 25964 44384
rect 25087 44353 25099 44356
rect 25041 44347 25099 44353
rect 25958 44344 25964 44356
rect 26016 44344 26022 44396
rect 15988 44288 16574 44316
rect 15988 44276 15994 44288
rect 19426 44276 19432 44328
rect 19484 44276 19490 44328
rect 21450 44276 21456 44328
rect 21508 44276 21514 44328
rect 22094 44276 22100 44328
rect 22152 44316 22158 44328
rect 23477 44319 23535 44325
rect 23477 44316 23489 44319
rect 22152 44288 23489 44316
rect 22152 44276 22158 44288
rect 23477 44285 23489 44288
rect 23523 44285 23535 44319
rect 23477 44279 23535 44285
rect 23750 44276 23756 44328
rect 23808 44276 23814 44328
rect 25317 44319 25375 44325
rect 25317 44285 25329 44319
rect 25363 44316 25375 44319
rect 25498 44316 25504 44328
rect 25363 44288 25504 44316
rect 25363 44285 25375 44288
rect 25317 44279 25375 44285
rect 25498 44276 25504 44288
rect 25556 44276 25562 44328
rect 14550 44248 14556 44260
rect 14384 44220 14556 44248
rect 14550 44208 14556 44220
rect 14608 44208 14614 44260
rect 14921 44251 14979 44257
rect 14921 44217 14933 44251
rect 14967 44248 14979 44251
rect 15378 44248 15384 44260
rect 14967 44220 15384 44248
rect 14967 44217 14979 44220
rect 14921 44211 14979 44217
rect 15378 44208 15384 44220
rect 15436 44208 15442 44260
rect 20806 44208 20812 44260
rect 20864 44248 20870 44260
rect 22005 44251 22063 44257
rect 22005 44248 22017 44251
rect 20864 44220 22017 44248
rect 20864 44208 20870 44220
rect 22005 44217 22017 44220
rect 22051 44217 22063 44251
rect 22005 44211 22063 44217
rect 13541 44183 13599 44189
rect 13541 44149 13553 44183
rect 13587 44180 13599 44183
rect 14182 44180 14188 44192
rect 13587 44152 14188 44180
rect 13587 44149 13599 44152
rect 13541 44143 13599 44149
rect 14182 44140 14188 44152
rect 14240 44140 14246 44192
rect 19058 44140 19064 44192
rect 19116 44180 19122 44192
rect 19797 44183 19855 44189
rect 19797 44180 19809 44183
rect 19116 44152 19809 44180
rect 19116 44140 19122 44152
rect 19797 44149 19809 44152
rect 19843 44180 19855 44183
rect 21082 44180 21088 44192
rect 19843 44152 21088 44180
rect 19843 44149 19855 44152
rect 19797 44143 19855 44149
rect 21082 44140 21088 44152
rect 21140 44180 21146 44192
rect 21269 44183 21327 44189
rect 21269 44180 21281 44183
rect 21140 44152 21281 44180
rect 21140 44140 21146 44152
rect 21269 44149 21281 44152
rect 21315 44149 21327 44183
rect 21269 44143 21327 44149
rect 1104 44090 25852 44112
rect 1104 44038 2950 44090
rect 3002 44038 3014 44090
rect 3066 44038 3078 44090
rect 3130 44038 3142 44090
rect 3194 44038 3206 44090
rect 3258 44038 12950 44090
rect 13002 44038 13014 44090
rect 13066 44038 13078 44090
rect 13130 44038 13142 44090
rect 13194 44038 13206 44090
rect 13258 44038 22950 44090
rect 23002 44038 23014 44090
rect 23066 44038 23078 44090
rect 23130 44038 23142 44090
rect 23194 44038 23206 44090
rect 23258 44038 25852 44090
rect 1104 44016 25852 44038
rect 9122 43936 9128 43988
rect 9180 43976 9186 43988
rect 10505 43979 10563 43985
rect 10505 43976 10517 43979
rect 9180 43948 10517 43976
rect 9180 43936 9186 43948
rect 10505 43945 10517 43948
rect 10551 43945 10563 43979
rect 10505 43939 10563 43945
rect 20898 43936 20904 43988
rect 20956 43976 20962 43988
rect 21177 43979 21235 43985
rect 21177 43976 21189 43979
rect 20956 43948 21189 43976
rect 20956 43936 20962 43948
rect 21177 43945 21189 43948
rect 21223 43945 21235 43979
rect 21177 43939 21235 43945
rect 22005 43979 22063 43985
rect 22005 43945 22017 43979
rect 22051 43976 22063 43979
rect 22094 43976 22100 43988
rect 22051 43948 22100 43976
rect 22051 43945 22063 43948
rect 22005 43939 22063 43945
rect 22094 43936 22100 43948
rect 22152 43936 22158 43988
rect 24121 43979 24179 43985
rect 24121 43945 24133 43979
rect 24167 43976 24179 43979
rect 24210 43976 24216 43988
rect 24167 43948 24216 43976
rect 24167 43945 24179 43948
rect 24121 43939 24179 43945
rect 24210 43936 24216 43948
rect 24268 43936 24274 43988
rect 24762 43936 24768 43988
rect 24820 43976 24826 43988
rect 25041 43979 25099 43985
rect 25041 43976 25053 43979
rect 24820 43948 25053 43976
rect 24820 43936 24826 43948
rect 25041 43945 25053 43948
rect 25087 43945 25099 43979
rect 25041 43939 25099 43945
rect 6178 43868 6184 43920
rect 6236 43908 6242 43920
rect 6365 43911 6423 43917
rect 6365 43908 6377 43911
rect 6236 43880 6377 43908
rect 6236 43868 6242 43880
rect 6365 43877 6377 43880
rect 6411 43877 6423 43911
rect 6365 43871 6423 43877
rect 7834 43868 7840 43920
rect 7892 43908 7898 43920
rect 8297 43911 8355 43917
rect 8297 43908 8309 43911
rect 7892 43880 8309 43908
rect 7892 43868 7898 43880
rect 8297 43877 8309 43880
rect 8343 43877 8355 43911
rect 8297 43871 8355 43877
rect 9490 43868 9496 43920
rect 9548 43908 9554 43920
rect 9677 43911 9735 43917
rect 9677 43908 9689 43911
rect 9548 43880 9689 43908
rect 9548 43868 9554 43880
rect 9677 43877 9689 43880
rect 9723 43877 9735 43911
rect 24581 43911 24639 43917
rect 24581 43908 24593 43911
rect 9677 43871 9735 43877
rect 23676 43880 24593 43908
rect 9033 43843 9091 43849
rect 9033 43809 9045 43843
rect 9079 43840 9091 43843
rect 14918 43840 14924 43852
rect 9079 43812 14924 43840
rect 9079 43809 9091 43812
rect 9033 43803 9091 43809
rect 1302 43732 1308 43784
rect 1360 43772 1366 43784
rect 1581 43775 1639 43781
rect 1581 43772 1593 43775
rect 1360 43744 1593 43772
rect 1360 43732 1366 43744
rect 1581 43741 1593 43744
rect 1627 43772 1639 43775
rect 2041 43775 2099 43781
rect 2041 43772 2053 43775
rect 1627 43744 2053 43772
rect 1627 43741 1639 43744
rect 1581 43735 1639 43741
rect 2041 43741 2053 43744
rect 2087 43741 2099 43775
rect 2041 43735 2099 43741
rect 8481 43775 8539 43781
rect 8481 43741 8493 43775
rect 8527 43772 8539 43775
rect 9048 43772 9076 43803
rect 14918 43800 14924 43812
rect 14976 43800 14982 43852
rect 15470 43800 15476 43852
rect 15528 43840 15534 43852
rect 15841 43843 15899 43849
rect 15841 43840 15853 43843
rect 15528 43812 15853 43840
rect 15528 43800 15534 43812
rect 15841 43809 15853 43812
rect 15887 43809 15899 43843
rect 15841 43803 15899 43809
rect 18598 43800 18604 43852
rect 18656 43840 18662 43852
rect 23676 43840 23704 43880
rect 24581 43877 24593 43880
rect 24627 43877 24639 43911
rect 24581 43871 24639 43877
rect 18656 43812 23704 43840
rect 18656 43800 18662 43812
rect 23750 43800 23756 43852
rect 23808 43840 23814 43852
rect 25038 43840 25044 43852
rect 23808 43812 25044 43840
rect 23808 43800 23814 43812
rect 25038 43800 25044 43812
rect 25096 43800 25102 43852
rect 8527 43744 9076 43772
rect 9401 43775 9459 43781
rect 8527 43741 8539 43744
rect 8481 43735 8539 43741
rect 9401 43741 9413 43775
rect 9447 43772 9459 43775
rect 9861 43775 9919 43781
rect 9861 43772 9873 43775
rect 9447 43744 9873 43772
rect 9447 43741 9459 43744
rect 9401 43735 9459 43741
rect 9861 43741 9873 43744
rect 9907 43772 9919 43775
rect 10502 43772 10508 43784
rect 9907 43744 10508 43772
rect 9907 43741 9919 43744
rect 9861 43735 9919 43741
rect 10502 43732 10508 43744
rect 10560 43732 10566 43784
rect 10686 43732 10692 43784
rect 10744 43772 10750 43784
rect 11790 43772 11796 43784
rect 10744 43744 11796 43772
rect 10744 43732 10750 43744
rect 11790 43732 11796 43744
rect 11848 43732 11854 43784
rect 19426 43732 19432 43784
rect 19484 43732 19490 43784
rect 20806 43732 20812 43784
rect 20864 43772 20870 43784
rect 21082 43772 21088 43784
rect 20864 43744 21088 43772
rect 20864 43732 20870 43744
rect 21082 43732 21088 43744
rect 21140 43772 21146 43784
rect 21453 43775 21511 43781
rect 21453 43772 21465 43775
rect 21140 43744 21465 43772
rect 21140 43732 21146 43744
rect 21453 43741 21465 43744
rect 21499 43772 21511 43775
rect 22002 43772 22008 43784
rect 21499 43744 22008 43772
rect 21499 43741 21511 43744
rect 21453 43735 21511 43741
rect 22002 43732 22008 43744
rect 22060 43772 22066 43784
rect 22060 43744 22402 43772
rect 22060 43732 22066 43744
rect 24762 43732 24768 43784
rect 24820 43732 24826 43784
rect 6549 43707 6607 43713
rect 6549 43673 6561 43707
rect 6595 43673 6607 43707
rect 6549 43667 6607 43673
rect 10597 43707 10655 43713
rect 10597 43673 10609 43707
rect 10643 43704 10655 43707
rect 11057 43707 11115 43713
rect 11057 43704 11069 43707
rect 10643 43676 11069 43704
rect 10643 43673 10655 43676
rect 10597 43667 10655 43673
rect 11057 43673 11069 43676
rect 11103 43704 11115 43707
rect 11698 43704 11704 43716
rect 11103 43676 11704 43704
rect 11103 43673 11115 43676
rect 11057 43667 11115 43673
rect 1762 43596 1768 43648
rect 1820 43596 1826 43648
rect 6564 43636 6592 43667
rect 11698 43664 11704 43676
rect 11756 43664 11762 43716
rect 12069 43707 12127 43713
rect 12069 43673 12081 43707
rect 12115 43704 12127 43707
rect 12342 43704 12348 43716
rect 12115 43676 12348 43704
rect 12115 43673 12127 43676
rect 12069 43667 12127 43673
rect 12342 43664 12348 43676
rect 12400 43664 12406 43716
rect 13294 43676 13768 43704
rect 13740 43648 13768 43676
rect 15838 43664 15844 43716
rect 15896 43704 15902 43716
rect 16117 43707 16175 43713
rect 16117 43704 16129 43707
rect 15896 43676 16129 43704
rect 15896 43664 15902 43676
rect 16117 43673 16129 43676
rect 16163 43673 16175 43707
rect 17494 43704 17500 43716
rect 17342 43676 17500 43704
rect 16117 43667 16175 43673
rect 17494 43664 17500 43676
rect 17552 43704 17558 43716
rect 17957 43707 18015 43713
rect 17957 43704 17969 43707
rect 17552 43676 17969 43704
rect 17552 43664 17558 43676
rect 17957 43673 17969 43676
rect 18003 43704 18015 43707
rect 18046 43704 18052 43716
rect 18003 43676 18052 43704
rect 18003 43673 18015 43676
rect 17957 43667 18015 43673
rect 18046 43664 18052 43676
rect 18104 43664 18110 43716
rect 19705 43707 19763 43713
rect 19705 43673 19717 43707
rect 19751 43704 19763 43707
rect 19978 43704 19984 43716
rect 19751 43676 19984 43704
rect 19751 43673 19763 43676
rect 19705 43667 19763 43673
rect 19978 43664 19984 43676
rect 20036 43664 20042 43716
rect 23477 43707 23535 43713
rect 23477 43673 23489 43707
rect 23523 43704 23535 43707
rect 23750 43704 23756 43716
rect 23523 43676 23756 43704
rect 23523 43673 23535 43676
rect 23477 43667 23535 43673
rect 23750 43664 23756 43676
rect 23808 43664 23814 43716
rect 7009 43639 7067 43645
rect 7009 43636 7021 43639
rect 6564 43608 7021 43636
rect 7009 43605 7021 43608
rect 7055 43636 7067 43639
rect 9122 43636 9128 43648
rect 7055 43608 9128 43636
rect 7055 43605 7067 43608
rect 7009 43599 7067 43605
rect 9122 43596 9128 43608
rect 9180 43596 9186 43648
rect 10778 43596 10784 43648
rect 10836 43636 10842 43648
rect 11241 43639 11299 43645
rect 11241 43636 11253 43639
rect 10836 43608 11253 43636
rect 10836 43596 10842 43608
rect 11241 43605 11253 43608
rect 11287 43605 11299 43639
rect 11241 43599 11299 43605
rect 13541 43639 13599 43645
rect 13541 43605 13553 43639
rect 13587 43636 13599 43639
rect 13630 43636 13636 43648
rect 13587 43608 13636 43636
rect 13587 43605 13599 43608
rect 13541 43599 13599 43605
rect 13630 43596 13636 43608
rect 13688 43596 13694 43648
rect 13722 43596 13728 43648
rect 13780 43636 13786 43648
rect 14093 43639 14151 43645
rect 14093 43636 14105 43639
rect 13780 43608 14105 43636
rect 13780 43596 13786 43608
rect 14093 43605 14105 43608
rect 14139 43605 14151 43639
rect 14093 43599 14151 43605
rect 17586 43596 17592 43648
rect 17644 43596 17650 43648
rect 25498 43596 25504 43648
rect 25556 43596 25562 43648
rect 1104 43546 25852 43568
rect 1104 43494 7950 43546
rect 8002 43494 8014 43546
rect 8066 43494 8078 43546
rect 8130 43494 8142 43546
rect 8194 43494 8206 43546
rect 8258 43494 17950 43546
rect 18002 43494 18014 43546
rect 18066 43494 18078 43546
rect 18130 43494 18142 43546
rect 18194 43494 18206 43546
rect 18258 43494 25852 43546
rect 1104 43472 25852 43494
rect 1762 43392 1768 43444
rect 1820 43432 1826 43444
rect 2041 43435 2099 43441
rect 2041 43432 2053 43435
rect 1820 43404 2053 43432
rect 1820 43392 1826 43404
rect 2041 43401 2053 43404
rect 2087 43401 2099 43435
rect 2041 43395 2099 43401
rect 5721 43435 5779 43441
rect 5721 43401 5733 43435
rect 5767 43432 5779 43435
rect 6546 43432 6552 43444
rect 5767 43404 6552 43432
rect 5767 43401 5779 43404
rect 5721 43395 5779 43401
rect 6546 43392 6552 43404
rect 6604 43392 6610 43444
rect 8662 43392 8668 43444
rect 8720 43392 8726 43444
rect 12158 43392 12164 43444
rect 12216 43432 12222 43444
rect 12253 43435 12311 43441
rect 12253 43432 12265 43435
rect 12216 43404 12265 43432
rect 12216 43392 12222 43404
rect 12253 43401 12265 43404
rect 12299 43401 12311 43435
rect 12253 43395 12311 43401
rect 17126 43392 17132 43444
rect 17184 43432 17190 43444
rect 17313 43435 17371 43441
rect 17313 43432 17325 43435
rect 17184 43404 17325 43432
rect 17184 43392 17190 43404
rect 17313 43401 17325 43404
rect 17359 43401 17371 43435
rect 17313 43395 17371 43401
rect 17957 43435 18015 43441
rect 17957 43401 17969 43435
rect 18003 43432 18015 43435
rect 19886 43432 19892 43444
rect 18003 43404 19892 43432
rect 18003 43401 18015 43404
rect 17957 43395 18015 43401
rect 10042 43364 10048 43376
rect 9706 43336 10048 43364
rect 10042 43324 10048 43336
rect 10100 43364 10106 43376
rect 10778 43364 10784 43376
rect 10100 43336 10784 43364
rect 10100 43324 10106 43336
rect 10778 43324 10784 43336
rect 10836 43324 10842 43376
rect 17221 43367 17279 43373
rect 17221 43333 17233 43367
rect 17267 43364 17279 43367
rect 17972 43364 18000 43395
rect 19886 43392 19892 43404
rect 19944 43392 19950 43444
rect 22002 43392 22008 43444
rect 22060 43432 22066 43444
rect 22060 43404 23612 43432
rect 22060 43392 22066 43404
rect 17267 43336 18000 43364
rect 17267 43333 17279 43336
rect 17221 43327 17279 43333
rect 22278 43324 22284 43376
rect 22336 43364 22342 43376
rect 22554 43364 22560 43376
rect 22336 43336 22560 43364
rect 22336 43324 22342 43336
rect 22554 43324 22560 43336
rect 22612 43324 22618 43376
rect 23584 43364 23612 43404
rect 23750 43392 23756 43444
rect 23808 43432 23814 43444
rect 24394 43432 24400 43444
rect 23808 43404 24400 43432
rect 23808 43392 23814 43404
rect 24394 43392 24400 43404
rect 24452 43392 24458 43444
rect 23658 43364 23664 43376
rect 23506 43336 23664 43364
rect 23658 43324 23664 43336
rect 23716 43364 23722 43376
rect 24210 43364 24216 43376
rect 23716 43336 24216 43364
rect 23716 43324 23722 43336
rect 24210 43324 24216 43336
rect 24268 43364 24274 43376
rect 24305 43367 24363 43373
rect 24305 43364 24317 43367
rect 24268 43336 24317 43364
rect 24268 43324 24274 43336
rect 24305 43333 24317 43336
rect 24351 43333 24363 43367
rect 24305 43327 24363 43333
rect 2225 43299 2283 43305
rect 2225 43265 2237 43299
rect 2271 43296 2283 43299
rect 2501 43299 2559 43305
rect 2501 43296 2513 43299
rect 2271 43268 2513 43296
rect 2271 43265 2283 43268
rect 2225 43259 2283 43265
rect 2501 43265 2513 43268
rect 2547 43296 2559 43299
rect 4982 43296 4988 43308
rect 2547 43268 4988 43296
rect 2547 43265 2559 43268
rect 2501 43259 2559 43265
rect 4982 43256 4988 43268
rect 5040 43256 5046 43308
rect 5166 43256 5172 43308
rect 5224 43296 5230 43308
rect 5537 43299 5595 43305
rect 5537 43296 5549 43299
rect 5224 43268 5549 43296
rect 5224 43256 5230 43268
rect 5537 43265 5549 43268
rect 5583 43265 5595 43299
rect 5537 43259 5595 43265
rect 10413 43299 10471 43305
rect 10413 43265 10425 43299
rect 10459 43296 10471 43299
rect 10686 43296 10692 43308
rect 10459 43268 10692 43296
rect 10459 43265 10471 43268
rect 10413 43259 10471 43265
rect 10686 43256 10692 43268
rect 10744 43256 10750 43308
rect 12621 43299 12679 43305
rect 12621 43265 12633 43299
rect 12667 43296 12679 43299
rect 15654 43296 15660 43308
rect 12667 43268 15660 43296
rect 12667 43265 12679 43268
rect 12621 43259 12679 43265
rect 15654 43256 15660 43268
rect 15712 43256 15718 43308
rect 25317 43299 25375 43305
rect 25317 43265 25329 43299
rect 25363 43296 25375 43299
rect 25406 43296 25412 43308
rect 25363 43268 25412 43296
rect 25363 43265 25375 43268
rect 25317 43259 25375 43265
rect 25406 43256 25412 43268
rect 25464 43256 25470 43308
rect 10137 43231 10195 43237
rect 10137 43197 10149 43231
rect 10183 43228 10195 43231
rect 10778 43228 10784 43240
rect 10183 43200 10784 43228
rect 10183 43197 10195 43200
rect 10137 43191 10195 43197
rect 10778 43188 10784 43200
rect 10836 43188 10842 43240
rect 11054 43188 11060 43240
rect 11112 43228 11118 43240
rect 12713 43231 12771 43237
rect 12713 43228 12725 43231
rect 11112 43200 12725 43228
rect 11112 43188 11118 43200
rect 12713 43197 12725 43200
rect 12759 43197 12771 43231
rect 12713 43191 12771 43197
rect 12805 43231 12863 43237
rect 12805 43197 12817 43231
rect 12851 43197 12863 43231
rect 12805 43191 12863 43197
rect 17405 43231 17463 43237
rect 17405 43197 17417 43231
rect 17451 43197 17463 43231
rect 17405 43191 17463 43197
rect 11882 43120 11888 43172
rect 11940 43160 11946 43172
rect 12820 43160 12848 43191
rect 11940 43132 12848 43160
rect 11940 43120 11946 43132
rect 14090 43120 14096 43172
rect 14148 43160 14154 43172
rect 17420 43160 17448 43191
rect 22002 43188 22008 43240
rect 22060 43188 22066 43240
rect 14148 43132 17448 43160
rect 14148 43120 14154 43132
rect 8205 43095 8263 43101
rect 8205 43061 8217 43095
rect 8251 43092 8263 43095
rect 8478 43092 8484 43104
rect 8251 43064 8484 43092
rect 8251 43061 8263 43064
rect 8205 43055 8263 43061
rect 8478 43052 8484 43064
rect 8536 43052 8542 43104
rect 16666 43052 16672 43104
rect 16724 43092 16730 43104
rect 16853 43095 16911 43101
rect 16853 43092 16865 43095
rect 16724 43064 16865 43092
rect 16724 43052 16730 43064
rect 16853 43061 16865 43064
rect 16899 43061 16911 43095
rect 16853 43055 16911 43061
rect 25133 43095 25191 43101
rect 25133 43061 25145 43095
rect 25179 43092 25191 43095
rect 25222 43092 25228 43104
rect 25179 43064 25228 43092
rect 25179 43061 25191 43064
rect 25133 43055 25191 43061
rect 25222 43052 25228 43064
rect 25280 43052 25286 43104
rect 1104 43002 25852 43024
rect 1104 42950 2950 43002
rect 3002 42950 3014 43002
rect 3066 42950 3078 43002
rect 3130 42950 3142 43002
rect 3194 42950 3206 43002
rect 3258 42950 12950 43002
rect 13002 42950 13014 43002
rect 13066 42950 13078 43002
rect 13130 42950 13142 43002
rect 13194 42950 13206 43002
rect 13258 42950 22950 43002
rect 23002 42950 23014 43002
rect 23066 42950 23078 43002
rect 23130 42950 23142 43002
rect 23194 42950 23206 43002
rect 23258 42950 25852 43002
rect 1104 42928 25852 42950
rect 12710 42848 12716 42900
rect 12768 42888 12774 42900
rect 14534 42891 14592 42897
rect 14534 42888 14546 42891
rect 12768 42860 14546 42888
rect 12768 42848 12774 42860
rect 14534 42857 14546 42860
rect 14580 42888 14592 42891
rect 17402 42888 17408 42900
rect 14580 42860 17408 42888
rect 14580 42857 14592 42860
rect 14534 42851 14592 42857
rect 17402 42848 17408 42860
rect 17460 42848 17466 42900
rect 15838 42780 15844 42832
rect 15896 42820 15902 42832
rect 16850 42820 16856 42832
rect 15896 42792 16856 42820
rect 15896 42780 15902 42792
rect 16850 42780 16856 42792
rect 16908 42820 16914 42832
rect 16908 42792 18092 42820
rect 16908 42780 16914 42792
rect 4154 42712 4160 42764
rect 4212 42712 4218 42764
rect 6273 42755 6331 42761
rect 6273 42721 6285 42755
rect 6319 42752 6331 42755
rect 6362 42752 6368 42764
rect 6319 42724 6368 42752
rect 6319 42721 6331 42724
rect 6273 42715 6331 42721
rect 6362 42712 6368 42724
rect 6420 42712 6426 42764
rect 8294 42712 8300 42764
rect 8352 42712 8358 42764
rect 9125 42755 9183 42761
rect 9125 42721 9137 42755
rect 9171 42752 9183 42755
rect 9214 42752 9220 42764
rect 9171 42724 9220 42752
rect 9171 42721 9183 42724
rect 9125 42715 9183 42721
rect 9214 42712 9220 42724
rect 9272 42752 9278 42764
rect 9493 42755 9551 42761
rect 9493 42752 9505 42755
rect 9272 42724 9505 42752
rect 9272 42712 9278 42724
rect 9493 42721 9505 42724
rect 9539 42721 9551 42755
rect 9493 42715 9551 42721
rect 12526 42712 12532 42764
rect 12584 42712 12590 42764
rect 14274 42712 14280 42764
rect 14332 42712 14338 42764
rect 18064 42761 18092 42792
rect 25130 42780 25136 42832
rect 25188 42820 25194 42832
rect 25406 42820 25412 42832
rect 25188 42792 25412 42820
rect 25188 42780 25194 42792
rect 25406 42780 25412 42792
rect 25464 42780 25470 42832
rect 18049 42755 18107 42761
rect 18049 42721 18061 42755
rect 18095 42721 18107 42755
rect 18049 42715 18107 42721
rect 7009 42687 7067 42693
rect 7009 42653 7021 42687
rect 7055 42684 7067 42687
rect 7558 42684 7564 42696
rect 7055 42656 7564 42684
rect 7055 42653 7067 42656
rect 7009 42647 7067 42653
rect 7558 42644 7564 42656
rect 7616 42644 7622 42696
rect 7653 42687 7711 42693
rect 7653 42653 7665 42687
rect 7699 42653 7711 42687
rect 7653 42647 7711 42653
rect 4341 42619 4399 42625
rect 4341 42585 4353 42619
rect 4387 42585 4399 42619
rect 4341 42579 4399 42585
rect 5997 42619 6055 42625
rect 5997 42585 6009 42619
rect 6043 42616 6055 42619
rect 6454 42616 6460 42628
rect 6043 42588 6460 42616
rect 6043 42585 6055 42588
rect 5997 42579 6055 42585
rect 4356 42548 4384 42579
rect 6454 42576 6460 42588
rect 6512 42576 6518 42628
rect 7668 42616 7696 42647
rect 8478 42644 8484 42696
rect 8536 42684 8542 42696
rect 9030 42684 9036 42696
rect 8536 42656 9036 42684
rect 8536 42644 8542 42656
rect 9030 42644 9036 42656
rect 9088 42644 9094 42696
rect 9674 42644 9680 42696
rect 9732 42684 9738 42696
rect 9769 42687 9827 42693
rect 9769 42684 9781 42687
rect 9732 42656 9781 42684
rect 9732 42644 9738 42656
rect 9769 42653 9781 42656
rect 9815 42653 9827 42687
rect 9769 42647 9827 42653
rect 11238 42644 11244 42696
rect 11296 42684 11302 42696
rect 11790 42684 11796 42696
rect 11296 42656 11796 42684
rect 11296 42644 11302 42656
rect 11790 42644 11796 42656
rect 11848 42684 11854 42696
rect 14292 42684 14320 42712
rect 11848 42656 14320 42684
rect 17957 42687 18015 42693
rect 11848 42644 11854 42656
rect 17957 42653 17969 42687
rect 18003 42684 18015 42687
rect 18322 42684 18328 42696
rect 18003 42656 18328 42684
rect 18003 42653 18015 42656
rect 17957 42647 18015 42653
rect 18322 42644 18328 42656
rect 18380 42644 18386 42696
rect 21174 42644 21180 42696
rect 21232 42684 21238 42696
rect 22002 42684 22008 42696
rect 21232 42656 22008 42684
rect 21232 42644 21238 42656
rect 22002 42644 22008 42656
rect 22060 42684 22066 42696
rect 22278 42684 22284 42696
rect 22060 42656 22284 42684
rect 22060 42644 22066 42656
rect 22278 42644 22284 42656
rect 22336 42644 22342 42696
rect 23658 42644 23664 42696
rect 23716 42644 23722 42696
rect 24765 42687 24823 42693
rect 24765 42653 24777 42687
rect 24811 42684 24823 42687
rect 24811 42656 24900 42684
rect 24811 42653 24823 42656
rect 24765 42647 24823 42653
rect 9490 42616 9496 42628
rect 7668 42588 9496 42616
rect 9490 42576 9496 42588
rect 9548 42576 9554 42628
rect 10962 42576 10968 42628
rect 11020 42616 11026 42628
rect 11020 42588 12020 42616
rect 11020 42576 11026 42588
rect 4801 42551 4859 42557
rect 4801 42548 4813 42551
rect 4356 42520 4813 42548
rect 4801 42517 4813 42520
rect 4847 42548 4859 42551
rect 6822 42548 6828 42560
rect 4847 42520 6828 42548
rect 4847 42517 4859 42520
rect 4801 42511 4859 42517
rect 6822 42508 6828 42520
rect 6880 42508 6886 42560
rect 7193 42551 7251 42557
rect 7193 42517 7205 42551
rect 7239 42548 7251 42551
rect 7374 42548 7380 42560
rect 7239 42520 7380 42548
rect 7239 42517 7251 42520
rect 7193 42511 7251 42517
rect 7374 42508 7380 42520
rect 7432 42508 7438 42560
rect 7650 42508 7656 42560
rect 7708 42548 7714 42560
rect 7837 42551 7895 42557
rect 7837 42548 7849 42551
rect 7708 42520 7849 42548
rect 7708 42508 7714 42520
rect 7837 42517 7849 42520
rect 7883 42517 7895 42551
rect 7837 42511 7895 42517
rect 9677 42551 9735 42557
rect 9677 42517 9689 42551
rect 9723 42548 9735 42551
rect 9858 42548 9864 42560
rect 9723 42520 9864 42548
rect 9723 42517 9735 42520
rect 9677 42511 9735 42517
rect 9858 42508 9864 42520
rect 9916 42508 9922 42560
rect 10137 42551 10195 42557
rect 10137 42517 10149 42551
rect 10183 42548 10195 42551
rect 11054 42548 11060 42560
rect 10183 42520 11060 42548
rect 10183 42517 10195 42520
rect 10137 42511 10195 42517
rect 11054 42508 11060 42520
rect 11112 42508 11118 42560
rect 11992 42557 12020 42588
rect 13722 42576 13728 42628
rect 13780 42616 13786 42628
rect 15010 42616 15016 42628
rect 13780 42588 15016 42616
rect 13780 42576 13786 42588
rect 15010 42576 15016 42588
rect 15068 42576 15074 42628
rect 20470 42588 20576 42616
rect 20548 42560 20576 42588
rect 20898 42576 20904 42628
rect 20956 42576 20962 42628
rect 21729 42619 21787 42625
rect 21729 42616 21741 42619
rect 21008 42588 21741 42616
rect 11977 42551 12035 42557
rect 11977 42517 11989 42551
rect 12023 42517 12035 42551
rect 11977 42511 12035 42517
rect 12066 42508 12072 42560
rect 12124 42548 12130 42560
rect 12345 42551 12403 42557
rect 12345 42548 12357 42551
rect 12124 42520 12357 42548
rect 12124 42508 12130 42520
rect 12345 42517 12357 42520
rect 12391 42517 12403 42551
rect 12345 42511 12403 42517
rect 12434 42508 12440 42560
rect 12492 42508 12498 42560
rect 15562 42508 15568 42560
rect 15620 42548 15626 42560
rect 16025 42551 16083 42557
rect 16025 42548 16037 42551
rect 15620 42520 16037 42548
rect 15620 42508 15626 42520
rect 16025 42517 16037 42520
rect 16071 42517 16083 42551
rect 16025 42511 16083 42517
rect 16298 42508 16304 42560
rect 16356 42508 16362 42560
rect 17497 42551 17555 42557
rect 17497 42517 17509 42551
rect 17543 42548 17555 42551
rect 17678 42548 17684 42560
rect 17543 42520 17684 42548
rect 17543 42517 17555 42520
rect 17497 42511 17555 42517
rect 17678 42508 17684 42520
rect 17736 42508 17742 42560
rect 17862 42508 17868 42560
rect 17920 42548 17926 42560
rect 18509 42551 18567 42557
rect 18509 42548 18521 42551
rect 17920 42520 18521 42548
rect 17920 42508 17926 42520
rect 18509 42517 18521 42520
rect 18555 42517 18567 42551
rect 18509 42511 18567 42517
rect 19334 42508 19340 42560
rect 19392 42548 19398 42560
rect 19429 42551 19487 42557
rect 19429 42548 19441 42551
rect 19392 42520 19441 42548
rect 19392 42508 19398 42520
rect 19429 42517 19441 42520
rect 19475 42517 19487 42551
rect 19429 42511 19487 42517
rect 20530 42508 20536 42560
rect 20588 42548 20594 42560
rect 20806 42548 20812 42560
rect 20588 42520 20812 42548
rect 20588 42508 20594 42520
rect 20806 42508 20812 42520
rect 20864 42548 20870 42560
rect 21008 42548 21036 42588
rect 21729 42585 21741 42588
rect 21775 42585 21787 42619
rect 21729 42579 21787 42585
rect 22554 42576 22560 42628
rect 22612 42576 22618 42628
rect 24872 42560 24900 42656
rect 20864 42520 21036 42548
rect 20864 42508 20870 42520
rect 21266 42508 21272 42560
rect 21324 42548 21330 42560
rect 21545 42551 21603 42557
rect 21545 42548 21557 42551
rect 21324 42520 21557 42548
rect 21324 42508 21330 42520
rect 21545 42517 21557 42520
rect 21591 42517 21603 42551
rect 21545 42511 21603 42517
rect 24029 42551 24087 42557
rect 24029 42517 24041 42551
rect 24075 42548 24087 42551
rect 24486 42548 24492 42560
rect 24075 42520 24492 42548
rect 24075 42517 24087 42520
rect 24029 42511 24087 42517
rect 24486 42508 24492 42520
rect 24544 42508 24550 42560
rect 24578 42508 24584 42560
rect 24636 42508 24642 42560
rect 24854 42508 24860 42560
rect 24912 42548 24918 42560
rect 25041 42551 25099 42557
rect 25041 42548 25053 42551
rect 24912 42520 25053 42548
rect 24912 42508 24918 42520
rect 25041 42517 25053 42520
rect 25087 42517 25099 42551
rect 25041 42511 25099 42517
rect 25498 42508 25504 42560
rect 25556 42508 25562 42560
rect 1104 42458 25852 42480
rect 1104 42406 7950 42458
rect 8002 42406 8014 42458
rect 8066 42406 8078 42458
rect 8130 42406 8142 42458
rect 8194 42406 8206 42458
rect 8258 42406 17950 42458
rect 18002 42406 18014 42458
rect 18066 42406 18078 42458
rect 18130 42406 18142 42458
rect 18194 42406 18206 42458
rect 18258 42406 25852 42458
rect 1104 42384 25852 42406
rect 6914 42304 6920 42356
rect 6972 42344 6978 42356
rect 7374 42344 7380 42356
rect 6972 42316 7380 42344
rect 6972 42304 6978 42316
rect 7374 42304 7380 42316
rect 7432 42304 7438 42356
rect 9398 42344 9404 42356
rect 7944 42316 9404 42344
rect 3694 42236 3700 42288
rect 3752 42236 3758 42288
rect 7944 42276 7972 42316
rect 9398 42304 9404 42316
rect 9456 42304 9462 42356
rect 9953 42347 10011 42353
rect 9953 42313 9965 42347
rect 9999 42344 10011 42347
rect 10042 42344 10048 42356
rect 9999 42316 10048 42344
rect 9999 42313 10011 42316
rect 9953 42307 10011 42313
rect 10042 42304 10048 42316
rect 10100 42344 10106 42356
rect 10962 42344 10968 42356
rect 10100 42316 10968 42344
rect 10100 42304 10106 42316
rect 10962 42304 10968 42316
rect 11020 42304 11026 42356
rect 11514 42304 11520 42356
rect 11572 42344 11578 42356
rect 11793 42347 11851 42353
rect 11793 42344 11805 42347
rect 11572 42316 11805 42344
rect 11572 42304 11578 42316
rect 11793 42313 11805 42316
rect 11839 42313 11851 42347
rect 11793 42307 11851 42313
rect 12434 42304 12440 42356
rect 12492 42344 12498 42356
rect 16758 42344 16764 42356
rect 12492 42316 16764 42344
rect 12492 42304 12498 42316
rect 16758 42304 16764 42316
rect 16816 42304 16822 42356
rect 19426 42344 19432 42356
rect 18432 42316 19432 42344
rect 18432 42288 18460 42316
rect 19426 42304 19432 42316
rect 19484 42304 19490 42356
rect 22281 42347 22339 42353
rect 22281 42313 22293 42347
rect 22327 42344 22339 42347
rect 22830 42344 22836 42356
rect 22327 42316 22836 42344
rect 22327 42313 22339 42316
rect 22281 42307 22339 42313
rect 22830 42304 22836 42316
rect 22888 42304 22894 42356
rect 23293 42347 23351 42353
rect 23293 42313 23305 42347
rect 23339 42313 23351 42347
rect 23842 42344 23848 42356
rect 23293 42307 23351 42313
rect 23676 42316 23848 42344
rect 7852 42248 7972 42276
rect 3881 42211 3939 42217
rect 3881 42177 3893 42211
rect 3927 42208 3939 42211
rect 4338 42208 4344 42220
rect 3927 42180 4344 42208
rect 3927 42177 3939 42180
rect 3881 42171 3939 42177
rect 4338 42168 4344 42180
rect 4396 42168 4402 42220
rect 7852 42217 7880 42248
rect 8570 42236 8576 42288
rect 8628 42236 8634 42288
rect 12161 42279 12219 42285
rect 12161 42245 12173 42279
rect 12207 42276 12219 42279
rect 12342 42276 12348 42288
rect 12207 42248 12348 42276
rect 12207 42245 12219 42248
rect 12161 42239 12219 42245
rect 12342 42236 12348 42248
rect 12400 42236 12406 42288
rect 13722 42236 13728 42288
rect 13780 42276 13786 42288
rect 13780 42248 13938 42276
rect 13780 42236 13786 42248
rect 15010 42236 15016 42288
rect 15068 42276 15074 42288
rect 15657 42279 15715 42285
rect 15657 42276 15669 42279
rect 15068 42248 15669 42276
rect 15068 42236 15074 42248
rect 15657 42245 15669 42248
rect 15703 42276 15715 42279
rect 16298 42276 16304 42288
rect 15703 42248 16304 42276
rect 15703 42245 15715 42248
rect 15657 42239 15715 42245
rect 16298 42236 16304 42248
rect 16356 42236 16362 42288
rect 18414 42276 18420 42288
rect 17880 42248 18420 42276
rect 7837 42211 7895 42217
rect 7837 42177 7849 42211
rect 7883 42177 7895 42211
rect 7837 42171 7895 42177
rect 12253 42211 12311 42217
rect 12253 42177 12265 42211
rect 12299 42208 12311 42211
rect 13814 42208 13820 42220
rect 12299 42180 13820 42208
rect 12299 42177 12311 42180
rect 12253 42171 12311 42177
rect 13814 42168 13820 42180
rect 13872 42168 13878 42220
rect 15381 42211 15439 42217
rect 15381 42177 15393 42211
rect 15427 42208 15439 42211
rect 15470 42208 15476 42220
rect 15427 42180 15476 42208
rect 15427 42177 15439 42180
rect 15381 42171 15439 42177
rect 15470 42168 15476 42180
rect 15528 42208 15534 42220
rect 17880 42217 17908 42248
rect 18414 42236 18420 42248
rect 18472 42236 18478 42288
rect 20717 42279 20775 42285
rect 20717 42245 20729 42279
rect 20763 42276 20775 42279
rect 21174 42276 21180 42288
rect 20763 42248 21180 42276
rect 20763 42245 20775 42248
rect 20717 42239 20775 42245
rect 21174 42236 21180 42248
rect 21232 42236 21238 42288
rect 22738 42236 22744 42288
rect 22796 42276 22802 42288
rect 23308 42276 23336 42307
rect 22796 42248 23336 42276
rect 22796 42236 22802 42248
rect 23676 42220 23704 42316
rect 23842 42304 23848 42316
rect 23900 42344 23906 42356
rect 25317 42347 25375 42353
rect 25317 42344 25329 42347
rect 23900 42316 25329 42344
rect 23900 42304 23906 42316
rect 25317 42313 25329 42316
rect 25363 42313 25375 42347
rect 25317 42307 25375 42313
rect 24486 42236 24492 42288
rect 24544 42276 24550 42288
rect 24670 42276 24676 42288
rect 24544 42248 24676 42276
rect 24544 42236 24550 42248
rect 24670 42236 24676 42248
rect 24728 42276 24734 42288
rect 24765 42279 24823 42285
rect 24765 42276 24777 42279
rect 24728 42248 24777 42276
rect 24728 42236 24734 42248
rect 24765 42245 24777 42248
rect 24811 42245 24823 42279
rect 24765 42239 24823 42245
rect 17865 42211 17923 42217
rect 17865 42208 17877 42211
rect 15528 42180 17877 42208
rect 15528 42168 15534 42180
rect 17865 42177 17877 42180
rect 17911 42177 17923 42211
rect 17865 42171 17923 42177
rect 19242 42168 19248 42220
rect 19300 42208 19306 42220
rect 19300 42180 20024 42208
rect 19300 42168 19306 42180
rect 8113 42143 8171 42149
rect 8113 42109 8125 42143
rect 8159 42140 8171 42143
rect 8478 42140 8484 42152
rect 8159 42112 8484 42140
rect 8159 42109 8171 42112
rect 8113 42103 8171 42109
rect 8478 42100 8484 42112
rect 8536 42100 8542 42152
rect 11146 42100 11152 42152
rect 11204 42140 11210 42152
rect 12345 42143 12403 42149
rect 12345 42140 12357 42143
rect 11204 42112 12357 42140
rect 11204 42100 11210 42112
rect 12345 42109 12357 42112
rect 12391 42109 12403 42143
rect 12345 42103 12403 42109
rect 15105 42143 15163 42149
rect 15105 42109 15117 42143
rect 15151 42140 15163 42143
rect 15562 42140 15568 42152
rect 15151 42112 15568 42140
rect 15151 42109 15163 42112
rect 15105 42103 15163 42109
rect 15562 42100 15568 42112
rect 15620 42100 15626 42152
rect 18141 42143 18199 42149
rect 18141 42109 18153 42143
rect 18187 42140 18199 42143
rect 19150 42140 19156 42152
rect 18187 42112 19156 42140
rect 18187 42109 18199 42112
rect 18141 42103 18199 42109
rect 19150 42100 19156 42112
rect 19208 42100 19214 42152
rect 9585 42075 9643 42081
rect 9585 42041 9597 42075
rect 9631 42072 9643 42075
rect 11514 42072 11520 42084
rect 9631 42044 11520 42072
rect 9631 42041 9643 42044
rect 9585 42035 9643 42041
rect 11514 42032 11520 42044
rect 11572 42032 11578 42084
rect 19996 42081 20024 42180
rect 21082 42168 21088 42220
rect 21140 42208 21146 42220
rect 21453 42211 21511 42217
rect 21453 42208 21465 42211
rect 21140 42180 21465 42208
rect 21140 42168 21146 42180
rect 21453 42177 21465 42180
rect 21499 42177 21511 42211
rect 21453 42171 21511 42177
rect 22370 42168 22376 42220
rect 22428 42168 22434 42220
rect 23658 42168 23664 42220
rect 23716 42168 23722 42220
rect 22186 42100 22192 42152
rect 22244 42140 22250 42152
rect 22554 42140 22560 42152
rect 22244 42112 22560 42140
rect 22244 42100 22250 42112
rect 22554 42100 22560 42112
rect 22612 42100 22618 42152
rect 25038 42100 25044 42152
rect 25096 42100 25102 42152
rect 19981 42075 20039 42081
rect 19981 42041 19993 42075
rect 20027 42072 20039 42075
rect 20530 42072 20536 42084
rect 20027 42044 20536 42072
rect 20027 42041 20039 42044
rect 19981 42035 20039 42041
rect 20530 42032 20536 42044
rect 20588 42032 20594 42084
rect 22741 42075 22799 42081
rect 22741 42041 22753 42075
rect 22787 42072 22799 42075
rect 22787 42044 23796 42072
rect 22787 42041 22799 42044
rect 22741 42035 22799 42041
rect 4338 41964 4344 42016
rect 4396 41964 4402 42016
rect 8662 41964 8668 42016
rect 8720 42004 8726 42016
rect 11422 42004 11428 42016
rect 8720 41976 11428 42004
rect 8720 41964 8726 41976
rect 11422 41964 11428 41976
rect 11480 41964 11486 42016
rect 13633 42007 13691 42013
rect 13633 41973 13645 42007
rect 13679 42004 13691 42007
rect 14550 42004 14556 42016
rect 13679 41976 14556 42004
rect 13679 41973 13691 41976
rect 13633 41967 13691 41973
rect 14550 41964 14556 41976
rect 14608 41964 14614 42016
rect 19610 41964 19616 42016
rect 19668 41964 19674 42016
rect 20257 42007 20315 42013
rect 20257 41973 20269 42007
rect 20303 42004 20315 42007
rect 21082 42004 21088 42016
rect 20303 41976 21088 42004
rect 20303 41973 20315 41976
rect 20257 41967 20315 41973
rect 21082 41964 21088 41976
rect 21140 41964 21146 42016
rect 23768 42004 23796 42044
rect 25130 42004 25136 42016
rect 23768 41976 25136 42004
rect 25130 41964 25136 41976
rect 25188 41964 25194 42016
rect 1104 41914 25852 41936
rect 1104 41862 2950 41914
rect 3002 41862 3014 41914
rect 3066 41862 3078 41914
rect 3130 41862 3142 41914
rect 3194 41862 3206 41914
rect 3258 41862 12950 41914
rect 13002 41862 13014 41914
rect 13066 41862 13078 41914
rect 13130 41862 13142 41914
rect 13194 41862 13206 41914
rect 13258 41862 22950 41914
rect 23002 41862 23014 41914
rect 23066 41862 23078 41914
rect 23130 41862 23142 41914
rect 23194 41862 23206 41914
rect 23258 41862 25852 41914
rect 1104 41840 25852 41862
rect 4430 41760 4436 41812
rect 4488 41760 4494 41812
rect 5350 41760 5356 41812
rect 5408 41760 5414 41812
rect 7282 41760 7288 41812
rect 7340 41800 7346 41812
rect 7837 41803 7895 41809
rect 7837 41800 7849 41803
rect 7340 41772 7849 41800
rect 7340 41760 7346 41772
rect 7837 41769 7849 41772
rect 7883 41769 7895 41803
rect 7837 41763 7895 41769
rect 16206 41760 16212 41812
rect 16264 41800 16270 41812
rect 17313 41803 17371 41809
rect 17313 41800 17325 41803
rect 16264 41772 17325 41800
rect 16264 41760 16270 41772
rect 8478 41624 8484 41676
rect 8536 41624 8542 41676
rect 11238 41624 11244 41676
rect 11296 41624 11302 41676
rect 11514 41624 11520 41676
rect 11572 41624 11578 41676
rect 15197 41667 15255 41673
rect 15197 41633 15209 41667
rect 15243 41664 15255 41667
rect 15470 41664 15476 41676
rect 15243 41636 15476 41664
rect 15243 41633 15255 41636
rect 15197 41627 15255 41633
rect 15470 41624 15476 41636
rect 15528 41624 15534 41676
rect 16500 41664 16528 41772
rect 17313 41769 17325 41772
rect 17359 41800 17371 41803
rect 17494 41800 17500 41812
rect 17359 41772 17500 41800
rect 17359 41769 17371 41772
rect 17313 41763 17371 41769
rect 17494 41760 17500 41772
rect 17552 41800 17558 41812
rect 19242 41800 19248 41812
rect 17552 41772 19248 41800
rect 17552 41760 17558 41772
rect 19242 41760 19248 41772
rect 19300 41760 19306 41812
rect 21266 41760 21272 41812
rect 21324 41800 21330 41812
rect 23566 41800 23572 41812
rect 21324 41772 23572 41800
rect 21324 41760 21330 41772
rect 23566 41760 23572 41772
rect 23624 41760 23630 41812
rect 16945 41735 17003 41741
rect 16945 41701 16957 41735
rect 16991 41732 17003 41735
rect 19058 41732 19064 41744
rect 16991 41704 19064 41732
rect 16991 41701 17003 41704
rect 16945 41695 17003 41701
rect 19058 41692 19064 41704
rect 19116 41692 19122 41744
rect 19334 41692 19340 41744
rect 19392 41732 19398 41744
rect 21453 41735 21511 41741
rect 19392 41704 20024 41732
rect 19392 41692 19398 41704
rect 16500 41636 16620 41664
rect 4525 41599 4583 41605
rect 4525 41565 4537 41599
rect 4571 41596 4583 41599
rect 4985 41599 5043 41605
rect 4985 41596 4997 41599
rect 4571 41568 4997 41596
rect 4571 41565 4583 41568
rect 4525 41559 4583 41565
rect 4985 41565 4997 41568
rect 5031 41596 5043 41599
rect 6638 41596 6644 41608
rect 5031 41568 6644 41596
rect 5031 41565 5043 41568
rect 4985 41559 5043 41565
rect 6638 41556 6644 41568
rect 6696 41556 6702 41608
rect 8205 41599 8263 41605
rect 8205 41565 8217 41599
rect 8251 41596 8263 41599
rect 8294 41596 8300 41608
rect 8251 41568 8300 41596
rect 8251 41565 8263 41568
rect 8205 41559 8263 41565
rect 8294 41556 8300 41568
rect 8352 41556 8358 41608
rect 13262 41596 13268 41608
rect 12650 41568 13268 41596
rect 13262 41556 13268 41568
rect 13320 41596 13326 41608
rect 13722 41596 13728 41608
rect 13320 41568 13728 41596
rect 13320 41556 13326 41568
rect 13722 41556 13728 41568
rect 13780 41556 13786 41608
rect 16592 41582 16620 41636
rect 18414 41624 18420 41676
rect 18472 41664 18478 41676
rect 18693 41667 18751 41673
rect 18693 41664 18705 41667
rect 18472 41636 18705 41664
rect 18472 41624 18478 41636
rect 18693 41633 18705 41636
rect 18739 41633 18751 41667
rect 18693 41627 18751 41633
rect 19702 41624 19708 41676
rect 19760 41664 19766 41676
rect 19996 41673 20024 41704
rect 21453 41701 21465 41735
rect 21499 41732 21511 41735
rect 23198 41732 23204 41744
rect 21499 41704 23204 41732
rect 21499 41701 21511 41704
rect 21453 41695 21511 41701
rect 23198 41692 23204 41704
rect 23256 41692 23262 41744
rect 24394 41692 24400 41744
rect 24452 41732 24458 41744
rect 24452 41704 25176 41732
rect 24452 41692 24458 41704
rect 19889 41667 19947 41673
rect 19889 41664 19901 41667
rect 19760 41636 19901 41664
rect 19760 41624 19766 41636
rect 19889 41633 19901 41636
rect 19935 41633 19947 41667
rect 19889 41627 19947 41633
rect 19981 41667 20039 41673
rect 19981 41633 19993 41667
rect 20027 41633 20039 41667
rect 19981 41627 20039 41633
rect 20806 41624 20812 41676
rect 20864 41624 20870 41676
rect 20990 41624 20996 41676
rect 21048 41624 21054 41676
rect 22094 41624 22100 41676
rect 22152 41624 22158 41676
rect 23382 41624 23388 41676
rect 23440 41624 23446 41676
rect 23658 41624 23664 41676
rect 23716 41664 23722 41676
rect 25148 41673 25176 41704
rect 25133 41667 25191 41673
rect 23716 41636 24992 41664
rect 23716 41624 23722 41636
rect 17681 41599 17739 41605
rect 17681 41565 17693 41599
rect 17727 41596 17739 41599
rect 17957 41599 18015 41605
rect 17957 41596 17969 41599
rect 17727 41568 17969 41596
rect 17727 41565 17739 41568
rect 17681 41559 17739 41565
rect 17957 41565 17969 41568
rect 18003 41596 18015 41599
rect 21082 41596 21088 41608
rect 18003 41568 21088 41596
rect 18003 41565 18015 41568
rect 17957 41559 18015 41565
rect 21082 41556 21088 41568
rect 21140 41556 21146 41608
rect 21910 41556 21916 41608
rect 21968 41596 21974 41608
rect 23400 41596 23428 41624
rect 21968 41568 23428 41596
rect 21968 41556 21974 41568
rect 23750 41556 23756 41608
rect 23808 41556 23814 41608
rect 24029 41599 24087 41605
rect 24029 41565 24041 41599
rect 24075 41596 24087 41599
rect 24762 41596 24768 41608
rect 24075 41568 24768 41596
rect 24075 41565 24087 41568
rect 24029 41559 24087 41565
rect 24762 41556 24768 41568
rect 24820 41556 24826 41608
rect 24964 41605 24992 41636
rect 25133 41633 25145 41667
rect 25179 41633 25191 41667
rect 25133 41627 25191 41633
rect 24949 41599 25007 41605
rect 24949 41565 24961 41599
rect 24995 41565 25007 41599
rect 24949 41559 25007 41565
rect 1670 41488 1676 41540
rect 1728 41528 1734 41540
rect 2133 41531 2191 41537
rect 2133 41528 2145 41531
rect 1728 41500 2145 41528
rect 1728 41488 1734 41500
rect 2133 41497 2145 41500
rect 2179 41497 2191 41531
rect 2133 41491 2191 41497
rect 5445 41531 5503 41537
rect 5445 41497 5457 41531
rect 5491 41497 5503 41531
rect 15473 41531 15531 41537
rect 15473 41528 15485 41531
rect 5445 41491 5503 41497
rect 13004 41500 15485 41528
rect 1765 41463 1823 41469
rect 1765 41429 1777 41463
rect 1811 41460 1823 41463
rect 3602 41460 3608 41472
rect 1811 41432 3608 41460
rect 1811 41429 1823 41432
rect 1765 41423 1823 41429
rect 3602 41420 3608 41432
rect 3660 41420 3666 41472
rect 5460 41460 5488 41491
rect 5905 41463 5963 41469
rect 5905 41460 5917 41463
rect 5460 41432 5917 41460
rect 5905 41429 5917 41432
rect 5951 41460 5963 41463
rect 6270 41460 6276 41472
rect 5951 41432 6276 41460
rect 5951 41429 5963 41432
rect 5905 41423 5963 41429
rect 6270 41420 6276 41432
rect 6328 41420 6334 41472
rect 8297 41463 8355 41469
rect 8297 41429 8309 41463
rect 8343 41460 8355 41463
rect 9582 41460 9588 41472
rect 8343 41432 9588 41460
rect 8343 41429 8355 41432
rect 8297 41423 8355 41429
rect 9582 41420 9588 41432
rect 9640 41420 9646 41472
rect 12526 41420 12532 41472
rect 12584 41460 12590 41472
rect 13004 41469 13032 41500
rect 15473 41497 15485 41500
rect 15519 41497 15531 41531
rect 15473 41491 15531 41497
rect 22281 41531 22339 41537
rect 22281 41497 22293 41531
rect 22327 41528 22339 41531
rect 22327 41500 24624 41528
rect 22327 41497 22339 41500
rect 22281 41491 22339 41497
rect 12989 41463 13047 41469
rect 12989 41460 13001 41463
rect 12584 41432 13001 41460
rect 12584 41420 12590 41432
rect 12989 41429 13001 41432
rect 13035 41429 13047 41463
rect 12989 41423 13047 41429
rect 13262 41420 13268 41472
rect 13320 41420 13326 41472
rect 19426 41420 19432 41472
rect 19484 41420 19490 41472
rect 19518 41420 19524 41472
rect 19576 41460 19582 41472
rect 19797 41463 19855 41469
rect 19797 41460 19809 41463
rect 19576 41432 19809 41460
rect 19576 41420 19582 41432
rect 19797 41429 19809 41432
rect 19843 41429 19855 41463
rect 19797 41423 19855 41429
rect 21085 41463 21143 41469
rect 21085 41429 21097 41463
rect 21131 41460 21143 41463
rect 21174 41460 21180 41472
rect 21131 41432 21180 41460
rect 21131 41429 21143 41432
rect 21085 41423 21143 41429
rect 21174 41420 21180 41432
rect 21232 41420 21238 41472
rect 22373 41463 22431 41469
rect 22373 41429 22385 41463
rect 22419 41460 22431 41463
rect 22646 41460 22652 41472
rect 22419 41432 22652 41460
rect 22419 41429 22431 41432
rect 22373 41423 22431 41429
rect 22646 41420 22652 41432
rect 22704 41420 22710 41472
rect 22741 41463 22799 41469
rect 22741 41429 22753 41463
rect 22787 41460 22799 41463
rect 23474 41460 23480 41472
rect 22787 41432 23480 41460
rect 22787 41429 22799 41432
rect 22741 41423 22799 41429
rect 23474 41420 23480 41432
rect 23532 41420 23538 41472
rect 24596 41469 24624 41500
rect 24581 41463 24639 41469
rect 24581 41429 24593 41463
rect 24627 41429 24639 41463
rect 24581 41423 24639 41429
rect 24946 41420 24952 41472
rect 25004 41460 25010 41472
rect 25041 41463 25099 41469
rect 25041 41460 25053 41463
rect 25004 41432 25053 41460
rect 25004 41420 25010 41432
rect 25041 41429 25053 41432
rect 25087 41429 25099 41463
rect 25041 41423 25099 41429
rect 1104 41370 25852 41392
rect 1104 41318 7950 41370
rect 8002 41318 8014 41370
rect 8066 41318 8078 41370
rect 8130 41318 8142 41370
rect 8194 41318 8206 41370
rect 8258 41318 17950 41370
rect 18002 41318 18014 41370
rect 18066 41318 18078 41370
rect 18130 41318 18142 41370
rect 18194 41318 18206 41370
rect 18258 41318 25852 41370
rect 1104 41296 25852 41318
rect 3970 41216 3976 41268
rect 4028 41216 4034 41268
rect 4522 41216 4528 41268
rect 4580 41256 4586 41268
rect 7558 41256 7564 41268
rect 4580 41228 7564 41256
rect 4580 41216 4586 41228
rect 7558 41216 7564 41228
rect 7616 41256 7622 41268
rect 8297 41259 8355 41265
rect 7616 41228 8248 41256
rect 7616 41216 7622 41228
rect 7098 41148 7104 41200
rect 7156 41188 7162 41200
rect 8220 41188 8248 41228
rect 8297 41225 8309 41259
rect 8343 41256 8355 41259
rect 8478 41256 8484 41268
rect 8343 41228 8484 41256
rect 8343 41225 8355 41228
rect 8297 41219 8355 41225
rect 8478 41216 8484 41228
rect 8536 41216 8542 41268
rect 9674 41256 9680 41268
rect 9646 41216 9680 41256
rect 9732 41256 9738 41268
rect 12250 41256 12256 41268
rect 9732 41228 12256 41256
rect 9732 41216 9738 41228
rect 12250 41216 12256 41228
rect 12308 41216 12314 41268
rect 12437 41259 12495 41265
rect 12437 41225 12449 41259
rect 12483 41256 12495 41259
rect 12618 41256 12624 41268
rect 12483 41228 12624 41256
rect 12483 41225 12495 41228
rect 12437 41219 12495 41225
rect 12618 41216 12624 41228
rect 12676 41216 12682 41268
rect 12805 41259 12863 41265
rect 12805 41225 12817 41259
rect 12851 41256 12863 41259
rect 13262 41256 13268 41268
rect 12851 41228 13268 41256
rect 12851 41225 12863 41228
rect 12805 41219 12863 41225
rect 9646 41188 9674 41216
rect 10962 41188 10968 41200
rect 7156 41160 7314 41188
rect 8220 41160 9674 41188
rect 10902 41160 10968 41188
rect 7156 41148 7162 41160
rect 10962 41148 10968 41160
rect 11020 41188 11026 41200
rect 12820 41188 12848 41219
rect 13262 41216 13268 41228
rect 13320 41256 13326 41268
rect 15381 41259 15439 41265
rect 15381 41256 15393 41259
rect 13320 41228 15393 41256
rect 13320 41216 13326 41228
rect 11020 41160 12848 41188
rect 11020 41148 11026 41160
rect 14366 41148 14372 41200
rect 14424 41188 14430 41200
rect 14476 41188 14504 41228
rect 15381 41225 15393 41228
rect 15427 41225 15439 41259
rect 15381 41219 15439 41225
rect 17310 41216 17316 41268
rect 17368 41216 17374 41268
rect 19334 41256 19340 41268
rect 18708 41228 19340 41256
rect 14424 41160 14504 41188
rect 14424 41148 14430 41160
rect 14550 41148 14556 41200
rect 14608 41188 14614 41200
rect 14829 41191 14887 41197
rect 14829 41188 14841 41191
rect 14608 41160 14841 41188
rect 14608 41148 14614 41160
rect 14829 41157 14841 41160
rect 14875 41157 14887 41191
rect 14829 41151 14887 41157
rect 16206 41148 16212 41200
rect 16264 41188 16270 41200
rect 18708 41197 18736 41228
rect 19334 41216 19340 41228
rect 19392 41216 19398 41268
rect 22002 41216 22008 41268
rect 22060 41256 22066 41268
rect 22554 41256 22560 41268
rect 22060 41228 22560 41256
rect 22060 41216 22066 41228
rect 22554 41216 22560 41228
rect 22612 41216 22618 41268
rect 22738 41216 22744 41268
rect 22796 41216 22802 41268
rect 23842 41216 23848 41268
rect 23900 41256 23906 41268
rect 23900 41228 24348 41256
rect 23900 41216 23906 41228
rect 18693 41191 18751 41197
rect 18693 41188 18705 41191
rect 16264 41160 18705 41188
rect 16264 41148 16270 41160
rect 18693 41157 18705 41160
rect 18739 41157 18751 41191
rect 18693 41151 18751 41157
rect 24210 41148 24216 41200
rect 24268 41188 24274 41200
rect 24320 41188 24348 41228
rect 25225 41191 25283 41197
rect 25225 41188 25237 41191
rect 24268 41160 25237 41188
rect 24268 41148 24274 41160
rect 25225 41157 25237 41160
rect 25271 41157 25283 41191
rect 25225 41151 25283 41157
rect 4065 41123 4123 41129
rect 4065 41089 4077 41123
rect 4111 41120 4123 41123
rect 4246 41120 4252 41132
rect 4111 41092 4252 41120
rect 4111 41089 4123 41092
rect 4065 41083 4123 41089
rect 4246 41080 4252 41092
rect 4304 41080 4310 41132
rect 12069 41123 12127 41129
rect 12069 41120 12081 41123
rect 11072 41092 12081 41120
rect 6362 41012 6368 41064
rect 6420 41052 6426 41064
rect 6549 41055 6607 41061
rect 6549 41052 6561 41055
rect 6420 41024 6561 41052
rect 6420 41012 6426 41024
rect 6549 41021 6561 41024
rect 6595 41021 6607 41055
rect 6549 41015 6607 41021
rect 6825 41055 6883 41061
rect 6825 41021 6837 41055
rect 6871 41052 6883 41055
rect 7834 41052 7840 41064
rect 6871 41024 7840 41052
rect 6871 41021 6883 41024
rect 6825 41015 6883 41021
rect 7834 41012 7840 41024
rect 7892 41012 7898 41064
rect 9398 41012 9404 41064
rect 9456 41012 9462 41064
rect 9677 41055 9735 41061
rect 9677 41021 9689 41055
rect 9723 41052 9735 41055
rect 9723 41024 10824 41052
rect 9723 41021 9735 41024
rect 9677 41015 9735 41021
rect 10796 40984 10824 41024
rect 10870 41012 10876 41064
rect 10928 41052 10934 41064
rect 11072 41052 11100 41092
rect 12069 41089 12081 41092
rect 12115 41089 12127 41123
rect 12069 41083 12127 41089
rect 15105 41123 15163 41129
rect 15105 41089 15117 41123
rect 15151 41120 15163 41123
rect 15470 41120 15476 41132
rect 15151 41092 15476 41120
rect 15151 41089 15163 41092
rect 15105 41083 15163 41089
rect 15470 41080 15476 41092
rect 15528 41080 15534 41132
rect 17218 41080 17224 41132
rect 17276 41080 17282 41132
rect 18414 41080 18420 41132
rect 18472 41080 18478 41132
rect 22373 41123 22431 41129
rect 10928 41024 11100 41052
rect 10928 41012 10934 41024
rect 11882 41012 11888 41064
rect 11940 41012 11946 41064
rect 11977 41055 12035 41061
rect 11977 41021 11989 41055
rect 12023 41052 12035 41055
rect 14826 41052 14832 41064
rect 12023 41024 14832 41052
rect 12023 41021 12035 41024
rect 11977 41015 12035 41021
rect 14826 41012 14832 41024
rect 14884 41012 14890 41064
rect 17402 41012 17408 41064
rect 17460 41012 17466 41064
rect 19812 41052 19840 41106
rect 22373 41089 22385 41123
rect 22419 41120 22431 41123
rect 23382 41120 23388 41132
rect 22419 41092 23388 41120
rect 22419 41089 22431 41092
rect 22373 41083 22431 41089
rect 23382 41080 23388 41092
rect 23440 41080 23446 41132
rect 20530 41052 20536 41064
rect 19812 41024 20536 41052
rect 20530 41012 20536 41024
rect 20588 41052 20594 41064
rect 21358 41052 21364 41064
rect 20588 41024 21364 41052
rect 20588 41012 20594 41024
rect 21358 41012 21364 41024
rect 21416 41012 21422 41064
rect 21453 41055 21511 41061
rect 21453 41021 21465 41055
rect 21499 41052 21511 41055
rect 21726 41052 21732 41064
rect 21499 41024 21732 41052
rect 21499 41021 21511 41024
rect 21453 41015 21511 41021
rect 21726 41012 21732 41024
rect 21784 41012 21790 41064
rect 22186 41012 22192 41064
rect 22244 41012 22250 41064
rect 22281 41055 22339 41061
rect 22281 41021 22293 41055
rect 22327 41052 22339 41055
rect 22554 41052 22560 41064
rect 22327 41024 22560 41052
rect 22327 41021 22339 41024
rect 22281 41015 22339 41021
rect 22554 41012 22560 41024
rect 22612 41012 22618 41064
rect 24118 41012 24124 41064
rect 24176 41052 24182 41064
rect 24673 41055 24731 41061
rect 24673 41052 24685 41055
rect 24176 41024 24685 41052
rect 24176 41012 24182 41024
rect 24673 41021 24685 41024
rect 24719 41021 24731 41055
rect 24673 41015 24731 41021
rect 24946 41012 24952 41064
rect 25004 41012 25010 41064
rect 11330 40984 11336 40996
rect 10796 40956 11336 40984
rect 11330 40944 11336 40956
rect 11388 40944 11394 40996
rect 21542 40984 21548 40996
rect 19904 40956 21548 40984
rect 4246 40876 4252 40928
rect 4304 40916 4310 40928
rect 4433 40919 4491 40925
rect 4433 40916 4445 40919
rect 4304 40888 4445 40916
rect 4304 40876 4310 40888
rect 4433 40885 4445 40888
rect 4479 40885 4491 40919
rect 4433 40879 4491 40885
rect 8570 40876 8576 40928
rect 8628 40876 8634 40928
rect 11146 40876 11152 40928
rect 11204 40916 11210 40928
rect 11882 40916 11888 40928
rect 11204 40888 11888 40916
rect 11204 40876 11210 40888
rect 11882 40876 11888 40888
rect 11940 40876 11946 40928
rect 13357 40919 13415 40925
rect 13357 40885 13369 40919
rect 13403 40916 13415 40919
rect 13630 40916 13636 40928
rect 13403 40888 13636 40916
rect 13403 40885 13415 40888
rect 13357 40879 13415 40885
rect 13630 40876 13636 40888
rect 13688 40876 13694 40928
rect 13814 40876 13820 40928
rect 13872 40916 13878 40928
rect 14458 40916 14464 40928
rect 13872 40888 14464 40916
rect 13872 40876 13878 40888
rect 14458 40876 14464 40888
rect 14516 40876 14522 40928
rect 16850 40876 16856 40928
rect 16908 40876 16914 40928
rect 17218 40876 17224 40928
rect 17276 40916 17282 40928
rect 17865 40919 17923 40925
rect 17865 40916 17877 40919
rect 17276 40888 17877 40916
rect 17276 40876 17282 40888
rect 17865 40885 17877 40888
rect 17911 40916 17923 40919
rect 19904 40916 19932 40956
rect 21542 40944 21548 40956
rect 21600 40944 21606 40996
rect 22204 40984 22232 41012
rect 23201 40987 23259 40993
rect 23201 40984 23213 40987
rect 22204 40956 23213 40984
rect 23201 40953 23213 40956
rect 23247 40953 23259 40987
rect 26050 40984 26056 40996
rect 23201 40947 23259 40953
rect 24872 40956 26056 40984
rect 17911 40888 19932 40916
rect 17911 40885 17923 40888
rect 17865 40879 17923 40885
rect 19978 40876 19984 40928
rect 20036 40916 20042 40928
rect 20165 40919 20223 40925
rect 20165 40916 20177 40919
rect 20036 40888 20177 40916
rect 20036 40876 20042 40888
rect 20165 40885 20177 40888
rect 20211 40885 20223 40919
rect 20165 40879 20223 40885
rect 20530 40876 20536 40928
rect 20588 40916 20594 40928
rect 24872 40916 24900 40956
rect 26050 40944 26056 40956
rect 26108 40944 26114 40996
rect 20588 40888 24900 40916
rect 20588 40876 20594 40888
rect 25314 40876 25320 40928
rect 25372 40916 25378 40928
rect 25409 40919 25467 40925
rect 25409 40916 25421 40919
rect 25372 40888 25421 40916
rect 25372 40876 25378 40888
rect 25409 40885 25421 40888
rect 25455 40885 25467 40919
rect 25409 40879 25467 40885
rect 1104 40826 25852 40848
rect 1104 40774 2950 40826
rect 3002 40774 3014 40826
rect 3066 40774 3078 40826
rect 3130 40774 3142 40826
rect 3194 40774 3206 40826
rect 3258 40774 12950 40826
rect 13002 40774 13014 40826
rect 13066 40774 13078 40826
rect 13130 40774 13142 40826
rect 13194 40774 13206 40826
rect 13258 40774 22950 40826
rect 23002 40774 23014 40826
rect 23066 40774 23078 40826
rect 23130 40774 23142 40826
rect 23194 40774 23206 40826
rect 23258 40774 25852 40826
rect 1104 40752 25852 40774
rect 8570 40672 8576 40724
rect 8628 40712 8634 40724
rect 9858 40712 9864 40724
rect 8628 40684 9864 40712
rect 8628 40672 8634 40684
rect 9858 40672 9864 40684
rect 9916 40672 9922 40724
rect 14185 40715 14243 40721
rect 14185 40681 14197 40715
rect 14231 40712 14243 40715
rect 14366 40712 14372 40724
rect 14231 40684 14372 40712
rect 14231 40681 14243 40684
rect 14185 40675 14243 40681
rect 14366 40672 14372 40684
rect 14424 40672 14430 40724
rect 15654 40672 15660 40724
rect 15712 40712 15718 40724
rect 17405 40715 17463 40721
rect 17405 40712 17417 40715
rect 15712 40684 17417 40712
rect 15712 40672 15718 40684
rect 17405 40681 17417 40684
rect 17451 40681 17463 40715
rect 17405 40675 17463 40681
rect 17494 40672 17500 40724
rect 17552 40712 17558 40724
rect 25133 40715 25191 40721
rect 25133 40712 25145 40715
rect 17552 40684 25145 40712
rect 17552 40672 17558 40684
rect 25133 40681 25145 40684
rect 25179 40681 25191 40715
rect 25133 40675 25191 40681
rect 2961 40647 3019 40653
rect 2961 40613 2973 40647
rect 3007 40644 3019 40647
rect 3326 40644 3332 40656
rect 3007 40616 3332 40644
rect 3007 40613 3019 40616
rect 2961 40607 3019 40613
rect 3326 40604 3332 40616
rect 3384 40604 3390 40656
rect 13004 40616 14412 40644
rect 7834 40536 7840 40588
rect 7892 40576 7898 40588
rect 8113 40579 8171 40585
rect 8113 40576 8125 40579
rect 7892 40548 8125 40576
rect 7892 40536 7898 40548
rect 8113 40545 8125 40548
rect 8159 40545 8171 40579
rect 8113 40539 8171 40545
rect 11238 40536 11244 40588
rect 11296 40576 11302 40588
rect 12069 40579 12127 40585
rect 12069 40576 12081 40579
rect 11296 40548 12081 40576
rect 11296 40536 11302 40548
rect 12069 40545 12081 40548
rect 12115 40576 12127 40579
rect 12158 40576 12164 40588
rect 12115 40548 12164 40576
rect 12115 40545 12127 40548
rect 12069 40539 12127 40545
rect 12158 40536 12164 40548
rect 12216 40536 12222 40588
rect 5902 40468 5908 40520
rect 5960 40508 5966 40520
rect 6362 40508 6368 40520
rect 5960 40480 6368 40508
rect 5960 40468 5966 40480
rect 6362 40468 6368 40480
rect 6420 40468 6426 40520
rect 13004 40508 13032 40616
rect 13081 40579 13139 40585
rect 13081 40545 13093 40579
rect 13127 40576 13139 40579
rect 13446 40576 13452 40588
rect 13127 40548 13452 40576
rect 13127 40545 13139 40548
rect 13081 40539 13139 40545
rect 13446 40536 13452 40548
rect 13504 40536 13510 40588
rect 13173 40511 13231 40517
rect 13173 40508 13185 40511
rect 13004 40480 13185 40508
rect 13173 40477 13185 40480
rect 13219 40477 13231 40511
rect 13173 40471 13231 40477
rect 13265 40511 13323 40517
rect 13265 40477 13277 40511
rect 13311 40508 13323 40511
rect 13354 40508 13360 40520
rect 13311 40480 13360 40508
rect 13311 40477 13323 40480
rect 13265 40471 13323 40477
rect 13354 40468 13360 40480
rect 13412 40468 13418 40520
rect 13630 40468 13636 40520
rect 13688 40468 13694 40520
rect 2777 40443 2835 40449
rect 2777 40409 2789 40443
rect 2823 40409 2835 40443
rect 2777 40403 2835 40409
rect 6641 40443 6699 40449
rect 6641 40409 6653 40443
rect 6687 40440 6699 40443
rect 6730 40440 6736 40452
rect 6687 40412 6736 40440
rect 6687 40409 6699 40412
rect 6641 40403 6699 40409
rect 2792 40372 2820 40403
rect 6730 40400 6736 40412
rect 6788 40400 6794 40452
rect 7098 40440 7104 40452
rect 6840 40412 7104 40440
rect 3329 40375 3387 40381
rect 3329 40372 3341 40375
rect 2792 40344 3341 40372
rect 3329 40341 3341 40344
rect 3375 40372 3387 40375
rect 4154 40372 4160 40384
rect 3375 40344 4160 40372
rect 3375 40341 3387 40344
rect 3329 40335 3387 40341
rect 4154 40332 4160 40344
rect 4212 40332 4218 40384
rect 6546 40332 6552 40384
rect 6604 40372 6610 40384
rect 6840 40372 6868 40412
rect 7098 40400 7104 40412
rect 7156 40400 7162 40452
rect 11333 40443 11391 40449
rect 11333 40409 11345 40443
rect 11379 40440 11391 40443
rect 13648 40440 13676 40468
rect 14384 40449 14412 40616
rect 17862 40604 17868 40656
rect 17920 40644 17926 40656
rect 20809 40647 20867 40653
rect 20809 40644 20821 40647
rect 17920 40616 20821 40644
rect 17920 40604 17926 40616
rect 20809 40613 20821 40616
rect 20855 40644 20867 40647
rect 20990 40644 20996 40656
rect 20855 40616 20996 40644
rect 20855 40613 20867 40616
rect 20809 40607 20867 40613
rect 20990 40604 20996 40616
rect 21048 40644 21054 40656
rect 21634 40644 21640 40656
rect 21048 40616 21640 40644
rect 21048 40604 21054 40616
rect 21634 40604 21640 40616
rect 21692 40604 21698 40656
rect 23937 40647 23995 40653
rect 23937 40613 23949 40647
rect 23983 40644 23995 40647
rect 24210 40644 24216 40656
rect 23983 40616 24216 40644
rect 23983 40613 23995 40616
rect 23937 40607 23995 40613
rect 24210 40604 24216 40616
rect 24268 40604 24274 40656
rect 24489 40647 24547 40653
rect 24489 40613 24501 40647
rect 24535 40644 24547 40647
rect 24762 40644 24768 40656
rect 24535 40616 24768 40644
rect 24535 40613 24547 40616
rect 24489 40607 24547 40613
rect 24762 40604 24768 40616
rect 24820 40604 24826 40656
rect 16022 40536 16028 40588
rect 16080 40536 16086 40588
rect 16117 40579 16175 40585
rect 16117 40545 16129 40579
rect 16163 40576 16175 40579
rect 16666 40576 16672 40588
rect 16163 40548 16672 40576
rect 16163 40545 16175 40548
rect 16117 40539 16175 40545
rect 16666 40536 16672 40548
rect 16724 40536 16730 40588
rect 17129 40579 17187 40585
rect 17129 40545 17141 40579
rect 17175 40576 17187 40579
rect 17957 40579 18015 40585
rect 17957 40576 17969 40579
rect 17175 40548 17969 40576
rect 17175 40545 17187 40548
rect 17129 40539 17187 40545
rect 17957 40545 17969 40548
rect 18003 40545 18015 40579
rect 17957 40539 18015 40545
rect 15654 40468 15660 40520
rect 15712 40508 15718 40520
rect 17144 40508 17172 40539
rect 19150 40536 19156 40588
rect 19208 40576 19214 40588
rect 19521 40579 19579 40585
rect 19521 40576 19533 40579
rect 19208 40548 19533 40576
rect 19208 40536 19214 40548
rect 19521 40545 19533 40548
rect 19567 40545 19579 40579
rect 19521 40539 19579 40545
rect 19705 40579 19763 40585
rect 19705 40545 19717 40579
rect 19751 40576 19763 40579
rect 20070 40576 20076 40588
rect 19751 40548 20076 40576
rect 19751 40545 19763 40548
rect 19705 40539 19763 40545
rect 20070 40536 20076 40548
rect 20128 40536 20134 40588
rect 20533 40579 20591 40585
rect 20533 40545 20545 40579
rect 20579 40576 20591 40579
rect 20714 40576 20720 40588
rect 20579 40548 20720 40576
rect 20579 40545 20591 40548
rect 20533 40539 20591 40545
rect 15712 40480 17172 40508
rect 19797 40511 19855 40517
rect 15712 40468 15718 40480
rect 19797 40477 19809 40511
rect 19843 40508 19855 40511
rect 20548 40508 20576 40539
rect 20714 40536 20720 40548
rect 20772 40576 20778 40588
rect 21450 40576 21456 40588
rect 20772 40548 21456 40576
rect 20772 40536 20778 40548
rect 21450 40536 21456 40548
rect 21508 40536 21514 40588
rect 22278 40536 22284 40588
rect 22336 40576 22342 40588
rect 22925 40579 22983 40585
rect 22925 40576 22937 40579
rect 22336 40548 22937 40576
rect 22336 40536 22342 40548
rect 22925 40545 22937 40548
rect 22971 40576 22983 40579
rect 24946 40576 24952 40588
rect 22971 40548 24952 40576
rect 22971 40545 22983 40548
rect 22925 40539 22983 40545
rect 24946 40536 24952 40548
rect 25004 40536 25010 40588
rect 19843 40480 20576 40508
rect 19843 40477 19855 40480
rect 19797 40471 19855 40477
rect 23382 40468 23388 40520
rect 23440 40468 23446 40520
rect 25317 40511 25375 40517
rect 25317 40508 25329 40511
rect 24872 40480 25329 40508
rect 11379 40412 11413 40440
rect 13372 40412 13676 40440
rect 14369 40443 14427 40449
rect 11379 40409 11391 40412
rect 11333 40403 11391 40409
rect 8389 40375 8447 40381
rect 8389 40372 8401 40375
rect 6604 40344 8401 40372
rect 6604 40332 6610 40344
rect 8389 40341 8401 40344
rect 8435 40372 8447 40375
rect 8570 40372 8576 40384
rect 8435 40344 8576 40372
rect 8435 40341 8447 40344
rect 8389 40335 8447 40341
rect 8570 40332 8576 40344
rect 8628 40332 8634 40384
rect 10226 40332 10232 40384
rect 10284 40372 10290 40384
rect 11348 40372 11376 40403
rect 13372 40384 13400 40412
rect 14369 40409 14381 40443
rect 14415 40440 14427 40443
rect 16390 40440 16396 40452
rect 14415 40412 16396 40440
rect 14415 40409 14427 40412
rect 14369 40403 14427 40409
rect 16390 40400 16396 40412
rect 16448 40400 16454 40452
rect 17773 40443 17831 40449
rect 17773 40409 17785 40443
rect 17819 40440 17831 40443
rect 18690 40440 18696 40452
rect 17819 40412 18696 40440
rect 17819 40409 17831 40412
rect 17773 40403 17831 40409
rect 18690 40400 18696 40412
rect 18748 40400 18754 40452
rect 21358 40400 21364 40452
rect 21416 40440 21422 40452
rect 22649 40443 22707 40449
rect 21416 40412 21482 40440
rect 21416 40400 21422 40412
rect 22649 40409 22661 40443
rect 22695 40440 22707 40443
rect 22695 40412 22876 40440
rect 22695 40409 22707 40412
rect 22649 40403 22707 40409
rect 22848 40384 22876 40412
rect 12529 40375 12587 40381
rect 12529 40372 12541 40375
rect 10284 40344 12541 40372
rect 10284 40332 10290 40344
rect 12529 40341 12541 40344
rect 12575 40341 12587 40375
rect 12529 40335 12587 40341
rect 13354 40332 13360 40384
rect 13412 40332 13418 40384
rect 13633 40375 13691 40381
rect 13633 40341 13645 40375
rect 13679 40372 13691 40375
rect 13998 40372 14004 40384
rect 13679 40344 14004 40372
rect 13679 40341 13691 40344
rect 13633 40335 13691 40341
rect 13998 40332 14004 40344
rect 14056 40332 14062 40384
rect 15470 40332 15476 40384
rect 15528 40372 15534 40384
rect 16209 40375 16267 40381
rect 16209 40372 16221 40375
rect 15528 40344 16221 40372
rect 15528 40332 15534 40344
rect 16209 40341 16221 40344
rect 16255 40341 16267 40375
rect 16209 40335 16267 40341
rect 16577 40375 16635 40381
rect 16577 40341 16589 40375
rect 16623 40372 16635 40375
rect 16666 40372 16672 40384
rect 16623 40344 16672 40372
rect 16623 40341 16635 40344
rect 16577 40335 16635 40341
rect 16666 40332 16672 40344
rect 16724 40332 16730 40384
rect 17865 40375 17923 40381
rect 17865 40341 17877 40375
rect 17911 40372 17923 40375
rect 18322 40372 18328 40384
rect 17911 40344 18328 40372
rect 17911 40341 17923 40344
rect 17865 40335 17923 40341
rect 18322 40332 18328 40344
rect 18380 40372 18386 40384
rect 18598 40372 18604 40384
rect 18380 40344 18604 40372
rect 18380 40332 18386 40344
rect 18598 40332 18604 40344
rect 18656 40332 18662 40384
rect 20162 40332 20168 40384
rect 20220 40332 20226 40384
rect 21177 40375 21235 40381
rect 21177 40341 21189 40375
rect 21223 40372 21235 40375
rect 21634 40372 21640 40384
rect 21223 40344 21640 40372
rect 21223 40341 21235 40344
rect 21177 40335 21235 40341
rect 21634 40332 21640 40344
rect 21692 40332 21698 40384
rect 22830 40332 22836 40384
rect 22888 40332 22894 40384
rect 24210 40332 24216 40384
rect 24268 40332 24274 40384
rect 24762 40332 24768 40384
rect 24820 40372 24826 40384
rect 24872 40381 24900 40480
rect 25317 40477 25329 40480
rect 25363 40477 25375 40511
rect 25317 40471 25375 40477
rect 24857 40375 24915 40381
rect 24857 40372 24869 40375
rect 24820 40344 24869 40372
rect 24820 40332 24826 40344
rect 24857 40341 24869 40344
rect 24903 40341 24915 40375
rect 24857 40335 24915 40341
rect 1104 40282 25852 40304
rect 1104 40230 7950 40282
rect 8002 40230 8014 40282
rect 8066 40230 8078 40282
rect 8130 40230 8142 40282
rect 8194 40230 8206 40282
rect 8258 40230 17950 40282
rect 18002 40230 18014 40282
rect 18066 40230 18078 40282
rect 18130 40230 18142 40282
rect 18194 40230 18206 40282
rect 18258 40230 25852 40282
rect 1104 40208 25852 40230
rect 7558 40128 7564 40180
rect 7616 40168 7622 40180
rect 8113 40171 8171 40177
rect 8113 40168 8125 40171
rect 7616 40140 8125 40168
rect 7616 40128 7622 40140
rect 8113 40137 8125 40140
rect 8159 40137 8171 40171
rect 8113 40131 8171 40137
rect 8481 40171 8539 40177
rect 8481 40137 8493 40171
rect 8527 40168 8539 40171
rect 10042 40168 10048 40180
rect 8527 40140 10048 40168
rect 8527 40137 8539 40140
rect 8481 40131 8539 40137
rect 10042 40128 10048 40140
rect 10100 40128 10106 40180
rect 14274 40168 14280 40180
rect 10244 40140 14280 40168
rect 6362 40060 6368 40112
rect 6420 40100 6426 40112
rect 9033 40103 9091 40109
rect 9033 40100 9045 40103
rect 6420 40072 9045 40100
rect 6420 40060 6426 40072
rect 9033 40069 9045 40072
rect 9079 40100 9091 40103
rect 9398 40100 9404 40112
rect 9079 40072 9404 40100
rect 9079 40069 9091 40072
rect 9033 40063 9091 40069
rect 9398 40060 9404 40072
rect 9456 40060 9462 40112
rect 10244 40100 10272 40140
rect 14274 40128 14280 40140
rect 14332 40168 14338 40180
rect 14829 40171 14887 40177
rect 14829 40168 14841 40171
rect 14332 40140 14841 40168
rect 14332 40128 14338 40140
rect 14829 40137 14841 40140
rect 14875 40137 14887 40171
rect 14829 40131 14887 40137
rect 15565 40171 15623 40177
rect 15565 40137 15577 40171
rect 15611 40168 15623 40171
rect 20346 40168 20352 40180
rect 15611 40140 20352 40168
rect 15611 40137 15623 40140
rect 15565 40131 15623 40137
rect 13722 40100 13728 40112
rect 9784 40072 10272 40100
rect 13662 40072 13728 40100
rect 4062 39992 4068 40044
rect 4120 40032 4126 40044
rect 7377 40035 7435 40041
rect 7377 40032 7389 40035
rect 4120 40004 7389 40032
rect 4120 39992 4126 40004
rect 7377 40001 7389 40004
rect 7423 40032 7435 40035
rect 8021 40035 8079 40041
rect 8021 40032 8033 40035
rect 7423 40004 8033 40032
rect 7423 40001 7435 40004
rect 7377 39995 7435 40001
rect 8021 40001 8033 40004
rect 8067 40001 8079 40035
rect 9416 40032 9444 40060
rect 9674 40032 9680 40044
rect 9416 40004 9680 40032
rect 8021 39995 8079 40001
rect 7098 39924 7104 39976
rect 7156 39964 7162 39976
rect 7837 39967 7895 39973
rect 7837 39964 7849 39967
rect 7156 39936 7849 39964
rect 7156 39924 7162 39936
rect 7837 39933 7849 39936
rect 7883 39933 7895 39967
rect 8036 39964 8064 39995
rect 9674 39992 9680 40004
rect 9732 39992 9738 40044
rect 9784 39964 9812 40072
rect 13722 40060 13728 40072
rect 13780 40100 13786 40112
rect 14366 40100 14372 40112
rect 13780 40072 14372 40100
rect 13780 40060 13786 40072
rect 14366 40060 14372 40072
rect 14424 40060 14430 40112
rect 14844 40100 14872 40131
rect 20346 40128 20352 40140
rect 20404 40168 20410 40180
rect 20530 40168 20536 40180
rect 20404 40140 20536 40168
rect 20404 40128 20410 40140
rect 20530 40128 20536 40140
rect 20588 40128 20594 40180
rect 20990 40128 20996 40180
rect 21048 40128 21054 40180
rect 21453 40171 21511 40177
rect 21453 40137 21465 40171
rect 21499 40137 21511 40171
rect 21453 40131 21511 40137
rect 15657 40103 15715 40109
rect 15657 40100 15669 40103
rect 14844 40072 15669 40100
rect 15657 40069 15669 40072
rect 15703 40069 15715 40103
rect 15657 40063 15715 40069
rect 16390 40060 16396 40112
rect 16448 40100 16454 40112
rect 16942 40100 16948 40112
rect 16448 40072 16948 40100
rect 16448 40060 16454 40072
rect 16942 40060 16948 40072
rect 17000 40060 17006 40112
rect 21085 40103 21143 40109
rect 21085 40069 21097 40103
rect 21131 40069 21143 40103
rect 21468 40100 21496 40131
rect 21726 40128 21732 40180
rect 21784 40168 21790 40180
rect 22373 40171 22431 40177
rect 22373 40168 22385 40171
rect 21784 40140 22385 40168
rect 21784 40128 21790 40140
rect 22373 40137 22385 40140
rect 22419 40137 22431 40171
rect 22373 40131 22431 40137
rect 22646 40128 22652 40180
rect 22704 40168 22710 40180
rect 22741 40171 22799 40177
rect 22741 40168 22753 40171
rect 22704 40140 22753 40168
rect 22704 40128 22710 40140
rect 22741 40137 22753 40140
rect 22787 40137 22799 40171
rect 22741 40131 22799 40137
rect 23658 40100 23664 40112
rect 21468 40072 23664 40100
rect 21085 40063 21143 40069
rect 9861 40035 9919 40041
rect 9861 40001 9873 40035
rect 9907 40032 9919 40035
rect 10226 40032 10232 40044
rect 9907 40004 10232 40032
rect 9907 40001 9919 40004
rect 9861 39995 9919 40001
rect 10226 39992 10232 40004
rect 10284 39992 10290 40044
rect 12158 39992 12164 40044
rect 12216 39992 12222 40044
rect 21100 40032 21128 40063
rect 23658 40060 23664 40072
rect 23716 40060 23722 40112
rect 21818 40032 21824 40044
rect 14292 40004 15884 40032
rect 8036 39936 9812 39964
rect 7837 39927 7895 39933
rect 12434 39924 12440 39976
rect 12492 39964 12498 39976
rect 13814 39964 13820 39976
rect 12492 39936 13820 39964
rect 12492 39924 12498 39936
rect 13814 39924 13820 39936
rect 13872 39964 13878 39976
rect 14292 39964 14320 40004
rect 13872 39936 14320 39964
rect 13872 39924 13878 39936
rect 14366 39924 14372 39976
rect 14424 39924 14430 39976
rect 15856 39973 15884 40004
rect 19812 40004 21824 40032
rect 15841 39967 15899 39973
rect 15841 39933 15853 39967
rect 15887 39964 15899 39967
rect 16942 39964 16948 39976
rect 15887 39936 16948 39964
rect 15887 39933 15899 39936
rect 15841 39927 15899 39933
rect 16942 39924 16948 39936
rect 17000 39924 17006 39976
rect 7374 39788 7380 39840
rect 7432 39828 7438 39840
rect 8202 39828 8208 39840
rect 7432 39800 8208 39828
rect 7432 39788 7438 39800
rect 8202 39788 8208 39800
rect 8260 39788 8266 39840
rect 10226 39788 10232 39840
rect 10284 39788 10290 39840
rect 11330 39788 11336 39840
rect 11388 39828 11394 39840
rect 11790 39828 11796 39840
rect 11388 39800 11796 39828
rect 11388 39788 11394 39800
rect 11790 39788 11796 39800
rect 11848 39828 11854 39840
rect 13906 39828 13912 39840
rect 11848 39800 13912 39828
rect 11848 39788 11854 39800
rect 13906 39788 13912 39800
rect 13964 39788 13970 39840
rect 15194 39788 15200 39840
rect 15252 39788 15258 39840
rect 19702 39788 19708 39840
rect 19760 39828 19766 39840
rect 19812 39828 19840 40004
rect 21818 39992 21824 40004
rect 21876 39992 21882 40044
rect 24578 40032 24584 40044
rect 22204 40004 24584 40032
rect 20714 39924 20720 39976
rect 20772 39964 20778 39976
rect 20809 39967 20867 39973
rect 20809 39964 20821 39967
rect 20772 39936 20821 39964
rect 20772 39924 20778 39936
rect 20809 39933 20821 39936
rect 20855 39964 20867 39967
rect 22002 39964 22008 39976
rect 20855 39936 22008 39964
rect 20855 39933 20867 39936
rect 20809 39927 20867 39933
rect 22002 39924 22008 39936
rect 22060 39924 22066 39976
rect 22204 39973 22232 40004
rect 24578 39992 24584 40004
rect 24636 39992 24642 40044
rect 22189 39967 22247 39973
rect 22189 39933 22201 39967
rect 22235 39933 22247 39967
rect 22189 39927 22247 39933
rect 22281 39967 22339 39973
rect 22281 39933 22293 39967
rect 22327 39933 22339 39967
rect 22281 39927 22339 39933
rect 19886 39856 19892 39908
rect 19944 39896 19950 39908
rect 20070 39896 20076 39908
rect 19944 39868 20076 39896
rect 19944 39856 19950 39868
rect 20070 39856 20076 39868
rect 20128 39896 20134 39908
rect 20349 39899 20407 39905
rect 20349 39896 20361 39899
rect 20128 39868 20361 39896
rect 20128 39856 20134 39868
rect 20349 39865 20361 39868
rect 20395 39865 20407 39899
rect 20349 39859 20407 39865
rect 20165 39831 20223 39837
rect 20165 39828 20177 39831
rect 19760 39800 20177 39828
rect 19760 39788 19766 39800
rect 20165 39797 20177 39800
rect 20211 39797 20223 39831
rect 20165 39791 20223 39797
rect 20438 39788 20444 39840
rect 20496 39828 20502 39840
rect 22296 39828 22324 39927
rect 22646 39924 22652 39976
rect 22704 39964 22710 39976
rect 23566 39964 23572 39976
rect 22704 39936 23572 39964
rect 22704 39924 22710 39936
rect 23566 39924 23572 39936
rect 23624 39924 23630 39976
rect 23658 39924 23664 39976
rect 23716 39964 23722 39976
rect 23753 39967 23811 39973
rect 23753 39964 23765 39967
rect 23716 39936 23765 39964
rect 23716 39924 23722 39936
rect 23753 39933 23765 39936
rect 23799 39933 23811 39967
rect 23753 39927 23811 39933
rect 24029 39967 24087 39973
rect 24029 39933 24041 39967
rect 24075 39964 24087 39967
rect 24210 39964 24216 39976
rect 24075 39936 24216 39964
rect 24075 39933 24087 39936
rect 24029 39927 24087 39933
rect 24210 39924 24216 39936
rect 24268 39964 24274 39976
rect 24946 39964 24952 39976
rect 24268 39936 24952 39964
rect 24268 39924 24274 39936
rect 24946 39924 24952 39936
rect 25004 39924 25010 39976
rect 25038 39924 25044 39976
rect 25096 39924 25102 39976
rect 25314 39924 25320 39976
rect 25372 39924 25378 39976
rect 20496 39800 22324 39828
rect 20496 39788 20502 39800
rect 1104 39738 25852 39760
rect 1104 39686 2950 39738
rect 3002 39686 3014 39738
rect 3066 39686 3078 39738
rect 3130 39686 3142 39738
rect 3194 39686 3206 39738
rect 3258 39686 12950 39738
rect 13002 39686 13014 39738
rect 13066 39686 13078 39738
rect 13130 39686 13142 39738
rect 13194 39686 13206 39738
rect 13258 39686 22950 39738
rect 23002 39686 23014 39738
rect 23066 39686 23078 39738
rect 23130 39686 23142 39738
rect 23194 39686 23206 39738
rect 23258 39686 25852 39738
rect 1104 39664 25852 39686
rect 8386 39584 8392 39636
rect 8444 39584 8450 39636
rect 14277 39627 14335 39633
rect 8496 39596 12112 39624
rect 6730 39516 6736 39568
rect 6788 39556 6794 39568
rect 8496 39556 8524 39596
rect 6788 39528 8524 39556
rect 6788 39516 6794 39528
rect 9858 39516 9864 39568
rect 9916 39556 9922 39568
rect 12084 39556 12112 39596
rect 14277 39593 14289 39627
rect 14323 39624 14335 39627
rect 14458 39624 14464 39636
rect 14323 39596 14464 39624
rect 14323 39593 14335 39596
rect 14277 39587 14335 39593
rect 14458 39584 14464 39596
rect 14516 39584 14522 39636
rect 19518 39584 19524 39636
rect 19576 39584 19582 39636
rect 20806 39584 20812 39636
rect 20864 39624 20870 39636
rect 20990 39624 20996 39636
rect 20864 39596 20996 39624
rect 20864 39584 20870 39596
rect 20990 39584 20996 39596
rect 21048 39584 21054 39636
rect 22738 39584 22744 39636
rect 22796 39624 22802 39636
rect 23198 39624 23204 39636
rect 22796 39596 23204 39624
rect 22796 39584 22802 39596
rect 23198 39584 23204 39596
rect 23256 39584 23262 39636
rect 23382 39584 23388 39636
rect 23440 39624 23446 39636
rect 23569 39627 23627 39633
rect 23569 39624 23581 39627
rect 23440 39596 23581 39624
rect 23440 39584 23446 39596
rect 23569 39593 23581 39596
rect 23615 39593 23627 39627
rect 23569 39587 23627 39593
rect 9916 39528 10824 39556
rect 12084 39528 12434 39556
rect 9916 39516 9922 39528
rect 6914 39448 6920 39500
rect 6972 39488 6978 39500
rect 7745 39491 7803 39497
rect 7745 39488 7757 39491
rect 6972 39460 7757 39488
rect 6972 39448 6978 39460
rect 7745 39457 7757 39460
rect 7791 39457 7803 39491
rect 9217 39491 9275 39497
rect 9217 39488 9229 39491
rect 7745 39451 7803 39457
rect 8128 39460 9229 39488
rect 7374 39380 7380 39432
rect 7432 39420 7438 39432
rect 8128 39420 8156 39460
rect 9217 39457 9229 39460
rect 9263 39457 9275 39491
rect 9217 39451 9275 39457
rect 10413 39491 10471 39497
rect 10413 39457 10425 39491
rect 10459 39488 10471 39491
rect 10686 39488 10692 39500
rect 10459 39460 10692 39488
rect 10459 39457 10471 39460
rect 10413 39451 10471 39457
rect 10686 39448 10692 39460
rect 10744 39448 10750 39500
rect 7432 39392 8156 39420
rect 7432 39380 7438 39392
rect 8202 39380 8208 39432
rect 8260 39420 8266 39432
rect 8665 39423 8723 39429
rect 8665 39420 8677 39423
rect 8260 39392 8677 39420
rect 8260 39380 8266 39392
rect 8665 39389 8677 39392
rect 8711 39420 8723 39423
rect 9493 39423 9551 39429
rect 9493 39420 9505 39423
rect 8711 39392 9505 39420
rect 8711 39389 8723 39392
rect 8665 39383 8723 39389
rect 9493 39389 9505 39392
rect 9539 39420 9551 39423
rect 9539 39392 10640 39420
rect 10796 39406 10824 39528
rect 11882 39448 11888 39500
rect 11940 39448 11946 39500
rect 12158 39448 12164 39500
rect 12216 39448 12222 39500
rect 12406 39488 12434 39528
rect 13630 39516 13636 39568
rect 13688 39556 13694 39568
rect 15749 39559 15807 39565
rect 15749 39556 15761 39559
rect 13688 39528 15761 39556
rect 13688 39516 13694 39528
rect 15749 39525 15761 39528
rect 15795 39525 15807 39559
rect 18414 39556 18420 39568
rect 15749 39519 15807 39525
rect 16132 39528 18420 39556
rect 13173 39491 13231 39497
rect 13173 39488 13185 39491
rect 12406 39460 13185 39488
rect 13173 39457 13185 39460
rect 13219 39457 13231 39491
rect 13173 39451 13231 39457
rect 13906 39448 13912 39500
rect 13964 39488 13970 39500
rect 14829 39491 14887 39497
rect 14829 39488 14841 39491
rect 13964 39460 14841 39488
rect 13964 39448 13970 39460
rect 14829 39457 14841 39460
rect 14875 39457 14887 39491
rect 14829 39451 14887 39457
rect 9539 39389 9551 39392
rect 9493 39383 9551 39389
rect 7929 39355 7987 39361
rect 7929 39321 7941 39355
rect 7975 39352 7987 39355
rect 9306 39352 9312 39364
rect 7975 39324 9312 39352
rect 7975 39321 7987 39324
rect 7929 39315 7987 39321
rect 9306 39312 9312 39324
rect 9364 39312 9370 39364
rect 9401 39355 9459 39361
rect 9401 39321 9413 39355
rect 9447 39352 9459 39355
rect 9950 39352 9956 39364
rect 9447 39324 9956 39352
rect 9447 39321 9459 39324
rect 9401 39315 9459 39321
rect 9950 39312 9956 39324
rect 10008 39352 10014 39364
rect 10502 39352 10508 39364
rect 10008 39324 10508 39352
rect 10008 39312 10014 39324
rect 10502 39312 10508 39324
rect 10560 39312 10566 39364
rect 8021 39287 8079 39293
rect 8021 39253 8033 39287
rect 8067 39284 8079 39287
rect 8478 39284 8484 39296
rect 8067 39256 8484 39284
rect 8067 39253 8079 39256
rect 8021 39247 8079 39253
rect 8478 39244 8484 39256
rect 8536 39244 8542 39296
rect 9858 39244 9864 39296
rect 9916 39244 9922 39296
rect 10612 39284 10640 39392
rect 12250 39380 12256 39432
rect 12308 39420 12314 39432
rect 13081 39423 13139 39429
rect 13081 39420 13093 39423
rect 12308 39392 13093 39420
rect 12308 39380 12314 39392
rect 13081 39389 13093 39392
rect 13127 39389 13139 39423
rect 13081 39383 13139 39389
rect 14737 39423 14795 39429
rect 14737 39389 14749 39423
rect 14783 39420 14795 39423
rect 15194 39420 15200 39432
rect 14783 39392 15200 39420
rect 14783 39389 14795 39392
rect 14737 39383 14795 39389
rect 15194 39380 15200 39392
rect 15252 39380 15258 39432
rect 12989 39355 13047 39361
rect 12989 39321 13001 39355
rect 13035 39352 13047 39355
rect 16132 39352 16160 39528
rect 18414 39516 18420 39528
rect 18472 39556 18478 39568
rect 25038 39556 25044 39568
rect 18472 39528 25044 39556
rect 18472 39516 18478 39528
rect 25038 39516 25044 39528
rect 25096 39516 25102 39568
rect 16393 39491 16451 39497
rect 16393 39457 16405 39491
rect 16439 39457 16451 39491
rect 16393 39451 16451 39457
rect 16408 39420 16436 39451
rect 17586 39448 17592 39500
rect 17644 39448 17650 39500
rect 17678 39448 17684 39500
rect 17736 39448 17742 39500
rect 20165 39491 20223 39497
rect 20165 39457 20177 39491
rect 20211 39488 20223 39491
rect 20806 39488 20812 39500
rect 20211 39460 20812 39488
rect 20211 39457 20223 39460
rect 20165 39451 20223 39457
rect 20806 39448 20812 39460
rect 20864 39448 20870 39500
rect 20901 39491 20959 39497
rect 20901 39457 20913 39491
rect 20947 39457 20959 39491
rect 20901 39451 20959 39457
rect 18782 39420 18788 39432
rect 16408 39392 18788 39420
rect 18782 39380 18788 39392
rect 18840 39380 18846 39432
rect 20916 39420 20944 39451
rect 21634 39448 21640 39500
rect 21692 39488 21698 39500
rect 22465 39491 22523 39497
rect 22465 39488 22477 39491
rect 21692 39460 22477 39488
rect 21692 39448 21698 39460
rect 22465 39457 22477 39460
rect 22511 39457 22523 39491
rect 22465 39451 22523 39457
rect 23017 39491 23075 39497
rect 23017 39457 23029 39491
rect 23063 39488 23075 39491
rect 23063 39460 24164 39488
rect 23063 39457 23075 39460
rect 23017 39451 23075 39457
rect 22830 39420 22836 39432
rect 20916 39392 22836 39420
rect 22830 39380 22836 39392
rect 22888 39380 22894 39432
rect 13035 39324 16160 39352
rect 16209 39355 16267 39361
rect 13035 39321 13047 39324
rect 12989 39315 13047 39321
rect 16209 39321 16221 39355
rect 16255 39352 16267 39355
rect 19242 39352 19248 39364
rect 16255 39324 19248 39352
rect 16255 39321 16267 39324
rect 16209 39315 16267 39321
rect 19242 39312 19248 39324
rect 19300 39312 19306 39364
rect 20622 39352 20628 39364
rect 19904 39324 20628 39352
rect 19904 39296 19932 39324
rect 20622 39312 20628 39324
rect 20680 39352 20686 39364
rect 21085 39355 21143 39361
rect 21085 39352 21097 39355
rect 20680 39324 21097 39352
rect 20680 39312 20686 39324
rect 21085 39321 21097 39324
rect 21131 39321 21143 39355
rect 22281 39355 22339 39361
rect 22281 39352 22293 39355
rect 21085 39315 21143 39321
rect 21468 39324 22293 39352
rect 11238 39284 11244 39296
rect 10612 39256 11244 39284
rect 11238 39244 11244 39256
rect 11296 39244 11302 39296
rect 12618 39244 12624 39296
rect 12676 39244 12682 39296
rect 14642 39244 14648 39296
rect 14700 39244 14706 39296
rect 15930 39244 15936 39296
rect 15988 39284 15994 39296
rect 16117 39287 16175 39293
rect 16117 39284 16129 39287
rect 15988 39256 16129 39284
rect 15988 39244 15994 39256
rect 16117 39253 16129 39256
rect 16163 39253 16175 39287
rect 16117 39247 16175 39253
rect 16574 39244 16580 39296
rect 16632 39284 16638 39296
rect 17773 39287 17831 39293
rect 17773 39284 17785 39287
rect 16632 39256 17785 39284
rect 16632 39244 16638 39256
rect 17773 39253 17785 39256
rect 17819 39253 17831 39287
rect 17773 39247 17831 39253
rect 18141 39287 18199 39293
rect 18141 39253 18153 39287
rect 18187 39284 18199 39287
rect 19794 39284 19800 39296
rect 18187 39256 19800 39284
rect 18187 39253 18199 39256
rect 18141 39247 18199 39253
rect 19794 39244 19800 39256
rect 19852 39244 19858 39296
rect 19886 39244 19892 39296
rect 19944 39244 19950 39296
rect 19981 39287 20039 39293
rect 19981 39253 19993 39287
rect 20027 39284 20039 39287
rect 20070 39284 20076 39296
rect 20027 39256 20076 39284
rect 20027 39253 20039 39256
rect 19981 39247 20039 39253
rect 20070 39244 20076 39256
rect 20128 39284 20134 39296
rect 21468 39293 21496 39324
rect 22281 39321 22293 39324
rect 22327 39321 22339 39355
rect 22281 39315 22339 39321
rect 22373 39355 22431 39361
rect 22373 39321 22385 39355
rect 22419 39352 22431 39355
rect 22462 39352 22468 39364
rect 22419 39324 22468 39352
rect 22419 39321 22431 39324
rect 22373 39315 22431 39321
rect 22462 39312 22468 39324
rect 22520 39312 22526 39364
rect 20993 39287 21051 39293
rect 20993 39284 21005 39287
rect 20128 39256 21005 39284
rect 20128 39244 20134 39256
rect 20993 39253 21005 39256
rect 21039 39253 21051 39287
rect 20993 39247 21051 39253
rect 21453 39287 21511 39293
rect 21453 39253 21465 39287
rect 21499 39253 21511 39287
rect 21453 39247 21511 39253
rect 21910 39244 21916 39296
rect 21968 39244 21974 39296
rect 22094 39244 22100 39296
rect 22152 39284 22158 39296
rect 23032 39284 23060 39451
rect 23382 39380 23388 39432
rect 23440 39420 23446 39432
rect 24029 39423 24087 39429
rect 24029 39420 24041 39423
rect 23440 39392 24041 39420
rect 23440 39380 23446 39392
rect 24029 39389 24041 39392
rect 24075 39389 24087 39423
rect 24136 39420 24164 39460
rect 24670 39448 24676 39500
rect 24728 39488 24734 39500
rect 25133 39491 25191 39497
rect 25133 39488 25145 39491
rect 24728 39460 25145 39488
rect 24728 39448 24734 39460
rect 25133 39457 25145 39460
rect 25179 39457 25191 39491
rect 25133 39451 25191 39457
rect 25406 39420 25412 39432
rect 24136 39392 25412 39420
rect 24029 39383 24087 39389
rect 25406 39380 25412 39392
rect 25464 39380 25470 39432
rect 23198 39312 23204 39364
rect 23256 39352 23262 39364
rect 24949 39355 25007 39361
rect 24949 39352 24961 39355
rect 23256 39324 24961 39352
rect 23256 39312 23262 39324
rect 24949 39321 24961 39324
rect 24995 39321 25007 39355
rect 24949 39315 25007 39321
rect 25041 39355 25099 39361
rect 25041 39321 25053 39355
rect 25087 39352 25099 39355
rect 25130 39352 25136 39364
rect 25087 39324 25136 39352
rect 25087 39321 25099 39324
rect 25041 39315 25099 39321
rect 25130 39312 25136 39324
rect 25188 39312 25194 39364
rect 22152 39256 23060 39284
rect 23845 39287 23903 39293
rect 22152 39244 22158 39256
rect 23845 39253 23857 39287
rect 23891 39284 23903 39287
rect 24026 39284 24032 39296
rect 23891 39256 24032 39284
rect 23891 39253 23903 39256
rect 23845 39247 23903 39253
rect 24026 39244 24032 39256
rect 24084 39244 24090 39296
rect 24581 39287 24639 39293
rect 24581 39253 24593 39287
rect 24627 39284 24639 39287
rect 24670 39284 24676 39296
rect 24627 39256 24676 39284
rect 24627 39253 24639 39256
rect 24581 39247 24639 39253
rect 24670 39244 24676 39256
rect 24728 39244 24734 39296
rect 1104 39194 25852 39216
rect 1104 39142 7950 39194
rect 8002 39142 8014 39194
rect 8066 39142 8078 39194
rect 8130 39142 8142 39194
rect 8194 39142 8206 39194
rect 8258 39142 17950 39194
rect 18002 39142 18014 39194
rect 18066 39142 18078 39194
rect 18130 39142 18142 39194
rect 18194 39142 18206 39194
rect 18258 39142 25852 39194
rect 1104 39120 25852 39142
rect 5997 39083 6055 39089
rect 4908 39052 5948 39080
rect 4908 39012 4936 39052
rect 4982 39012 4988 39024
rect 4908 38984 4988 39012
rect 4982 38972 4988 38984
rect 5040 38972 5046 39024
rect 5920 39012 5948 39052
rect 5997 39049 6009 39083
rect 6043 39080 6055 39083
rect 6730 39080 6736 39092
rect 6043 39052 6736 39080
rect 6043 39049 6055 39052
rect 5997 39043 6055 39049
rect 6730 39040 6736 39052
rect 6788 39040 6794 39092
rect 9766 39040 9772 39092
rect 9824 39040 9830 39092
rect 12342 39040 12348 39092
rect 12400 39080 12406 39092
rect 12529 39083 12587 39089
rect 12529 39080 12541 39083
rect 12400 39052 12541 39080
rect 12400 39040 12406 39052
rect 12529 39049 12541 39052
rect 12575 39049 12587 39083
rect 12529 39043 12587 39049
rect 12894 39040 12900 39092
rect 12952 39080 12958 39092
rect 13722 39080 13728 39092
rect 12952 39052 13728 39080
rect 12952 39040 12958 39052
rect 13722 39040 13728 39052
rect 13780 39040 13786 39092
rect 14093 39083 14151 39089
rect 14093 39049 14105 39083
rect 14139 39080 14151 39083
rect 14366 39080 14372 39092
rect 14139 39052 14372 39080
rect 14139 39049 14151 39052
rect 14093 39043 14151 39049
rect 14366 39040 14372 39052
rect 14424 39040 14430 39092
rect 14461 39083 14519 39089
rect 14461 39049 14473 39083
rect 14507 39080 14519 39083
rect 15470 39080 15476 39092
rect 14507 39052 15476 39080
rect 14507 39049 14519 39052
rect 14461 39043 14519 39049
rect 15470 39040 15476 39052
rect 15528 39040 15534 39092
rect 15749 39083 15807 39089
rect 15749 39049 15761 39083
rect 15795 39080 15807 39083
rect 16850 39080 16856 39092
rect 15795 39052 16856 39080
rect 15795 39049 15807 39052
rect 15749 39043 15807 39049
rect 16850 39040 16856 39052
rect 16908 39040 16914 39092
rect 17586 39040 17592 39092
rect 17644 39080 17650 39092
rect 17862 39080 17868 39092
rect 17644 39052 17868 39080
rect 17644 39040 17650 39052
rect 17862 39040 17868 39052
rect 17920 39040 17926 39092
rect 20162 39040 20168 39092
rect 20220 39040 20226 39092
rect 20622 39040 20628 39092
rect 20680 39080 20686 39092
rect 21085 39083 21143 39089
rect 21085 39080 21097 39083
rect 20680 39052 21097 39080
rect 20680 39040 20686 39052
rect 21085 39049 21097 39052
rect 21131 39080 21143 39083
rect 23477 39083 23535 39089
rect 23477 39080 23489 39083
rect 21131 39052 21864 39080
rect 21131 39049 21143 39052
rect 21085 39043 21143 39049
rect 6365 39015 6423 39021
rect 6365 39012 6377 39015
rect 5920 38984 6377 39012
rect 6365 38981 6377 38984
rect 6411 39012 6423 39015
rect 6546 39012 6552 39024
rect 6411 38984 6552 39012
rect 6411 38981 6423 38984
rect 6365 38975 6423 38981
rect 6546 38972 6552 38984
rect 6604 38972 6610 39024
rect 10137 39015 10195 39021
rect 10137 38981 10149 39015
rect 10183 39012 10195 39015
rect 10318 39012 10324 39024
rect 10183 38984 10324 39012
rect 10183 38981 10195 38984
rect 10137 38975 10195 38981
rect 10318 38972 10324 38984
rect 10376 38972 10382 39024
rect 10502 38972 10508 39024
rect 10560 39012 10566 39024
rect 14734 39012 14740 39024
rect 10560 38984 14740 39012
rect 10560 38972 10566 38984
rect 14734 38972 14740 38984
rect 14792 38972 14798 39024
rect 18598 38972 18604 39024
rect 18656 38972 18662 39024
rect 19058 38972 19064 39024
rect 19116 39012 19122 39024
rect 20257 39015 20315 39021
rect 20257 39012 20269 39015
rect 19116 38984 20269 39012
rect 19116 38972 19122 38984
rect 20257 38981 20269 38984
rect 20303 38981 20315 39015
rect 20257 38975 20315 38981
rect 1210 38904 1216 38956
rect 1268 38944 1274 38956
rect 1581 38947 1639 38953
rect 1581 38944 1593 38947
rect 1268 38916 1593 38944
rect 1268 38904 1274 38916
rect 1581 38913 1593 38916
rect 1627 38944 1639 38947
rect 2041 38947 2099 38953
rect 2041 38944 2053 38947
rect 1627 38916 2053 38944
rect 1627 38913 1639 38916
rect 1581 38907 1639 38913
rect 2041 38913 2053 38916
rect 2087 38913 2099 38947
rect 2041 38907 2099 38913
rect 12158 38904 12164 38956
rect 12216 38904 12222 38956
rect 14090 38944 14096 38956
rect 13924 38916 14096 38944
rect 4249 38879 4307 38885
rect 4249 38845 4261 38879
rect 4295 38845 4307 38879
rect 4249 38839 4307 38845
rect 4525 38879 4583 38885
rect 4525 38845 4537 38879
rect 4571 38876 4583 38879
rect 4982 38876 4988 38888
rect 4571 38848 4988 38876
rect 4571 38845 4583 38848
rect 4525 38839 4583 38845
rect 1765 38743 1823 38749
rect 1765 38709 1777 38743
rect 1811 38740 1823 38743
rect 3970 38740 3976 38752
rect 1811 38712 3976 38740
rect 1811 38709 1823 38712
rect 1765 38703 1823 38709
rect 3970 38700 3976 38712
rect 4028 38700 4034 38752
rect 4264 38740 4292 38839
rect 4982 38836 4988 38848
rect 5040 38836 5046 38888
rect 8570 38836 8576 38888
rect 8628 38836 8634 38888
rect 10229 38879 10287 38885
rect 10229 38845 10241 38879
rect 10275 38845 10287 38879
rect 10229 38839 10287 38845
rect 10244 38808 10272 38839
rect 10410 38836 10416 38888
rect 10468 38836 10474 38888
rect 10965 38879 11023 38885
rect 10965 38845 10977 38879
rect 11011 38876 11023 38879
rect 11054 38876 11060 38888
rect 11011 38848 11060 38876
rect 11011 38845 11023 38848
rect 10965 38839 11023 38845
rect 11054 38836 11060 38848
rect 11112 38836 11118 38888
rect 11790 38836 11796 38888
rect 11848 38876 11854 38888
rect 11885 38879 11943 38885
rect 11885 38876 11897 38879
rect 11848 38848 11897 38876
rect 11848 38836 11854 38848
rect 11885 38845 11897 38848
rect 11931 38845 11943 38879
rect 11885 38839 11943 38845
rect 11974 38836 11980 38888
rect 12032 38876 12038 38888
rect 12069 38879 12127 38885
rect 12069 38876 12081 38879
rect 12032 38848 12081 38876
rect 12032 38836 12038 38848
rect 12069 38845 12081 38848
rect 12115 38845 12127 38879
rect 12069 38839 12127 38845
rect 12250 38836 12256 38888
rect 12308 38876 12314 38888
rect 13924 38885 13952 38916
rect 14090 38904 14096 38916
rect 14148 38904 14154 38956
rect 15194 38904 15200 38956
rect 15252 38944 15258 38956
rect 15841 38947 15899 38953
rect 15841 38944 15853 38947
rect 15252 38916 15853 38944
rect 15252 38904 15258 38916
rect 15841 38913 15853 38916
rect 15887 38913 15899 38947
rect 20993 38947 21051 38953
rect 20993 38944 21005 38947
rect 15841 38907 15899 38913
rect 20088 38916 21005 38944
rect 13909 38879 13967 38885
rect 12308 38848 13216 38876
rect 12308 38836 12314 38848
rect 12434 38808 12440 38820
rect 10244 38780 12440 38808
rect 12434 38768 12440 38780
rect 12492 38768 12498 38820
rect 5902 38740 5908 38752
rect 4264 38712 5908 38740
rect 5902 38700 5908 38712
rect 5960 38700 5966 38752
rect 11330 38700 11336 38752
rect 11388 38740 11394 38752
rect 12250 38740 12256 38752
rect 11388 38712 12256 38740
rect 11388 38700 11394 38712
rect 12250 38700 12256 38712
rect 12308 38700 12314 38752
rect 12342 38700 12348 38752
rect 12400 38740 12406 38752
rect 12894 38740 12900 38752
rect 12400 38712 12900 38740
rect 12400 38700 12406 38712
rect 12894 38700 12900 38712
rect 12952 38700 12958 38752
rect 13188 38740 13216 38848
rect 13909 38845 13921 38879
rect 13955 38845 13967 38879
rect 13909 38839 13967 38845
rect 14001 38879 14059 38885
rect 14001 38845 14013 38879
rect 14047 38845 14059 38879
rect 14001 38839 14059 38845
rect 13357 38743 13415 38749
rect 13357 38740 13369 38743
rect 13188 38712 13369 38740
rect 13357 38709 13369 38712
rect 13403 38740 13415 38743
rect 14016 38740 14044 38839
rect 15562 38836 15568 38888
rect 15620 38836 15626 38888
rect 18598 38836 18604 38888
rect 18656 38876 18662 38888
rect 19429 38879 19487 38885
rect 18656 38848 19380 38876
rect 18656 38836 18662 38848
rect 17310 38768 17316 38820
rect 17368 38808 17374 38820
rect 17681 38811 17739 38817
rect 17681 38808 17693 38811
rect 17368 38780 17693 38808
rect 17368 38768 17374 38780
rect 17681 38777 17693 38780
rect 17727 38777 17739 38811
rect 19352 38808 19380 38848
rect 19429 38845 19441 38879
rect 19475 38876 19487 38879
rect 19518 38876 19524 38888
rect 19475 38848 19524 38876
rect 19475 38845 19487 38848
rect 19429 38839 19487 38845
rect 19518 38836 19524 38848
rect 19576 38836 19582 38888
rect 19610 38836 19616 38888
rect 19668 38876 19674 38888
rect 19981 38879 20039 38885
rect 19981 38876 19993 38879
rect 19668 38848 19993 38876
rect 19668 38836 19674 38848
rect 19981 38845 19993 38848
rect 20027 38845 20039 38879
rect 19981 38839 20039 38845
rect 20088 38808 20116 38916
rect 20993 38913 21005 38916
rect 21039 38944 21051 38947
rect 21358 38944 21364 38956
rect 21039 38916 21364 38944
rect 21039 38913 21051 38916
rect 20993 38907 21051 38913
rect 21358 38904 21364 38916
rect 21416 38904 21422 38956
rect 21836 38944 21864 39052
rect 22066 39052 23489 39080
rect 22066 39024 22094 39052
rect 23477 39049 23489 39052
rect 23523 39049 23535 39083
rect 23477 39043 23535 39049
rect 22002 38972 22008 39024
rect 22060 38984 22094 39024
rect 22465 39015 22523 39021
rect 22060 38972 22066 38984
rect 22465 38981 22477 39015
rect 22511 39012 22523 39015
rect 22646 39012 22652 39024
rect 22511 38984 22652 39012
rect 22511 38981 22523 38984
rect 22465 38975 22523 38981
rect 22646 38972 22652 38984
rect 22704 38972 22710 39024
rect 24302 38972 24308 39024
rect 24360 38972 24366 39024
rect 24949 39015 25007 39021
rect 24949 38981 24961 39015
rect 24995 39012 25007 39015
rect 25038 39012 25044 39024
rect 24995 38984 25044 39012
rect 24995 38981 25007 38984
rect 24949 38975 25007 38981
rect 25038 38972 25044 38984
rect 25096 38972 25102 39024
rect 22094 38944 22100 38956
rect 21836 38916 22100 38944
rect 22094 38904 22100 38916
rect 22152 38904 22158 38956
rect 22373 38947 22431 38953
rect 22373 38913 22385 38947
rect 22419 38913 22431 38947
rect 22373 38907 22431 38913
rect 20162 38836 20168 38888
rect 20220 38876 20226 38888
rect 21545 38879 21603 38885
rect 21545 38876 21557 38879
rect 20220 38848 21557 38876
rect 20220 38836 20226 38848
rect 21545 38845 21557 38848
rect 21591 38845 21603 38879
rect 21545 38839 21603 38845
rect 21818 38836 21824 38888
rect 21876 38876 21882 38888
rect 22002 38876 22008 38888
rect 21876 38848 22008 38876
rect 21876 38836 21882 38848
rect 22002 38836 22008 38848
rect 22060 38836 22066 38888
rect 22388 38876 22416 38907
rect 22462 38876 22468 38888
rect 22388 38848 22468 38876
rect 22462 38836 22468 38848
rect 22520 38836 22526 38888
rect 22557 38879 22615 38885
rect 22557 38845 22569 38879
rect 22603 38845 22615 38879
rect 22557 38839 22615 38845
rect 25225 38879 25283 38885
rect 25225 38845 25237 38879
rect 25271 38845 25283 38879
rect 25225 38839 25283 38845
rect 22572 38808 22600 38839
rect 19352 38780 20116 38808
rect 20456 38780 22600 38808
rect 17681 38771 17739 38777
rect 13403 38712 14044 38740
rect 13403 38709 13415 38712
rect 13357 38703 13415 38709
rect 14918 38700 14924 38752
rect 14976 38740 14982 38752
rect 15197 38743 15255 38749
rect 15197 38740 15209 38743
rect 14976 38712 15209 38740
rect 14976 38700 14982 38712
rect 15197 38709 15209 38712
rect 15243 38740 15255 38743
rect 15286 38740 15292 38752
rect 15243 38712 15292 38740
rect 15243 38709 15255 38712
rect 15197 38703 15255 38709
rect 15286 38700 15292 38712
rect 15344 38700 15350 38752
rect 16209 38743 16267 38749
rect 16209 38709 16221 38743
rect 16255 38740 16267 38743
rect 17402 38740 17408 38752
rect 16255 38712 17408 38740
rect 16255 38709 16267 38712
rect 16209 38703 16267 38709
rect 17402 38700 17408 38712
rect 17460 38700 17466 38752
rect 18966 38700 18972 38752
rect 19024 38740 19030 38752
rect 19165 38743 19223 38749
rect 19165 38740 19177 38743
rect 19024 38712 19177 38740
rect 19024 38700 19030 38712
rect 19165 38709 19177 38712
rect 19211 38740 19223 38743
rect 20456 38740 20484 38780
rect 23382 38768 23388 38820
rect 23440 38808 23446 38820
rect 23440 38780 23612 38808
rect 23440 38768 23446 38780
rect 19211 38712 20484 38740
rect 19211 38709 19223 38712
rect 19165 38703 19223 38709
rect 20530 38700 20536 38752
rect 20588 38740 20594 38752
rect 20625 38743 20683 38749
rect 20625 38740 20637 38743
rect 20588 38712 20637 38740
rect 20588 38700 20594 38712
rect 20625 38709 20637 38712
rect 20671 38709 20683 38743
rect 20625 38703 20683 38709
rect 22002 38700 22008 38752
rect 22060 38700 22066 38752
rect 22094 38700 22100 38752
rect 22152 38740 22158 38752
rect 22370 38740 22376 38752
rect 22152 38712 22376 38740
rect 22152 38700 22158 38712
rect 22370 38700 22376 38712
rect 22428 38740 22434 38752
rect 23017 38743 23075 38749
rect 23017 38740 23029 38743
rect 22428 38712 23029 38740
rect 22428 38700 22434 38712
rect 23017 38709 23029 38712
rect 23063 38709 23075 38743
rect 23584 38740 23612 38780
rect 25240 38740 25268 38839
rect 23584 38712 25268 38740
rect 23017 38703 23075 38709
rect 1104 38650 25852 38672
rect 1104 38598 2950 38650
rect 3002 38598 3014 38650
rect 3066 38598 3078 38650
rect 3130 38598 3142 38650
rect 3194 38598 3206 38650
rect 3258 38598 12950 38650
rect 13002 38598 13014 38650
rect 13066 38598 13078 38650
rect 13130 38598 13142 38650
rect 13194 38598 13206 38650
rect 13258 38598 22950 38650
rect 23002 38598 23014 38650
rect 23066 38598 23078 38650
rect 23130 38598 23142 38650
rect 23194 38598 23206 38650
rect 23258 38598 25852 38650
rect 1104 38576 25852 38598
rect 4893 38539 4951 38545
rect 4893 38505 4905 38539
rect 4939 38536 4951 38539
rect 6914 38536 6920 38548
rect 4939 38508 6920 38536
rect 4939 38505 4951 38508
rect 4893 38499 4951 38505
rect 6914 38496 6920 38508
rect 6972 38496 6978 38548
rect 8294 38496 8300 38548
rect 8352 38536 8358 38548
rect 8573 38539 8631 38545
rect 8573 38536 8585 38539
rect 8352 38508 8585 38536
rect 8352 38496 8358 38508
rect 8573 38505 8585 38508
rect 8619 38505 8631 38539
rect 8573 38499 8631 38505
rect 9306 38496 9312 38548
rect 9364 38536 9370 38548
rect 9493 38539 9551 38545
rect 9493 38536 9505 38539
rect 9364 38508 9505 38536
rect 9364 38496 9370 38508
rect 9493 38505 9505 38508
rect 9539 38505 9551 38539
rect 11330 38536 11336 38548
rect 9493 38499 9551 38505
rect 9600 38508 11336 38536
rect 8110 38428 8116 38480
rect 8168 38468 8174 38480
rect 9600 38468 9628 38508
rect 11330 38496 11336 38508
rect 11388 38496 11394 38548
rect 11425 38539 11483 38545
rect 11425 38505 11437 38539
rect 11471 38536 11483 38539
rect 12066 38536 12072 38548
rect 11471 38508 12072 38536
rect 11471 38505 11483 38508
rect 11425 38499 11483 38505
rect 12066 38496 12072 38508
rect 12124 38496 12130 38548
rect 12710 38496 12716 38548
rect 12768 38536 12774 38548
rect 12986 38536 12992 38548
rect 12768 38508 12992 38536
rect 12768 38496 12774 38508
rect 12986 38496 12992 38508
rect 13044 38496 13050 38548
rect 16393 38539 16451 38545
rect 16393 38505 16405 38539
rect 16439 38536 16451 38539
rect 16574 38536 16580 38548
rect 16439 38508 16580 38536
rect 16439 38505 16451 38508
rect 16393 38499 16451 38505
rect 16574 38496 16580 38508
rect 16632 38496 16638 38548
rect 16758 38496 16764 38548
rect 16816 38536 16822 38548
rect 16853 38539 16911 38545
rect 16853 38536 16865 38539
rect 16816 38508 16865 38536
rect 16816 38496 16822 38508
rect 16853 38505 16865 38508
rect 16899 38505 16911 38539
rect 16853 38499 16911 38505
rect 20165 38539 20223 38545
rect 20165 38505 20177 38539
rect 20211 38536 20223 38539
rect 22738 38536 22744 38548
rect 20211 38508 22744 38536
rect 20211 38505 20223 38508
rect 20165 38499 20223 38505
rect 22738 38496 22744 38508
rect 22796 38496 22802 38548
rect 25958 38536 25964 38548
rect 23124 38508 25964 38536
rect 11977 38471 12035 38477
rect 11977 38468 11989 38471
rect 8168 38440 9628 38468
rect 9784 38440 11989 38468
rect 8168 38428 8174 38440
rect 5902 38360 5908 38412
rect 5960 38400 5966 38412
rect 6641 38403 6699 38409
rect 6641 38400 6653 38403
rect 5960 38372 6653 38400
rect 5960 38360 5966 38372
rect 6641 38369 6653 38372
rect 6687 38369 6699 38403
rect 6641 38363 6699 38369
rect 7834 38360 7840 38412
rect 7892 38400 7898 38412
rect 8021 38403 8079 38409
rect 8021 38400 8033 38403
rect 7892 38372 8033 38400
rect 7892 38360 7898 38372
rect 8021 38369 8033 38372
rect 8067 38400 8079 38403
rect 8067 38372 8892 38400
rect 8067 38369 8079 38372
rect 8021 38363 8079 38369
rect 7190 38292 7196 38344
rect 7248 38332 7254 38344
rect 7561 38335 7619 38341
rect 7561 38332 7573 38335
rect 7248 38304 7573 38332
rect 7248 38292 7254 38304
rect 7561 38301 7573 38304
rect 7607 38332 7619 38335
rect 8110 38332 8116 38344
rect 7607 38304 8116 38332
rect 7607 38301 7619 38304
rect 7561 38295 7619 38301
rect 8110 38292 8116 38304
rect 8168 38292 8174 38344
rect 8205 38335 8263 38341
rect 8205 38301 8217 38335
rect 8251 38332 8263 38335
rect 8570 38332 8576 38344
rect 8251 38304 8576 38332
rect 8251 38301 8263 38304
rect 8205 38295 8263 38301
rect 8570 38292 8576 38304
rect 8628 38292 8634 38344
rect 8864 38332 8892 38372
rect 9582 38360 9588 38412
rect 9640 38400 9646 38412
rect 9784 38400 9812 38440
rect 11977 38437 11989 38440
rect 12023 38437 12035 38471
rect 22922 38468 22928 38480
rect 11977 38431 12035 38437
rect 12084 38440 17448 38468
rect 9640 38372 9812 38400
rect 9640 38360 9646 38372
rect 9858 38360 9864 38412
rect 9916 38400 9922 38412
rect 9953 38403 10011 38409
rect 9953 38400 9965 38403
rect 9916 38372 9965 38400
rect 9916 38360 9922 38372
rect 9953 38369 9965 38372
rect 9999 38369 10011 38403
rect 9953 38363 10011 38369
rect 10134 38360 10140 38412
rect 10192 38360 10198 38412
rect 10873 38403 10931 38409
rect 10873 38369 10885 38403
rect 10919 38400 10931 38403
rect 11514 38400 11520 38412
rect 10919 38372 11520 38400
rect 10919 38369 10931 38372
rect 10873 38363 10931 38369
rect 11514 38360 11520 38372
rect 11572 38400 11578 38412
rect 12084 38400 12112 38440
rect 12529 38403 12587 38409
rect 12529 38400 12541 38403
rect 11572 38372 12112 38400
rect 12406 38372 12541 38400
rect 11572 38360 11578 38372
rect 8864 38304 10272 38332
rect 5934 38236 6040 38264
rect 6012 38196 6040 38236
rect 6086 38224 6092 38276
rect 6144 38264 6150 38276
rect 6365 38267 6423 38273
rect 6365 38264 6377 38267
rect 6144 38236 6377 38264
rect 6144 38224 6150 38236
rect 6365 38233 6377 38236
rect 6411 38264 6423 38267
rect 10134 38264 10140 38276
rect 6411 38236 10140 38264
rect 6411 38233 6423 38236
rect 6365 38227 6423 38233
rect 10134 38224 10140 38236
rect 10192 38224 10198 38276
rect 10244 38264 10272 38304
rect 11054 38292 11060 38344
rect 11112 38292 11118 38344
rect 12406 38332 12434 38372
rect 12529 38369 12541 38372
rect 12575 38369 12587 38403
rect 12529 38363 12587 38369
rect 15105 38403 15163 38409
rect 15105 38369 15117 38403
rect 15151 38400 15163 38403
rect 15562 38400 15568 38412
rect 15151 38372 15568 38400
rect 15151 38369 15163 38372
rect 15105 38363 15163 38369
rect 15562 38360 15568 38372
rect 15620 38360 15626 38412
rect 15838 38360 15844 38412
rect 15896 38360 15902 38412
rect 17420 38409 17448 38440
rect 18432 38440 22928 38468
rect 17405 38403 17463 38409
rect 17405 38369 17417 38403
rect 17451 38369 17463 38403
rect 17405 38363 17463 38369
rect 11164 38304 12434 38332
rect 14829 38335 14887 38341
rect 11164 38264 11192 38304
rect 14829 38301 14841 38335
rect 14875 38332 14887 38335
rect 18432 38332 18460 38440
rect 22922 38428 22928 38440
rect 22980 38468 22986 38480
rect 23124 38468 23152 38508
rect 25958 38496 25964 38508
rect 26016 38496 26022 38548
rect 25130 38468 25136 38480
rect 22980 38440 23152 38468
rect 23216 38440 25136 38468
rect 22980 38428 22986 38440
rect 19613 38403 19671 38409
rect 19613 38369 19625 38403
rect 19659 38400 19671 38403
rect 19978 38400 19984 38412
rect 19659 38372 19984 38400
rect 19659 38369 19671 38372
rect 19613 38363 19671 38369
rect 19978 38360 19984 38372
rect 20036 38360 20042 38412
rect 22094 38360 22100 38412
rect 22152 38400 22158 38412
rect 22646 38400 22652 38412
rect 22152 38372 22652 38400
rect 22152 38360 22158 38372
rect 22646 38360 22652 38372
rect 22704 38360 22710 38412
rect 23216 38409 23244 38440
rect 25130 38428 25136 38440
rect 25188 38428 25194 38480
rect 23201 38403 23259 38409
rect 23201 38369 23213 38403
rect 23247 38369 23259 38403
rect 23201 38363 23259 38369
rect 23290 38360 23296 38412
rect 23348 38360 23354 38412
rect 14875 38304 18460 38332
rect 14875 38301 14887 38304
rect 14829 38295 14887 38301
rect 19426 38292 19432 38344
rect 19484 38332 19490 38344
rect 19705 38335 19763 38341
rect 19705 38332 19717 38335
rect 19484 38304 19717 38332
rect 19484 38292 19490 38304
rect 19705 38301 19717 38304
rect 19751 38301 19763 38335
rect 19705 38295 19763 38301
rect 22278 38292 22284 38344
rect 22336 38332 22342 38344
rect 23382 38332 23388 38344
rect 22336 38304 23388 38332
rect 22336 38292 22342 38304
rect 23382 38292 23388 38304
rect 23440 38292 23446 38344
rect 24857 38335 24915 38341
rect 24857 38301 24869 38335
rect 24903 38332 24915 38335
rect 25317 38335 25375 38341
rect 25317 38332 25329 38335
rect 24903 38304 25329 38332
rect 24903 38301 24915 38304
rect 24857 38295 24915 38301
rect 25317 38301 25329 38304
rect 25363 38332 25375 38335
rect 25406 38332 25412 38344
rect 25363 38304 25412 38332
rect 25363 38301 25375 38304
rect 25317 38295 25375 38301
rect 25406 38292 25412 38304
rect 25464 38292 25470 38344
rect 10244 38236 11192 38264
rect 11238 38224 11244 38276
rect 11296 38264 11302 38276
rect 12066 38264 12072 38276
rect 11296 38236 12072 38264
rect 11296 38224 11302 38236
rect 12066 38224 12072 38236
rect 12124 38264 12130 38276
rect 14093 38267 14151 38273
rect 14093 38264 14105 38267
rect 12124 38236 14105 38264
rect 12124 38224 12130 38236
rect 14093 38233 14105 38236
rect 14139 38264 14151 38267
rect 14921 38267 14979 38273
rect 14921 38264 14933 38267
rect 14139 38236 14933 38264
rect 14139 38233 14151 38236
rect 14093 38227 14151 38233
rect 14921 38233 14933 38236
rect 14967 38233 14979 38267
rect 14921 38227 14979 38233
rect 15286 38224 15292 38276
rect 15344 38264 15350 38276
rect 15933 38267 15991 38273
rect 15933 38264 15945 38267
rect 15344 38236 15945 38264
rect 15344 38224 15350 38236
rect 15933 38233 15945 38236
rect 15979 38233 15991 38267
rect 15933 38227 15991 38233
rect 17313 38267 17371 38273
rect 17313 38233 17325 38267
rect 17359 38264 17371 38267
rect 17494 38264 17500 38276
rect 17359 38236 17500 38264
rect 17359 38233 17371 38236
rect 17313 38227 17371 38233
rect 17494 38224 17500 38236
rect 17552 38224 17558 38276
rect 21453 38267 21511 38273
rect 21453 38233 21465 38267
rect 21499 38233 21511 38267
rect 21453 38227 21511 38233
rect 6546 38196 6552 38208
rect 6012 38168 6552 38196
rect 6546 38156 6552 38168
rect 6604 38196 6610 38208
rect 6917 38199 6975 38205
rect 6917 38196 6929 38199
rect 6604 38168 6929 38196
rect 6604 38156 6610 38168
rect 6917 38165 6929 38168
rect 6963 38196 6975 38199
rect 8294 38196 8300 38208
rect 6963 38168 8300 38196
rect 6963 38165 6975 38168
rect 6917 38159 6975 38165
rect 8294 38156 8300 38168
rect 8352 38156 8358 38208
rect 9858 38156 9864 38208
rect 9916 38156 9922 38208
rect 10962 38156 10968 38208
rect 11020 38156 11026 38208
rect 12250 38156 12256 38208
rect 12308 38196 12314 38208
rect 12345 38199 12403 38205
rect 12345 38196 12357 38199
rect 12308 38168 12357 38196
rect 12308 38156 12314 38168
rect 12345 38165 12357 38168
rect 12391 38165 12403 38199
rect 12345 38159 12403 38165
rect 12437 38199 12495 38205
rect 12437 38165 12449 38199
rect 12483 38196 12495 38199
rect 12618 38196 12624 38208
rect 12483 38168 12624 38196
rect 12483 38165 12495 38168
rect 12437 38159 12495 38165
rect 12618 38156 12624 38168
rect 12676 38156 12682 38208
rect 14458 38156 14464 38208
rect 14516 38156 14522 38208
rect 16025 38199 16083 38205
rect 16025 38165 16037 38199
rect 16071 38196 16083 38199
rect 16114 38196 16120 38208
rect 16071 38168 16120 38196
rect 16071 38165 16083 38168
rect 16025 38159 16083 38165
rect 16114 38156 16120 38168
rect 16172 38156 16178 38208
rect 16482 38156 16488 38208
rect 16540 38196 16546 38208
rect 17221 38199 17279 38205
rect 17221 38196 17233 38199
rect 16540 38168 17233 38196
rect 16540 38156 16546 38168
rect 17221 38165 17233 38168
rect 17267 38165 17279 38199
rect 17221 38159 17279 38165
rect 18598 38156 18604 38208
rect 18656 38196 18662 38208
rect 18877 38199 18935 38205
rect 18877 38196 18889 38199
rect 18656 38168 18889 38196
rect 18656 38156 18662 38168
rect 18877 38165 18889 38168
rect 18923 38165 18935 38199
rect 18877 38159 18935 38165
rect 19334 38156 19340 38208
rect 19392 38196 19398 38208
rect 19797 38199 19855 38205
rect 19797 38196 19809 38199
rect 19392 38168 19809 38196
rect 19392 38156 19398 38168
rect 19797 38165 19809 38168
rect 19843 38165 19855 38199
rect 19797 38159 19855 38165
rect 20714 38156 20720 38208
rect 20772 38196 20778 38208
rect 21082 38196 21088 38208
rect 20772 38168 21088 38196
rect 20772 38156 20778 38168
rect 21082 38156 21088 38168
rect 21140 38196 21146 38208
rect 21468 38196 21496 38227
rect 22462 38224 22468 38276
rect 22520 38264 22526 38276
rect 22520 38236 25176 38264
rect 22520 38224 22526 38236
rect 21140 38168 21496 38196
rect 21140 38156 21146 38168
rect 21542 38156 21548 38208
rect 21600 38196 21606 38208
rect 22649 38199 22707 38205
rect 22649 38196 22661 38199
rect 21600 38168 22661 38196
rect 21600 38156 21606 38168
rect 22649 38165 22661 38168
rect 22695 38165 22707 38199
rect 22649 38159 22707 38165
rect 22830 38156 22836 38208
rect 22888 38196 22894 38208
rect 23385 38199 23443 38205
rect 23385 38196 23397 38199
rect 22888 38168 23397 38196
rect 22888 38156 22894 38168
rect 23385 38165 23397 38168
rect 23431 38165 23443 38199
rect 23385 38159 23443 38165
rect 23750 38156 23756 38208
rect 23808 38156 23814 38208
rect 24486 38156 24492 38208
rect 24544 38156 24550 38208
rect 24673 38199 24731 38205
rect 24673 38165 24685 38199
rect 24719 38196 24731 38199
rect 24762 38196 24768 38208
rect 24719 38168 24768 38196
rect 24719 38165 24731 38168
rect 24673 38159 24731 38165
rect 24762 38156 24768 38168
rect 24820 38156 24826 38208
rect 25148 38205 25176 38236
rect 25133 38199 25191 38205
rect 25133 38165 25145 38199
rect 25179 38165 25191 38199
rect 25133 38159 25191 38165
rect 1104 38106 25852 38128
rect 1104 38054 7950 38106
rect 8002 38054 8014 38106
rect 8066 38054 8078 38106
rect 8130 38054 8142 38106
rect 8194 38054 8206 38106
rect 8258 38054 17950 38106
rect 18002 38054 18014 38106
rect 18066 38054 18078 38106
rect 18130 38054 18142 38106
rect 18194 38054 18206 38106
rect 18258 38054 25852 38106
rect 1104 38032 25852 38054
rect 10870 37952 10876 38004
rect 10928 37952 10934 38004
rect 12158 37952 12164 38004
rect 12216 37992 12222 38004
rect 12253 37995 12311 38001
rect 12253 37992 12265 37995
rect 12216 37964 12265 37992
rect 12216 37952 12222 37964
rect 12253 37961 12265 37964
rect 12299 37961 12311 37995
rect 12253 37955 12311 37961
rect 12894 37952 12900 38004
rect 12952 37992 12958 38004
rect 13173 37995 13231 38001
rect 13173 37992 13185 37995
rect 12952 37964 13185 37992
rect 12952 37952 12958 37964
rect 13173 37961 13185 37964
rect 13219 37961 13231 37995
rect 13173 37955 13231 37961
rect 13633 37995 13691 38001
rect 13633 37961 13645 37995
rect 13679 37992 13691 37995
rect 15194 37992 15200 38004
rect 13679 37964 15200 37992
rect 13679 37961 13691 37964
rect 13633 37955 13691 37961
rect 15194 37952 15200 37964
rect 15252 37952 15258 38004
rect 15378 37952 15384 38004
rect 15436 37952 15442 38004
rect 16114 37952 16120 38004
rect 16172 37952 16178 38004
rect 19518 37992 19524 38004
rect 17052 37964 19524 37992
rect 9306 37884 9312 37936
rect 9364 37924 9370 37936
rect 9401 37927 9459 37933
rect 9401 37924 9413 37927
rect 9364 37896 9413 37924
rect 9364 37884 9370 37896
rect 9401 37893 9413 37896
rect 9447 37924 9459 37927
rect 10410 37924 10416 37936
rect 9447 37896 10416 37924
rect 9447 37893 9459 37896
rect 9401 37887 9459 37893
rect 10410 37884 10416 37896
rect 10468 37884 10474 37936
rect 10686 37884 10692 37936
rect 10744 37924 10750 37936
rect 15562 37924 15568 37936
rect 10744 37896 15568 37924
rect 10744 37884 10750 37896
rect 15562 37884 15568 37896
rect 15620 37884 15626 37936
rect 8294 37816 8300 37868
rect 8352 37816 8358 37868
rect 9674 37816 9680 37868
rect 9732 37816 9738 37868
rect 10502 37816 10508 37868
rect 10560 37816 10566 37868
rect 13265 37859 13323 37865
rect 10888 37828 13216 37856
rect 7374 37748 7380 37800
rect 7432 37788 7438 37800
rect 7653 37791 7711 37797
rect 7653 37788 7665 37791
rect 7432 37760 7665 37788
rect 7432 37748 7438 37760
rect 7653 37757 7665 37760
rect 7699 37757 7711 37791
rect 7653 37751 7711 37757
rect 9398 37748 9404 37800
rect 9456 37788 9462 37800
rect 10229 37791 10287 37797
rect 10229 37788 10241 37791
rect 9456 37760 10241 37788
rect 9456 37748 9462 37760
rect 10229 37757 10241 37760
rect 10275 37757 10287 37791
rect 10229 37751 10287 37757
rect 10244 37720 10272 37751
rect 10410 37748 10416 37800
rect 10468 37748 10474 37800
rect 10888 37732 10916 37828
rect 12986 37748 12992 37800
rect 13044 37748 13050 37800
rect 13188 37788 13216 37828
rect 13265 37825 13277 37859
rect 13311 37856 13323 37859
rect 14093 37859 14151 37865
rect 14093 37856 14105 37859
rect 13311 37828 14105 37856
rect 13311 37825 13323 37828
rect 13265 37819 13323 37825
rect 14093 37825 14105 37828
rect 14139 37825 14151 37859
rect 14093 37819 14151 37825
rect 15194 37816 15200 37868
rect 15252 37856 15258 37868
rect 17052 37865 17080 37964
rect 19518 37952 19524 37964
rect 19576 37952 19582 38004
rect 22005 37995 22063 38001
rect 22005 37961 22017 37995
rect 22051 37992 22063 37995
rect 22186 37992 22192 38004
rect 22051 37964 22192 37992
rect 22051 37961 22063 37964
rect 22005 37955 22063 37961
rect 22186 37952 22192 37964
rect 22244 37952 22250 38004
rect 22370 37952 22376 38004
rect 22428 37952 22434 38004
rect 18598 37924 18604 37936
rect 18538 37896 18604 37924
rect 18598 37884 18604 37896
rect 18656 37884 18662 37936
rect 20625 37927 20683 37933
rect 20625 37893 20637 37927
rect 20671 37924 20683 37927
rect 22094 37924 22100 37936
rect 20671 37896 22100 37924
rect 20671 37893 20683 37896
rect 20625 37887 20683 37893
rect 22094 37884 22100 37896
rect 22152 37884 22158 37936
rect 22465 37927 22523 37933
rect 22465 37924 22477 37927
rect 22296 37896 22477 37924
rect 15289 37859 15347 37865
rect 15289 37856 15301 37859
rect 15252 37828 15301 37856
rect 15252 37816 15258 37828
rect 15289 37825 15301 37828
rect 15335 37856 15347 37859
rect 16669 37859 16727 37865
rect 16669 37856 16681 37859
rect 15335 37828 16681 37856
rect 15335 37825 15347 37828
rect 15289 37819 15347 37825
rect 16669 37825 16681 37828
rect 16715 37825 16727 37859
rect 16669 37819 16727 37825
rect 17037 37859 17095 37865
rect 17037 37825 17049 37859
rect 17083 37825 17095 37859
rect 19150 37856 19156 37868
rect 17037 37819 17095 37825
rect 18708 37828 19156 37856
rect 13188 37760 13308 37788
rect 10870 37720 10876 37732
rect 10244 37692 10876 37720
rect 10870 37680 10876 37692
rect 10928 37680 10934 37732
rect 12802 37720 12808 37732
rect 11164 37692 12808 37720
rect 7466 37612 7472 37664
rect 7524 37652 7530 37664
rect 10962 37652 10968 37664
rect 7524 37624 10968 37652
rect 7524 37612 7530 37624
rect 10962 37612 10968 37624
rect 11020 37652 11026 37664
rect 11164 37661 11192 37692
rect 12802 37680 12808 37692
rect 12860 37680 12866 37732
rect 13280 37720 13308 37760
rect 13354 37748 13360 37800
rect 13412 37788 13418 37800
rect 13722 37788 13728 37800
rect 13412 37760 13728 37788
rect 13412 37748 13418 37760
rect 13722 37748 13728 37760
rect 13780 37788 13786 37800
rect 15473 37791 15531 37797
rect 15473 37788 15485 37791
rect 13780 37760 15485 37788
rect 13780 37748 13786 37760
rect 15473 37757 15485 37760
rect 15519 37757 15531 37791
rect 15473 37751 15531 37757
rect 15654 37720 15660 37732
rect 13280 37692 15660 37720
rect 15654 37680 15660 37692
rect 15712 37680 15718 37732
rect 11149 37655 11207 37661
rect 11149 37652 11161 37655
rect 11020 37624 11161 37652
rect 11020 37612 11026 37624
rect 11149 37621 11161 37624
rect 11195 37621 11207 37655
rect 11149 37615 11207 37621
rect 11514 37612 11520 37664
rect 11572 37652 11578 37664
rect 12342 37652 12348 37664
rect 11572 37624 12348 37652
rect 11572 37612 11578 37624
rect 12342 37612 12348 37624
rect 12400 37612 12406 37664
rect 14918 37612 14924 37664
rect 14976 37612 14982 37664
rect 16684 37652 16712 37819
rect 17310 37748 17316 37800
rect 17368 37748 17374 37800
rect 18046 37748 18052 37800
rect 18104 37788 18110 37800
rect 18708 37788 18736 37828
rect 19150 37816 19156 37828
rect 19208 37816 19214 37868
rect 19886 37816 19892 37868
rect 19944 37856 19950 37868
rect 20533 37859 20591 37865
rect 20533 37856 20545 37859
rect 19944 37828 20545 37856
rect 19944 37816 19950 37828
rect 20533 37825 20545 37828
rect 20579 37825 20591 37859
rect 20533 37819 20591 37825
rect 21542 37816 21548 37868
rect 21600 37856 21606 37868
rect 22296 37856 22324 37896
rect 22465 37893 22477 37896
rect 22511 37893 22523 37927
rect 23382 37924 23388 37936
rect 22465 37887 22523 37893
rect 23216 37896 23388 37924
rect 23216 37865 23244 37896
rect 23382 37884 23388 37896
rect 23440 37884 23446 37936
rect 21600 37828 22324 37856
rect 23201 37859 23259 37865
rect 21600 37816 21606 37828
rect 23201 37825 23213 37859
rect 23247 37825 23259 37859
rect 23201 37819 23259 37825
rect 18104 37760 18736 37788
rect 18104 37748 18110 37760
rect 18782 37748 18788 37800
rect 18840 37748 18846 37800
rect 19426 37748 19432 37800
rect 19484 37748 19490 37800
rect 20441 37791 20499 37797
rect 20441 37757 20453 37791
rect 20487 37757 20499 37791
rect 20441 37751 20499 37757
rect 19702 37720 19708 37732
rect 18340 37692 19708 37720
rect 18340 37652 18368 37692
rect 19702 37680 19708 37692
rect 19760 37680 19766 37732
rect 20456 37720 20484 37751
rect 20806 37748 20812 37800
rect 20864 37788 20870 37800
rect 22649 37791 22707 37797
rect 22649 37788 22661 37791
rect 20864 37760 22661 37788
rect 20864 37748 20870 37760
rect 22649 37757 22661 37760
rect 22695 37788 22707 37791
rect 23842 37788 23848 37800
rect 22695 37760 23848 37788
rect 22695 37757 22707 37760
rect 22649 37751 22707 37757
rect 23842 37748 23848 37760
rect 23900 37788 23906 37800
rect 24118 37788 24124 37800
rect 23900 37760 24124 37788
rect 23900 37748 23906 37760
rect 24118 37748 24124 37760
rect 24176 37748 24182 37800
rect 20622 37720 20628 37732
rect 20456 37692 20628 37720
rect 20622 37680 20628 37692
rect 20680 37680 20686 37732
rect 20993 37723 21051 37729
rect 20993 37689 21005 37723
rect 21039 37720 21051 37723
rect 22462 37720 22468 37732
rect 21039 37692 22468 37720
rect 21039 37689 21051 37692
rect 20993 37683 21051 37689
rect 22462 37680 22468 37692
rect 22520 37680 22526 37732
rect 24486 37680 24492 37732
rect 24544 37720 24550 37732
rect 24596 37720 24624 37842
rect 25409 37723 25467 37729
rect 25409 37720 25421 37723
rect 24544 37692 25421 37720
rect 24544 37680 24550 37692
rect 25409 37689 25421 37692
rect 25455 37689 25467 37723
rect 25409 37683 25467 37689
rect 16684 37624 18368 37652
rect 18414 37612 18420 37664
rect 18472 37652 18478 37664
rect 19061 37655 19119 37661
rect 19061 37652 19073 37655
rect 18472 37624 19073 37652
rect 18472 37612 18478 37624
rect 19061 37621 19073 37624
rect 19107 37621 19119 37655
rect 19061 37615 19119 37621
rect 19886 37612 19892 37664
rect 19944 37612 19950 37664
rect 22646 37612 22652 37664
rect 22704 37652 22710 37664
rect 22922 37652 22928 37664
rect 22704 37624 22928 37652
rect 22704 37612 22710 37624
rect 22922 37612 22928 37624
rect 22980 37612 22986 37664
rect 23474 37661 23480 37664
rect 23464 37655 23480 37661
rect 23464 37621 23476 37655
rect 23464 37615 23480 37621
rect 23474 37612 23480 37615
rect 23532 37612 23538 37664
rect 24949 37655 25007 37661
rect 24949 37621 24961 37655
rect 24995 37652 25007 37655
rect 25130 37652 25136 37664
rect 24995 37624 25136 37652
rect 24995 37621 25007 37624
rect 24949 37615 25007 37621
rect 25130 37612 25136 37624
rect 25188 37612 25194 37664
rect 25314 37612 25320 37664
rect 25372 37612 25378 37664
rect 1104 37562 25852 37584
rect 1104 37510 2950 37562
rect 3002 37510 3014 37562
rect 3066 37510 3078 37562
rect 3130 37510 3142 37562
rect 3194 37510 3206 37562
rect 3258 37510 12950 37562
rect 13002 37510 13014 37562
rect 13066 37510 13078 37562
rect 13130 37510 13142 37562
rect 13194 37510 13206 37562
rect 13258 37510 22950 37562
rect 23002 37510 23014 37562
rect 23066 37510 23078 37562
rect 23130 37510 23142 37562
rect 23194 37510 23206 37562
rect 23258 37510 25852 37562
rect 1104 37488 25852 37510
rect 5902 37408 5908 37460
rect 5960 37448 5966 37460
rect 7466 37448 7472 37460
rect 5960 37420 7472 37448
rect 5960 37408 5966 37420
rect 7466 37408 7472 37420
rect 7524 37408 7530 37460
rect 8294 37408 8300 37460
rect 8352 37448 8358 37460
rect 8941 37451 8999 37457
rect 8941 37448 8953 37451
rect 8352 37420 8953 37448
rect 8352 37408 8358 37420
rect 8941 37417 8953 37420
rect 8987 37417 8999 37451
rect 8941 37411 8999 37417
rect 8956 37380 8984 37411
rect 9122 37408 9128 37460
rect 9180 37448 9186 37460
rect 9309 37451 9367 37457
rect 9309 37448 9321 37451
rect 9180 37420 9321 37448
rect 9180 37408 9186 37420
rect 9309 37417 9321 37420
rect 9355 37448 9367 37451
rect 10410 37448 10416 37460
rect 9355 37420 10416 37448
rect 9355 37417 9367 37420
rect 9309 37411 9367 37417
rect 10410 37408 10416 37420
rect 10468 37408 10474 37460
rect 10778 37408 10784 37460
rect 10836 37448 10842 37460
rect 12618 37448 12624 37460
rect 10836 37420 12624 37448
rect 10836 37408 10842 37420
rect 12618 37408 12624 37420
rect 12676 37408 12682 37460
rect 12802 37408 12808 37460
rect 12860 37408 12866 37460
rect 20898 37448 20904 37460
rect 18340 37420 20904 37448
rect 9401 37383 9459 37389
rect 9401 37380 9413 37383
rect 8956 37352 9413 37380
rect 9401 37349 9413 37352
rect 9447 37349 9459 37383
rect 18046 37380 18052 37392
rect 9401 37343 9459 37349
rect 17696 37352 18052 37380
rect 5537 37315 5595 37321
rect 5537 37281 5549 37315
rect 5583 37312 5595 37315
rect 6914 37312 6920 37324
rect 5583 37284 6920 37312
rect 5583 37281 5595 37284
rect 5537 37275 5595 37281
rect 6914 37272 6920 37284
rect 6972 37272 6978 37324
rect 7190 37272 7196 37324
rect 7248 37312 7254 37324
rect 8297 37315 8355 37321
rect 8297 37312 8309 37315
rect 7248 37284 8309 37312
rect 7248 37272 7254 37284
rect 8297 37281 8309 37284
rect 8343 37281 8355 37315
rect 8297 37275 8355 37281
rect 10413 37315 10471 37321
rect 10413 37281 10425 37315
rect 10459 37312 10471 37315
rect 10778 37312 10784 37324
rect 10459 37284 10784 37312
rect 10459 37281 10471 37284
rect 10413 37275 10471 37281
rect 10778 37272 10784 37284
rect 10836 37272 10842 37324
rect 10870 37272 10876 37324
rect 10928 37272 10934 37324
rect 11422 37272 11428 37324
rect 11480 37312 11486 37324
rect 11885 37315 11943 37321
rect 11885 37312 11897 37315
rect 11480 37284 11897 37312
rect 11480 37272 11486 37284
rect 11885 37281 11897 37284
rect 11931 37281 11943 37315
rect 11885 37275 11943 37281
rect 12066 37272 12072 37324
rect 12124 37312 12130 37324
rect 12437 37315 12495 37321
rect 12437 37312 12449 37315
rect 12124 37284 12449 37312
rect 12124 37272 12130 37284
rect 12437 37281 12449 37284
rect 12483 37281 12495 37315
rect 12437 37275 12495 37281
rect 12618 37272 12624 37324
rect 12676 37312 12682 37324
rect 15565 37315 15623 37321
rect 15565 37312 15577 37315
rect 12676 37284 15577 37312
rect 12676 37272 12682 37284
rect 15565 37281 15577 37284
rect 15611 37312 15623 37315
rect 15838 37312 15844 37324
rect 15611 37284 15844 37312
rect 15611 37281 15623 37284
rect 15565 37275 15623 37281
rect 15838 37272 15844 37284
rect 15896 37272 15902 37324
rect 16669 37315 16727 37321
rect 16669 37281 16681 37315
rect 16715 37312 16727 37315
rect 17696 37312 17724 37352
rect 18046 37340 18052 37352
rect 18104 37340 18110 37392
rect 16715 37284 17724 37312
rect 16715 37281 16727 37284
rect 16669 37275 16727 37281
rect 17770 37272 17776 37324
rect 17828 37272 17834 37324
rect 18340 37321 18368 37420
rect 20898 37408 20904 37420
rect 20956 37408 20962 37460
rect 20990 37408 20996 37460
rect 21048 37448 21054 37460
rect 21048 37420 23796 37448
rect 21048 37408 21054 37420
rect 23768 37380 23796 37420
rect 23842 37408 23848 37460
rect 23900 37448 23906 37460
rect 25498 37448 25504 37460
rect 23900 37420 25504 37448
rect 23900 37408 23906 37420
rect 25498 37408 25504 37420
rect 25556 37408 25562 37460
rect 25682 37380 25688 37392
rect 23768 37352 25688 37380
rect 25682 37340 25688 37352
rect 25740 37340 25746 37392
rect 18325 37315 18383 37321
rect 18325 37281 18337 37315
rect 18371 37281 18383 37315
rect 18325 37275 18383 37281
rect 18414 37272 18420 37324
rect 18472 37272 18478 37324
rect 21453 37315 21511 37321
rect 21453 37281 21465 37315
rect 21499 37312 21511 37315
rect 22278 37312 22284 37324
rect 21499 37284 22284 37312
rect 21499 37281 21511 37284
rect 21453 37275 21511 37281
rect 22278 37272 22284 37284
rect 22336 37272 22342 37324
rect 23569 37315 23627 37321
rect 23569 37281 23581 37315
rect 23615 37312 23627 37315
rect 24394 37312 24400 37324
rect 23615 37284 24400 37312
rect 23615 37281 23627 37284
rect 23569 37275 23627 37281
rect 5258 37204 5264 37256
rect 5316 37204 5322 37256
rect 8113 37247 8171 37253
rect 8113 37213 8125 37247
rect 8159 37244 8171 37247
rect 9950 37244 9956 37256
rect 8159 37216 9956 37244
rect 8159 37213 8171 37216
rect 8113 37207 8171 37213
rect 9950 37204 9956 37216
rect 10008 37204 10014 37256
rect 10042 37204 10048 37256
rect 10100 37244 10106 37256
rect 10229 37247 10287 37253
rect 10229 37244 10241 37247
rect 10100 37216 10241 37244
rect 10100 37204 10106 37216
rect 10229 37213 10241 37216
rect 10275 37213 10287 37247
rect 10229 37207 10287 37213
rect 11701 37247 11759 37253
rect 11701 37213 11713 37247
rect 11747 37244 11759 37247
rect 15286 37244 15292 37256
rect 11747 37216 15292 37244
rect 11747 37213 11759 37216
rect 11701 37207 11759 37213
rect 15286 37204 15292 37216
rect 15344 37204 15350 37256
rect 16853 37247 16911 37253
rect 16853 37213 16865 37247
rect 16899 37244 16911 37247
rect 19426 37244 19432 37256
rect 16899 37216 19432 37244
rect 16899 37213 16911 37216
rect 16853 37207 16911 37213
rect 19426 37204 19432 37216
rect 19484 37204 19490 37256
rect 19518 37204 19524 37256
rect 19576 37204 19582 37256
rect 23584 37244 23612 37275
rect 24394 37272 24400 37284
rect 24452 37312 24458 37324
rect 24673 37315 24731 37321
rect 24673 37312 24685 37315
rect 24452 37284 24685 37312
rect 24452 37272 24458 37284
rect 24673 37281 24685 37284
rect 24719 37281 24731 37315
rect 24673 37275 24731 37281
rect 22862 37216 23612 37244
rect 24029 37247 24087 37253
rect 24029 37213 24041 37247
rect 24075 37244 24087 37247
rect 24075 37216 24532 37244
rect 24075 37213 24087 37216
rect 24029 37207 24087 37213
rect 6546 37136 6552 37188
rect 6604 37136 6610 37188
rect 7098 37136 7104 37188
rect 7156 37176 7162 37188
rect 7285 37179 7343 37185
rect 7285 37176 7297 37179
rect 7156 37148 7297 37176
rect 7156 37136 7162 37148
rect 7285 37145 7297 37148
rect 7331 37145 7343 37179
rect 7285 37139 7343 37145
rect 8205 37179 8263 37185
rect 8205 37145 8217 37179
rect 8251 37176 8263 37179
rect 10137 37179 10195 37185
rect 8251 37148 9812 37176
rect 8251 37145 8263 37148
rect 8205 37139 8263 37145
rect 7742 37068 7748 37120
rect 7800 37068 7806 37120
rect 9784 37117 9812 37148
rect 10137 37145 10149 37179
rect 10183 37176 10195 37179
rect 11238 37176 11244 37188
rect 10183 37148 11244 37176
rect 10183 37145 10195 37148
rect 10137 37139 10195 37145
rect 11238 37136 11244 37148
rect 11296 37136 11302 37188
rect 11793 37179 11851 37185
rect 11793 37145 11805 37179
rect 11839 37176 11851 37179
rect 15381 37179 15439 37185
rect 11839 37148 15056 37176
rect 11839 37145 11851 37148
rect 11793 37139 11851 37145
rect 9769 37111 9827 37117
rect 9769 37077 9781 37111
rect 9815 37077 9827 37111
rect 9769 37071 9827 37077
rect 10870 37068 10876 37120
rect 10928 37108 10934 37120
rect 15028 37117 15056 37148
rect 15381 37145 15393 37179
rect 15427 37176 15439 37179
rect 17494 37176 17500 37188
rect 15427 37148 17500 37176
rect 15427 37145 15439 37148
rect 15381 37139 15439 37145
rect 17494 37136 17500 37148
rect 17552 37136 17558 37188
rect 17954 37136 17960 37188
rect 18012 37176 18018 37188
rect 18509 37179 18567 37185
rect 18509 37176 18521 37179
rect 18012 37148 18521 37176
rect 18012 37136 18018 37148
rect 18509 37145 18521 37148
rect 18555 37145 18567 37179
rect 19058 37176 19064 37188
rect 18509 37139 18567 37145
rect 18708 37148 19064 37176
rect 11333 37111 11391 37117
rect 11333 37108 11345 37111
rect 10928 37080 11345 37108
rect 10928 37068 10934 37080
rect 11333 37077 11345 37080
rect 11379 37077 11391 37111
rect 11333 37071 11391 37077
rect 15013 37111 15071 37117
rect 15013 37077 15025 37111
rect 15059 37077 15071 37111
rect 15013 37071 15071 37077
rect 15470 37068 15476 37120
rect 15528 37108 15534 37120
rect 16022 37108 16028 37120
rect 15528 37080 16028 37108
rect 15528 37068 15534 37080
rect 16022 37068 16028 37080
rect 16080 37068 16086 37120
rect 16298 37068 16304 37120
rect 16356 37108 16362 37120
rect 16761 37111 16819 37117
rect 16761 37108 16773 37111
rect 16356 37080 16773 37108
rect 16356 37068 16362 37080
rect 16761 37077 16773 37080
rect 16807 37077 16819 37111
rect 16761 37071 16819 37077
rect 17221 37111 17279 37117
rect 17221 37077 17233 37111
rect 17267 37108 17279 37111
rect 18708 37108 18736 37148
rect 19058 37136 19064 37148
rect 19116 37136 19122 37188
rect 20349 37179 20407 37185
rect 20349 37145 20361 37179
rect 20395 37176 20407 37179
rect 20714 37176 20720 37188
rect 20395 37148 20720 37176
rect 20395 37145 20407 37148
rect 20349 37139 20407 37145
rect 20714 37136 20720 37148
rect 20772 37136 20778 37188
rect 21634 37136 21640 37188
rect 21692 37176 21698 37188
rect 24504 37185 24532 37216
rect 25314 37204 25320 37256
rect 25372 37204 25378 37256
rect 21729 37179 21787 37185
rect 21729 37176 21741 37179
rect 21692 37148 21741 37176
rect 21692 37136 21698 37148
rect 21729 37145 21741 37148
rect 21775 37145 21787 37179
rect 21729 37139 21787 37145
rect 24489 37179 24547 37185
rect 24489 37145 24501 37179
rect 24535 37176 24547 37179
rect 24946 37176 24952 37188
rect 24535 37148 24952 37176
rect 24535 37145 24547 37148
rect 24489 37139 24547 37145
rect 24946 37136 24952 37148
rect 25004 37136 25010 37188
rect 17267 37080 18736 37108
rect 18877 37111 18935 37117
rect 17267 37077 17279 37080
rect 17221 37071 17279 37077
rect 18877 37077 18889 37111
rect 18923 37108 18935 37111
rect 20438 37108 20444 37120
rect 18923 37080 20444 37108
rect 18923 37077 18935 37080
rect 18877 37071 18935 37077
rect 20438 37068 20444 37080
rect 20496 37068 20502 37120
rect 23014 37068 23020 37120
rect 23072 37108 23078 37120
rect 23201 37111 23259 37117
rect 23201 37108 23213 37111
rect 23072 37080 23213 37108
rect 23072 37068 23078 37080
rect 23201 37077 23213 37080
rect 23247 37077 23259 37111
rect 23201 37071 23259 37077
rect 23842 37068 23848 37120
rect 23900 37068 23906 37120
rect 24118 37068 24124 37120
rect 24176 37108 24182 37120
rect 25133 37111 25191 37117
rect 25133 37108 25145 37111
rect 24176 37080 25145 37108
rect 24176 37068 24182 37080
rect 25133 37077 25145 37080
rect 25179 37077 25191 37111
rect 25133 37071 25191 37077
rect 1104 37018 25852 37040
rect 1104 36966 7950 37018
rect 8002 36966 8014 37018
rect 8066 36966 8078 37018
rect 8130 36966 8142 37018
rect 8194 36966 8206 37018
rect 8258 36966 17950 37018
rect 18002 36966 18014 37018
rect 18066 36966 18078 37018
rect 18130 36966 18142 37018
rect 18194 36966 18206 37018
rect 18258 36966 25852 37018
rect 1104 36944 25852 36966
rect 5166 36864 5172 36916
rect 5224 36864 5230 36916
rect 5629 36907 5687 36913
rect 5629 36873 5641 36907
rect 5675 36904 5687 36907
rect 9122 36904 9128 36916
rect 5675 36876 9128 36904
rect 5675 36873 5687 36876
rect 5629 36867 5687 36873
rect 9122 36864 9128 36876
rect 9180 36864 9186 36916
rect 9306 36864 9312 36916
rect 9364 36864 9370 36916
rect 9490 36864 9496 36916
rect 9548 36904 9554 36916
rect 9769 36907 9827 36913
rect 9769 36904 9781 36907
rect 9548 36876 9781 36904
rect 9548 36864 9554 36876
rect 9769 36873 9781 36876
rect 9815 36873 9827 36907
rect 9769 36867 9827 36873
rect 10502 36864 10508 36916
rect 10560 36904 10566 36916
rect 10965 36907 11023 36913
rect 10965 36904 10977 36907
rect 10560 36876 10977 36904
rect 10560 36864 10566 36876
rect 10965 36873 10977 36876
rect 11011 36873 11023 36907
rect 10965 36867 11023 36873
rect 12066 36864 12072 36916
rect 12124 36864 12130 36916
rect 12158 36864 12164 36916
rect 12216 36864 12222 36916
rect 12434 36864 12440 36916
rect 12492 36904 12498 36916
rect 12989 36907 13047 36913
rect 12989 36904 13001 36907
rect 12492 36876 13001 36904
rect 12492 36864 12498 36876
rect 12989 36873 13001 36876
rect 13035 36873 13047 36907
rect 12989 36867 13047 36873
rect 13449 36907 13507 36913
rect 13449 36873 13461 36907
rect 13495 36904 13507 36907
rect 14458 36904 14464 36916
rect 13495 36876 14464 36904
rect 13495 36873 13507 36876
rect 13449 36867 13507 36873
rect 14458 36864 14464 36876
rect 14516 36864 14522 36916
rect 15286 36864 15292 36916
rect 15344 36864 15350 36916
rect 15749 36907 15807 36913
rect 15749 36873 15761 36907
rect 15795 36904 15807 36907
rect 16482 36904 16488 36916
rect 15795 36876 16488 36904
rect 15795 36873 15807 36876
rect 15749 36867 15807 36873
rect 16482 36864 16488 36876
rect 16540 36904 16546 36916
rect 18230 36904 18236 36916
rect 16540 36876 18236 36904
rect 16540 36864 16546 36876
rect 18230 36864 18236 36876
rect 18288 36864 18294 36916
rect 18322 36864 18328 36916
rect 18380 36904 18386 36916
rect 18417 36907 18475 36913
rect 18417 36904 18429 36907
rect 18380 36876 18429 36904
rect 18380 36864 18386 36876
rect 18417 36873 18429 36876
rect 18463 36873 18475 36907
rect 18417 36867 18475 36873
rect 19242 36864 19248 36916
rect 19300 36904 19306 36916
rect 19705 36907 19763 36913
rect 19705 36904 19717 36907
rect 19300 36876 19717 36904
rect 19300 36864 19306 36876
rect 19705 36873 19717 36876
rect 19751 36873 19763 36907
rect 19705 36867 19763 36873
rect 20165 36907 20223 36913
rect 20165 36873 20177 36907
rect 20211 36904 20223 36907
rect 22002 36904 22008 36916
rect 20211 36876 22008 36904
rect 20211 36873 20223 36876
rect 20165 36867 20223 36873
rect 22002 36864 22008 36876
rect 22060 36864 22066 36916
rect 23842 36904 23848 36916
rect 22940 36876 23848 36904
rect 8294 36796 8300 36848
rect 8352 36796 8358 36848
rect 13357 36839 13415 36845
rect 13357 36805 13369 36839
rect 13403 36836 13415 36839
rect 13538 36836 13544 36848
rect 13403 36808 13544 36836
rect 13403 36805 13415 36808
rect 13357 36799 13415 36805
rect 13538 36796 13544 36808
rect 13596 36796 13602 36848
rect 15378 36796 15384 36848
rect 15436 36836 15442 36848
rect 16298 36836 16304 36848
rect 15436 36808 16304 36836
rect 15436 36796 15442 36808
rect 16298 36796 16304 36808
rect 16356 36796 16362 36848
rect 17310 36796 17316 36848
rect 17368 36836 17374 36848
rect 17368 36808 19288 36836
rect 17368 36796 17374 36808
rect 1302 36728 1308 36780
rect 1360 36768 1366 36780
rect 1581 36771 1639 36777
rect 1581 36768 1593 36771
rect 1360 36740 1593 36768
rect 1360 36728 1366 36740
rect 1581 36737 1593 36740
rect 1627 36768 1639 36771
rect 2041 36771 2099 36777
rect 2041 36768 2053 36771
rect 1627 36740 2053 36768
rect 1627 36737 1639 36740
rect 1581 36731 1639 36737
rect 2041 36737 2053 36740
rect 2087 36737 2099 36771
rect 2041 36731 2099 36737
rect 5350 36728 5356 36780
rect 5408 36768 5414 36780
rect 5537 36771 5595 36777
rect 5537 36768 5549 36771
rect 5408 36740 5549 36768
rect 5408 36728 5414 36740
rect 5537 36737 5549 36740
rect 5583 36737 5595 36771
rect 5537 36731 5595 36737
rect 10134 36728 10140 36780
rect 10192 36728 10198 36780
rect 10229 36771 10287 36777
rect 10229 36737 10241 36771
rect 10275 36768 10287 36771
rect 10962 36768 10968 36780
rect 10275 36740 10968 36768
rect 10275 36737 10287 36740
rect 10229 36731 10287 36737
rect 10962 36728 10968 36740
rect 11020 36728 11026 36780
rect 14829 36771 14887 36777
rect 14829 36737 14841 36771
rect 14875 36768 14887 36771
rect 15657 36771 15715 36777
rect 15657 36768 15669 36771
rect 14875 36740 15669 36768
rect 14875 36737 14887 36740
rect 14829 36731 14887 36737
rect 15657 36737 15669 36740
rect 15703 36737 15715 36771
rect 16758 36768 16764 36780
rect 15657 36731 15715 36737
rect 15856 36740 16764 36768
rect 15856 36712 15884 36740
rect 16758 36728 16764 36740
rect 16816 36728 16822 36780
rect 19058 36768 19064 36780
rect 18248 36740 19064 36768
rect 5721 36703 5779 36709
rect 5721 36669 5733 36703
rect 5767 36669 5779 36703
rect 5721 36663 5779 36669
rect 4982 36592 4988 36644
rect 5040 36632 5046 36644
rect 5736 36632 5764 36663
rect 7558 36660 7564 36712
rect 7616 36660 7622 36712
rect 7837 36703 7895 36709
rect 7837 36669 7849 36703
rect 7883 36700 7895 36703
rect 9398 36700 9404 36712
rect 7883 36672 9404 36700
rect 7883 36669 7895 36672
rect 7837 36663 7895 36669
rect 9398 36660 9404 36672
rect 9456 36660 9462 36712
rect 9490 36660 9496 36712
rect 9548 36700 9554 36712
rect 10321 36703 10379 36709
rect 10321 36700 10333 36703
rect 9548 36672 10333 36700
rect 9548 36660 9554 36672
rect 10321 36669 10333 36672
rect 10367 36669 10379 36703
rect 10321 36663 10379 36669
rect 11606 36660 11612 36712
rect 11664 36700 11670 36712
rect 12253 36703 12311 36709
rect 12253 36700 12265 36703
rect 11664 36672 12265 36700
rect 11664 36660 11670 36672
rect 12253 36669 12265 36672
rect 12299 36669 12311 36703
rect 12253 36663 12311 36669
rect 13541 36703 13599 36709
rect 13541 36669 13553 36703
rect 13587 36669 13599 36703
rect 13541 36663 13599 36669
rect 5040 36604 5764 36632
rect 5040 36592 5046 36604
rect 11238 36592 11244 36644
rect 11296 36632 11302 36644
rect 11296 36604 11836 36632
rect 11296 36592 11302 36604
rect 1765 36567 1823 36573
rect 1765 36533 1777 36567
rect 1811 36564 1823 36567
rect 1946 36564 1952 36576
rect 1811 36536 1952 36564
rect 1811 36533 1823 36536
rect 1765 36527 1823 36533
rect 1946 36524 1952 36536
rect 2004 36524 2010 36576
rect 9582 36524 9588 36576
rect 9640 36564 9646 36576
rect 11701 36567 11759 36573
rect 11701 36564 11713 36567
rect 9640 36536 11713 36564
rect 9640 36524 9646 36536
rect 11701 36533 11713 36536
rect 11747 36533 11759 36567
rect 11808 36564 11836 36604
rect 11882 36592 11888 36644
rect 11940 36632 11946 36644
rect 13556 36632 13584 36663
rect 15838 36660 15844 36712
rect 15896 36660 15902 36712
rect 16298 36660 16304 36712
rect 16356 36700 16362 36712
rect 18248 36709 18276 36740
rect 19058 36728 19064 36740
rect 19116 36728 19122 36780
rect 16853 36703 16911 36709
rect 16853 36700 16865 36703
rect 16356 36672 16865 36700
rect 16356 36660 16362 36672
rect 16853 36669 16865 36672
rect 16899 36669 16911 36703
rect 16853 36663 16911 36669
rect 18233 36703 18291 36709
rect 18233 36669 18245 36703
rect 18279 36669 18291 36703
rect 18233 36663 18291 36669
rect 18325 36703 18383 36709
rect 18325 36669 18337 36703
rect 18371 36700 18383 36703
rect 18506 36700 18512 36712
rect 18371 36672 18512 36700
rect 18371 36669 18383 36672
rect 18325 36663 18383 36669
rect 18506 36660 18512 36672
rect 18564 36700 18570 36712
rect 19150 36700 19156 36712
rect 18564 36672 19156 36700
rect 18564 36660 18570 36672
rect 19150 36660 19156 36672
rect 19208 36660 19214 36712
rect 19260 36700 19288 36808
rect 19426 36796 19432 36848
rect 19484 36836 19490 36848
rect 22940 36836 22968 36876
rect 23842 36864 23848 36876
rect 23900 36864 23906 36916
rect 19484 36808 22968 36836
rect 19484 36796 19490 36808
rect 23014 36796 23020 36848
rect 23072 36796 23078 36848
rect 24394 36836 24400 36848
rect 24242 36808 24400 36836
rect 24394 36796 24400 36808
rect 24452 36796 24458 36848
rect 20073 36771 20131 36777
rect 20073 36737 20085 36771
rect 20119 36768 20131 36771
rect 22186 36768 22192 36780
rect 20119 36740 22192 36768
rect 20119 36737 20131 36740
rect 20073 36731 20131 36737
rect 22186 36728 22192 36740
rect 22244 36728 22250 36780
rect 22278 36728 22284 36780
rect 22336 36768 22342 36780
rect 22741 36771 22799 36777
rect 22741 36768 22753 36771
rect 22336 36740 22753 36768
rect 22336 36728 22342 36740
rect 22741 36737 22753 36740
rect 22787 36737 22799 36771
rect 22741 36731 22799 36737
rect 24762 36728 24768 36780
rect 24820 36768 24826 36780
rect 25317 36771 25375 36777
rect 25317 36768 25329 36771
rect 24820 36740 25329 36768
rect 24820 36728 24826 36740
rect 25317 36737 25329 36740
rect 25363 36737 25375 36771
rect 25317 36731 25375 36737
rect 20257 36703 20315 36709
rect 20257 36700 20269 36703
rect 19260 36672 20269 36700
rect 20257 36669 20269 36672
rect 20303 36669 20315 36703
rect 20257 36663 20315 36669
rect 21726 36660 21732 36712
rect 21784 36700 21790 36712
rect 23014 36700 23020 36712
rect 21784 36672 23020 36700
rect 21784 36660 21790 36672
rect 23014 36660 23020 36672
rect 23072 36660 23078 36712
rect 11940 36604 13584 36632
rect 11940 36592 11946 36604
rect 15194 36592 15200 36644
rect 15252 36632 15258 36644
rect 19337 36635 19395 36641
rect 19337 36632 19349 36635
rect 15252 36604 19349 36632
rect 15252 36592 15258 36604
rect 19337 36601 19349 36604
rect 19383 36632 19395 36635
rect 20714 36632 20720 36644
rect 19383 36604 20720 36632
rect 19383 36601 19395 36604
rect 19337 36595 19395 36601
rect 20714 36592 20720 36604
rect 20772 36592 20778 36644
rect 25133 36635 25191 36641
rect 25133 36632 25145 36635
rect 24044 36604 25145 36632
rect 16850 36564 16856 36576
rect 11808 36536 16856 36564
rect 11701 36527 11759 36533
rect 16850 36524 16856 36536
rect 16908 36524 16914 36576
rect 18506 36524 18512 36576
rect 18564 36564 18570 36576
rect 18785 36567 18843 36573
rect 18785 36564 18797 36567
rect 18564 36536 18797 36564
rect 18564 36524 18570 36536
rect 18785 36533 18797 36536
rect 18831 36533 18843 36567
rect 18785 36527 18843 36533
rect 19150 36524 19156 36576
rect 19208 36524 19214 36576
rect 23198 36524 23204 36576
rect 23256 36564 23262 36576
rect 24044 36564 24072 36604
rect 25133 36601 25145 36604
rect 25179 36601 25191 36635
rect 25133 36595 25191 36601
rect 23256 36536 24072 36564
rect 23256 36524 23262 36536
rect 24486 36524 24492 36576
rect 24544 36524 24550 36576
rect 1104 36474 25852 36496
rect 1104 36422 2950 36474
rect 3002 36422 3014 36474
rect 3066 36422 3078 36474
rect 3130 36422 3142 36474
rect 3194 36422 3206 36474
rect 3258 36422 12950 36474
rect 13002 36422 13014 36474
rect 13066 36422 13078 36474
rect 13130 36422 13142 36474
rect 13194 36422 13206 36474
rect 13258 36422 22950 36474
rect 23002 36422 23014 36474
rect 23066 36422 23078 36474
rect 23130 36422 23142 36474
rect 23194 36422 23206 36474
rect 23258 36422 25852 36474
rect 1104 36400 25852 36422
rect 6086 36320 6092 36372
rect 6144 36320 6150 36372
rect 8205 36363 8263 36369
rect 8205 36329 8217 36363
rect 8251 36360 8263 36363
rect 8294 36360 8300 36372
rect 8251 36332 8300 36360
rect 8251 36329 8263 36332
rect 8205 36323 8263 36329
rect 8294 36320 8300 36332
rect 8352 36360 8358 36372
rect 9306 36360 9312 36372
rect 8352 36332 9312 36360
rect 8352 36320 8358 36332
rect 9306 36320 9312 36332
rect 9364 36320 9370 36372
rect 15381 36363 15439 36369
rect 15381 36329 15393 36363
rect 15427 36360 15439 36363
rect 15654 36360 15660 36372
rect 15427 36332 15660 36360
rect 15427 36329 15439 36332
rect 15381 36323 15439 36329
rect 15654 36320 15660 36332
rect 15712 36320 15718 36372
rect 16669 36363 16727 36369
rect 16669 36329 16681 36363
rect 16715 36360 16727 36363
rect 19334 36360 19340 36372
rect 16715 36332 19340 36360
rect 16715 36329 16727 36332
rect 16669 36323 16727 36329
rect 19334 36320 19340 36332
rect 19392 36320 19398 36372
rect 19610 36320 19616 36372
rect 19668 36360 19674 36372
rect 20438 36360 20444 36372
rect 19668 36332 20444 36360
rect 19668 36320 19674 36332
rect 20438 36320 20444 36332
rect 20496 36320 20502 36372
rect 21818 36360 21824 36372
rect 20640 36332 21824 36360
rect 9030 36252 9036 36304
rect 9088 36292 9094 36304
rect 15565 36295 15623 36301
rect 15565 36292 15577 36295
rect 9088 36264 15577 36292
rect 9088 36252 9094 36264
rect 15565 36261 15577 36264
rect 15611 36292 15623 36295
rect 15611 36264 16252 36292
rect 15611 36261 15623 36264
rect 15565 36255 15623 36261
rect 7006 36184 7012 36236
rect 7064 36224 7070 36236
rect 7558 36224 7564 36236
rect 7064 36196 7564 36224
rect 7064 36184 7070 36196
rect 7558 36184 7564 36196
rect 7616 36224 7622 36236
rect 7837 36227 7895 36233
rect 7837 36224 7849 36227
rect 7616 36196 7849 36224
rect 7616 36184 7622 36196
rect 7837 36193 7849 36196
rect 7883 36224 7895 36227
rect 9217 36227 9275 36233
rect 9217 36224 9229 36227
rect 7883 36196 9229 36224
rect 7883 36193 7895 36196
rect 7837 36187 7895 36193
rect 9217 36193 9229 36196
rect 9263 36193 9275 36227
rect 9217 36187 9275 36193
rect 10502 36184 10508 36236
rect 10560 36184 10566 36236
rect 14921 36227 14979 36233
rect 14921 36193 14933 36227
rect 14967 36224 14979 36227
rect 15010 36224 15016 36236
rect 14967 36196 15016 36224
rect 14967 36193 14979 36196
rect 14921 36187 14979 36193
rect 15010 36184 15016 36196
rect 15068 36184 15074 36236
rect 16022 36184 16028 36236
rect 16080 36184 16086 36236
rect 8757 36159 8815 36165
rect 8757 36125 8769 36159
rect 8803 36156 8815 36159
rect 10045 36159 10103 36165
rect 10045 36156 10057 36159
rect 8803 36128 10057 36156
rect 8803 36125 8815 36128
rect 8757 36119 8815 36125
rect 10045 36125 10057 36128
rect 10091 36156 10103 36159
rect 10226 36156 10232 36168
rect 10091 36128 10232 36156
rect 10091 36125 10103 36128
rect 10045 36119 10103 36125
rect 10226 36116 10232 36128
rect 10284 36156 10290 36168
rect 12161 36159 12219 36165
rect 12161 36156 12173 36159
rect 10284 36128 12173 36156
rect 10284 36116 10290 36128
rect 12161 36125 12173 36128
rect 12207 36156 12219 36159
rect 12437 36159 12495 36165
rect 12437 36156 12449 36159
rect 12207 36128 12449 36156
rect 12207 36125 12219 36128
rect 12161 36119 12219 36125
rect 12437 36125 12449 36128
rect 12483 36156 12495 36159
rect 15194 36156 15200 36168
rect 12483 36128 15200 36156
rect 12483 36125 12495 36128
rect 12437 36119 12495 36125
rect 15194 36116 15200 36128
rect 15252 36116 15258 36168
rect 16224 36165 16252 36264
rect 17126 36252 17132 36304
rect 17184 36252 17190 36304
rect 17218 36252 17224 36304
rect 17276 36292 17282 36304
rect 20640 36292 20668 36332
rect 21818 36320 21824 36332
rect 21876 36320 21882 36372
rect 22189 36363 22247 36369
rect 22189 36329 22201 36363
rect 22235 36360 22247 36363
rect 22830 36360 22836 36372
rect 22235 36332 22836 36360
rect 22235 36329 22247 36332
rect 22189 36323 22247 36329
rect 22830 36320 22836 36332
rect 22888 36320 22894 36372
rect 23474 36360 23480 36372
rect 23400 36332 23480 36360
rect 17276 36264 20668 36292
rect 20717 36295 20775 36301
rect 17276 36252 17282 36264
rect 20717 36261 20729 36295
rect 20763 36292 20775 36295
rect 22554 36292 22560 36304
rect 20763 36264 22560 36292
rect 20763 36261 20775 36264
rect 20717 36255 20775 36261
rect 22554 36252 22560 36264
rect 22612 36252 22618 36304
rect 17681 36227 17739 36233
rect 17681 36224 17693 36227
rect 16408 36196 17693 36224
rect 16209 36159 16267 36165
rect 16209 36125 16221 36159
rect 16255 36125 16267 36159
rect 16209 36119 16267 36125
rect 16298 36116 16304 36168
rect 16356 36116 16362 36168
rect 6546 36048 6552 36100
rect 6604 36048 6610 36100
rect 7561 36091 7619 36097
rect 7561 36057 7573 36091
rect 7607 36057 7619 36091
rect 7561 36051 7619 36057
rect 7374 35980 7380 36032
rect 7432 36020 7438 36032
rect 7576 36020 7604 36051
rect 9674 36048 9680 36100
rect 9732 36088 9738 36100
rect 10870 36088 10876 36100
rect 9732 36060 10876 36088
rect 9732 36048 9738 36060
rect 10870 36048 10876 36060
rect 10928 36048 10934 36100
rect 11146 36048 11152 36100
rect 11204 36088 11210 36100
rect 11333 36091 11391 36097
rect 11333 36088 11345 36091
rect 11204 36060 11345 36088
rect 11204 36048 11210 36060
rect 11333 36057 11345 36060
rect 11379 36057 11391 36091
rect 16408 36088 16436 36196
rect 17681 36193 17693 36196
rect 17727 36193 17739 36227
rect 20165 36227 20223 36233
rect 17681 36187 17739 36193
rect 18340 36196 20116 36224
rect 17586 36116 17592 36168
rect 17644 36116 17650 36168
rect 11333 36051 11391 36057
rect 12820 36060 16436 36088
rect 17497 36091 17555 36097
rect 12820 36020 12848 36060
rect 17497 36057 17509 36091
rect 17543 36088 17555 36091
rect 18340 36088 18368 36196
rect 18690 36116 18696 36168
rect 18748 36156 18754 36168
rect 19426 36156 19432 36168
rect 18748 36128 19432 36156
rect 18748 36116 18754 36128
rect 19426 36116 19432 36128
rect 19484 36116 19490 36168
rect 17543 36060 18368 36088
rect 20088 36088 20116 36196
rect 20165 36193 20177 36227
rect 20211 36224 20223 36227
rect 20806 36224 20812 36236
rect 20211 36196 20812 36224
rect 20211 36193 20223 36196
rect 20165 36187 20223 36193
rect 20806 36184 20812 36196
rect 20864 36184 20870 36236
rect 21082 36184 21088 36236
rect 21140 36224 21146 36236
rect 21545 36227 21603 36233
rect 21545 36224 21557 36227
rect 21140 36196 21557 36224
rect 21140 36184 21146 36196
rect 21545 36193 21557 36196
rect 21591 36224 21603 36227
rect 23400 36224 23428 36332
rect 23474 36320 23480 36332
rect 23532 36360 23538 36372
rect 24486 36360 24492 36372
rect 23532 36332 24492 36360
rect 23532 36320 23538 36332
rect 24486 36320 24492 36332
rect 24544 36320 24550 36372
rect 23842 36292 23848 36304
rect 23492 36264 23848 36292
rect 23492 36233 23520 36264
rect 23842 36252 23848 36264
rect 23900 36292 23906 36304
rect 25038 36292 25044 36304
rect 23900 36264 25044 36292
rect 23900 36252 23906 36264
rect 25038 36252 25044 36264
rect 25096 36252 25102 36304
rect 21591 36196 23428 36224
rect 23477 36227 23535 36233
rect 21591 36193 21603 36196
rect 21545 36187 21603 36193
rect 23477 36193 23489 36227
rect 23523 36193 23535 36227
rect 23477 36187 23535 36193
rect 23569 36227 23627 36233
rect 23569 36193 23581 36227
rect 23615 36224 23627 36227
rect 23750 36224 23756 36236
rect 23615 36196 23756 36224
rect 23615 36193 23627 36196
rect 23569 36187 23627 36193
rect 23750 36184 23756 36196
rect 23808 36184 23814 36236
rect 20349 36159 20407 36165
rect 20349 36125 20361 36159
rect 20395 36156 20407 36159
rect 20438 36156 20444 36168
rect 20395 36128 20444 36156
rect 20395 36125 20407 36128
rect 20349 36119 20407 36125
rect 20438 36116 20444 36128
rect 20496 36116 20502 36168
rect 21450 36116 21456 36168
rect 21508 36156 21514 36168
rect 22465 36159 22523 36165
rect 22465 36156 22477 36159
rect 21508 36128 22477 36156
rect 21508 36116 21514 36128
rect 22465 36125 22477 36128
rect 22511 36125 22523 36159
rect 22465 36119 22523 36125
rect 24857 36159 24915 36165
rect 24857 36125 24869 36159
rect 24903 36156 24915 36159
rect 25314 36156 25320 36168
rect 24903 36128 25320 36156
rect 24903 36125 24915 36128
rect 24857 36119 24915 36125
rect 25314 36116 25320 36128
rect 25372 36116 25378 36168
rect 20898 36088 20904 36100
rect 20088 36060 20904 36088
rect 17543 36057 17555 36060
rect 17497 36051 17555 36057
rect 20898 36048 20904 36060
rect 20956 36088 20962 36100
rect 20956 36060 25176 36088
rect 20956 36048 20962 36060
rect 7432 35992 12848 36020
rect 7432 35980 7438 35992
rect 13354 35980 13360 36032
rect 13412 36020 13418 36032
rect 14277 36023 14335 36029
rect 14277 36020 14289 36023
rect 13412 35992 14289 36020
rect 13412 35980 13418 35992
rect 14277 35989 14289 35992
rect 14323 35989 14335 36023
rect 14277 35983 14335 35989
rect 14550 35980 14556 36032
rect 14608 36020 14614 36032
rect 14645 36023 14703 36029
rect 14645 36020 14657 36023
rect 14608 35992 14657 36020
rect 14608 35980 14614 35992
rect 14645 35989 14657 35992
rect 14691 35989 14703 36023
rect 14645 35983 14703 35989
rect 14734 35980 14740 36032
rect 14792 35980 14798 36032
rect 16574 35980 16580 36032
rect 16632 36020 16638 36032
rect 18414 36020 18420 36032
rect 16632 35992 18420 36020
rect 16632 35980 16638 35992
rect 18414 35980 18420 35992
rect 18472 36020 18478 36032
rect 20257 36023 20315 36029
rect 20257 36020 20269 36023
rect 18472 35992 20269 36020
rect 18472 35980 18478 35992
rect 20257 35989 20269 35992
rect 20303 36020 20315 36023
rect 20990 36020 20996 36032
rect 20303 35992 20996 36020
rect 20303 35989 20315 35992
rect 20257 35983 20315 35989
rect 20990 35980 20996 35992
rect 21048 35980 21054 36032
rect 21450 35980 21456 36032
rect 21508 36020 21514 36032
rect 21729 36023 21787 36029
rect 21729 36020 21741 36023
rect 21508 35992 21741 36020
rect 21508 35980 21514 35992
rect 21729 35989 21741 35992
rect 21775 35989 21787 36023
rect 21729 35983 21787 35989
rect 21818 35980 21824 36032
rect 21876 36020 21882 36032
rect 22094 36020 22100 36032
rect 21876 35992 22100 36020
rect 21876 35980 21882 35992
rect 22094 35980 22100 35992
rect 22152 36020 22158 36032
rect 22649 36023 22707 36029
rect 22649 36020 22661 36023
rect 22152 35992 22661 36020
rect 22152 35980 22158 35992
rect 22649 35989 22661 35992
rect 22695 35989 22707 36023
rect 22649 35983 22707 35989
rect 23106 35980 23112 36032
rect 23164 36020 23170 36032
rect 23290 36020 23296 36032
rect 23164 35992 23296 36020
rect 23164 35980 23170 35992
rect 23290 35980 23296 35992
rect 23348 35980 23354 36032
rect 23658 35980 23664 36032
rect 23716 35980 23722 36032
rect 24029 36023 24087 36029
rect 24029 35989 24041 36023
rect 24075 36020 24087 36023
rect 24578 36020 24584 36032
rect 24075 35992 24584 36020
rect 24075 35989 24087 35992
rect 24029 35983 24087 35989
rect 24578 35980 24584 35992
rect 24636 35980 24642 36032
rect 25148 36029 25176 36060
rect 25133 36023 25191 36029
rect 25133 35989 25145 36023
rect 25179 35989 25191 36023
rect 25133 35983 25191 35989
rect 1104 35930 25852 35952
rect 1104 35878 7950 35930
rect 8002 35878 8014 35930
rect 8066 35878 8078 35930
rect 8130 35878 8142 35930
rect 8194 35878 8206 35930
rect 8258 35878 17950 35930
rect 18002 35878 18014 35930
rect 18066 35878 18078 35930
rect 18130 35878 18142 35930
rect 18194 35878 18206 35930
rect 18258 35878 25852 35930
rect 1104 35856 25852 35878
rect 5997 35819 6055 35825
rect 5997 35785 6009 35819
rect 6043 35816 6055 35819
rect 7190 35816 7196 35828
rect 6043 35788 7196 35816
rect 6043 35785 6055 35788
rect 5997 35779 6055 35785
rect 7190 35776 7196 35788
rect 7248 35776 7254 35828
rect 9398 35776 9404 35828
rect 9456 35816 9462 35828
rect 11882 35816 11888 35828
rect 9456 35788 11888 35816
rect 9456 35776 9462 35788
rect 11882 35776 11888 35788
rect 11940 35776 11946 35828
rect 14182 35776 14188 35828
rect 14240 35816 14246 35828
rect 15565 35819 15623 35825
rect 15565 35816 15577 35819
rect 14240 35788 15577 35816
rect 14240 35776 14246 35788
rect 15565 35785 15577 35788
rect 15611 35785 15623 35819
rect 15565 35779 15623 35785
rect 16850 35776 16856 35828
rect 16908 35776 16914 35828
rect 17221 35819 17279 35825
rect 17221 35785 17233 35819
rect 17267 35816 17279 35819
rect 19702 35816 19708 35828
rect 17267 35788 19708 35816
rect 17267 35785 17279 35788
rect 17221 35779 17279 35785
rect 19702 35776 19708 35788
rect 19760 35776 19766 35828
rect 20254 35776 20260 35828
rect 20312 35816 20318 35828
rect 20806 35816 20812 35828
rect 20312 35788 20812 35816
rect 20312 35776 20318 35788
rect 20806 35776 20812 35788
rect 20864 35776 20870 35828
rect 23474 35776 23480 35828
rect 23532 35816 23538 35828
rect 23532 35788 25268 35816
rect 23532 35776 23538 35788
rect 6457 35751 6515 35757
rect 6457 35748 6469 35751
rect 5750 35720 6469 35748
rect 6457 35717 6469 35720
rect 6503 35748 6515 35751
rect 6546 35748 6552 35760
rect 6503 35720 6552 35748
rect 6503 35717 6515 35720
rect 6457 35711 6515 35717
rect 6546 35708 6552 35720
rect 6604 35708 6610 35760
rect 9306 35708 9312 35760
rect 9364 35748 9370 35760
rect 9364 35720 9706 35748
rect 9364 35708 9370 35720
rect 12158 35708 12164 35760
rect 12216 35708 12222 35760
rect 15010 35708 15016 35760
rect 15068 35748 15074 35760
rect 15378 35748 15384 35760
rect 15068 35720 15384 35748
rect 15068 35708 15074 35720
rect 15378 35708 15384 35720
rect 15436 35708 15442 35760
rect 15657 35751 15715 35757
rect 15657 35717 15669 35751
rect 15703 35748 15715 35751
rect 18874 35748 18880 35760
rect 15703 35720 18880 35748
rect 15703 35717 15715 35720
rect 15657 35711 15715 35717
rect 18874 35708 18880 35720
rect 18932 35708 18938 35760
rect 18966 35708 18972 35760
rect 19024 35708 19030 35760
rect 19610 35708 19616 35760
rect 19668 35708 19674 35760
rect 24394 35708 24400 35760
rect 24452 35708 24458 35760
rect 25240 35748 25268 35788
rect 25240 35720 25360 35748
rect 13814 35680 13820 35692
rect 13294 35666 13820 35680
rect 13280 35652 13820 35666
rect 4249 35615 4307 35621
rect 4249 35581 4261 35615
rect 4295 35612 4307 35615
rect 4295 35584 4384 35612
rect 4295 35581 4307 35584
rect 4249 35575 4307 35581
rect 4356 35476 4384 35584
rect 4522 35572 4528 35624
rect 4580 35572 4586 35624
rect 10226 35572 10232 35624
rect 10284 35612 10290 35624
rect 10873 35615 10931 35621
rect 10873 35612 10885 35615
rect 10284 35584 10885 35612
rect 10284 35572 10290 35584
rect 10873 35581 10885 35584
rect 10919 35581 10931 35615
rect 10873 35575 10931 35581
rect 11146 35572 11152 35624
rect 11204 35612 11210 35624
rect 11885 35615 11943 35621
rect 11885 35612 11897 35615
rect 11204 35584 11897 35612
rect 11204 35572 11210 35584
rect 11885 35581 11897 35584
rect 11931 35581 11943 35615
rect 13280 35612 13308 35652
rect 13814 35640 13820 35652
rect 13872 35640 13878 35692
rect 14366 35680 14372 35692
rect 13924 35652 14372 35680
rect 11885 35575 11943 35581
rect 11992 35584 13308 35612
rect 11992 35544 12020 35584
rect 13446 35572 13452 35624
rect 13504 35612 13510 35624
rect 13633 35615 13691 35621
rect 13633 35612 13645 35615
rect 13504 35584 13645 35612
rect 13504 35572 13510 35584
rect 13633 35581 13645 35584
rect 13679 35581 13691 35615
rect 13924 35612 13952 35652
rect 14366 35640 14372 35652
rect 14424 35680 14430 35692
rect 17313 35683 17371 35689
rect 14424 35652 15884 35680
rect 14424 35640 14430 35652
rect 13633 35575 13691 35581
rect 13740 35584 13952 35612
rect 11532 35516 12020 35544
rect 11532 35488 11560 35516
rect 5258 35476 5264 35488
rect 4356 35448 5264 35476
rect 5258 35436 5264 35448
rect 5316 35436 5322 35488
rect 10226 35436 10232 35488
rect 10284 35476 10290 35488
rect 10686 35476 10692 35488
rect 10284 35448 10692 35476
rect 10284 35436 10290 35448
rect 10686 35436 10692 35448
rect 10744 35436 10750 35488
rect 11238 35436 11244 35488
rect 11296 35476 11302 35488
rect 11514 35476 11520 35488
rect 11296 35448 11520 35476
rect 11296 35436 11302 35448
rect 11514 35436 11520 35448
rect 11572 35436 11578 35488
rect 11698 35436 11704 35488
rect 11756 35476 11762 35488
rect 13740 35476 13768 35584
rect 14734 35572 14740 35624
rect 14792 35572 14798 35624
rect 15654 35572 15660 35624
rect 15712 35612 15718 35624
rect 15749 35615 15807 35621
rect 15749 35612 15761 35615
rect 15712 35584 15761 35612
rect 15712 35572 15718 35584
rect 15749 35581 15761 35584
rect 15795 35581 15807 35615
rect 15856 35612 15884 35652
rect 17313 35649 17325 35683
rect 17359 35680 17371 35683
rect 17359 35652 18644 35680
rect 17359 35649 17371 35652
rect 17313 35643 17371 35649
rect 17405 35615 17463 35621
rect 17405 35612 17417 35615
rect 15856 35584 17417 35612
rect 15749 35575 15807 35581
rect 17405 35581 17417 35584
rect 17451 35581 17463 35615
rect 17405 35575 17463 35581
rect 14826 35504 14832 35556
rect 14884 35544 14890 35556
rect 15197 35547 15255 35553
rect 15197 35544 15209 35547
rect 14884 35516 15209 35544
rect 14884 35504 14890 35516
rect 15197 35513 15209 35516
rect 15243 35513 15255 35547
rect 18616 35544 18644 35652
rect 18690 35640 18696 35692
rect 18748 35640 18754 35692
rect 25332 35689 25360 35720
rect 25317 35683 25375 35689
rect 25317 35649 25329 35683
rect 25363 35649 25375 35683
rect 25317 35643 25375 35649
rect 19978 35612 19984 35624
rect 18800 35584 19984 35612
rect 18800 35544 18828 35584
rect 19978 35572 19984 35584
rect 20036 35612 20042 35624
rect 23569 35615 23627 35621
rect 20036 35584 22094 35612
rect 20036 35572 20042 35584
rect 20717 35547 20775 35553
rect 20717 35544 20729 35547
rect 18616 35516 18828 35544
rect 19996 35516 20729 35544
rect 15197 35507 15255 35513
rect 11756 35448 13768 35476
rect 11756 35436 11762 35448
rect 13814 35436 13820 35488
rect 13872 35476 13878 35488
rect 13909 35479 13967 35485
rect 13909 35476 13921 35479
rect 13872 35448 13921 35476
rect 13872 35436 13878 35448
rect 13909 35445 13921 35448
rect 13955 35445 13967 35479
rect 13909 35439 13967 35445
rect 18690 35436 18696 35488
rect 18748 35476 18754 35488
rect 19518 35476 19524 35488
rect 18748 35448 19524 35476
rect 18748 35436 18754 35448
rect 19518 35436 19524 35448
rect 19576 35436 19582 35488
rect 19610 35436 19616 35488
rect 19668 35476 19674 35488
rect 19996 35476 20024 35516
rect 20717 35513 20729 35516
rect 20763 35513 20775 35547
rect 22066 35544 22094 35584
rect 23569 35581 23581 35615
rect 23615 35612 23627 35615
rect 23842 35612 23848 35624
rect 23615 35584 23848 35612
rect 23615 35581 23627 35584
rect 23569 35575 23627 35581
rect 23842 35572 23848 35584
rect 23900 35572 23906 35624
rect 25038 35572 25044 35624
rect 25096 35572 25102 35624
rect 22066 35516 24072 35544
rect 20717 35507 20775 35513
rect 19668 35448 20024 35476
rect 19668 35436 19674 35448
rect 20346 35436 20352 35488
rect 20404 35476 20410 35488
rect 20441 35479 20499 35485
rect 20441 35476 20453 35479
rect 20404 35448 20453 35476
rect 20404 35436 20410 35448
rect 20441 35445 20453 35448
rect 20487 35445 20499 35479
rect 20441 35439 20499 35445
rect 22738 35436 22744 35488
rect 22796 35476 22802 35488
rect 23934 35476 23940 35488
rect 22796 35448 23940 35476
rect 22796 35436 22802 35448
rect 23934 35436 23940 35448
rect 23992 35436 23998 35488
rect 24044 35476 24072 35516
rect 25222 35476 25228 35488
rect 24044 35448 25228 35476
rect 25222 35436 25228 35448
rect 25280 35436 25286 35488
rect 1104 35386 25852 35408
rect 1104 35334 2950 35386
rect 3002 35334 3014 35386
rect 3066 35334 3078 35386
rect 3130 35334 3142 35386
rect 3194 35334 3206 35386
rect 3258 35334 12950 35386
rect 13002 35334 13014 35386
rect 13066 35334 13078 35386
rect 13130 35334 13142 35386
rect 13194 35334 13206 35386
rect 13258 35334 22950 35386
rect 23002 35334 23014 35386
rect 23066 35334 23078 35386
rect 23130 35334 23142 35386
rect 23194 35334 23206 35386
rect 23258 35334 25852 35386
rect 1104 35312 25852 35334
rect 4522 35232 4528 35284
rect 4580 35272 4586 35284
rect 5261 35275 5319 35281
rect 5261 35272 5273 35275
rect 4580 35244 5273 35272
rect 4580 35232 4586 35244
rect 5261 35241 5273 35244
rect 5307 35272 5319 35275
rect 5307 35244 7604 35272
rect 5307 35241 5319 35244
rect 5261 35235 5319 35241
rect 7576 35204 7604 35244
rect 7650 35232 7656 35284
rect 7708 35232 7714 35284
rect 10318 35232 10324 35284
rect 10376 35232 10382 35284
rect 13467 35275 13525 35281
rect 13467 35241 13479 35275
rect 13513 35272 13525 35275
rect 13722 35272 13728 35284
rect 13513 35244 13728 35272
rect 13513 35241 13525 35244
rect 13467 35235 13525 35241
rect 13722 35232 13728 35244
rect 13780 35232 13786 35284
rect 13998 35232 14004 35284
rect 14056 35272 14062 35284
rect 14461 35275 14519 35281
rect 14461 35272 14473 35275
rect 14056 35244 14473 35272
rect 14056 35232 14062 35244
rect 14461 35241 14473 35244
rect 14507 35241 14519 35275
rect 14461 35235 14519 35241
rect 15565 35275 15623 35281
rect 15565 35241 15577 35275
rect 15611 35272 15623 35275
rect 15930 35272 15936 35284
rect 15611 35244 15936 35272
rect 15611 35241 15623 35244
rect 15565 35235 15623 35241
rect 10778 35204 10784 35216
rect 7576 35176 10784 35204
rect 10778 35164 10784 35176
rect 10836 35164 10842 35216
rect 6086 35096 6092 35148
rect 6144 35136 6150 35148
rect 8205 35139 8263 35145
rect 8205 35136 8217 35139
rect 6144 35108 8217 35136
rect 6144 35096 6150 35108
rect 8205 35105 8217 35108
rect 8251 35105 8263 35139
rect 8205 35099 8263 35105
rect 9398 35096 9404 35148
rect 9456 35136 9462 35148
rect 9677 35139 9735 35145
rect 9677 35136 9689 35139
rect 9456 35108 9689 35136
rect 9456 35096 9462 35108
rect 9677 35105 9689 35108
rect 9723 35105 9735 35139
rect 11698 35136 11704 35148
rect 9677 35099 9735 35105
rect 9876 35108 11704 35136
rect 7006 35028 7012 35080
rect 7064 35028 7070 35080
rect 9876 35068 9904 35108
rect 11698 35096 11704 35108
rect 11756 35096 11762 35148
rect 11977 35139 12035 35145
rect 11977 35105 11989 35139
rect 12023 35136 12035 35139
rect 12158 35136 12164 35148
rect 12023 35108 12164 35136
rect 12023 35105 12035 35108
rect 11977 35099 12035 35105
rect 12158 35096 12164 35108
rect 12216 35136 12222 35148
rect 14090 35136 14096 35148
rect 12216 35108 14096 35136
rect 12216 35096 12222 35108
rect 14090 35096 14096 35108
rect 14148 35096 14154 35148
rect 7116 35040 9904 35068
rect 9953 35071 10011 35077
rect 7116 35012 7144 35040
rect 9953 35037 9965 35071
rect 9999 35068 10011 35071
rect 10502 35068 10508 35080
rect 9999 35040 10508 35068
rect 9999 35037 10011 35040
rect 9953 35031 10011 35037
rect 10502 35028 10508 35040
rect 10560 35028 10566 35080
rect 13722 35028 13728 35080
rect 13780 35028 13786 35080
rect 6733 35003 6791 35009
rect 6302 34972 6592 35000
rect 6564 34944 6592 34972
rect 6733 34969 6745 35003
rect 6779 35000 6791 35003
rect 7098 35000 7104 35012
rect 6779 34972 7104 35000
rect 6779 34969 6791 34972
rect 6733 34963 6791 34969
rect 7098 34960 7104 34972
rect 7156 34960 7162 35012
rect 13170 35000 13176 35012
rect 13018 34972 13176 35000
rect 13170 34960 13176 34972
rect 13228 35000 13234 35012
rect 13814 35000 13820 35012
rect 13228 34972 13820 35000
rect 13228 34960 13234 34972
rect 13814 34960 13820 34972
rect 13872 35000 13878 35012
rect 14093 35003 14151 35009
rect 14093 35000 14105 35003
rect 13872 34972 14105 35000
rect 13872 34960 13878 34972
rect 14093 34969 14105 34972
rect 14139 34969 14151 35003
rect 14476 35000 14504 35235
rect 15930 35232 15936 35244
rect 15988 35232 15994 35284
rect 16022 35232 16028 35284
rect 16080 35272 16086 35284
rect 22738 35272 22744 35284
rect 16080 35244 22744 35272
rect 16080 35232 16086 35244
rect 22738 35232 22744 35244
rect 22796 35232 22802 35284
rect 23477 35275 23535 35281
rect 23477 35241 23489 35275
rect 23523 35272 23535 35275
rect 23658 35272 23664 35284
rect 23523 35244 23664 35272
rect 23523 35241 23535 35244
rect 23477 35235 23535 35241
rect 23658 35232 23664 35244
rect 23716 35232 23722 35284
rect 14642 35164 14648 35216
rect 14700 35204 14706 35216
rect 18141 35207 18199 35213
rect 18141 35204 18153 35207
rect 14700 35176 18153 35204
rect 14700 35164 14706 35176
rect 18141 35173 18153 35176
rect 18187 35173 18199 35207
rect 18141 35167 18199 35173
rect 18782 35164 18788 35216
rect 18840 35204 18846 35216
rect 19610 35204 19616 35216
rect 18840 35176 19616 35204
rect 18840 35164 18846 35176
rect 19610 35164 19616 35176
rect 19668 35164 19674 35216
rect 20162 35164 20168 35216
rect 20220 35204 20226 35216
rect 24118 35204 24124 35216
rect 20220 35176 24124 35204
rect 20220 35164 20226 35176
rect 24118 35164 24124 35176
rect 24176 35164 24182 35216
rect 15013 35139 15071 35145
rect 15013 35105 15025 35139
rect 15059 35136 15071 35139
rect 17310 35136 17316 35148
rect 15059 35108 17316 35136
rect 15059 35105 15071 35108
rect 15013 35099 15071 35105
rect 17310 35096 17316 35108
rect 17368 35096 17374 35148
rect 18693 35139 18751 35145
rect 18693 35136 18705 35139
rect 17420 35108 18705 35136
rect 14734 35028 14740 35080
rect 14792 35068 14798 35080
rect 15197 35071 15255 35077
rect 15197 35068 15209 35071
rect 14792 35040 15209 35068
rect 14792 35028 14798 35040
rect 15197 35037 15209 35040
rect 15243 35037 15255 35071
rect 15197 35031 15255 35037
rect 16942 35028 16948 35080
rect 17000 35068 17006 35080
rect 17420 35068 17448 35108
rect 18693 35105 18705 35108
rect 18739 35105 18751 35139
rect 18693 35099 18751 35105
rect 18874 35096 18880 35148
rect 18932 35136 18938 35148
rect 20533 35139 20591 35145
rect 20533 35136 20545 35139
rect 18932 35108 19334 35136
rect 18932 35096 18938 35108
rect 17000 35040 17448 35068
rect 18509 35071 18567 35077
rect 17000 35028 17006 35040
rect 18509 35037 18521 35071
rect 18555 35068 18567 35071
rect 18598 35068 18604 35080
rect 18555 35040 18604 35068
rect 18555 35037 18567 35040
rect 18509 35031 18567 35037
rect 18598 35028 18604 35040
rect 18656 35028 18662 35080
rect 19306 35068 19334 35108
rect 20364 35108 20545 35136
rect 20364 35068 20392 35108
rect 20533 35105 20545 35108
rect 20579 35105 20591 35139
rect 20533 35099 20591 35105
rect 21726 35096 21732 35148
rect 21784 35096 21790 35148
rect 21821 35139 21879 35145
rect 21821 35105 21833 35139
rect 21867 35136 21879 35139
rect 21910 35136 21916 35148
rect 21867 35108 21916 35136
rect 21867 35105 21879 35108
rect 21821 35099 21879 35105
rect 21910 35096 21916 35108
rect 21968 35096 21974 35148
rect 22925 35139 22983 35145
rect 22925 35105 22937 35139
rect 22971 35136 22983 35139
rect 25038 35136 25044 35148
rect 22971 35108 25044 35136
rect 22971 35105 22983 35108
rect 22925 35099 22983 35105
rect 25038 35096 25044 35108
rect 25096 35096 25102 35148
rect 19306 35040 20392 35068
rect 20438 35028 20444 35080
rect 20496 35028 20502 35080
rect 22278 35028 22284 35080
rect 22336 35068 22342 35080
rect 24857 35071 24915 35077
rect 22336 35040 23152 35068
rect 22336 35028 22342 35040
rect 15105 35003 15163 35009
rect 15105 35000 15117 35003
rect 14476 34972 15117 35000
rect 14093 34963 14151 34969
rect 15105 34969 15117 34972
rect 15151 34969 15163 35003
rect 20162 35000 20168 35012
rect 15105 34963 15163 34969
rect 18616 34972 20168 35000
rect 6546 34892 6552 34944
rect 6604 34932 6610 34944
rect 7282 34932 7288 34944
rect 6604 34904 7288 34932
rect 6604 34892 6610 34904
rect 7282 34892 7288 34904
rect 7340 34892 7346 34944
rect 7834 34892 7840 34944
rect 7892 34932 7898 34944
rect 8021 34935 8079 34941
rect 8021 34932 8033 34935
rect 7892 34904 8033 34932
rect 7892 34892 7898 34904
rect 8021 34901 8033 34904
rect 8067 34901 8079 34935
rect 8021 34895 8079 34901
rect 8113 34935 8171 34941
rect 8113 34901 8125 34935
rect 8159 34932 8171 34935
rect 9030 34932 9036 34944
rect 8159 34904 9036 34932
rect 8159 34901 8171 34904
rect 8113 34895 8171 34901
rect 9030 34892 9036 34904
rect 9088 34892 9094 34944
rect 9858 34892 9864 34944
rect 9916 34892 9922 34944
rect 12158 34892 12164 34944
rect 12216 34932 12222 34944
rect 13998 34932 14004 34944
rect 12216 34904 14004 34932
rect 12216 34892 12222 34904
rect 13998 34892 14004 34904
rect 14056 34892 14062 34944
rect 18616 34941 18644 34972
rect 20162 34960 20168 34972
rect 20220 35000 20226 35012
rect 20349 35003 20407 35009
rect 20349 35000 20361 35003
rect 20220 34972 20361 35000
rect 20220 34960 20226 34972
rect 20349 34969 20361 34972
rect 20395 34969 20407 35003
rect 20456 35000 20484 35028
rect 23017 35003 23075 35009
rect 23017 35000 23029 35003
rect 20456 34972 23029 35000
rect 20349 34963 20407 34969
rect 23017 34969 23029 34972
rect 23063 34969 23075 35003
rect 23124 35000 23152 35040
rect 24857 35037 24869 35071
rect 24903 35068 24915 35071
rect 25317 35071 25375 35077
rect 25317 35068 25329 35071
rect 24903 35040 25329 35068
rect 24903 35037 24915 35040
rect 24857 35031 24915 35037
rect 25317 35037 25329 35040
rect 25363 35068 25375 35071
rect 25406 35068 25412 35080
rect 25363 35040 25412 35068
rect 25363 35037 25375 35040
rect 25317 35031 25375 35037
rect 25406 35028 25412 35040
rect 25464 35028 25470 35080
rect 23124 34972 25176 35000
rect 23017 34963 23075 34969
rect 18601 34935 18659 34941
rect 18601 34901 18613 34935
rect 18647 34901 18659 34935
rect 18601 34895 18659 34901
rect 18690 34892 18696 34944
rect 18748 34932 18754 34944
rect 19981 34935 20039 34941
rect 19981 34932 19993 34935
rect 18748 34904 19993 34932
rect 18748 34892 18754 34904
rect 19981 34901 19993 34904
rect 20027 34901 20039 34935
rect 19981 34895 20039 34901
rect 20254 34892 20260 34944
rect 20312 34932 20318 34944
rect 20441 34935 20499 34941
rect 20441 34932 20453 34935
rect 20312 34904 20453 34932
rect 20312 34892 20318 34904
rect 20441 34901 20453 34904
rect 20487 34901 20499 34935
rect 20441 34895 20499 34901
rect 20714 34892 20720 34944
rect 20772 34932 20778 34944
rect 21913 34935 21971 34941
rect 21913 34932 21925 34935
rect 20772 34904 21925 34932
rect 20772 34892 20778 34904
rect 21913 34901 21925 34904
rect 21959 34901 21971 34935
rect 21913 34895 21971 34901
rect 22281 34935 22339 34941
rect 22281 34901 22293 34935
rect 22327 34932 22339 34935
rect 22738 34932 22744 34944
rect 22327 34904 22744 34932
rect 22327 34901 22339 34904
rect 22281 34895 22339 34901
rect 22738 34892 22744 34904
rect 22796 34892 22802 34944
rect 23109 34935 23167 34941
rect 23109 34901 23121 34935
rect 23155 34932 23167 34935
rect 23198 34932 23204 34944
rect 23155 34904 23204 34932
rect 23155 34901 23167 34904
rect 23109 34895 23167 34901
rect 23198 34892 23204 34904
rect 23256 34892 23262 34944
rect 24394 34892 24400 34944
rect 24452 34932 24458 34944
rect 24673 34935 24731 34941
rect 24673 34932 24685 34935
rect 24452 34904 24685 34932
rect 24452 34892 24458 34904
rect 24673 34901 24685 34904
rect 24719 34932 24731 34935
rect 24762 34932 24768 34944
rect 24719 34904 24768 34932
rect 24719 34901 24731 34904
rect 24673 34895 24731 34901
rect 24762 34892 24768 34904
rect 24820 34892 24826 34944
rect 25148 34941 25176 34972
rect 25133 34935 25191 34941
rect 25133 34901 25145 34935
rect 25179 34901 25191 34935
rect 25133 34895 25191 34901
rect 1104 34842 25852 34864
rect 1104 34790 7950 34842
rect 8002 34790 8014 34842
rect 8066 34790 8078 34842
rect 8130 34790 8142 34842
rect 8194 34790 8206 34842
rect 8258 34790 17950 34842
rect 18002 34790 18014 34842
rect 18066 34790 18078 34842
rect 18130 34790 18142 34842
rect 18194 34790 18206 34842
rect 18258 34790 25852 34842
rect 1104 34768 25852 34790
rect 1765 34731 1823 34737
rect 1765 34697 1777 34731
rect 1811 34728 1823 34731
rect 2682 34728 2688 34740
rect 1811 34700 2688 34728
rect 1811 34697 1823 34700
rect 1765 34691 1823 34697
rect 2682 34688 2688 34700
rect 2740 34688 2746 34740
rect 3513 34731 3571 34737
rect 3513 34697 3525 34731
rect 3559 34728 3571 34731
rect 4982 34728 4988 34740
rect 3559 34700 4988 34728
rect 3559 34697 3571 34700
rect 3513 34691 3571 34697
rect 4982 34688 4988 34700
rect 5040 34688 5046 34740
rect 5629 34731 5687 34737
rect 5629 34697 5641 34731
rect 5675 34728 5687 34731
rect 5810 34728 5816 34740
rect 5675 34700 5816 34728
rect 5675 34697 5687 34700
rect 5629 34691 5687 34697
rect 5644 34660 5672 34691
rect 5810 34688 5816 34700
rect 5868 34728 5874 34740
rect 6546 34728 6552 34740
rect 5868 34700 6552 34728
rect 5868 34688 5874 34700
rect 6546 34688 6552 34700
rect 6604 34688 6610 34740
rect 7190 34688 7196 34740
rect 7248 34688 7254 34740
rect 8478 34688 8484 34740
rect 8536 34728 8542 34740
rect 9033 34731 9091 34737
rect 9033 34728 9045 34731
rect 8536 34700 9045 34728
rect 8536 34688 8542 34700
rect 9033 34697 9045 34700
rect 9079 34697 9091 34731
rect 9401 34731 9459 34737
rect 9401 34728 9413 34731
rect 9033 34691 9091 34697
rect 9140 34700 9413 34728
rect 4554 34632 5672 34660
rect 7009 34663 7067 34669
rect 7009 34629 7021 34663
rect 7055 34660 7067 34663
rect 7208 34660 7236 34688
rect 7055 34632 7236 34660
rect 7055 34629 7067 34632
rect 7009 34623 7067 34629
rect 7282 34620 7288 34672
rect 7340 34660 7346 34672
rect 9140 34660 9168 34700
rect 9401 34697 9413 34700
rect 9447 34697 9459 34731
rect 9401 34691 9459 34697
rect 11146 34688 11152 34740
rect 11204 34728 11210 34740
rect 13722 34728 13728 34740
rect 11204 34700 13728 34728
rect 11204 34688 11210 34700
rect 9766 34660 9772 34672
rect 7340 34632 7498 34660
rect 8312 34632 9168 34660
rect 9416 34632 9772 34660
rect 7340 34620 7346 34632
rect 1578 34552 1584 34604
rect 1636 34592 1642 34604
rect 2041 34595 2099 34601
rect 2041 34592 2053 34595
rect 1636 34564 2053 34592
rect 1636 34552 1642 34564
rect 2041 34561 2053 34564
rect 2087 34561 2099 34595
rect 2041 34555 2099 34561
rect 5258 34484 5264 34536
rect 5316 34524 5322 34536
rect 6730 34524 6736 34536
rect 5316 34496 6736 34524
rect 5316 34484 5322 34496
rect 6730 34484 6736 34496
rect 6788 34524 6794 34536
rect 7006 34524 7012 34536
rect 6788 34496 7012 34524
rect 6788 34484 6794 34496
rect 7006 34484 7012 34496
rect 7064 34484 7070 34536
rect 7650 34484 7656 34536
rect 7708 34524 7714 34536
rect 8312 34524 8340 34632
rect 9416 34592 9444 34632
rect 9766 34620 9772 34632
rect 9824 34620 9830 34672
rect 13170 34660 13176 34672
rect 12742 34632 13176 34660
rect 13170 34620 13176 34632
rect 13228 34620 13234 34672
rect 13464 34601 13492 34700
rect 13722 34688 13728 34700
rect 13780 34688 13786 34740
rect 13998 34688 14004 34740
rect 14056 34728 14062 34740
rect 14093 34731 14151 34737
rect 14093 34728 14105 34731
rect 14056 34700 14105 34728
rect 14056 34688 14062 34700
rect 14093 34697 14105 34700
rect 14139 34697 14151 34731
rect 14093 34691 14151 34697
rect 14461 34731 14519 34737
rect 14461 34697 14473 34731
rect 14507 34728 14519 34731
rect 16022 34728 16028 34740
rect 14507 34700 16028 34728
rect 14507 34697 14519 34700
rect 14461 34691 14519 34697
rect 16022 34688 16028 34700
rect 16080 34688 16086 34740
rect 16850 34688 16856 34740
rect 16908 34728 16914 34740
rect 16908 34700 18644 34728
rect 16908 34688 16914 34700
rect 13817 34663 13875 34669
rect 13817 34629 13829 34663
rect 13863 34660 13875 34663
rect 14274 34660 14280 34672
rect 13863 34632 14280 34660
rect 13863 34629 13875 34632
rect 13817 34623 13875 34629
rect 14274 34620 14280 34632
rect 14332 34660 14338 34672
rect 14553 34663 14611 34669
rect 14553 34660 14565 34663
rect 14332 34632 14565 34660
rect 14332 34620 14338 34632
rect 14553 34629 14565 34632
rect 14599 34629 14611 34663
rect 18230 34660 18236 34672
rect 17894 34632 18236 34660
rect 14553 34623 14611 34629
rect 18230 34620 18236 34632
rect 18288 34620 18294 34672
rect 18616 34660 18644 34700
rect 18966 34688 18972 34740
rect 19024 34728 19030 34740
rect 19429 34731 19487 34737
rect 19429 34728 19441 34731
rect 19024 34700 19441 34728
rect 19024 34688 19030 34700
rect 19429 34697 19441 34700
rect 19475 34728 19487 34731
rect 19475 34700 22324 34728
rect 19475 34697 19487 34700
rect 19429 34691 19487 34697
rect 19334 34660 19340 34672
rect 18616 34632 19340 34660
rect 18616 34601 18644 34632
rect 19334 34620 19340 34632
rect 19392 34660 19398 34672
rect 19518 34660 19524 34672
rect 19392 34632 19524 34660
rect 19392 34620 19398 34632
rect 19518 34620 19524 34632
rect 19576 34620 19582 34672
rect 7708 34496 8340 34524
rect 8496 34564 9444 34592
rect 9493 34595 9551 34601
rect 7708 34484 7714 34496
rect 8496 34465 8524 34564
rect 9493 34561 9505 34595
rect 9539 34592 9551 34595
rect 13449 34595 13507 34601
rect 9539 34564 11744 34592
rect 9539 34561 9551 34564
rect 9493 34555 9551 34561
rect 9677 34527 9735 34533
rect 9677 34493 9689 34527
rect 9723 34524 9735 34527
rect 10042 34524 10048 34536
rect 9723 34496 10048 34524
rect 9723 34493 9735 34496
rect 9677 34487 9735 34493
rect 10042 34484 10048 34496
rect 10100 34484 10106 34536
rect 11716 34524 11744 34564
rect 13449 34561 13461 34595
rect 13495 34561 13507 34595
rect 13449 34555 13507 34561
rect 18601 34595 18659 34601
rect 18601 34561 18613 34595
rect 18647 34561 18659 34595
rect 18601 34555 18659 34561
rect 19058 34552 19064 34604
rect 19116 34592 19122 34604
rect 19242 34592 19248 34604
rect 19116 34564 19248 34592
rect 19116 34552 19122 34564
rect 19242 34552 19248 34564
rect 19300 34592 19306 34604
rect 19300 34564 19656 34592
rect 19300 34552 19306 34564
rect 12802 34524 12808 34536
rect 11716 34496 12808 34524
rect 12802 34484 12808 34496
rect 12860 34484 12866 34536
rect 13173 34527 13231 34533
rect 13173 34493 13185 34527
rect 13219 34524 13231 34527
rect 14645 34527 14703 34533
rect 13219 34496 13492 34524
rect 13219 34493 13231 34496
rect 13173 34487 13231 34493
rect 13464 34468 13492 34496
rect 14645 34493 14657 34527
rect 14691 34493 14703 34527
rect 14645 34487 14703 34493
rect 8481 34459 8539 34465
rect 8481 34425 8493 34459
rect 8527 34425 8539 34459
rect 8481 34419 8539 34425
rect 13446 34416 13452 34468
rect 13504 34416 13510 34468
rect 4982 34348 4988 34400
rect 5040 34397 5046 34400
rect 5040 34391 5055 34397
rect 5043 34357 5055 34391
rect 5040 34351 5055 34357
rect 5040 34348 5046 34351
rect 11698 34348 11704 34400
rect 11756 34348 11762 34400
rect 14550 34348 14556 34400
rect 14608 34388 14614 34400
rect 14660 34388 14688 34487
rect 16758 34484 16764 34536
rect 16816 34524 16822 34536
rect 16853 34527 16911 34533
rect 16853 34524 16865 34527
rect 16816 34496 16865 34524
rect 16816 34484 16822 34496
rect 16853 34493 16865 34496
rect 16899 34493 16911 34527
rect 16853 34487 16911 34493
rect 18325 34527 18383 34533
rect 18325 34493 18337 34527
rect 18371 34524 18383 34527
rect 18371 34496 18552 34524
rect 18371 34493 18383 34496
rect 18325 34487 18383 34493
rect 18524 34456 18552 34496
rect 19426 34484 19432 34536
rect 19484 34524 19490 34536
rect 19628 34533 19656 34564
rect 19702 34552 19708 34604
rect 19760 34592 19766 34604
rect 22296 34592 22324 34700
rect 22370 34688 22376 34740
rect 22428 34688 22434 34740
rect 22462 34688 22468 34740
rect 22520 34688 22526 34740
rect 23198 34688 23204 34740
rect 23256 34688 23262 34740
rect 25222 34592 25228 34604
rect 19760 34564 22094 34592
rect 22296 34564 25228 34592
rect 19760 34552 19766 34564
rect 19521 34527 19579 34533
rect 19521 34524 19533 34527
rect 19484 34496 19533 34524
rect 19484 34484 19490 34496
rect 19521 34493 19533 34496
rect 19567 34493 19579 34527
rect 19521 34487 19579 34493
rect 19613 34527 19671 34533
rect 19613 34493 19625 34527
rect 19659 34493 19671 34527
rect 19613 34487 19671 34493
rect 20254 34484 20260 34536
rect 20312 34484 20318 34536
rect 22066 34524 22094 34564
rect 25222 34552 25228 34564
rect 25280 34552 25286 34604
rect 25314 34552 25320 34604
rect 25372 34552 25378 34604
rect 22278 34524 22284 34536
rect 22066 34496 22284 34524
rect 22278 34484 22284 34496
rect 22336 34484 22342 34536
rect 22557 34527 22615 34533
rect 22557 34493 22569 34527
rect 22603 34493 22615 34527
rect 22557 34487 22615 34493
rect 20162 34456 20168 34468
rect 18524 34428 20168 34456
rect 20162 34416 20168 34428
rect 20220 34416 20226 34468
rect 22572 34456 22600 34487
rect 23658 34484 23664 34536
rect 23716 34524 23722 34536
rect 23716 34496 25176 34524
rect 23716 34484 23722 34496
rect 25148 34465 25176 34496
rect 22480 34428 22600 34456
rect 25133 34459 25191 34465
rect 22480 34400 22508 34428
rect 25133 34425 25145 34459
rect 25179 34425 25191 34459
rect 25133 34419 25191 34425
rect 14608 34360 14688 34388
rect 14608 34348 14614 34360
rect 19058 34348 19064 34400
rect 19116 34348 19122 34400
rect 22002 34348 22008 34400
rect 22060 34348 22066 34400
rect 22462 34348 22468 34400
rect 22520 34348 22526 34400
rect 1104 34298 25852 34320
rect 1104 34246 2950 34298
rect 3002 34246 3014 34298
rect 3066 34246 3078 34298
rect 3130 34246 3142 34298
rect 3194 34246 3206 34298
rect 3258 34246 12950 34298
rect 13002 34246 13014 34298
rect 13066 34246 13078 34298
rect 13130 34246 13142 34298
rect 13194 34246 13206 34298
rect 13258 34246 22950 34298
rect 23002 34246 23014 34298
rect 23066 34246 23078 34298
rect 23130 34246 23142 34298
rect 23194 34246 23206 34298
rect 23258 34246 25852 34298
rect 1104 34224 25852 34246
rect 7009 34187 7067 34193
rect 7009 34153 7021 34187
rect 7055 34184 7067 34187
rect 7282 34184 7288 34196
rect 7055 34156 7288 34184
rect 7055 34153 7067 34156
rect 7009 34147 7067 34153
rect 7282 34144 7288 34156
rect 7340 34184 7346 34196
rect 8478 34184 8484 34196
rect 7340 34156 8484 34184
rect 7340 34144 7346 34156
rect 8478 34144 8484 34156
rect 8536 34184 8542 34196
rect 8665 34187 8723 34193
rect 8665 34184 8677 34187
rect 8536 34156 8677 34184
rect 8536 34144 8542 34156
rect 8665 34153 8677 34156
rect 8711 34153 8723 34187
rect 8665 34147 8723 34153
rect 9122 34144 9128 34196
rect 9180 34144 9186 34196
rect 10962 34144 10968 34196
rect 11020 34184 11026 34196
rect 12253 34187 12311 34193
rect 12253 34184 12265 34187
rect 11020 34156 12265 34184
rect 11020 34144 11026 34156
rect 12253 34153 12265 34156
rect 12299 34153 12311 34187
rect 12253 34147 12311 34153
rect 20165 34187 20223 34193
rect 20165 34153 20177 34187
rect 20211 34184 20223 34187
rect 20714 34184 20720 34196
rect 20211 34156 20720 34184
rect 20211 34153 20223 34156
rect 20165 34147 20223 34153
rect 20714 34144 20720 34156
rect 20772 34144 20778 34196
rect 21634 34184 21640 34196
rect 20916 34156 21640 34184
rect 20916 34116 20944 34156
rect 21634 34144 21640 34156
rect 21692 34144 21698 34196
rect 6564 34088 9720 34116
rect 4706 34008 4712 34060
rect 4764 34048 4770 34060
rect 4893 34051 4951 34057
rect 4893 34048 4905 34051
rect 4764 34020 4905 34048
rect 4764 34008 4770 34020
rect 4893 34017 4905 34020
rect 4939 34048 4951 34051
rect 4982 34048 4988 34060
rect 4939 34020 4988 34048
rect 4939 34017 4951 34020
rect 4893 34011 4951 34017
rect 4982 34008 4988 34020
rect 5040 34048 5046 34060
rect 6564 34048 6592 34088
rect 5040 34020 6592 34048
rect 5040 34008 5046 34020
rect 9582 34008 9588 34060
rect 9640 34008 9646 34060
rect 9692 34057 9720 34088
rect 19628 34088 20944 34116
rect 19628 34057 19656 34088
rect 9677 34051 9735 34057
rect 9677 34017 9689 34051
rect 9723 34017 9735 34051
rect 12805 34051 12863 34057
rect 12805 34048 12817 34051
rect 9677 34011 9735 34017
rect 12406 34020 12817 34048
rect 6641 33983 6699 33989
rect 6641 33949 6653 33983
rect 6687 33980 6699 33983
rect 6730 33980 6736 33992
rect 6687 33952 6736 33980
rect 6687 33949 6699 33952
rect 6641 33943 6699 33949
rect 6730 33940 6736 33952
rect 6788 33980 6794 33992
rect 7742 33980 7748 33992
rect 6788 33952 7748 33980
rect 6788 33940 6794 33952
rect 7742 33940 7748 33952
rect 7800 33940 7806 33992
rect 9214 33940 9220 33992
rect 9272 33980 9278 33992
rect 12406 33980 12434 34020
rect 12805 34017 12817 34020
rect 12851 34017 12863 34051
rect 12805 34011 12863 34017
rect 19613 34051 19671 34057
rect 19613 34017 19625 34051
rect 19659 34017 19671 34051
rect 19613 34011 19671 34017
rect 20809 34051 20867 34057
rect 20809 34017 20821 34051
rect 20855 34048 20867 34051
rect 22278 34048 22284 34060
rect 20855 34020 22284 34048
rect 20855 34017 20867 34020
rect 20809 34011 20867 34017
rect 22278 34008 22284 34020
rect 22336 34048 22342 34060
rect 23474 34048 23480 34060
rect 22336 34020 23480 34048
rect 22336 34008 22342 34020
rect 23474 34008 23480 34020
rect 23532 34008 23538 34060
rect 9272 33952 12434 33980
rect 12713 33983 12771 33989
rect 9272 33940 9278 33952
rect 12713 33949 12725 33983
rect 12759 33980 12771 33983
rect 13354 33980 13360 33992
rect 12759 33952 13360 33980
rect 12759 33949 12771 33952
rect 12713 33943 12771 33949
rect 13354 33940 13360 33952
rect 13412 33940 13418 33992
rect 19797 33983 19855 33989
rect 19797 33949 19809 33983
rect 19843 33980 19855 33983
rect 20254 33980 20260 33992
rect 19843 33952 20260 33980
rect 19843 33949 19855 33952
rect 19797 33943 19855 33949
rect 20254 33940 20260 33952
rect 20312 33940 20318 33992
rect 23566 33940 23572 33992
rect 23624 33940 23630 33992
rect 24581 33983 24639 33989
rect 24581 33949 24593 33983
rect 24627 33980 24639 33983
rect 24670 33980 24676 33992
rect 24627 33952 24676 33980
rect 24627 33949 24639 33952
rect 24581 33943 24639 33949
rect 24670 33940 24676 33952
rect 24728 33940 24734 33992
rect 5810 33872 5816 33924
rect 5868 33872 5874 33924
rect 6365 33915 6423 33921
rect 6365 33881 6377 33915
rect 6411 33912 6423 33915
rect 7282 33912 7288 33924
rect 6411 33884 7288 33912
rect 6411 33881 6423 33884
rect 6365 33875 6423 33881
rect 7282 33872 7288 33884
rect 7340 33872 7346 33924
rect 12621 33915 12679 33921
rect 12621 33881 12633 33915
rect 12667 33912 12679 33915
rect 15654 33912 15660 33924
rect 12667 33884 15660 33912
rect 12667 33881 12679 33884
rect 12621 33875 12679 33881
rect 15654 33872 15660 33884
rect 15712 33872 15718 33924
rect 19518 33872 19524 33924
rect 19576 33912 19582 33924
rect 20622 33912 20628 33924
rect 19576 33884 20628 33912
rect 19576 33872 19582 33884
rect 20622 33872 20628 33884
rect 20680 33912 20686 33924
rect 21085 33915 21143 33921
rect 21085 33912 21097 33915
rect 20680 33884 21097 33912
rect 20680 33872 20686 33884
rect 21085 33881 21097 33884
rect 21131 33881 21143 33915
rect 22646 33912 22652 33924
rect 22310 33884 22652 33912
rect 21085 33875 21143 33881
rect 22646 33872 22652 33884
rect 22704 33912 22710 33924
rect 22925 33915 22983 33921
rect 22925 33912 22937 33915
rect 22704 33884 22937 33912
rect 22704 33872 22710 33884
rect 22925 33881 22937 33884
rect 22971 33912 22983 33915
rect 24854 33912 24860 33924
rect 22971 33884 24860 33912
rect 22971 33881 22983 33884
rect 22925 33875 22983 33881
rect 24854 33872 24860 33884
rect 24912 33912 24918 33924
rect 25409 33915 25467 33921
rect 25409 33912 25421 33915
rect 24912 33884 25421 33912
rect 24912 33872 24918 33884
rect 25409 33881 25421 33884
rect 25455 33881 25467 33915
rect 25409 33875 25467 33881
rect 9493 33847 9551 33853
rect 9493 33813 9505 33847
rect 9539 33844 9551 33847
rect 12342 33844 12348 33856
rect 9539 33816 12348 33844
rect 9539 33813 9551 33816
rect 9493 33807 9551 33813
rect 12342 33804 12348 33816
rect 12400 33804 12406 33856
rect 13633 33847 13691 33853
rect 13633 33813 13645 33847
rect 13679 33844 13691 33847
rect 13722 33844 13728 33856
rect 13679 33816 13728 33844
rect 13679 33813 13691 33816
rect 13633 33807 13691 33813
rect 13722 33804 13728 33816
rect 13780 33804 13786 33856
rect 18230 33804 18236 33856
rect 18288 33844 18294 33856
rect 18782 33844 18788 33856
rect 18288 33816 18788 33844
rect 18288 33804 18294 33816
rect 18782 33804 18788 33816
rect 18840 33804 18846 33856
rect 18966 33804 18972 33856
rect 19024 33844 19030 33856
rect 19705 33847 19763 33853
rect 19705 33844 19717 33847
rect 19024 33816 19717 33844
rect 19024 33804 19030 33816
rect 19705 33813 19717 33816
rect 19751 33813 19763 33847
rect 19705 33807 19763 33813
rect 22462 33804 22468 33856
rect 22520 33844 22526 33856
rect 22557 33847 22615 33853
rect 22557 33844 22569 33847
rect 22520 33816 22569 33844
rect 22520 33804 22526 33816
rect 22557 33813 22569 33816
rect 22603 33813 22615 33847
rect 22557 33807 22615 33813
rect 23753 33847 23811 33853
rect 23753 33813 23765 33847
rect 23799 33844 23811 33847
rect 24394 33844 24400 33856
rect 23799 33816 24400 33844
rect 23799 33813 23811 33816
rect 23753 33807 23811 33813
rect 24394 33804 24400 33816
rect 24452 33804 24458 33856
rect 24670 33804 24676 33856
rect 24728 33844 24734 33856
rect 24765 33847 24823 33853
rect 24765 33844 24777 33847
rect 24728 33816 24777 33844
rect 24728 33804 24734 33816
rect 24765 33813 24777 33816
rect 24811 33813 24823 33847
rect 24765 33807 24823 33813
rect 25314 33804 25320 33856
rect 25372 33804 25378 33856
rect 1104 33754 25852 33776
rect 1104 33702 7950 33754
rect 8002 33702 8014 33754
rect 8066 33702 8078 33754
rect 8130 33702 8142 33754
rect 8194 33702 8206 33754
rect 8258 33702 17950 33754
rect 18002 33702 18014 33754
rect 18066 33702 18078 33754
rect 18130 33702 18142 33754
rect 18194 33702 18206 33754
rect 18258 33702 25852 33754
rect 1104 33680 25852 33702
rect 7558 33600 7564 33652
rect 7616 33640 7622 33652
rect 7616 33612 9352 33640
rect 7616 33600 7622 33612
rect 8478 33532 8484 33584
rect 8536 33532 8542 33584
rect 9324 33572 9352 33612
rect 9490 33600 9496 33652
rect 9548 33600 9554 33652
rect 9950 33600 9956 33652
rect 10008 33600 10014 33652
rect 11885 33643 11943 33649
rect 11885 33609 11897 33643
rect 11931 33640 11943 33643
rect 11974 33640 11980 33652
rect 11931 33612 11980 33640
rect 11931 33609 11943 33612
rect 11885 33603 11943 33609
rect 11974 33600 11980 33612
rect 12032 33600 12038 33652
rect 12250 33600 12256 33652
rect 12308 33640 12314 33652
rect 13814 33640 13820 33652
rect 12308 33612 13820 33640
rect 12308 33600 12314 33612
rect 13814 33600 13820 33612
rect 13872 33600 13878 33652
rect 13906 33600 13912 33652
rect 13964 33600 13970 33652
rect 14918 33600 14924 33652
rect 14976 33600 14982 33652
rect 18601 33643 18659 33649
rect 18601 33609 18613 33643
rect 18647 33640 18659 33643
rect 19610 33640 19616 33652
rect 18647 33612 19616 33640
rect 18647 33609 18659 33612
rect 18601 33603 18659 33609
rect 19610 33600 19616 33612
rect 19668 33600 19674 33652
rect 21910 33600 21916 33652
rect 21968 33640 21974 33652
rect 22373 33643 22431 33649
rect 22373 33640 22385 33643
rect 21968 33612 22385 33640
rect 21968 33600 21974 33612
rect 22373 33609 22385 33612
rect 22419 33640 22431 33643
rect 22646 33640 22652 33652
rect 22419 33612 22652 33640
rect 22419 33609 22431 33612
rect 22373 33603 22431 33609
rect 22646 33600 22652 33612
rect 22704 33600 22710 33652
rect 25225 33643 25283 33649
rect 25225 33609 25237 33643
rect 25271 33640 25283 33643
rect 25498 33640 25504 33652
rect 25271 33612 25504 33640
rect 25271 33609 25283 33612
rect 25225 33603 25283 33609
rect 25498 33600 25504 33612
rect 25556 33600 25562 33652
rect 10321 33575 10379 33581
rect 10321 33572 10333 33575
rect 9324 33544 10333 33572
rect 10321 33541 10333 33544
rect 10367 33541 10379 33575
rect 10321 33535 10379 33541
rect 10686 33532 10692 33584
rect 10744 33572 10750 33584
rect 11698 33572 11704 33584
rect 10744 33544 11704 33572
rect 10744 33532 10750 33544
rect 11698 33532 11704 33544
rect 11756 33572 11762 33584
rect 11756 33544 14044 33572
rect 11756 33532 11762 33544
rect 9766 33464 9772 33516
rect 9824 33504 9830 33516
rect 9950 33504 9956 33516
rect 9824 33476 9956 33504
rect 9824 33464 9830 33476
rect 9950 33464 9956 33476
rect 10008 33464 10014 33516
rect 11882 33504 11888 33516
rect 11256 33476 11888 33504
rect 7742 33396 7748 33448
rect 7800 33396 7806 33448
rect 8021 33439 8079 33445
rect 8021 33405 8033 33439
rect 8067 33436 8079 33439
rect 9214 33436 9220 33448
rect 8067 33408 9220 33436
rect 8067 33405 8079 33408
rect 8021 33399 8079 33405
rect 9214 33396 9220 33408
rect 9272 33396 9278 33448
rect 10410 33396 10416 33448
rect 10468 33396 10474 33448
rect 10597 33439 10655 33445
rect 10597 33405 10609 33439
rect 10643 33436 10655 33439
rect 10778 33436 10784 33448
rect 10643 33408 10784 33436
rect 10643 33405 10655 33408
rect 10597 33399 10655 33405
rect 10778 33396 10784 33408
rect 10836 33396 10842 33448
rect 9030 33328 9036 33380
rect 9088 33368 9094 33380
rect 9490 33368 9496 33380
rect 9088 33340 9496 33368
rect 9088 33328 9094 33340
rect 9490 33328 9496 33340
rect 9548 33328 9554 33380
rect 6454 33260 6460 33312
rect 6512 33300 6518 33312
rect 11256 33309 11284 33476
rect 11882 33464 11888 33476
rect 11940 33504 11946 33516
rect 12253 33507 12311 33513
rect 12253 33504 12265 33507
rect 11940 33476 12265 33504
rect 11940 33464 11946 33476
rect 12253 33473 12265 33476
rect 12299 33473 12311 33507
rect 12253 33467 12311 33473
rect 13817 33507 13875 33513
rect 13817 33473 13829 33507
rect 13863 33504 13875 33507
rect 13906 33504 13912 33516
rect 13863 33476 13912 33504
rect 13863 33473 13875 33476
rect 13817 33467 13875 33473
rect 13906 33464 13912 33476
rect 13964 33464 13970 33516
rect 11514 33396 11520 33448
rect 11572 33436 11578 33448
rect 11609 33439 11667 33445
rect 11609 33436 11621 33439
rect 11572 33408 11621 33436
rect 11572 33396 11578 33408
rect 11609 33405 11621 33408
rect 11655 33436 11667 33439
rect 12066 33436 12072 33448
rect 11655 33408 12072 33436
rect 11655 33405 11667 33408
rect 11609 33399 11667 33405
rect 12066 33396 12072 33408
rect 12124 33436 12130 33448
rect 12345 33439 12403 33445
rect 12345 33436 12357 33439
rect 12124 33408 12357 33436
rect 12124 33396 12130 33408
rect 12345 33405 12357 33408
rect 12391 33405 12403 33439
rect 12345 33399 12403 33405
rect 12526 33396 12532 33448
rect 12584 33396 12590 33448
rect 14016 33445 14044 33544
rect 15562 33532 15568 33584
rect 15620 33572 15626 33584
rect 15620 33544 18828 33572
rect 15620 33532 15626 33544
rect 15010 33464 15016 33516
rect 15068 33464 15074 33516
rect 14001 33439 14059 33445
rect 14001 33405 14013 33439
rect 14047 33405 14059 33439
rect 14001 33399 14059 33405
rect 14090 33396 14096 33448
rect 14148 33436 14154 33448
rect 18800 33445 18828 33544
rect 23474 33464 23480 33516
rect 23532 33464 23538 33516
rect 24854 33464 24860 33516
rect 24912 33464 24918 33516
rect 14737 33439 14795 33445
rect 14737 33436 14749 33439
rect 14148 33408 14749 33436
rect 14148 33396 14154 33408
rect 14737 33405 14749 33408
rect 14783 33405 14795 33439
rect 14737 33399 14795 33405
rect 18693 33439 18751 33445
rect 18693 33405 18705 33439
rect 18739 33405 18751 33439
rect 18693 33399 18751 33405
rect 18785 33439 18843 33445
rect 18785 33405 18797 33439
rect 18831 33405 18843 33439
rect 18785 33399 18843 33405
rect 13538 33328 13544 33380
rect 13596 33368 13602 33380
rect 18233 33371 18291 33377
rect 18233 33368 18245 33371
rect 13596 33340 18245 33368
rect 13596 33328 13602 33340
rect 18233 33337 18245 33340
rect 18279 33337 18291 33371
rect 18708 33368 18736 33399
rect 23750 33396 23756 33448
rect 23808 33396 23814 33448
rect 23290 33368 23296 33380
rect 18708 33340 23296 33368
rect 18233 33331 18291 33337
rect 23290 33328 23296 33340
rect 23348 33328 23354 33380
rect 11241 33303 11299 33309
rect 11241 33300 11253 33303
rect 6512 33272 11253 33300
rect 6512 33260 6518 33272
rect 11241 33269 11253 33272
rect 11287 33269 11299 33303
rect 11241 33263 11299 33269
rect 13446 33260 13452 33312
rect 13504 33260 13510 33312
rect 15381 33303 15439 33309
rect 15381 33269 15393 33303
rect 15427 33300 15439 33303
rect 16022 33300 16028 33312
rect 15427 33272 16028 33300
rect 15427 33269 15439 33272
rect 15381 33263 15439 33269
rect 16022 33260 16028 33272
rect 16080 33260 16086 33312
rect 1104 33210 25852 33232
rect 1104 33158 2950 33210
rect 3002 33158 3014 33210
rect 3066 33158 3078 33210
rect 3130 33158 3142 33210
rect 3194 33158 3206 33210
rect 3258 33158 12950 33210
rect 13002 33158 13014 33210
rect 13066 33158 13078 33210
rect 13130 33158 13142 33210
rect 13194 33158 13206 33210
rect 13258 33158 22950 33210
rect 23002 33158 23014 33210
rect 23066 33158 23078 33210
rect 23130 33158 23142 33210
rect 23194 33158 23206 33210
rect 23258 33158 25852 33210
rect 1104 33136 25852 33158
rect 7282 33056 7288 33108
rect 7340 33096 7346 33108
rect 9306 33096 9312 33108
rect 7340 33068 9312 33096
rect 7340 33056 7346 33068
rect 9306 33056 9312 33068
rect 9364 33056 9370 33108
rect 9490 33056 9496 33108
rect 9548 33096 9554 33108
rect 9861 33099 9919 33105
rect 9548 33068 9812 33096
rect 9548 33056 9554 33068
rect 9784 33028 9812 33068
rect 9861 33065 9873 33099
rect 9907 33096 9919 33099
rect 10134 33096 10140 33108
rect 9907 33068 10140 33096
rect 9907 33065 9919 33068
rect 9861 33059 9919 33065
rect 10134 33056 10140 33068
rect 10192 33056 10198 33108
rect 13633 33099 13691 33105
rect 13633 33065 13645 33099
rect 13679 33096 13691 33099
rect 15010 33096 15016 33108
rect 13679 33068 15016 33096
rect 13679 33065 13691 33068
rect 13633 33059 13691 33065
rect 15010 33056 15016 33068
rect 15068 33056 15074 33108
rect 16942 33056 16948 33108
rect 17000 33096 17006 33108
rect 17678 33096 17684 33108
rect 17000 33068 17684 33096
rect 17000 33056 17006 33068
rect 17678 33056 17684 33068
rect 17736 33056 17742 33108
rect 18601 33099 18659 33105
rect 18601 33065 18613 33099
rect 18647 33096 18659 33099
rect 19518 33096 19524 33108
rect 18647 33068 19524 33096
rect 18647 33065 18659 33068
rect 18601 33059 18659 33065
rect 19518 33056 19524 33068
rect 19576 33056 19582 33108
rect 19705 33099 19763 33105
rect 19705 33065 19717 33099
rect 19751 33096 19763 33099
rect 21726 33096 21732 33108
rect 19751 33068 21732 33096
rect 19751 33065 19763 33068
rect 19705 33059 19763 33065
rect 21726 33056 21732 33068
rect 21784 33056 21790 33108
rect 22554 33056 22560 33108
rect 22612 33096 22618 33108
rect 23106 33096 23112 33108
rect 22612 33068 23112 33096
rect 22612 33056 22618 33068
rect 23106 33056 23112 33068
rect 23164 33056 23170 33108
rect 11701 33031 11759 33037
rect 11701 33028 11713 33031
rect 9784 33000 11713 33028
rect 11701 32997 11713 33000
rect 11747 32997 11759 33031
rect 11701 32991 11759 32997
rect 16666 32988 16672 33040
rect 16724 33028 16730 33040
rect 16724 33000 16988 33028
rect 16724 32988 16730 33000
rect 5537 32963 5595 32969
rect 5537 32929 5549 32963
rect 5583 32960 5595 32963
rect 7742 32960 7748 32972
rect 5583 32932 7748 32960
rect 5583 32929 5595 32932
rect 5537 32923 5595 32929
rect 7742 32920 7748 32932
rect 7800 32920 7806 32972
rect 9214 32920 9220 32972
rect 9272 32920 9278 32972
rect 9306 32920 9312 32972
rect 9364 32960 9370 32972
rect 11606 32960 11612 32972
rect 9364 32932 11612 32960
rect 9364 32920 9370 32932
rect 11606 32920 11612 32932
rect 11664 32920 11670 32972
rect 12158 32920 12164 32972
rect 12216 32920 12222 32972
rect 12253 32963 12311 32969
rect 12253 32929 12265 32963
rect 12299 32929 12311 32963
rect 12253 32923 12311 32929
rect 13081 32963 13139 32969
rect 13081 32929 13093 32963
rect 13127 32960 13139 32963
rect 13630 32960 13636 32972
rect 13127 32932 13636 32960
rect 13127 32929 13139 32932
rect 13081 32923 13139 32929
rect 8294 32852 8300 32904
rect 8352 32892 8358 32904
rect 12268 32892 12296 32923
rect 13630 32920 13636 32932
rect 13688 32920 13694 32972
rect 16850 32920 16856 32972
rect 16908 32920 16914 32972
rect 16960 32960 16988 33000
rect 18322 32988 18328 33040
rect 18380 33028 18386 33040
rect 18380 33000 19656 33028
rect 18380 32988 18386 33000
rect 19628 32960 19656 33000
rect 20162 32988 20168 33040
rect 20220 33028 20226 33040
rect 20441 33031 20499 33037
rect 20441 33028 20453 33031
rect 20220 33000 20453 33028
rect 20220 32988 20226 33000
rect 20441 32997 20453 33000
rect 20487 32997 20499 33031
rect 20441 32991 20499 32997
rect 20714 32960 20720 32972
rect 16960 32932 19564 32960
rect 19628 32932 20720 32960
rect 8352 32864 12296 32892
rect 8352 32852 8358 32864
rect 12710 32852 12716 32904
rect 12768 32892 12774 32904
rect 13173 32895 13231 32901
rect 13173 32892 13185 32895
rect 12768 32864 13185 32892
rect 12768 32852 12774 32864
rect 13173 32861 13185 32864
rect 13219 32861 13231 32895
rect 13173 32855 13231 32861
rect 14550 32852 14556 32904
rect 14608 32892 14614 32904
rect 15102 32892 15108 32904
rect 14608 32864 15108 32892
rect 14608 32852 14614 32864
rect 15102 32852 15108 32864
rect 15160 32852 15166 32904
rect 19536 32901 19564 32932
rect 20714 32920 20720 32932
rect 20772 32920 20778 32972
rect 21910 32960 21916 32972
rect 20824 32932 21916 32960
rect 19521 32895 19579 32901
rect 19521 32861 19533 32895
rect 19567 32861 19579 32895
rect 19521 32855 19579 32861
rect 5813 32827 5871 32833
rect 5813 32793 5825 32827
rect 5859 32824 5871 32827
rect 6086 32824 6092 32836
rect 5859 32796 6092 32824
rect 5859 32793 5871 32796
rect 5813 32787 5871 32793
rect 6086 32784 6092 32796
rect 6144 32784 6150 32836
rect 7098 32824 7104 32836
rect 7038 32796 7104 32824
rect 7098 32784 7104 32796
rect 7156 32824 7162 32836
rect 7653 32827 7711 32833
rect 7653 32824 7665 32827
rect 7156 32796 7665 32824
rect 7156 32784 7162 32796
rect 7653 32793 7665 32796
rect 7699 32824 7711 32827
rect 8478 32824 8484 32836
rect 7699 32796 8484 32824
rect 7699 32793 7711 32796
rect 7653 32787 7711 32793
rect 8478 32784 8484 32796
rect 8536 32784 8542 32836
rect 9401 32827 9459 32833
rect 9401 32793 9413 32827
rect 9447 32824 9459 32827
rect 9766 32824 9772 32836
rect 9447 32796 9772 32824
rect 9447 32793 9459 32796
rect 9401 32787 9459 32793
rect 9766 32784 9772 32796
rect 9824 32784 9830 32836
rect 12069 32827 12127 32833
rect 12069 32793 12081 32827
rect 12115 32824 12127 32827
rect 15746 32824 15752 32836
rect 12115 32796 15752 32824
rect 12115 32793 12127 32796
rect 12069 32787 12127 32793
rect 15746 32784 15752 32796
rect 15804 32784 15810 32836
rect 16114 32784 16120 32836
rect 16172 32824 16178 32836
rect 17129 32827 17187 32833
rect 17129 32824 17141 32827
rect 16172 32796 17141 32824
rect 16172 32784 16178 32796
rect 17129 32793 17141 32796
rect 17175 32793 17187 32827
rect 17129 32787 17187 32793
rect 17512 32796 17618 32824
rect 9490 32716 9496 32768
rect 9548 32716 9554 32768
rect 9582 32716 9588 32768
rect 9640 32756 9646 32768
rect 10137 32759 10195 32765
rect 10137 32756 10149 32759
rect 9640 32728 10149 32756
rect 9640 32716 9646 32728
rect 10137 32725 10149 32728
rect 10183 32725 10195 32759
rect 10137 32719 10195 32725
rect 13265 32759 13323 32765
rect 13265 32725 13277 32759
rect 13311 32756 13323 32759
rect 13354 32756 13360 32768
rect 13311 32728 13360 32756
rect 13311 32725 13323 32728
rect 13265 32719 13323 32725
rect 13354 32716 13360 32728
rect 13412 32716 13418 32768
rect 13998 32716 14004 32768
rect 14056 32756 14062 32768
rect 14277 32759 14335 32765
rect 14277 32756 14289 32759
rect 14056 32728 14289 32756
rect 14056 32716 14062 32728
rect 14277 32725 14289 32728
rect 14323 32725 14335 32759
rect 14277 32719 14335 32725
rect 16206 32716 16212 32768
rect 16264 32756 16270 32768
rect 16301 32759 16359 32765
rect 16301 32756 16313 32759
rect 16264 32728 16313 32756
rect 16264 32716 16270 32728
rect 16301 32725 16313 32728
rect 16347 32756 16359 32759
rect 17512 32756 17540 32796
rect 18138 32756 18144 32768
rect 16347 32728 18144 32756
rect 16347 32725 16359 32728
rect 16301 32719 16359 32725
rect 18138 32716 18144 32728
rect 18196 32756 18202 32768
rect 18782 32756 18788 32768
rect 18196 32728 18788 32756
rect 18196 32716 18202 32728
rect 18782 32716 18788 32728
rect 18840 32756 18846 32768
rect 18877 32759 18935 32765
rect 18877 32756 18889 32759
rect 18840 32728 18889 32756
rect 18840 32716 18846 32728
rect 18877 32725 18889 32728
rect 18923 32756 18935 32759
rect 20824 32756 20852 32932
rect 21910 32920 21916 32932
rect 21968 32920 21974 32972
rect 22189 32963 22247 32969
rect 22189 32929 22201 32963
rect 22235 32960 22247 32963
rect 22278 32960 22284 32972
rect 22235 32932 22284 32960
rect 22235 32929 22247 32932
rect 22189 32923 22247 32929
rect 22278 32920 22284 32932
rect 22336 32960 22342 32972
rect 22554 32960 22560 32972
rect 22336 32932 22560 32960
rect 22336 32920 22342 32932
rect 22554 32920 22560 32932
rect 22612 32920 22618 32972
rect 22830 32920 22836 32972
rect 22888 32960 22894 32972
rect 23201 32963 23259 32969
rect 23201 32960 23213 32963
rect 22888 32932 23213 32960
rect 22888 32920 22894 32932
rect 23201 32929 23213 32932
rect 23247 32929 23259 32963
rect 23201 32923 23259 32929
rect 23017 32895 23075 32901
rect 23017 32861 23029 32895
rect 23063 32892 23075 32895
rect 23290 32892 23296 32904
rect 23063 32864 23296 32892
rect 23063 32861 23075 32864
rect 23017 32855 23075 32861
rect 23290 32852 23296 32864
rect 23348 32852 23354 32904
rect 24857 32895 24915 32901
rect 24857 32861 24869 32895
rect 24903 32892 24915 32895
rect 25314 32892 25320 32904
rect 24903 32864 25320 32892
rect 24903 32861 24915 32864
rect 24857 32855 24915 32861
rect 25314 32852 25320 32864
rect 25372 32852 25378 32904
rect 21913 32827 21971 32833
rect 21913 32793 21925 32827
rect 21959 32824 21971 32827
rect 22462 32824 22468 32836
rect 21959 32796 22468 32824
rect 21959 32793 21971 32796
rect 21913 32787 21971 32793
rect 22462 32784 22468 32796
rect 22520 32824 22526 32836
rect 23198 32824 23204 32836
rect 22520 32796 23204 32824
rect 22520 32784 22526 32796
rect 23198 32784 23204 32796
rect 23256 32784 23262 32836
rect 18923 32728 20852 32756
rect 18923 32725 18935 32728
rect 18877 32719 18935 32725
rect 22646 32716 22652 32768
rect 22704 32716 22710 32768
rect 23106 32716 23112 32768
rect 23164 32716 23170 32768
rect 23658 32716 23664 32768
rect 23716 32756 23722 32768
rect 25133 32759 25191 32765
rect 25133 32756 25145 32759
rect 23716 32728 25145 32756
rect 23716 32716 23722 32728
rect 25133 32725 25145 32728
rect 25179 32725 25191 32759
rect 25133 32719 25191 32725
rect 1104 32666 25852 32688
rect 1104 32614 7950 32666
rect 8002 32614 8014 32666
rect 8066 32614 8078 32666
rect 8130 32614 8142 32666
rect 8194 32614 8206 32666
rect 8258 32614 17950 32666
rect 18002 32614 18014 32666
rect 18066 32614 18078 32666
rect 18130 32614 18142 32666
rect 18194 32614 18206 32666
rect 18258 32614 25852 32666
rect 1104 32592 25852 32614
rect 7098 32512 7104 32564
rect 7156 32512 7162 32564
rect 8665 32555 8723 32561
rect 8665 32521 8677 32555
rect 8711 32552 8723 32555
rect 9490 32552 9496 32564
rect 8711 32524 9496 32552
rect 8711 32521 8723 32524
rect 8665 32515 8723 32521
rect 9490 32512 9496 32524
rect 9548 32512 9554 32564
rect 9582 32512 9588 32564
rect 9640 32552 9646 32564
rect 11238 32552 11244 32564
rect 9640 32524 11244 32552
rect 9640 32512 9646 32524
rect 11238 32512 11244 32524
rect 11296 32512 11302 32564
rect 12710 32512 12716 32564
rect 12768 32512 12774 32564
rect 13354 32512 13360 32564
rect 13412 32512 13418 32564
rect 14918 32512 14924 32564
rect 14976 32552 14982 32564
rect 18049 32555 18107 32561
rect 18049 32552 18061 32555
rect 14976 32524 18061 32552
rect 14976 32512 14982 32524
rect 18049 32521 18061 32524
rect 18095 32521 18107 32555
rect 18049 32515 18107 32521
rect 18417 32555 18475 32561
rect 18417 32521 18429 32555
rect 18463 32552 18475 32555
rect 19058 32552 19064 32564
rect 18463 32524 19064 32552
rect 18463 32521 18475 32524
rect 18417 32515 18475 32521
rect 19058 32512 19064 32524
rect 19116 32512 19122 32564
rect 19613 32555 19671 32561
rect 19613 32521 19625 32555
rect 19659 32552 19671 32555
rect 19702 32552 19708 32564
rect 19659 32524 19708 32552
rect 19659 32521 19671 32524
rect 19613 32515 19671 32521
rect 19702 32512 19708 32524
rect 19760 32512 19766 32564
rect 20898 32512 20904 32564
rect 20956 32552 20962 32564
rect 20993 32555 21051 32561
rect 20993 32552 21005 32555
rect 20956 32524 21005 32552
rect 20956 32512 20962 32524
rect 20993 32521 21005 32524
rect 21039 32521 21051 32555
rect 20993 32515 21051 32521
rect 21085 32555 21143 32561
rect 21085 32521 21097 32555
rect 21131 32552 21143 32555
rect 21266 32552 21272 32564
rect 21131 32524 21272 32552
rect 21131 32521 21143 32524
rect 21085 32515 21143 32521
rect 21266 32512 21272 32524
rect 21324 32512 21330 32564
rect 22094 32512 22100 32564
rect 22152 32552 22158 32564
rect 22649 32555 22707 32561
rect 22649 32552 22661 32555
rect 22152 32524 22661 32552
rect 22152 32512 22158 32524
rect 22649 32521 22661 32524
rect 22695 32521 22707 32555
rect 25130 32552 25136 32564
rect 22649 32515 22707 32521
rect 22848 32524 25136 32552
rect 8478 32444 8484 32496
rect 8536 32484 8542 32496
rect 9600 32484 9628 32512
rect 8536 32456 9890 32484
rect 8536 32444 8542 32456
rect 13722 32444 13728 32496
rect 13780 32484 13786 32496
rect 13780 32456 14766 32484
rect 13780 32444 13786 32456
rect 17034 32444 17040 32496
rect 17092 32484 17098 32496
rect 17221 32487 17279 32493
rect 17221 32484 17233 32487
rect 17092 32456 17233 32484
rect 17092 32444 17098 32456
rect 17221 32453 17233 32456
rect 17267 32453 17279 32487
rect 17221 32447 17279 32453
rect 18506 32444 18512 32496
rect 18564 32444 18570 32496
rect 19794 32444 19800 32496
rect 19852 32484 19858 32496
rect 19852 32456 22048 32484
rect 19852 32444 19858 32456
rect 1302 32376 1308 32428
rect 1360 32416 1366 32428
rect 1581 32419 1639 32425
rect 1581 32416 1593 32419
rect 1360 32388 1593 32416
rect 1360 32376 1366 32388
rect 1581 32385 1593 32388
rect 1627 32416 1639 32419
rect 2041 32419 2099 32425
rect 2041 32416 2053 32419
rect 1627 32388 2053 32416
rect 1627 32385 1639 32388
rect 1581 32379 1639 32385
rect 2041 32385 2053 32388
rect 2087 32385 2099 32419
rect 2041 32379 2099 32385
rect 16209 32419 16267 32425
rect 16209 32385 16221 32419
rect 16255 32416 16267 32419
rect 16850 32416 16856 32428
rect 16255 32388 16856 32416
rect 16255 32385 16267 32388
rect 16209 32379 16267 32385
rect 16850 32376 16856 32388
rect 16908 32376 16914 32428
rect 18874 32416 18880 32428
rect 17052 32388 18880 32416
rect 4982 32308 4988 32360
rect 5040 32308 5046 32360
rect 7466 32308 7472 32360
rect 7524 32308 7530 32360
rect 7742 32308 7748 32360
rect 7800 32348 7806 32360
rect 9122 32348 9128 32360
rect 7800 32320 9128 32348
rect 7800 32308 7806 32320
rect 9122 32308 9128 32320
rect 9180 32308 9186 32360
rect 9398 32308 9404 32360
rect 9456 32308 9462 32360
rect 11790 32308 11796 32360
rect 11848 32348 11854 32360
rect 12526 32348 12532 32360
rect 11848 32320 12532 32348
rect 11848 32308 11854 32320
rect 12526 32308 12532 32320
rect 12584 32308 12590 32360
rect 13722 32308 13728 32360
rect 13780 32348 13786 32360
rect 14458 32348 14464 32360
rect 13780 32320 14464 32348
rect 13780 32308 13786 32320
rect 14458 32308 14464 32320
rect 14516 32308 14522 32360
rect 14550 32308 14556 32360
rect 14608 32308 14614 32360
rect 15930 32308 15936 32360
rect 15988 32308 15994 32360
rect 17052 32357 17080 32388
rect 18874 32376 18880 32388
rect 18932 32376 18938 32428
rect 19705 32419 19763 32425
rect 19705 32385 19717 32419
rect 19751 32416 19763 32419
rect 19978 32416 19984 32428
rect 19751 32388 19984 32416
rect 19751 32385 19763 32388
rect 19705 32379 19763 32385
rect 19978 32376 19984 32388
rect 20036 32376 20042 32428
rect 22020 32425 22048 32456
rect 22005 32419 22063 32425
rect 22005 32385 22017 32419
rect 22051 32385 22063 32419
rect 22005 32379 22063 32385
rect 17037 32351 17095 32357
rect 17037 32317 17049 32351
rect 17083 32317 17095 32351
rect 17037 32311 17095 32317
rect 17129 32351 17187 32357
rect 17129 32317 17141 32351
rect 17175 32317 17187 32351
rect 18601 32351 18659 32357
rect 18601 32348 18613 32351
rect 17129 32311 17187 32317
rect 17236 32320 18613 32348
rect 6914 32240 6920 32292
rect 6972 32280 6978 32292
rect 7760 32280 7788 32308
rect 14568 32280 14596 32308
rect 6972 32252 7788 32280
rect 10888 32252 14596 32280
rect 6972 32240 6978 32252
rect 1765 32215 1823 32221
rect 1765 32181 1777 32215
rect 1811 32212 1823 32215
rect 2590 32212 2596 32224
rect 1811 32184 2596 32212
rect 1811 32181 1823 32184
rect 1765 32175 1823 32181
rect 2590 32172 2596 32184
rect 2648 32172 2654 32224
rect 9582 32172 9588 32224
rect 9640 32212 9646 32224
rect 10888 32221 10916 32252
rect 16942 32240 16948 32292
rect 17000 32280 17006 32292
rect 17144 32280 17172 32311
rect 17000 32252 17172 32280
rect 17000 32240 17006 32252
rect 10873 32215 10931 32221
rect 10873 32212 10885 32215
rect 9640 32184 10885 32212
rect 9640 32172 9646 32184
rect 10873 32181 10885 32184
rect 10919 32181 10931 32215
rect 10873 32175 10931 32181
rect 11790 32172 11796 32224
rect 11848 32212 11854 32224
rect 12710 32212 12716 32224
rect 11848 32184 12716 32212
rect 11848 32172 11854 32184
rect 12710 32172 12716 32184
rect 12768 32172 12774 32224
rect 14461 32215 14519 32221
rect 14461 32181 14473 32215
rect 14507 32212 14519 32215
rect 14550 32212 14556 32224
rect 14507 32184 14556 32212
rect 14507 32181 14519 32184
rect 14461 32175 14519 32181
rect 14550 32172 14556 32184
rect 14608 32212 14614 32224
rect 17236 32212 17264 32320
rect 18601 32317 18613 32320
rect 18647 32317 18659 32351
rect 18601 32311 18659 32317
rect 19797 32351 19855 32357
rect 19797 32317 19809 32351
rect 19843 32317 19855 32351
rect 19797 32311 19855 32317
rect 17310 32240 17316 32292
rect 17368 32280 17374 32292
rect 17368 32252 17724 32280
rect 17368 32240 17374 32252
rect 14608 32184 17264 32212
rect 14608 32172 14614 32184
rect 17586 32172 17592 32224
rect 17644 32172 17650 32224
rect 17696 32212 17724 32252
rect 17862 32240 17868 32292
rect 17920 32280 17926 32292
rect 19245 32283 19303 32289
rect 19245 32280 19257 32283
rect 17920 32252 19257 32280
rect 17920 32240 17926 32252
rect 19245 32249 19257 32252
rect 19291 32249 19303 32283
rect 19245 32243 19303 32249
rect 19812 32212 19840 32311
rect 21174 32308 21180 32360
rect 21232 32308 21238 32360
rect 22370 32308 22376 32360
rect 22428 32348 22434 32360
rect 22848 32348 22876 32524
rect 25130 32512 25136 32524
rect 25188 32512 25194 32564
rect 22922 32444 22928 32496
rect 22980 32484 22986 32496
rect 22980 32456 23888 32484
rect 22980 32444 22986 32456
rect 23017 32419 23075 32425
rect 23017 32385 23029 32419
rect 23063 32416 23075 32419
rect 23290 32416 23296 32428
rect 23063 32388 23296 32416
rect 23063 32385 23075 32388
rect 23017 32379 23075 32385
rect 23290 32376 23296 32388
rect 23348 32376 23354 32428
rect 23860 32425 23888 32456
rect 23845 32419 23903 32425
rect 23845 32385 23857 32419
rect 23891 32385 23903 32419
rect 23845 32379 23903 32385
rect 24857 32419 24915 32425
rect 24857 32385 24869 32419
rect 24903 32416 24915 32419
rect 25314 32416 25320 32428
rect 24903 32388 25320 32416
rect 24903 32385 24915 32388
rect 24857 32379 24915 32385
rect 25314 32376 25320 32388
rect 25372 32376 25378 32428
rect 23109 32351 23167 32357
rect 23109 32348 23121 32351
rect 22428 32320 23121 32348
rect 22428 32308 22434 32320
rect 23109 32317 23121 32320
rect 23155 32317 23167 32351
rect 23109 32311 23167 32317
rect 23198 32308 23204 32360
rect 23256 32308 23262 32360
rect 19978 32240 19984 32292
rect 20036 32280 20042 32292
rect 25133 32283 25191 32289
rect 25133 32280 25145 32283
rect 20036 32252 25145 32280
rect 20036 32240 20042 32252
rect 25133 32249 25145 32252
rect 25179 32249 25191 32283
rect 25133 32243 25191 32249
rect 17696 32184 19840 32212
rect 20622 32172 20628 32224
rect 20680 32172 20686 32224
rect 22189 32215 22247 32221
rect 22189 32181 22201 32215
rect 22235 32212 22247 32215
rect 23934 32212 23940 32224
rect 22235 32184 23940 32212
rect 22235 32181 22247 32184
rect 22189 32175 22247 32181
rect 23934 32172 23940 32184
rect 23992 32172 23998 32224
rect 24029 32215 24087 32221
rect 24029 32181 24041 32215
rect 24075 32212 24087 32215
rect 24486 32212 24492 32224
rect 24075 32184 24492 32212
rect 24075 32181 24087 32184
rect 24029 32175 24087 32181
rect 24486 32172 24492 32184
rect 24544 32172 24550 32224
rect 1104 32122 25852 32144
rect 1104 32070 2950 32122
rect 3002 32070 3014 32122
rect 3066 32070 3078 32122
rect 3130 32070 3142 32122
rect 3194 32070 3206 32122
rect 3258 32070 12950 32122
rect 13002 32070 13014 32122
rect 13066 32070 13078 32122
rect 13130 32070 13142 32122
rect 13194 32070 13206 32122
rect 13258 32070 22950 32122
rect 23002 32070 23014 32122
rect 23066 32070 23078 32122
rect 23130 32070 23142 32122
rect 23194 32070 23206 32122
rect 23258 32070 25852 32122
rect 1104 32048 25852 32070
rect 5169 32011 5227 32017
rect 5169 31977 5181 32011
rect 5215 32008 5227 32011
rect 6086 32008 6092 32020
rect 5215 31980 6092 32008
rect 5215 31977 5227 31980
rect 5169 31971 5227 31977
rect 6086 31968 6092 31980
rect 6144 31968 6150 32020
rect 7282 31968 7288 32020
rect 7340 32008 7346 32020
rect 10778 32008 10784 32020
rect 7340 31980 10784 32008
rect 7340 31968 7346 31980
rect 10778 31968 10784 31980
rect 10836 31968 10842 32020
rect 11238 31968 11244 32020
rect 11296 31968 11302 32020
rect 12342 31968 12348 32020
rect 12400 31968 12406 32020
rect 15197 32011 15255 32017
rect 15197 31977 15209 32011
rect 15243 32008 15255 32011
rect 15930 32008 15936 32020
rect 15243 31980 15936 32008
rect 15243 31977 15255 31980
rect 15197 31971 15255 31977
rect 15930 31968 15936 31980
rect 15988 32008 15994 32020
rect 15988 31980 17632 32008
rect 15988 31968 15994 31980
rect 7834 31900 7840 31952
rect 7892 31940 7898 31952
rect 8205 31943 8263 31949
rect 8205 31940 8217 31943
rect 7892 31912 8217 31940
rect 7892 31900 7898 31912
rect 8205 31909 8217 31912
rect 8251 31909 8263 31943
rect 17604 31940 17632 31980
rect 17678 31968 17684 32020
rect 17736 31968 17742 32020
rect 19794 32008 19800 32020
rect 19628 31980 19800 32008
rect 19242 31940 19248 31952
rect 8205 31903 8263 31909
rect 16868 31912 17540 31940
rect 17604 31912 19248 31940
rect 6641 31875 6699 31881
rect 6641 31841 6653 31875
rect 6687 31872 6699 31875
rect 7653 31875 7711 31881
rect 7653 31872 7665 31875
rect 6687 31844 7665 31872
rect 6687 31841 6699 31844
rect 6641 31835 6699 31841
rect 7576 31816 7604 31844
rect 7653 31841 7665 31844
rect 7699 31872 7711 31875
rect 8294 31872 8300 31884
rect 7699 31844 8300 31872
rect 7699 31841 7711 31844
rect 7653 31835 7711 31841
rect 8294 31832 8300 31844
rect 8352 31832 8358 31884
rect 9125 31875 9183 31881
rect 9125 31841 9137 31875
rect 9171 31872 9183 31875
rect 9214 31872 9220 31884
rect 9171 31844 9220 31872
rect 9171 31841 9183 31844
rect 9125 31835 9183 31841
rect 9214 31832 9220 31844
rect 9272 31832 9278 31884
rect 11606 31832 11612 31884
rect 11664 31872 11670 31884
rect 12897 31875 12955 31881
rect 12897 31872 12909 31875
rect 11664 31844 12909 31872
rect 11664 31832 11670 31844
rect 12897 31841 12909 31844
rect 12943 31841 12955 31875
rect 16868 31872 16896 31912
rect 12897 31835 12955 31841
rect 15488 31844 16896 31872
rect 6914 31764 6920 31816
rect 6972 31764 6978 31816
rect 7558 31764 7564 31816
rect 7616 31764 7622 31816
rect 7745 31807 7803 31813
rect 7745 31773 7757 31807
rect 7791 31804 7803 31807
rect 9030 31804 9036 31816
rect 7791 31776 9036 31804
rect 7791 31773 7803 31776
rect 7745 31767 7803 31773
rect 9030 31764 9036 31776
rect 9088 31764 9094 31816
rect 9490 31764 9496 31816
rect 9548 31764 9554 31816
rect 10873 31807 10931 31813
rect 10873 31773 10885 31807
rect 10919 31804 10931 31807
rect 10962 31804 10968 31816
rect 10919 31776 10968 31804
rect 10919 31773 10931 31776
rect 10873 31767 10931 31773
rect 10962 31764 10968 31776
rect 11020 31764 11026 31816
rect 12069 31807 12127 31813
rect 12069 31773 12081 31807
rect 12115 31804 12127 31807
rect 12805 31807 12863 31813
rect 12115 31776 12756 31804
rect 12115 31773 12127 31776
rect 12069 31767 12127 31773
rect 12728 31748 12756 31776
rect 12805 31773 12817 31807
rect 12851 31804 12863 31807
rect 15488 31804 15516 31844
rect 16942 31832 16948 31884
rect 17000 31832 17006 31884
rect 17034 31832 17040 31884
rect 17092 31872 17098 31884
rect 17405 31875 17463 31881
rect 17405 31872 17417 31875
rect 17092 31844 17417 31872
rect 17092 31832 17098 31844
rect 17405 31841 17417 31844
rect 17451 31841 17463 31875
rect 17405 31835 17463 31841
rect 12851 31776 15516 31804
rect 17512 31804 17540 31912
rect 19242 31900 19248 31912
rect 19300 31900 19306 31952
rect 19628 31804 19656 31980
rect 19794 31968 19800 31980
rect 19852 32008 19858 32020
rect 19978 32008 19984 32020
rect 19852 31980 19984 32008
rect 19852 31968 19858 31980
rect 19978 31968 19984 31980
rect 20036 31968 20042 32020
rect 20257 32011 20315 32017
rect 20257 31977 20269 32011
rect 20303 32008 20315 32011
rect 20438 32008 20444 32020
rect 20303 31980 20444 32008
rect 20303 31977 20315 31980
rect 20257 31971 20315 31977
rect 20438 31968 20444 31980
rect 20496 31968 20502 32020
rect 20714 31968 20720 32020
rect 20772 32008 20778 32020
rect 25133 32011 25191 32017
rect 25133 32008 25145 32011
rect 20772 31980 25145 32008
rect 20772 31968 20778 31980
rect 25133 31977 25145 31980
rect 25179 31977 25191 32011
rect 25133 31971 25191 31977
rect 21082 31940 21088 31952
rect 19720 31912 21088 31940
rect 19720 31881 19748 31912
rect 21082 31900 21088 31912
rect 21140 31900 21146 31952
rect 21453 31943 21511 31949
rect 21453 31909 21465 31943
rect 21499 31940 21511 31943
rect 22278 31940 22284 31952
rect 21499 31912 22284 31940
rect 21499 31909 21511 31912
rect 21453 31903 21511 31909
rect 22278 31900 22284 31912
rect 22336 31900 22342 31952
rect 22370 31900 22376 31952
rect 22428 31940 22434 31952
rect 22649 31943 22707 31949
rect 22649 31940 22661 31943
rect 22428 31912 22661 31940
rect 22428 31900 22434 31912
rect 22649 31909 22661 31912
rect 22695 31909 22707 31943
rect 22649 31903 22707 31909
rect 22738 31900 22744 31952
rect 22796 31940 22802 31952
rect 23382 31940 23388 31952
rect 22796 31912 23388 31940
rect 22796 31900 22802 31912
rect 23382 31900 23388 31912
rect 23440 31900 23446 31952
rect 23845 31943 23903 31949
rect 23845 31909 23857 31943
rect 23891 31940 23903 31943
rect 25590 31940 25596 31952
rect 23891 31912 25596 31940
rect 23891 31909 23903 31912
rect 23845 31903 23903 31909
rect 19705 31875 19763 31881
rect 19705 31841 19717 31875
rect 19751 31841 19763 31875
rect 19705 31835 19763 31841
rect 19797 31875 19855 31881
rect 19797 31841 19809 31875
rect 19843 31872 19855 31875
rect 19843 31844 19932 31872
rect 19843 31841 19855 31844
rect 19797 31835 19855 31841
rect 17512 31776 19656 31804
rect 12851 31773 12863 31776
rect 12805 31767 12863 31773
rect 7098 31736 7104 31748
rect 6210 31708 7104 31736
rect 7098 31696 7104 31708
rect 7156 31696 7162 31748
rect 10594 31696 10600 31748
rect 10652 31696 10658 31748
rect 12710 31736 12716 31748
rect 12671 31708 12716 31736
rect 12710 31696 12716 31708
rect 12768 31736 12774 31748
rect 13722 31736 13728 31748
rect 12768 31708 13728 31736
rect 12768 31696 12774 31708
rect 13722 31696 13728 31708
rect 13780 31696 13786 31748
rect 16206 31696 16212 31748
rect 16264 31696 16270 31748
rect 16666 31696 16672 31748
rect 16724 31696 16730 31748
rect 17313 31739 17371 31745
rect 17313 31705 17325 31739
rect 17359 31736 17371 31739
rect 18322 31736 18328 31748
rect 17359 31708 18328 31736
rect 17359 31705 17371 31708
rect 17313 31699 17371 31705
rect 18322 31696 18328 31708
rect 18380 31696 18386 31748
rect 19904 31736 19932 31844
rect 20346 31832 20352 31884
rect 20404 31872 20410 31884
rect 20809 31875 20867 31881
rect 20809 31872 20821 31875
rect 20404 31844 20821 31872
rect 20404 31832 20410 31844
rect 20809 31841 20821 31844
rect 20855 31872 20867 31875
rect 22005 31875 22063 31881
rect 22005 31872 22017 31875
rect 20855 31844 22017 31872
rect 20855 31841 20867 31844
rect 20809 31835 20867 31841
rect 22005 31841 22017 31844
rect 22051 31872 22063 31875
rect 22462 31872 22468 31884
rect 22051 31844 22468 31872
rect 22051 31841 22063 31844
rect 22005 31835 22063 31841
rect 22462 31832 22468 31844
rect 22520 31832 22526 31884
rect 23109 31875 23167 31881
rect 23109 31841 23121 31875
rect 23155 31872 23167 31875
rect 23290 31872 23296 31884
rect 23155 31844 23296 31872
rect 23155 31841 23167 31844
rect 23109 31835 23167 31841
rect 23290 31832 23296 31844
rect 23348 31832 23354 31884
rect 22186 31764 22192 31816
rect 22244 31804 22250 31816
rect 22738 31804 22744 31816
rect 22244 31776 22744 31804
rect 22244 31764 22250 31776
rect 22738 31764 22744 31776
rect 22796 31804 22802 31816
rect 23569 31807 23627 31813
rect 23569 31804 23581 31807
rect 22796 31776 23581 31804
rect 22796 31764 22802 31776
rect 23569 31773 23581 31776
rect 23615 31773 23627 31807
rect 23569 31767 23627 31773
rect 20438 31736 20444 31748
rect 19904 31708 20444 31736
rect 20438 31696 20444 31708
rect 20496 31736 20502 31748
rect 22281 31739 22339 31745
rect 22281 31736 22293 31739
rect 20496 31708 22293 31736
rect 20496 31696 20502 31708
rect 22281 31705 22293 31708
rect 22327 31736 22339 31739
rect 23860 31736 23888 31903
rect 25590 31900 25596 31912
rect 25648 31900 25654 31952
rect 24857 31807 24915 31813
rect 24857 31773 24869 31807
rect 24903 31804 24915 31807
rect 25317 31807 25375 31813
rect 25317 31804 25329 31807
rect 24903 31776 25329 31804
rect 24903 31773 24915 31776
rect 24857 31767 24915 31773
rect 25317 31773 25329 31776
rect 25363 31804 25375 31807
rect 25406 31804 25412 31816
rect 25363 31776 25412 31804
rect 25363 31773 25375 31776
rect 25317 31767 25375 31773
rect 25406 31764 25412 31776
rect 25464 31764 25470 31816
rect 22327 31708 23888 31736
rect 22327 31705 22339 31708
rect 22281 31699 22339 31705
rect 7834 31628 7840 31680
rect 7892 31628 7898 31680
rect 9950 31628 9956 31680
rect 10008 31668 10014 31680
rect 10612 31668 10640 31696
rect 10008 31640 10640 31668
rect 10008 31628 10014 31640
rect 14458 31628 14464 31680
rect 14516 31668 14522 31680
rect 18969 31671 19027 31677
rect 18969 31668 18981 31671
rect 14516 31640 18981 31668
rect 14516 31628 14522 31640
rect 18969 31637 18981 31640
rect 19015 31668 19027 31671
rect 19610 31668 19616 31680
rect 19015 31640 19616 31668
rect 19015 31637 19027 31640
rect 18969 31631 19027 31637
rect 19610 31628 19616 31640
rect 19668 31628 19674 31680
rect 19886 31628 19892 31680
rect 19944 31628 19950 31680
rect 20898 31628 20904 31680
rect 20956 31668 20962 31680
rect 20993 31671 21051 31677
rect 20993 31668 21005 31671
rect 20956 31640 21005 31668
rect 20956 31628 20962 31640
rect 20993 31637 21005 31640
rect 21039 31637 21051 31671
rect 20993 31631 21051 31637
rect 21085 31671 21143 31677
rect 21085 31637 21097 31671
rect 21131 31668 21143 31671
rect 21174 31668 21180 31680
rect 21131 31640 21180 31668
rect 21131 31637 21143 31640
rect 21085 31631 21143 31637
rect 21174 31628 21180 31640
rect 21232 31668 21238 31680
rect 21358 31668 21364 31680
rect 21232 31640 21364 31668
rect 21232 31628 21238 31640
rect 21358 31628 21364 31640
rect 21416 31628 21422 31680
rect 1104 31578 25852 31600
rect 1104 31526 7950 31578
rect 8002 31526 8014 31578
rect 8066 31526 8078 31578
rect 8130 31526 8142 31578
rect 8194 31526 8206 31578
rect 8258 31526 17950 31578
rect 18002 31526 18014 31578
rect 18066 31526 18078 31578
rect 18130 31526 18142 31578
rect 18194 31526 18206 31578
rect 18258 31526 25852 31578
rect 1104 31504 25852 31526
rect 4893 31467 4951 31473
rect 4893 31433 4905 31467
rect 4939 31464 4951 31467
rect 4982 31464 4988 31476
rect 4939 31436 4988 31464
rect 4939 31433 4951 31436
rect 4893 31427 4951 31433
rect 4982 31424 4988 31436
rect 5040 31424 5046 31476
rect 5261 31467 5319 31473
rect 5261 31433 5273 31467
rect 5307 31464 5319 31467
rect 5350 31464 5356 31476
rect 5307 31436 5356 31464
rect 5307 31433 5319 31436
rect 5261 31427 5319 31433
rect 5350 31424 5356 31436
rect 5408 31424 5414 31476
rect 7650 31424 7656 31476
rect 7708 31464 7714 31476
rect 7745 31467 7803 31473
rect 7745 31464 7757 31467
rect 7708 31436 7757 31464
rect 7708 31424 7714 31436
rect 7745 31433 7757 31436
rect 7791 31433 7803 31467
rect 7745 31427 7803 31433
rect 7834 31424 7840 31476
rect 7892 31464 7898 31476
rect 8205 31467 8263 31473
rect 8205 31464 8217 31467
rect 7892 31436 8217 31464
rect 7892 31424 7898 31436
rect 8205 31433 8217 31436
rect 8251 31433 8263 31467
rect 8205 31427 8263 31433
rect 9858 31424 9864 31476
rect 9916 31464 9922 31476
rect 10137 31467 10195 31473
rect 10137 31464 10149 31467
rect 9916 31436 10149 31464
rect 9916 31424 9922 31436
rect 10137 31433 10149 31436
rect 10183 31433 10195 31467
rect 10137 31427 10195 31433
rect 10226 31424 10232 31476
rect 10284 31464 10290 31476
rect 10502 31464 10508 31476
rect 10284 31436 10508 31464
rect 10284 31424 10290 31436
rect 10502 31424 10508 31436
rect 10560 31424 10566 31476
rect 10594 31424 10600 31476
rect 10652 31464 10658 31476
rect 15378 31464 15384 31476
rect 10652 31436 15384 31464
rect 10652 31424 10658 31436
rect 15378 31424 15384 31436
rect 15436 31464 15442 31476
rect 16850 31464 16856 31476
rect 15436 31436 16856 31464
rect 15436 31424 15442 31436
rect 16850 31424 16856 31436
rect 16908 31424 16914 31476
rect 17586 31424 17592 31476
rect 17644 31464 17650 31476
rect 17681 31467 17739 31473
rect 17681 31464 17693 31467
rect 17644 31436 17693 31464
rect 17644 31424 17650 31436
rect 17681 31433 17693 31436
rect 17727 31433 17739 31467
rect 17681 31427 17739 31433
rect 19610 31424 19616 31476
rect 19668 31464 19674 31476
rect 19886 31464 19892 31476
rect 19668 31436 19892 31464
rect 19668 31424 19674 31436
rect 19886 31424 19892 31436
rect 19944 31424 19950 31476
rect 20438 31424 20444 31476
rect 20496 31424 20502 31476
rect 20990 31424 20996 31476
rect 21048 31464 21054 31476
rect 23290 31464 23296 31476
rect 21048 31436 23296 31464
rect 21048 31424 21054 31436
rect 23290 31424 23296 31436
rect 23348 31424 23354 31476
rect 24213 31467 24271 31473
rect 24213 31433 24225 31467
rect 24259 31464 24271 31467
rect 24854 31464 24860 31476
rect 24259 31436 24860 31464
rect 24259 31433 24271 31436
rect 24213 31427 24271 31433
rect 24854 31424 24860 31436
rect 24912 31424 24918 31476
rect 17402 31356 17408 31408
rect 17460 31396 17466 31408
rect 17460 31368 19472 31396
rect 17460 31356 17466 31368
rect 6733 31331 6791 31337
rect 6733 31297 6745 31331
rect 6779 31328 6791 31331
rect 6822 31328 6828 31340
rect 6779 31300 6828 31328
rect 6779 31297 6791 31300
rect 6733 31291 6791 31297
rect 6822 31288 6828 31300
rect 6880 31328 6886 31340
rect 7098 31328 7104 31340
rect 6880 31300 7104 31328
rect 6880 31288 6886 31300
rect 7098 31288 7104 31300
rect 7156 31328 7162 31340
rect 7285 31331 7343 31337
rect 7285 31328 7297 31331
rect 7156 31300 7297 31328
rect 7156 31288 7162 31300
rect 7285 31297 7297 31300
rect 7331 31297 7343 31331
rect 7285 31291 7343 31297
rect 7377 31331 7435 31337
rect 7377 31297 7389 31331
rect 7423 31328 7435 31331
rect 8849 31331 8907 31337
rect 8849 31328 8861 31331
rect 7423 31300 8861 31328
rect 7423 31297 7435 31300
rect 7377 31291 7435 31297
rect 8849 31297 8861 31300
rect 8895 31297 8907 31331
rect 8849 31291 8907 31297
rect 10042 31288 10048 31340
rect 10100 31328 10106 31340
rect 10505 31331 10563 31337
rect 10505 31328 10517 31331
rect 10100 31300 10517 31328
rect 10100 31288 10106 31300
rect 10505 31297 10517 31300
rect 10551 31297 10563 31331
rect 10505 31291 10563 31297
rect 11238 31288 11244 31340
rect 11296 31328 11302 31340
rect 12250 31328 12256 31340
rect 11296 31300 12256 31328
rect 11296 31288 11302 31300
rect 12250 31288 12256 31300
rect 12308 31328 12314 31340
rect 12529 31331 12587 31337
rect 12529 31328 12541 31331
rect 12308 31300 12541 31328
rect 12308 31288 12314 31300
rect 12529 31297 12541 31300
rect 12575 31297 12587 31331
rect 12529 31291 12587 31297
rect 17589 31331 17647 31337
rect 17589 31297 17601 31331
rect 17635 31328 17647 31331
rect 18690 31328 18696 31340
rect 17635 31300 18696 31328
rect 17635 31297 17647 31300
rect 17589 31291 17647 31297
rect 18690 31288 18696 31300
rect 18748 31288 18754 31340
rect 19444 31337 19472 31368
rect 19429 31331 19487 31337
rect 19429 31297 19441 31331
rect 19475 31297 19487 31331
rect 19429 31291 19487 31297
rect 20530 31288 20536 31340
rect 20588 31328 20594 31340
rect 22005 31331 22063 31337
rect 22005 31328 22017 31331
rect 20588 31300 22017 31328
rect 20588 31288 20594 31300
rect 22005 31297 22017 31300
rect 22051 31297 22063 31331
rect 22005 31291 22063 31297
rect 23382 31288 23388 31340
rect 23440 31288 23446 31340
rect 25314 31288 25320 31340
rect 25372 31288 25378 31340
rect 4706 31220 4712 31272
rect 4764 31220 4770 31272
rect 4798 31220 4804 31272
rect 4856 31220 4862 31272
rect 7193 31263 7251 31269
rect 7193 31229 7205 31263
rect 7239 31229 7251 31263
rect 7193 31223 7251 31229
rect 4154 31152 4160 31204
rect 4212 31192 4218 31204
rect 4249 31195 4307 31201
rect 4249 31192 4261 31195
rect 4212 31164 4261 31192
rect 4212 31152 4218 31164
rect 4249 31161 4261 31164
rect 4295 31192 4307 31195
rect 4816 31192 4844 31220
rect 4295 31164 4844 31192
rect 7208 31192 7236 31223
rect 9858 31220 9864 31272
rect 9916 31260 9922 31272
rect 10594 31260 10600 31272
rect 9916 31232 10600 31260
rect 9916 31220 9922 31232
rect 10594 31220 10600 31232
rect 10652 31220 10658 31272
rect 10781 31263 10839 31269
rect 10781 31229 10793 31263
rect 10827 31260 10839 31263
rect 10870 31260 10876 31272
rect 10827 31232 10876 31260
rect 10827 31229 10839 31232
rect 10781 31223 10839 31229
rect 10870 31220 10876 31232
rect 10928 31220 10934 31272
rect 17770 31220 17776 31272
rect 17828 31220 17834 31272
rect 18046 31220 18052 31272
rect 18104 31260 18110 31272
rect 25041 31263 25099 31269
rect 25041 31260 25053 31263
rect 18104 31232 25053 31260
rect 18104 31220 18110 31232
rect 25041 31229 25053 31232
rect 25087 31229 25099 31263
rect 25041 31223 25099 31229
rect 7374 31192 7380 31204
rect 7208 31164 7380 31192
rect 4295 31161 4307 31164
rect 4249 31155 4307 31161
rect 7374 31152 7380 31164
rect 7432 31152 7438 31204
rect 19613 31195 19671 31201
rect 19613 31161 19625 31195
rect 19659 31192 19671 31195
rect 21266 31192 21272 31204
rect 19659 31164 21272 31192
rect 19659 31161 19671 31164
rect 19613 31155 19671 31161
rect 21266 31152 21272 31164
rect 21324 31152 21330 31204
rect 21358 31152 21364 31204
rect 21416 31192 21422 31204
rect 22465 31195 22523 31201
rect 22465 31192 22477 31195
rect 21416 31164 22477 31192
rect 21416 31152 21422 31164
rect 22465 31161 22477 31164
rect 22511 31161 22523 31195
rect 22465 31155 22523 31161
rect 23569 31195 23627 31201
rect 23569 31161 23581 31195
rect 23615 31192 23627 31195
rect 24302 31192 24308 31204
rect 23615 31164 24308 31192
rect 23615 31161 23627 31164
rect 23569 31155 23627 31161
rect 24302 31152 24308 31164
rect 24360 31152 24366 31204
rect 6362 31084 6368 31136
rect 6420 31124 6426 31136
rect 9677 31127 9735 31133
rect 9677 31124 9689 31127
rect 6420 31096 9689 31124
rect 6420 31084 6426 31096
rect 9677 31093 9689 31096
rect 9723 31124 9735 31127
rect 10042 31124 10048 31136
rect 9723 31096 10048 31124
rect 9723 31093 9735 31096
rect 9677 31087 9735 31093
rect 10042 31084 10048 31096
rect 10100 31084 10106 31136
rect 12526 31084 12532 31136
rect 12584 31124 12590 31136
rect 12897 31127 12955 31133
rect 12897 31124 12909 31127
rect 12584 31096 12909 31124
rect 12584 31084 12590 31096
rect 12897 31093 12909 31096
rect 12943 31124 12955 31127
rect 13354 31124 13360 31136
rect 12943 31096 13360 31124
rect 12943 31093 12955 31096
rect 12897 31087 12955 31093
rect 13354 31084 13360 31096
rect 13412 31084 13418 31136
rect 17218 31084 17224 31136
rect 17276 31084 17282 31136
rect 20898 31084 20904 31136
rect 20956 31124 20962 31136
rect 21545 31127 21603 31133
rect 21545 31124 21557 31127
rect 20956 31096 21557 31124
rect 20956 31084 20962 31096
rect 21545 31093 21557 31096
rect 21591 31124 21603 31127
rect 21634 31124 21640 31136
rect 21591 31096 21640 31124
rect 21591 31093 21603 31096
rect 21545 31087 21603 31093
rect 21634 31084 21640 31096
rect 21692 31084 21698 31136
rect 22189 31127 22247 31133
rect 22189 31093 22201 31127
rect 22235 31124 22247 31127
rect 25038 31124 25044 31136
rect 22235 31096 25044 31124
rect 22235 31093 22247 31096
rect 22189 31087 22247 31093
rect 25038 31084 25044 31096
rect 25096 31084 25102 31136
rect 1104 31034 25852 31056
rect 1104 30982 2950 31034
rect 3002 30982 3014 31034
rect 3066 30982 3078 31034
rect 3130 30982 3142 31034
rect 3194 30982 3206 31034
rect 3258 30982 12950 31034
rect 13002 30982 13014 31034
rect 13066 30982 13078 31034
rect 13130 30982 13142 31034
rect 13194 30982 13206 31034
rect 13258 30982 22950 31034
rect 23002 30982 23014 31034
rect 23066 30982 23078 31034
rect 23130 30982 23142 31034
rect 23194 30982 23206 31034
rect 23258 30982 25852 31034
rect 1104 30960 25852 30982
rect 7742 30880 7748 30932
rect 7800 30920 7806 30932
rect 7837 30923 7895 30929
rect 7837 30920 7849 30923
rect 7800 30892 7849 30920
rect 7800 30880 7806 30892
rect 7837 30889 7849 30892
rect 7883 30889 7895 30923
rect 7837 30883 7895 30889
rect 10778 30880 10784 30932
rect 10836 30920 10842 30932
rect 10836 30892 12434 30920
rect 10836 30880 10842 30892
rect 7282 30744 7288 30796
rect 7340 30744 7346 30796
rect 10689 30787 10747 30793
rect 10689 30753 10701 30787
rect 10735 30784 10747 30787
rect 10962 30784 10968 30796
rect 10735 30756 10968 30784
rect 10735 30753 10747 30756
rect 10689 30747 10747 30753
rect 10962 30744 10968 30756
rect 11020 30784 11026 30796
rect 12406 30784 12434 30892
rect 12802 30880 12808 30932
rect 12860 30920 12866 30932
rect 12989 30923 13047 30929
rect 12989 30920 13001 30923
rect 12860 30892 13001 30920
rect 12860 30880 12866 30892
rect 12989 30889 13001 30892
rect 13035 30889 13047 30923
rect 12989 30883 13047 30889
rect 17402 30880 17408 30932
rect 17460 30920 17466 30932
rect 21174 30920 21180 30932
rect 17460 30892 21180 30920
rect 17460 30880 17466 30892
rect 21174 30880 21180 30892
rect 21232 30880 21238 30932
rect 24854 30880 24860 30932
rect 24912 30920 24918 30932
rect 25225 30923 25283 30929
rect 25225 30920 25237 30923
rect 24912 30892 25237 30920
rect 24912 30880 24918 30892
rect 25225 30889 25237 30892
rect 25271 30889 25283 30923
rect 25225 30883 25283 30889
rect 25314 30880 25320 30932
rect 25372 30920 25378 30932
rect 25409 30923 25467 30929
rect 25409 30920 25421 30923
rect 25372 30892 25421 30920
rect 25372 30880 25378 30892
rect 25409 30889 25421 30892
rect 25455 30889 25467 30923
rect 25409 30883 25467 30889
rect 16482 30812 16488 30864
rect 16540 30852 16546 30864
rect 17678 30852 17684 30864
rect 16540 30824 17684 30852
rect 16540 30812 16546 30824
rect 17678 30812 17684 30824
rect 17736 30812 17742 30864
rect 13541 30787 13599 30793
rect 13541 30784 13553 30787
rect 11020 30756 12204 30784
rect 12406 30756 13553 30784
rect 11020 30744 11026 30756
rect 7466 30676 7472 30728
rect 7524 30676 7530 30728
rect 12176 30716 12204 30756
rect 13541 30753 13553 30756
rect 13587 30753 13599 30787
rect 13541 30747 13599 30753
rect 13814 30744 13820 30796
rect 13872 30784 13878 30796
rect 16669 30787 16727 30793
rect 13872 30756 16528 30784
rect 13872 30744 13878 30756
rect 14274 30716 14280 30728
rect 12176 30688 14280 30716
rect 14274 30676 14280 30688
rect 14332 30676 14338 30728
rect 16500 30716 16528 30756
rect 16669 30753 16681 30787
rect 16715 30784 16727 30787
rect 16942 30784 16948 30796
rect 16715 30756 16948 30784
rect 16715 30753 16727 30756
rect 16669 30747 16727 30753
rect 16942 30744 16948 30756
rect 17000 30784 17006 30796
rect 17310 30784 17316 30796
rect 17000 30756 17316 30784
rect 17000 30744 17006 30756
rect 17310 30744 17316 30756
rect 17368 30744 17374 30796
rect 18138 30744 18144 30796
rect 18196 30744 18202 30796
rect 18322 30744 18328 30796
rect 18380 30744 18386 30796
rect 20714 30744 20720 30796
rect 20772 30784 20778 30796
rect 20993 30787 21051 30793
rect 20993 30784 21005 30787
rect 20772 30756 21005 30784
rect 20772 30744 20778 30756
rect 20993 30753 21005 30756
rect 21039 30753 21051 30787
rect 20993 30747 21051 30753
rect 22281 30787 22339 30793
rect 22281 30753 22293 30787
rect 22327 30784 22339 30787
rect 22554 30784 22560 30796
rect 22327 30756 22560 30784
rect 22327 30753 22339 30756
rect 22281 30747 22339 30753
rect 22554 30744 22560 30756
rect 22612 30744 22618 30796
rect 18046 30716 18052 30728
rect 16500 30688 18052 30716
rect 18046 30676 18052 30688
rect 18104 30676 18110 30728
rect 19613 30719 19671 30725
rect 19613 30685 19625 30719
rect 19659 30716 19671 30719
rect 19978 30716 19984 30728
rect 19659 30688 19984 30716
rect 19659 30685 19671 30688
rect 19613 30679 19671 30685
rect 19978 30676 19984 30688
rect 20036 30716 20042 30728
rect 20806 30716 20812 30728
rect 20036 30688 20812 30716
rect 20036 30676 20042 30688
rect 20806 30676 20812 30688
rect 20864 30676 20870 30728
rect 20901 30719 20959 30725
rect 20901 30685 20913 30719
rect 20947 30716 20959 30719
rect 21542 30716 21548 30728
rect 20947 30688 21548 30716
rect 20947 30685 20959 30688
rect 20901 30679 20959 30685
rect 21542 30676 21548 30688
rect 21600 30676 21606 30728
rect 24578 30676 24584 30728
rect 24636 30676 24642 30728
rect 10686 30608 10692 30660
rect 10744 30648 10750 30660
rect 10965 30651 11023 30657
rect 10965 30648 10977 30651
rect 10744 30620 10977 30648
rect 10744 30608 10750 30620
rect 10965 30617 10977 30620
rect 11011 30617 11023 30651
rect 12250 30648 12256 30660
rect 12190 30620 12256 30648
rect 10965 30611 11023 30617
rect 12250 30608 12256 30620
rect 12308 30608 12314 30660
rect 13354 30608 13360 30660
rect 13412 30648 13418 30660
rect 14458 30648 14464 30660
rect 13412 30620 14464 30648
rect 13412 30608 13418 30620
rect 14458 30608 14464 30620
rect 14516 30608 14522 30660
rect 14550 30608 14556 30660
rect 14608 30608 14614 30660
rect 16114 30648 16120 30660
rect 15778 30620 16120 30648
rect 16114 30608 16120 30620
rect 16172 30608 16178 30660
rect 16761 30651 16819 30657
rect 16761 30617 16773 30651
rect 16807 30648 16819 30651
rect 16807 30620 18828 30648
rect 16807 30617 16819 30620
rect 16761 30611 16819 30617
rect 6638 30540 6644 30592
rect 6696 30580 6702 30592
rect 6825 30583 6883 30589
rect 6825 30580 6837 30583
rect 6696 30552 6837 30580
rect 6696 30540 6702 30552
rect 6825 30549 6837 30552
rect 6871 30580 6883 30583
rect 7006 30580 7012 30592
rect 6871 30552 7012 30580
rect 6871 30549 6883 30552
rect 6825 30543 6883 30549
rect 7006 30540 7012 30552
rect 7064 30580 7070 30592
rect 7377 30583 7435 30589
rect 7377 30580 7389 30583
rect 7064 30552 7389 30580
rect 7064 30540 7070 30552
rect 7377 30549 7389 30552
rect 7423 30549 7435 30583
rect 7377 30543 7435 30549
rect 12437 30583 12495 30589
rect 12437 30549 12449 30583
rect 12483 30580 12495 30583
rect 12802 30580 12808 30592
rect 12483 30552 12808 30580
rect 12483 30549 12495 30552
rect 12437 30543 12495 30549
rect 12802 30540 12808 30552
rect 12860 30540 12866 30592
rect 13449 30583 13507 30589
rect 13449 30549 13461 30583
rect 13495 30580 13507 30583
rect 13538 30580 13544 30592
rect 13495 30552 13544 30580
rect 13495 30549 13507 30552
rect 13449 30543 13507 30549
rect 13538 30540 13544 30552
rect 13596 30540 13602 30592
rect 16022 30540 16028 30592
rect 16080 30540 16086 30592
rect 16298 30540 16304 30592
rect 16356 30580 16362 30592
rect 16853 30583 16911 30589
rect 16853 30580 16865 30583
rect 16356 30552 16865 30580
rect 16356 30540 16362 30552
rect 16853 30549 16865 30552
rect 16899 30549 16911 30583
rect 16853 30543 16911 30549
rect 17221 30583 17279 30589
rect 17221 30549 17233 30583
rect 17267 30580 17279 30583
rect 17310 30580 17316 30592
rect 17267 30552 17316 30580
rect 17267 30549 17279 30552
rect 17221 30543 17279 30549
rect 17310 30540 17316 30552
rect 17368 30540 17374 30592
rect 17678 30540 17684 30592
rect 17736 30540 17742 30592
rect 18800 30589 18828 30620
rect 22462 30608 22468 30660
rect 22520 30648 22526 30660
rect 22557 30651 22615 30657
rect 22557 30648 22569 30651
rect 22520 30620 22569 30648
rect 22520 30608 22526 30620
rect 22557 30617 22569 30620
rect 22603 30617 22615 30651
rect 24854 30648 24860 30660
rect 23782 30620 24860 30648
rect 22557 30611 22615 30617
rect 24854 30608 24860 30620
rect 24912 30608 24918 30660
rect 18785 30583 18843 30589
rect 18785 30549 18797 30583
rect 18831 30580 18843 30583
rect 18966 30580 18972 30592
rect 18831 30552 18972 30580
rect 18831 30549 18843 30552
rect 18785 30543 18843 30549
rect 18966 30540 18972 30552
rect 19024 30540 19030 30592
rect 19426 30540 19432 30592
rect 19484 30540 19490 30592
rect 19610 30540 19616 30592
rect 19668 30580 19674 30592
rect 20441 30583 20499 30589
rect 20441 30580 20453 30583
rect 19668 30552 20453 30580
rect 19668 30540 19674 30552
rect 20441 30549 20453 30552
rect 20487 30549 20499 30583
rect 20441 30543 20499 30549
rect 20806 30540 20812 30592
rect 20864 30580 20870 30592
rect 23474 30580 23480 30592
rect 20864 30552 23480 30580
rect 20864 30540 20870 30552
rect 23474 30540 23480 30552
rect 23532 30540 23538 30592
rect 23566 30540 23572 30592
rect 23624 30580 23630 30592
rect 24029 30583 24087 30589
rect 24029 30580 24041 30583
rect 23624 30552 24041 30580
rect 23624 30540 23630 30552
rect 24029 30549 24041 30552
rect 24075 30580 24087 30583
rect 24578 30580 24584 30592
rect 24075 30552 24584 30580
rect 24075 30549 24087 30552
rect 24029 30543 24087 30549
rect 24578 30540 24584 30552
rect 24636 30540 24642 30592
rect 24762 30540 24768 30592
rect 24820 30540 24826 30592
rect 1104 30490 25852 30512
rect 1104 30438 7950 30490
rect 8002 30438 8014 30490
rect 8066 30438 8078 30490
rect 8130 30438 8142 30490
rect 8194 30438 8206 30490
rect 8258 30438 17950 30490
rect 18002 30438 18014 30490
rect 18066 30438 18078 30490
rect 18130 30438 18142 30490
rect 18194 30438 18206 30490
rect 18258 30438 25852 30490
rect 1104 30416 25852 30438
rect 7558 30336 7564 30388
rect 7616 30376 7622 30388
rect 7653 30379 7711 30385
rect 7653 30376 7665 30379
rect 7616 30348 7665 30376
rect 7616 30336 7622 30348
rect 7653 30345 7665 30348
rect 7699 30345 7711 30379
rect 15289 30379 15347 30385
rect 7653 30339 7711 30345
rect 9048 30348 9536 30376
rect 9048 30308 9076 30348
rect 8694 30280 9076 30308
rect 9122 30268 9128 30320
rect 9180 30308 9186 30320
rect 9180 30280 9444 30308
rect 9180 30268 9186 30280
rect 9416 30249 9444 30280
rect 9508 30252 9536 30348
rect 15289 30345 15301 30379
rect 15335 30376 15347 30379
rect 15838 30376 15844 30388
rect 15335 30348 15844 30376
rect 15335 30345 15347 30348
rect 15289 30339 15347 30345
rect 15838 30336 15844 30348
rect 15896 30336 15902 30388
rect 16114 30336 16120 30388
rect 16172 30336 16178 30388
rect 16298 30336 16304 30388
rect 16356 30376 16362 30388
rect 16482 30376 16488 30388
rect 16356 30348 16488 30376
rect 16356 30336 16362 30348
rect 16482 30336 16488 30348
rect 16540 30336 16546 30388
rect 17313 30379 17371 30385
rect 17313 30345 17325 30379
rect 17359 30345 17371 30379
rect 17313 30339 17371 30345
rect 17681 30379 17739 30385
rect 17681 30345 17693 30379
rect 17727 30376 17739 30379
rect 17727 30348 18552 30376
rect 17727 30345 17739 30348
rect 17681 30339 17739 30345
rect 10226 30268 10232 30320
rect 10284 30308 10290 30320
rect 12253 30311 12311 30317
rect 12253 30308 12265 30311
rect 10284 30280 12265 30308
rect 10284 30268 10290 30280
rect 12253 30277 12265 30280
rect 12299 30308 12311 30311
rect 12986 30308 12992 30320
rect 12299 30280 12992 30308
rect 12299 30277 12311 30280
rect 12253 30271 12311 30277
rect 12986 30268 12992 30280
rect 13044 30268 13050 30320
rect 15654 30268 15660 30320
rect 15712 30308 15718 30320
rect 17328 30308 17356 30339
rect 18524 30320 18552 30348
rect 19426 30336 19432 30388
rect 19484 30376 19490 30388
rect 20073 30379 20131 30385
rect 20073 30376 20085 30379
rect 19484 30348 20085 30376
rect 19484 30336 19490 30348
rect 20073 30345 20085 30348
rect 20119 30345 20131 30379
rect 24854 30376 24860 30388
rect 20073 30339 20131 30345
rect 22204 30348 22508 30376
rect 15712 30280 17356 30308
rect 15712 30268 15718 30280
rect 18506 30268 18512 30320
rect 18564 30268 18570 30320
rect 18969 30311 19027 30317
rect 18969 30277 18981 30311
rect 19015 30308 19027 30311
rect 22204 30308 22232 30348
rect 19015 30280 22232 30308
rect 19015 30277 19027 30280
rect 18969 30271 19027 30277
rect 22278 30268 22284 30320
rect 22336 30268 22342 30320
rect 22370 30268 22376 30320
rect 22428 30268 22434 30320
rect 22480 30308 22508 30348
rect 24596 30348 24860 30376
rect 23658 30308 23664 30320
rect 22480 30280 23664 30308
rect 23658 30268 23664 30280
rect 23716 30268 23722 30320
rect 24596 30308 24624 30348
rect 24854 30336 24860 30348
rect 24912 30336 24918 30388
rect 24518 30280 24624 30308
rect 9401 30243 9459 30249
rect 9401 30209 9413 30243
rect 9447 30209 9459 30243
rect 9401 30203 9459 30209
rect 9490 30200 9496 30252
rect 9548 30240 9554 30252
rect 9769 30243 9827 30249
rect 9769 30240 9781 30243
rect 9548 30212 9781 30240
rect 9548 30200 9554 30212
rect 9769 30209 9781 30212
rect 9815 30240 9827 30243
rect 11238 30240 11244 30252
rect 9815 30212 11244 30240
rect 9815 30209 9827 30212
rect 9769 30203 9827 30209
rect 11238 30200 11244 30212
rect 11296 30200 11302 30252
rect 13081 30243 13139 30249
rect 13081 30209 13093 30243
rect 13127 30240 13139 30243
rect 15010 30240 15016 30252
rect 13127 30212 15016 30240
rect 13127 30209 13139 30212
rect 13081 30203 13139 30209
rect 15010 30200 15016 30212
rect 15068 30200 15074 30252
rect 15197 30243 15255 30249
rect 15197 30209 15209 30243
rect 15243 30240 15255 30243
rect 16574 30240 16580 30252
rect 15243 30212 15516 30240
rect 15243 30209 15255 30212
rect 15197 30203 15255 30209
rect 9125 30175 9183 30181
rect 9125 30141 9137 30175
rect 9171 30172 9183 30175
rect 9582 30172 9588 30184
rect 9171 30144 9588 30172
rect 9171 30141 9183 30144
rect 9125 30135 9183 30141
rect 9582 30132 9588 30144
rect 9640 30132 9646 30184
rect 10962 30132 10968 30184
rect 11020 30172 11026 30184
rect 11701 30175 11759 30181
rect 11701 30172 11713 30175
rect 11020 30144 11713 30172
rect 11020 30132 11026 30144
rect 11701 30141 11713 30144
rect 11747 30141 11759 30175
rect 11701 30135 11759 30141
rect 13265 30175 13323 30181
rect 13265 30141 13277 30175
rect 13311 30172 13323 30175
rect 14366 30172 14372 30184
rect 13311 30144 14372 30172
rect 13311 30141 13323 30144
rect 13265 30135 13323 30141
rect 14366 30132 14372 30144
rect 14424 30132 14430 30184
rect 15378 30132 15384 30184
rect 15436 30132 15442 30184
rect 15488 30172 15516 30212
rect 15672 30212 16580 30240
rect 15672 30172 15700 30212
rect 16574 30200 16580 30212
rect 16632 30240 16638 30252
rect 16669 30243 16727 30249
rect 16669 30240 16681 30243
rect 16632 30212 16681 30240
rect 16632 30200 16638 30212
rect 16669 30209 16681 30212
rect 16715 30209 16727 30243
rect 16669 30203 16727 30209
rect 17773 30243 17831 30249
rect 17773 30209 17785 30243
rect 17819 30240 17831 30243
rect 17819 30212 18828 30240
rect 17819 30209 17831 30212
rect 17773 30203 17831 30209
rect 15488 30144 15700 30172
rect 15746 30132 15752 30184
rect 15804 30172 15810 30184
rect 15804 30144 16804 30172
rect 15804 30132 15810 30144
rect 10410 30064 10416 30116
rect 10468 30104 10474 30116
rect 12621 30107 12679 30113
rect 12621 30104 12633 30107
rect 10468 30076 12633 30104
rect 10468 30064 10474 30076
rect 12621 30073 12633 30076
rect 12667 30073 12679 30107
rect 16776 30104 16804 30144
rect 16850 30132 16856 30184
rect 16908 30172 16914 30184
rect 17865 30175 17923 30181
rect 17865 30172 17877 30175
rect 16908 30144 17877 30172
rect 16908 30132 16914 30144
rect 17865 30141 17877 30144
rect 17911 30141 17923 30175
rect 18800 30172 18828 30212
rect 18874 30200 18880 30252
rect 18932 30200 18938 30252
rect 23566 30240 23572 30252
rect 18984 30212 20116 30240
rect 18984 30172 19012 30212
rect 18800 30144 19012 30172
rect 17865 30135 17923 30141
rect 19058 30132 19064 30184
rect 19116 30132 19122 30184
rect 19889 30175 19947 30181
rect 19889 30141 19901 30175
rect 19935 30141 19947 30175
rect 19889 30135 19947 30141
rect 18509 30107 18567 30113
rect 18509 30104 18521 30107
rect 16776 30076 18521 30104
rect 12621 30067 12679 30073
rect 18509 30073 18521 30076
rect 18555 30073 18567 30107
rect 19904 30104 19932 30135
rect 19978 30132 19984 30184
rect 20036 30132 20042 30184
rect 20088 30172 20116 30212
rect 22204 30212 23572 30240
rect 22204 30184 22232 30212
rect 23566 30200 23572 30212
rect 23624 30200 23630 30252
rect 20806 30172 20812 30184
rect 20088 30144 20812 30172
rect 20806 30132 20812 30144
rect 20864 30132 20870 30184
rect 22186 30132 22192 30184
rect 22244 30132 22250 30184
rect 22830 30172 22836 30184
rect 22296 30144 22836 30172
rect 22296 30104 22324 30144
rect 22830 30132 22836 30144
rect 22888 30132 22894 30184
rect 23477 30175 23535 30181
rect 23477 30141 23489 30175
rect 23523 30172 23535 30175
rect 23750 30172 23756 30184
rect 23523 30144 23756 30172
rect 23523 30141 23535 30144
rect 23477 30135 23535 30141
rect 23750 30132 23756 30144
rect 23808 30132 23814 30184
rect 24578 30132 24584 30184
rect 24636 30172 24642 30184
rect 24949 30175 25007 30181
rect 24949 30172 24961 30175
rect 24636 30144 24961 30172
rect 24636 30132 24642 30144
rect 24949 30141 24961 30144
rect 24995 30141 25007 30175
rect 24949 30135 25007 30141
rect 25225 30175 25283 30181
rect 25225 30141 25237 30175
rect 25271 30141 25283 30175
rect 25225 30135 25283 30141
rect 19904 30076 22324 30104
rect 18509 30067 18567 30073
rect 22554 30064 22560 30116
rect 22612 30104 22618 30116
rect 22612 30076 23612 30104
rect 22612 30064 22618 30076
rect 14826 29996 14832 30048
rect 14884 29996 14890 30048
rect 15838 29996 15844 30048
rect 15896 30036 15902 30048
rect 15933 30039 15991 30045
rect 15933 30036 15945 30039
rect 15896 30008 15945 30036
rect 15896 29996 15902 30008
rect 15933 30005 15945 30008
rect 15979 30036 15991 30039
rect 16114 30036 16120 30048
rect 15979 30008 16120 30036
rect 15979 30005 15991 30008
rect 15933 29999 15991 30005
rect 16114 29996 16120 30008
rect 16172 29996 16178 30048
rect 16206 29996 16212 30048
rect 16264 30036 16270 30048
rect 16301 30039 16359 30045
rect 16301 30036 16313 30039
rect 16264 30008 16313 30036
rect 16264 29996 16270 30008
rect 16301 30005 16313 30008
rect 16347 30005 16359 30039
rect 16301 29999 16359 30005
rect 20438 29996 20444 30048
rect 20496 29996 20502 30048
rect 22741 30039 22799 30045
rect 22741 30005 22753 30039
rect 22787 30036 22799 30039
rect 23382 30036 23388 30048
rect 22787 30008 23388 30036
rect 22787 30005 22799 30008
rect 22741 29999 22799 30005
rect 23382 29996 23388 30008
rect 23440 29996 23446 30048
rect 23584 30036 23612 30076
rect 25240 30036 25268 30135
rect 23584 30008 25268 30036
rect 1104 29946 25852 29968
rect 1104 29894 2950 29946
rect 3002 29894 3014 29946
rect 3066 29894 3078 29946
rect 3130 29894 3142 29946
rect 3194 29894 3206 29946
rect 3258 29894 12950 29946
rect 13002 29894 13014 29946
rect 13066 29894 13078 29946
rect 13130 29894 13142 29946
rect 13194 29894 13206 29946
rect 13258 29894 22950 29946
rect 23002 29894 23014 29946
rect 23066 29894 23078 29946
rect 23130 29894 23142 29946
rect 23194 29894 23206 29946
rect 23258 29894 25852 29946
rect 1104 29872 25852 29894
rect 4338 29792 4344 29844
rect 4396 29832 4402 29844
rect 8481 29835 8539 29841
rect 8481 29832 8493 29835
rect 4396 29804 8493 29832
rect 4396 29792 4402 29804
rect 8481 29801 8493 29804
rect 8527 29801 8539 29835
rect 8481 29795 8539 29801
rect 1302 29656 1308 29708
rect 1360 29696 1366 29708
rect 2041 29699 2099 29705
rect 2041 29696 2053 29699
rect 1360 29668 2053 29696
rect 1360 29656 1366 29668
rect 2041 29665 2053 29668
rect 2087 29665 2099 29699
rect 2041 29659 2099 29665
rect 3970 29656 3976 29708
rect 4028 29656 4034 29708
rect 1762 29588 1768 29640
rect 1820 29588 1826 29640
rect 8496 29628 8524 29795
rect 9030 29792 9036 29844
rect 9088 29832 9094 29844
rect 9125 29835 9183 29841
rect 9125 29832 9137 29835
rect 9088 29804 9137 29832
rect 9088 29792 9094 29804
rect 9125 29801 9137 29804
rect 9171 29801 9183 29835
rect 9125 29795 9183 29801
rect 12802 29792 12808 29844
rect 12860 29832 12866 29844
rect 12860 29804 13032 29832
rect 12860 29792 12866 29804
rect 11333 29767 11391 29773
rect 11333 29733 11345 29767
rect 11379 29764 11391 29767
rect 11379 29736 12940 29764
rect 11379 29733 11391 29736
rect 11333 29727 11391 29733
rect 9582 29656 9588 29708
rect 9640 29696 9646 29708
rect 9677 29699 9735 29705
rect 9677 29696 9689 29699
rect 9640 29668 9689 29696
rect 9640 29656 9646 29668
rect 9677 29665 9689 29668
rect 9723 29665 9735 29699
rect 9677 29659 9735 29665
rect 10686 29656 10692 29708
rect 10744 29656 10750 29708
rect 10870 29656 10876 29708
rect 10928 29696 10934 29708
rect 12345 29699 12403 29705
rect 12345 29696 12357 29699
rect 10928 29668 12357 29696
rect 10928 29656 10934 29668
rect 12345 29665 12357 29668
rect 12391 29665 12403 29699
rect 12345 29659 12403 29665
rect 9398 29628 9404 29640
rect 8496 29600 9404 29628
rect 9398 29588 9404 29600
rect 9456 29628 9462 29640
rect 9493 29631 9551 29637
rect 9493 29628 9505 29631
rect 9456 29600 9505 29628
rect 9456 29588 9462 29600
rect 9493 29597 9505 29600
rect 9539 29597 9551 29631
rect 9493 29591 9551 29597
rect 10962 29588 10968 29640
rect 11020 29588 11026 29640
rect 12912 29628 12940 29736
rect 13004 29696 13032 29804
rect 15102 29792 15108 29844
rect 15160 29832 15166 29844
rect 19058 29832 19064 29844
rect 15160 29804 19064 29832
rect 15160 29792 15166 29804
rect 19058 29792 19064 29804
rect 19116 29792 19122 29844
rect 25130 29792 25136 29844
rect 25188 29792 25194 29844
rect 15010 29724 15016 29776
rect 15068 29764 15074 29776
rect 16482 29764 16488 29776
rect 15068 29736 16488 29764
rect 15068 29724 15074 29736
rect 16482 29724 16488 29736
rect 16540 29724 16546 29776
rect 17865 29767 17923 29773
rect 17865 29733 17877 29767
rect 17911 29764 17923 29767
rect 19242 29764 19248 29776
rect 17911 29736 19248 29764
rect 17911 29733 17923 29736
rect 17865 29727 17923 29733
rect 19242 29724 19248 29736
rect 19300 29724 19306 29776
rect 21174 29724 21180 29776
rect 21232 29764 21238 29776
rect 23750 29764 23756 29776
rect 21232 29736 22140 29764
rect 21232 29724 21238 29736
rect 13081 29699 13139 29705
rect 13081 29696 13093 29699
rect 13004 29668 13093 29696
rect 13081 29665 13093 29668
rect 13127 29665 13139 29699
rect 13081 29659 13139 29665
rect 13265 29699 13323 29705
rect 13265 29665 13277 29699
rect 13311 29696 13323 29699
rect 13446 29696 13452 29708
rect 13311 29668 13452 29696
rect 13311 29665 13323 29668
rect 13265 29659 13323 29665
rect 13446 29656 13452 29668
rect 13504 29656 13510 29708
rect 17313 29699 17371 29705
rect 17313 29665 17325 29699
rect 17359 29696 17371 29699
rect 17586 29696 17592 29708
rect 17359 29668 17592 29696
rect 17359 29665 17371 29668
rect 17313 29659 17371 29665
rect 17586 29656 17592 29668
rect 17644 29656 17650 29708
rect 18230 29656 18236 29708
rect 18288 29656 18294 29708
rect 19886 29656 19892 29708
rect 19944 29656 19950 29708
rect 19978 29656 19984 29708
rect 20036 29656 20042 29708
rect 20162 29656 20168 29708
rect 20220 29696 20226 29708
rect 22112 29705 22140 29736
rect 23308 29736 23756 29764
rect 21361 29699 21419 29705
rect 21361 29696 21373 29699
rect 20220 29668 21373 29696
rect 20220 29656 20226 29668
rect 21361 29665 21373 29668
rect 21407 29665 21419 29699
rect 21361 29659 21419 29665
rect 22097 29699 22155 29705
rect 22097 29665 22109 29699
rect 22143 29665 22155 29699
rect 22097 29659 22155 29665
rect 22278 29656 22284 29708
rect 22336 29656 22342 29708
rect 22462 29656 22468 29708
rect 22520 29696 22526 29708
rect 22738 29696 22744 29708
rect 22520 29668 22744 29696
rect 22520 29656 22526 29668
rect 22738 29656 22744 29668
rect 22796 29656 22802 29708
rect 23308 29705 23336 29736
rect 23750 29724 23756 29736
rect 23808 29724 23814 29776
rect 23293 29699 23351 29705
rect 23293 29665 23305 29699
rect 23339 29665 23351 29699
rect 23293 29659 23351 29665
rect 23382 29656 23388 29708
rect 23440 29696 23446 29708
rect 23477 29699 23535 29705
rect 23477 29696 23489 29699
rect 23440 29668 23489 29696
rect 23440 29656 23446 29668
rect 23477 29665 23489 29668
rect 23523 29665 23535 29699
rect 23477 29659 23535 29665
rect 13357 29631 13415 29637
rect 13357 29628 13369 29631
rect 12912 29600 13369 29628
rect 13357 29597 13369 29600
rect 13403 29597 13415 29631
rect 13357 29591 13415 29597
rect 17405 29631 17463 29637
rect 17405 29597 17417 29631
rect 17451 29628 17463 29631
rect 18248 29628 18276 29656
rect 17451 29600 18276 29628
rect 17451 29597 17463 29600
rect 17405 29591 17463 29597
rect 19794 29588 19800 29640
rect 19852 29588 19858 29640
rect 21269 29631 21327 29637
rect 21269 29597 21281 29631
rect 21315 29628 21327 29631
rect 22002 29628 22008 29640
rect 21315 29600 22008 29628
rect 21315 29597 21327 29600
rect 21269 29591 21327 29597
rect 22002 29588 22008 29600
rect 22060 29588 22066 29640
rect 22373 29631 22431 29637
rect 22373 29597 22385 29631
rect 22419 29628 22431 29631
rect 23658 29628 23664 29640
rect 22419 29600 23664 29628
rect 22419 29597 22431 29600
rect 22373 29591 22431 29597
rect 23658 29588 23664 29600
rect 23716 29588 23722 29640
rect 25314 29588 25320 29640
rect 25372 29588 25378 29640
rect 3510 29520 3516 29572
rect 3568 29560 3574 29572
rect 4157 29563 4215 29569
rect 4157 29560 4169 29563
rect 3568 29532 4169 29560
rect 3568 29520 3574 29532
rect 4157 29529 4169 29532
rect 4203 29529 4215 29563
rect 4157 29523 4215 29529
rect 5810 29520 5816 29572
rect 5868 29520 5874 29572
rect 8754 29520 8760 29572
rect 8812 29560 8818 29572
rect 9585 29563 9643 29569
rect 9585 29560 9597 29563
rect 8812 29532 9597 29560
rect 8812 29520 8818 29532
rect 9585 29529 9597 29532
rect 9631 29560 9643 29563
rect 12342 29560 12348 29572
rect 9631 29532 12348 29560
rect 9631 29529 9643 29532
rect 9585 29523 9643 29529
rect 12342 29520 12348 29532
rect 12400 29520 12406 29572
rect 12618 29520 12624 29572
rect 12676 29560 12682 29572
rect 16761 29563 16819 29569
rect 16761 29560 16773 29563
rect 12676 29532 16773 29560
rect 12676 29520 12682 29532
rect 16761 29529 16773 29532
rect 16807 29560 16819 29563
rect 17497 29563 17555 29569
rect 17497 29560 17509 29563
rect 16807 29532 17509 29560
rect 16807 29529 16819 29532
rect 16761 29523 16819 29529
rect 17497 29529 17509 29532
rect 17543 29529 17555 29563
rect 17497 29523 17555 29529
rect 21177 29563 21235 29569
rect 21177 29529 21189 29563
rect 21223 29560 21235 29563
rect 22094 29560 22100 29572
rect 21223 29532 22100 29560
rect 21223 29529 21235 29532
rect 21177 29523 21235 29529
rect 22094 29520 22100 29532
rect 22152 29520 22158 29572
rect 10134 29452 10140 29504
rect 10192 29492 10198 29504
rect 10229 29495 10287 29501
rect 10229 29492 10241 29495
rect 10192 29464 10241 29492
rect 10192 29452 10198 29464
rect 10229 29461 10241 29464
rect 10275 29492 10287 29495
rect 10318 29492 10324 29504
rect 10275 29464 10324 29492
rect 10275 29461 10287 29464
rect 10229 29455 10287 29461
rect 10318 29452 10324 29464
rect 10376 29492 10382 29504
rect 10873 29495 10931 29501
rect 10873 29492 10885 29495
rect 10376 29464 10885 29492
rect 10376 29452 10382 29464
rect 10873 29461 10885 29464
rect 10919 29461 10931 29495
rect 10873 29455 10931 29461
rect 10962 29452 10968 29504
rect 11020 29492 11026 29504
rect 11793 29495 11851 29501
rect 11793 29492 11805 29495
rect 11020 29464 11805 29492
rect 11020 29452 11026 29464
rect 11793 29461 11805 29464
rect 11839 29461 11851 29495
rect 11793 29455 11851 29461
rect 12158 29452 12164 29504
rect 12216 29452 12222 29504
rect 12250 29452 12256 29504
rect 12308 29492 12314 29504
rect 13078 29492 13084 29504
rect 12308 29464 13084 29492
rect 12308 29452 12314 29464
rect 13078 29452 13084 29464
rect 13136 29452 13142 29504
rect 13722 29452 13728 29504
rect 13780 29452 13786 29504
rect 19426 29452 19432 29504
rect 19484 29452 19490 29504
rect 20809 29495 20867 29501
rect 20809 29461 20821 29495
rect 20855 29492 20867 29495
rect 20990 29492 20996 29504
rect 20855 29464 20996 29492
rect 20855 29461 20867 29464
rect 20809 29455 20867 29461
rect 20990 29452 20996 29464
rect 21048 29452 21054 29504
rect 22738 29452 22744 29504
rect 22796 29452 22802 29504
rect 23566 29452 23572 29504
rect 23624 29452 23630 29504
rect 23934 29452 23940 29504
rect 23992 29452 23998 29504
rect 1104 29402 25852 29424
rect 1104 29350 7950 29402
rect 8002 29350 8014 29402
rect 8066 29350 8078 29402
rect 8130 29350 8142 29402
rect 8194 29350 8206 29402
rect 8258 29350 17950 29402
rect 18002 29350 18014 29402
rect 18066 29350 18078 29402
rect 18130 29350 18142 29402
rect 18194 29350 18206 29402
rect 18258 29350 25852 29402
rect 1104 29328 25852 29350
rect 8202 29248 8208 29300
rect 8260 29288 8266 29300
rect 10870 29288 10876 29300
rect 8260 29260 10876 29288
rect 8260 29248 8266 29260
rect 10870 29248 10876 29260
rect 10928 29248 10934 29300
rect 12158 29248 12164 29300
rect 12216 29288 12222 29300
rect 12894 29288 12900 29300
rect 12216 29260 12900 29288
rect 12216 29248 12222 29260
rect 12894 29248 12900 29260
rect 12952 29248 12958 29300
rect 13078 29248 13084 29300
rect 13136 29288 13142 29300
rect 14642 29288 14648 29300
rect 13136 29260 14648 29288
rect 13136 29248 13142 29260
rect 14642 29248 14648 29260
rect 14700 29288 14706 29300
rect 18414 29288 18420 29300
rect 14700 29260 18420 29288
rect 14700 29248 14706 29260
rect 18414 29248 18420 29260
rect 18472 29248 18478 29300
rect 19794 29288 19800 29300
rect 19260 29260 19800 29288
rect 9214 29180 9220 29232
rect 9272 29220 9278 29232
rect 9582 29220 9588 29232
rect 9272 29192 9588 29220
rect 9272 29180 9278 29192
rect 9582 29180 9588 29192
rect 9640 29220 9646 29232
rect 9640 29192 9996 29220
rect 9640 29180 9646 29192
rect 9968 29152 9996 29192
rect 10042 29180 10048 29232
rect 10100 29220 10106 29232
rect 10318 29220 10324 29232
rect 10100 29192 10324 29220
rect 10100 29180 10106 29192
rect 10318 29180 10324 29192
rect 10376 29180 10382 29232
rect 12253 29223 12311 29229
rect 12253 29189 12265 29223
rect 12299 29220 12311 29223
rect 13354 29220 13360 29232
rect 12299 29192 13360 29220
rect 12299 29189 12311 29192
rect 12253 29183 12311 29189
rect 13354 29180 13360 29192
rect 13412 29220 13418 29232
rect 16206 29220 16212 29232
rect 13412 29192 16212 29220
rect 13412 29180 13418 29192
rect 16206 29180 16212 29192
rect 16264 29180 16270 29232
rect 19260 29220 19288 29260
rect 19794 29248 19800 29260
rect 19852 29248 19858 29300
rect 25314 29248 25320 29300
rect 25372 29288 25378 29300
rect 25409 29291 25467 29297
rect 25409 29288 25421 29291
rect 25372 29260 25421 29288
rect 25372 29248 25378 29260
rect 25409 29257 25421 29260
rect 25455 29257 25467 29291
rect 25409 29251 25467 29257
rect 18814 29192 19288 29220
rect 19334 29180 19340 29232
rect 19392 29220 19398 29232
rect 19392 29192 19564 29220
rect 19392 29180 19398 29192
rect 10229 29155 10287 29161
rect 10229 29152 10241 29155
rect 9968 29124 10241 29152
rect 10229 29121 10241 29124
rect 10275 29121 10287 29155
rect 10229 29115 10287 29121
rect 12161 29155 12219 29161
rect 12161 29121 12173 29155
rect 12207 29152 12219 29155
rect 16301 29155 16359 29161
rect 12207 29124 13308 29152
rect 12207 29121 12219 29124
rect 12161 29115 12219 29121
rect 9950 29044 9956 29096
rect 10008 29044 10014 29096
rect 10042 29044 10048 29096
rect 10100 29084 10106 29096
rect 13280 29093 13308 29124
rect 16301 29121 16313 29155
rect 16347 29152 16359 29155
rect 16758 29152 16764 29164
rect 16347 29124 16764 29152
rect 16347 29121 16359 29124
rect 16301 29115 16359 29121
rect 16758 29112 16764 29124
rect 16816 29112 16822 29164
rect 19536 29161 19564 29192
rect 24670 29180 24676 29232
rect 24728 29220 24734 29232
rect 24765 29223 24823 29229
rect 24765 29220 24777 29223
rect 24728 29192 24777 29220
rect 24728 29180 24734 29192
rect 24765 29189 24777 29192
rect 24811 29189 24823 29223
rect 24765 29183 24823 29189
rect 19521 29155 19579 29161
rect 19521 29121 19533 29155
rect 19567 29121 19579 29155
rect 19521 29115 19579 29121
rect 23661 29155 23719 29161
rect 23661 29121 23673 29155
rect 23707 29152 23719 29155
rect 24118 29152 24124 29164
rect 23707 29124 24124 29152
rect 23707 29121 23719 29124
rect 23661 29115 23719 29121
rect 24118 29112 24124 29124
rect 24176 29112 24182 29164
rect 12345 29087 12403 29093
rect 12345 29084 12357 29087
rect 10100 29056 12357 29084
rect 10100 29044 10106 29056
rect 12345 29053 12357 29056
rect 12391 29053 12403 29087
rect 12345 29047 12403 29053
rect 13265 29087 13323 29093
rect 13265 29053 13277 29087
rect 13311 29084 13323 29087
rect 17494 29084 17500 29096
rect 13311 29056 17500 29084
rect 13311 29053 13323 29056
rect 13265 29047 13323 29053
rect 17494 29044 17500 29056
rect 17552 29044 17558 29096
rect 18782 29044 18788 29096
rect 18840 29084 18846 29096
rect 19245 29087 19303 29093
rect 19245 29084 19257 29087
rect 18840 29056 19257 29084
rect 18840 29044 18846 29056
rect 19245 29053 19257 29056
rect 19291 29053 19303 29087
rect 19245 29047 19303 29053
rect 19444 29056 22094 29084
rect 10410 28976 10416 29028
rect 10468 29016 10474 29028
rect 11793 29019 11851 29025
rect 11793 29016 11805 29019
rect 10468 28988 11805 29016
rect 10468 28976 10474 28988
rect 11793 28985 11805 28988
rect 11839 28985 11851 29019
rect 11793 28979 11851 28985
rect 12894 28976 12900 29028
rect 12952 29016 12958 29028
rect 15013 29019 15071 29025
rect 12952 28988 14964 29016
rect 12952 28976 12958 28988
rect 9695 28951 9753 28957
rect 9695 28917 9707 28951
rect 9741 28948 9753 28951
rect 9858 28948 9864 28960
rect 9741 28920 9864 28948
rect 9741 28917 9753 28920
rect 9695 28911 9753 28917
rect 9858 28908 9864 28920
rect 9916 28908 9922 28960
rect 12158 28908 12164 28960
rect 12216 28948 12222 28960
rect 13354 28948 13360 28960
rect 12216 28920 13360 28948
rect 12216 28908 12222 28920
rect 13354 28908 13360 28920
rect 13412 28908 13418 28960
rect 14936 28948 14964 28988
rect 15013 28985 15025 29019
rect 15059 29016 15071 29019
rect 15194 29016 15200 29028
rect 15059 28988 15200 29016
rect 15059 28985 15071 28988
rect 15013 28979 15071 28985
rect 15194 28976 15200 28988
rect 15252 28976 15258 29028
rect 15304 28988 16712 29016
rect 15304 28948 15332 28988
rect 14936 28920 15332 28948
rect 16684 28948 16712 28988
rect 16758 28976 16764 29028
rect 16816 28976 16822 29028
rect 17402 29016 17408 29028
rect 16868 28988 17408 29016
rect 16868 28948 16896 28988
rect 17402 28976 17408 28988
rect 17460 28976 17466 29028
rect 16684 28920 16896 28948
rect 17770 28908 17776 28960
rect 17828 28908 17834 28960
rect 18598 28908 18604 28960
rect 18656 28948 18662 28960
rect 19444 28948 19472 29056
rect 22066 29016 22094 29056
rect 22186 29044 22192 29096
rect 22244 29044 22250 29096
rect 23937 29019 23995 29025
rect 23937 29016 23949 29019
rect 22066 28988 23949 29016
rect 23937 28985 23949 28988
rect 23983 28985 23995 29019
rect 23937 28979 23995 28985
rect 24578 28976 24584 29028
rect 24636 28976 24642 29028
rect 18656 28920 19472 28948
rect 18656 28908 18662 28920
rect 1104 28858 25852 28880
rect 1104 28806 2950 28858
rect 3002 28806 3014 28858
rect 3066 28806 3078 28858
rect 3130 28806 3142 28858
rect 3194 28806 3206 28858
rect 3258 28806 12950 28858
rect 13002 28806 13014 28858
rect 13066 28806 13078 28858
rect 13130 28806 13142 28858
rect 13194 28806 13206 28858
rect 13258 28806 22950 28858
rect 23002 28806 23014 28858
rect 23066 28806 23078 28858
rect 23130 28806 23142 28858
rect 23194 28806 23206 28858
rect 23258 28806 25852 28858
rect 1104 28784 25852 28806
rect 4246 28704 4252 28756
rect 4304 28744 4310 28756
rect 7374 28744 7380 28756
rect 4304 28716 7380 28744
rect 4304 28704 4310 28716
rect 7374 28704 7380 28716
rect 7432 28744 7438 28756
rect 8481 28747 8539 28753
rect 8481 28744 8493 28747
rect 7432 28716 8493 28744
rect 7432 28704 7438 28716
rect 1946 28568 1952 28620
rect 2004 28608 2010 28620
rect 3973 28611 4031 28617
rect 3973 28608 3985 28611
rect 2004 28580 3985 28608
rect 2004 28568 2010 28580
rect 3973 28577 3985 28580
rect 4019 28577 4031 28611
rect 3973 28571 4031 28577
rect 8018 28568 8024 28620
rect 8076 28568 8082 28620
rect 4157 28475 4215 28481
rect 4157 28441 4169 28475
rect 4203 28441 4215 28475
rect 4157 28435 4215 28441
rect 4062 28364 4068 28416
rect 4120 28404 4126 28416
rect 4172 28404 4200 28435
rect 5718 28432 5724 28484
rect 5776 28472 5782 28484
rect 5813 28475 5871 28481
rect 5813 28472 5825 28475
rect 5776 28444 5825 28472
rect 5776 28432 5782 28444
rect 5813 28441 5825 28444
rect 5859 28441 5871 28475
rect 7466 28472 7472 28484
rect 7314 28444 7472 28472
rect 5813 28435 5871 28441
rect 7466 28432 7472 28444
rect 7524 28432 7530 28484
rect 7745 28475 7803 28481
rect 7745 28441 7757 28475
rect 7791 28472 7803 28475
rect 8202 28472 8208 28484
rect 7791 28444 8208 28472
rect 7791 28441 7803 28444
rect 7745 28435 7803 28441
rect 4120 28376 4200 28404
rect 6273 28407 6331 28413
rect 4120 28364 4126 28376
rect 6273 28373 6285 28407
rect 6319 28404 6331 28407
rect 6914 28404 6920 28416
rect 6319 28376 6920 28404
rect 6319 28373 6331 28376
rect 6273 28367 6331 28373
rect 6914 28364 6920 28376
rect 6972 28364 6978 28416
rect 7558 28364 7564 28416
rect 7616 28404 7622 28416
rect 7760 28404 7788 28435
rect 8202 28432 8208 28444
rect 8260 28432 8266 28484
rect 7616 28376 7788 28404
rect 8312 28404 8340 28716
rect 8481 28713 8493 28716
rect 8527 28713 8539 28747
rect 8481 28707 8539 28713
rect 9766 28704 9772 28756
rect 9824 28744 9830 28756
rect 9861 28747 9919 28753
rect 9861 28744 9873 28747
rect 9824 28716 9873 28744
rect 9824 28704 9830 28716
rect 9861 28713 9873 28716
rect 9907 28713 9919 28747
rect 9861 28707 9919 28713
rect 12618 28704 12624 28756
rect 12676 28744 12682 28756
rect 13449 28747 13507 28753
rect 13449 28744 13461 28747
rect 12676 28716 13461 28744
rect 12676 28704 12682 28716
rect 13449 28713 13461 28716
rect 13495 28713 13507 28747
rect 13449 28707 13507 28713
rect 14182 28704 14188 28756
rect 14240 28744 14246 28756
rect 16301 28747 16359 28753
rect 14240 28716 16252 28744
rect 14240 28704 14246 28716
rect 8389 28679 8447 28685
rect 8389 28645 8401 28679
rect 8435 28676 8447 28679
rect 8570 28676 8576 28688
rect 8435 28648 8576 28676
rect 8435 28645 8447 28648
rect 8389 28639 8447 28645
rect 8570 28636 8576 28648
rect 8628 28676 8634 28688
rect 9214 28676 9220 28688
rect 8628 28648 9220 28676
rect 8628 28636 8634 28648
rect 9214 28636 9220 28648
rect 9272 28636 9278 28688
rect 10778 28676 10784 28688
rect 9324 28648 10784 28676
rect 9324 28617 9352 28648
rect 10778 28636 10784 28648
rect 10836 28636 10842 28688
rect 16224 28676 16252 28716
rect 16301 28713 16313 28747
rect 16347 28744 16359 28747
rect 16666 28744 16672 28756
rect 16347 28716 16672 28744
rect 16347 28713 16359 28716
rect 16301 28707 16359 28713
rect 16666 28704 16672 28716
rect 16724 28704 16730 28756
rect 17586 28704 17592 28756
rect 17644 28744 17650 28756
rect 21082 28744 21088 28756
rect 17644 28716 21088 28744
rect 17644 28704 17650 28716
rect 21082 28704 21088 28716
rect 21140 28704 21146 28756
rect 22557 28747 22615 28753
rect 22557 28713 22569 28747
rect 22603 28744 22615 28747
rect 23566 28744 23572 28756
rect 22603 28716 23572 28744
rect 22603 28713 22615 28716
rect 22557 28707 22615 28713
rect 23566 28704 23572 28716
rect 23624 28704 23630 28756
rect 25133 28747 25191 28753
rect 25133 28713 25145 28747
rect 25179 28744 25191 28747
rect 25222 28744 25228 28756
rect 25179 28716 25228 28744
rect 25179 28713 25191 28716
rect 25133 28707 25191 28713
rect 25222 28704 25228 28716
rect 25280 28704 25286 28756
rect 16224 28648 19656 28676
rect 9309 28611 9367 28617
rect 9309 28577 9321 28611
rect 9355 28577 9367 28611
rect 9309 28571 9367 28577
rect 9950 28568 9956 28620
rect 10008 28608 10014 28620
rect 10962 28608 10968 28620
rect 10008 28580 10968 28608
rect 10008 28568 10014 28580
rect 10962 28568 10968 28580
rect 11020 28608 11026 28620
rect 11241 28611 11299 28617
rect 11241 28608 11253 28611
rect 11020 28580 11253 28608
rect 11020 28568 11026 28580
rect 11241 28577 11253 28580
rect 11287 28577 11299 28611
rect 11241 28571 11299 28577
rect 11517 28611 11575 28617
rect 11517 28577 11529 28611
rect 11563 28608 11575 28611
rect 12802 28608 12808 28620
rect 11563 28580 12808 28608
rect 11563 28577 11575 28580
rect 11517 28571 11575 28577
rect 12802 28568 12808 28580
rect 12860 28568 12866 28620
rect 12989 28611 13047 28617
rect 12989 28577 13001 28611
rect 13035 28608 13047 28611
rect 13630 28608 13636 28620
rect 13035 28580 13636 28608
rect 13035 28577 13047 28580
rect 12989 28571 13047 28577
rect 13630 28568 13636 28580
rect 13688 28568 13694 28620
rect 14274 28568 14280 28620
rect 14332 28608 14338 28620
rect 14553 28611 14611 28617
rect 14553 28608 14565 28611
rect 14332 28580 14565 28608
rect 14332 28568 14338 28580
rect 14553 28577 14565 28580
rect 14599 28577 14611 28611
rect 14553 28571 14611 28577
rect 14829 28611 14887 28617
rect 14829 28577 14841 28611
rect 14875 28608 14887 28611
rect 17589 28611 17647 28617
rect 17589 28608 17601 28611
rect 14875 28580 17601 28608
rect 14875 28577 14887 28580
rect 14829 28571 14887 28577
rect 17589 28577 17601 28580
rect 17635 28608 17647 28611
rect 17770 28608 17776 28620
rect 17635 28580 17776 28608
rect 17635 28577 17647 28580
rect 17589 28571 17647 28577
rect 17770 28568 17776 28580
rect 17828 28568 17834 28620
rect 19518 28568 19524 28620
rect 19576 28568 19582 28620
rect 19628 28608 19656 28648
rect 19702 28636 19708 28688
rect 19760 28676 19766 28688
rect 23845 28679 23903 28685
rect 23845 28676 23857 28679
rect 19760 28648 23857 28676
rect 19760 28636 19766 28648
rect 23845 28645 23857 28648
rect 23891 28645 23903 28679
rect 23845 28639 23903 28645
rect 20809 28611 20867 28617
rect 19628 28580 20760 28608
rect 8757 28543 8815 28549
rect 8757 28509 8769 28543
rect 8803 28540 8815 28543
rect 8938 28540 8944 28552
rect 8803 28512 8944 28540
rect 8803 28509 8815 28512
rect 8757 28503 8815 28509
rect 8938 28500 8944 28512
rect 8996 28540 9002 28552
rect 9401 28543 9459 28549
rect 9401 28540 9413 28543
rect 8996 28512 9413 28540
rect 8996 28500 9002 28512
rect 9401 28509 9413 28512
rect 9447 28540 9459 28543
rect 9490 28540 9496 28552
rect 9447 28512 9496 28540
rect 9447 28509 9459 28512
rect 9401 28503 9459 28509
rect 9490 28500 9496 28512
rect 9548 28500 9554 28552
rect 16574 28500 16580 28552
rect 16632 28540 16638 28552
rect 17126 28540 17132 28552
rect 16632 28512 17132 28540
rect 16632 28500 16638 28512
rect 17126 28500 17132 28512
rect 17184 28500 17190 28552
rect 19242 28500 19248 28552
rect 19300 28540 19306 28552
rect 19705 28543 19763 28549
rect 19705 28540 19717 28543
rect 19300 28512 19717 28540
rect 19300 28500 19306 28512
rect 19705 28509 19717 28512
rect 19751 28509 19763 28543
rect 19705 28503 19763 28509
rect 19797 28543 19855 28549
rect 19797 28509 19809 28543
rect 19843 28540 19855 28543
rect 20622 28540 20628 28552
rect 19843 28512 20628 28540
rect 19843 28509 19855 28512
rect 19797 28503 19855 28509
rect 20622 28500 20628 28512
rect 20680 28500 20686 28552
rect 20732 28540 20760 28580
rect 20809 28577 20821 28611
rect 20855 28608 20867 28611
rect 21174 28608 21180 28620
rect 20855 28580 21180 28608
rect 20855 28577 20867 28580
rect 20809 28571 20867 28577
rect 21174 28568 21180 28580
rect 21232 28568 21238 28620
rect 22005 28611 22063 28617
rect 22005 28577 22017 28611
rect 22051 28608 22063 28611
rect 22094 28608 22100 28620
rect 22051 28580 22100 28608
rect 22051 28577 22063 28580
rect 22005 28571 22063 28577
rect 22094 28568 22100 28580
rect 22152 28568 22158 28620
rect 24489 28611 24547 28617
rect 24489 28577 24501 28611
rect 24535 28608 24547 28611
rect 24670 28608 24676 28620
rect 24535 28580 24676 28608
rect 24535 28577 24547 28580
rect 24489 28571 24547 28577
rect 24670 28568 24676 28580
rect 24728 28568 24734 28620
rect 20732 28512 22140 28540
rect 12526 28432 12532 28484
rect 12584 28432 12590 28484
rect 17405 28475 17463 28481
rect 13832 28444 15318 28472
rect 13832 28416 13860 28444
rect 9493 28407 9551 28413
rect 9493 28404 9505 28407
rect 8312 28376 9505 28404
rect 7616 28364 7622 28376
rect 9493 28373 9505 28376
rect 9539 28373 9551 28407
rect 9493 28367 9551 28373
rect 13357 28407 13415 28413
rect 13357 28373 13369 28407
rect 13403 28404 13415 28407
rect 13814 28404 13820 28416
rect 13403 28376 13820 28404
rect 13403 28373 13415 28376
rect 13357 28367 13415 28373
rect 13814 28364 13820 28376
rect 13872 28364 13878 28416
rect 15212 28404 15240 28444
rect 17405 28441 17417 28475
rect 17451 28472 17463 28475
rect 18233 28475 18291 28481
rect 18233 28472 18245 28475
rect 17451 28444 18245 28472
rect 17451 28441 17463 28444
rect 17405 28435 17463 28441
rect 18233 28441 18245 28444
rect 18279 28441 18291 28475
rect 18233 28435 18291 28441
rect 20530 28432 20536 28484
rect 20588 28472 20594 28484
rect 22112 28481 22140 28512
rect 22186 28500 22192 28552
rect 22244 28500 22250 28552
rect 24029 28543 24087 28549
rect 24029 28509 24041 28543
rect 24075 28540 24087 28543
rect 25317 28543 25375 28549
rect 24075 28512 24716 28540
rect 24075 28509 24087 28512
rect 24029 28503 24087 28509
rect 20993 28475 21051 28481
rect 20993 28472 21005 28475
rect 20588 28444 21005 28472
rect 20588 28432 20594 28444
rect 20993 28441 21005 28444
rect 21039 28441 21051 28475
rect 20993 28435 21051 28441
rect 22097 28475 22155 28481
rect 22097 28441 22109 28475
rect 22143 28472 22155 28475
rect 22833 28475 22891 28481
rect 22833 28472 22845 28475
rect 22143 28444 22845 28472
rect 22143 28441 22155 28444
rect 22097 28435 22155 28441
rect 22833 28441 22845 28444
rect 22879 28441 22891 28475
rect 22833 28435 22891 28441
rect 16577 28407 16635 28413
rect 16577 28404 16589 28407
rect 15212 28376 16589 28404
rect 16577 28373 16589 28376
rect 16623 28373 16635 28407
rect 16577 28367 16635 28373
rect 17034 28364 17040 28416
rect 17092 28364 17098 28416
rect 17494 28364 17500 28416
rect 17552 28364 17558 28416
rect 18690 28364 18696 28416
rect 18748 28364 18754 28416
rect 19978 28364 19984 28416
rect 20036 28404 20042 28416
rect 20165 28407 20223 28413
rect 20165 28404 20177 28407
rect 20036 28376 20177 28404
rect 20036 28364 20042 28376
rect 20165 28373 20177 28376
rect 20211 28373 20223 28407
rect 20165 28367 20223 28373
rect 20898 28364 20904 28416
rect 20956 28364 20962 28416
rect 21358 28364 21364 28416
rect 21416 28364 21422 28416
rect 24688 28413 24716 28512
rect 25317 28509 25329 28543
rect 25363 28540 25375 28543
rect 25406 28540 25412 28552
rect 25363 28512 25412 28540
rect 25363 28509 25375 28512
rect 25317 28503 25375 28509
rect 25406 28500 25412 28512
rect 25464 28500 25470 28552
rect 24673 28407 24731 28413
rect 24673 28373 24685 28407
rect 24719 28404 24731 28407
rect 24854 28404 24860 28416
rect 24719 28376 24860 28404
rect 24719 28373 24731 28376
rect 24673 28367 24731 28373
rect 24854 28364 24860 28376
rect 24912 28364 24918 28416
rect 1104 28314 25852 28336
rect 1104 28262 7950 28314
rect 8002 28262 8014 28314
rect 8066 28262 8078 28314
rect 8130 28262 8142 28314
rect 8194 28262 8206 28314
rect 8258 28262 17950 28314
rect 18002 28262 18014 28314
rect 18066 28262 18078 28314
rect 18130 28262 18142 28314
rect 18194 28262 18206 28314
rect 18258 28262 25852 28314
rect 1104 28240 25852 28262
rect 7834 28200 7840 28212
rect 6564 28172 7840 28200
rect 6270 28024 6276 28076
rect 6328 28064 6334 28076
rect 6564 28073 6592 28172
rect 7834 28160 7840 28172
rect 7892 28160 7898 28212
rect 8570 28160 8576 28212
rect 8628 28160 8634 28212
rect 9217 28203 9275 28209
rect 9217 28169 9229 28203
rect 9263 28200 9275 28203
rect 9858 28200 9864 28212
rect 9263 28172 9864 28200
rect 9263 28169 9275 28172
rect 9217 28163 9275 28169
rect 9858 28160 9864 28172
rect 9916 28200 9922 28212
rect 11333 28203 11391 28209
rect 9916 28172 11100 28200
rect 9916 28160 9922 28172
rect 8588 28132 8616 28160
rect 8050 28104 9522 28132
rect 6549 28067 6607 28073
rect 6549 28064 6561 28067
rect 6328 28036 6561 28064
rect 6328 28024 6334 28036
rect 6549 28033 6561 28036
rect 6595 28033 6607 28067
rect 6549 28027 6607 28033
rect 10962 28024 10968 28076
rect 11020 28024 11026 28076
rect 11072 28064 11100 28172
rect 11333 28169 11345 28203
rect 11379 28200 11391 28203
rect 12526 28200 12532 28212
rect 11379 28172 12532 28200
rect 11379 28169 11391 28172
rect 11333 28163 11391 28169
rect 12526 28160 12532 28172
rect 12584 28160 12590 28212
rect 14645 28203 14703 28209
rect 14645 28169 14657 28203
rect 14691 28200 14703 28203
rect 15381 28203 15439 28209
rect 15381 28200 15393 28203
rect 14691 28172 15393 28200
rect 14691 28169 14703 28172
rect 14645 28163 14703 28169
rect 15381 28169 15393 28172
rect 15427 28200 15439 28203
rect 16574 28200 16580 28212
rect 15427 28172 16580 28200
rect 15427 28169 15439 28172
rect 15381 28163 15439 28169
rect 16574 28160 16580 28172
rect 16632 28160 16638 28212
rect 16853 28203 16911 28209
rect 16853 28169 16865 28203
rect 16899 28169 16911 28203
rect 16853 28163 16911 28169
rect 12253 28135 12311 28141
rect 12253 28101 12265 28135
rect 12299 28132 12311 28135
rect 12299 28104 13768 28132
rect 12299 28101 12311 28104
rect 12253 28095 12311 28101
rect 12618 28064 12624 28076
rect 11072 28036 12624 28064
rect 12618 28024 12624 28036
rect 12676 28024 12682 28076
rect 13740 28073 13768 28104
rect 16758 28092 16764 28144
rect 16816 28132 16822 28144
rect 16868 28132 16896 28163
rect 17310 28160 17316 28212
rect 17368 28160 17374 28212
rect 17494 28160 17500 28212
rect 17552 28200 17558 28212
rect 18049 28203 18107 28209
rect 18049 28200 18061 28203
rect 17552 28172 18061 28200
rect 17552 28160 17558 28172
rect 18049 28169 18061 28172
rect 18095 28169 18107 28203
rect 18049 28163 18107 28169
rect 18509 28203 18567 28209
rect 18509 28169 18521 28203
rect 18555 28200 18567 28203
rect 18598 28200 18604 28212
rect 18555 28172 18604 28200
rect 18555 28169 18567 28172
rect 18509 28163 18567 28169
rect 18598 28160 18604 28172
rect 18656 28160 18662 28212
rect 20438 28160 20444 28212
rect 20496 28200 20502 28212
rect 22281 28203 22339 28209
rect 22281 28200 22293 28203
rect 20496 28172 22293 28200
rect 20496 28160 20502 28172
rect 22281 28169 22293 28172
rect 22327 28169 22339 28203
rect 22281 28163 22339 28169
rect 22373 28203 22431 28209
rect 22373 28169 22385 28203
rect 22419 28200 22431 28203
rect 22646 28200 22652 28212
rect 22419 28172 22652 28200
rect 22419 28169 22431 28172
rect 22373 28163 22431 28169
rect 22646 28160 22652 28172
rect 22704 28160 22710 28212
rect 22741 28203 22799 28209
rect 22741 28169 22753 28203
rect 22787 28200 22799 28203
rect 22787 28172 25360 28200
rect 22787 28169 22799 28172
rect 22741 28163 22799 28169
rect 16816 28104 16896 28132
rect 17221 28135 17279 28141
rect 16816 28092 16822 28104
rect 17221 28101 17233 28135
rect 17267 28132 17279 28135
rect 17862 28132 17868 28144
rect 17267 28104 17868 28132
rect 17267 28101 17279 28104
rect 17221 28095 17279 28101
rect 17862 28092 17868 28104
rect 17920 28092 17926 28144
rect 17972 28104 19288 28132
rect 13725 28067 13783 28073
rect 13725 28033 13737 28067
rect 13771 28064 13783 28067
rect 13771 28036 14964 28064
rect 13771 28033 13783 28036
rect 13725 28027 13783 28033
rect 6825 27999 6883 28005
rect 6825 27965 6837 27999
rect 6871 27996 6883 27999
rect 6914 27996 6920 28008
rect 6871 27968 6920 27996
rect 6871 27965 6883 27968
rect 6825 27959 6883 27965
rect 6914 27956 6920 27968
rect 6972 27996 6978 28008
rect 7282 27996 7288 28008
rect 6972 27968 7288 27996
rect 6972 27956 6978 27968
rect 7282 27956 7288 27968
rect 7340 27956 7346 28008
rect 7834 27956 7840 28008
rect 7892 27996 7898 28008
rect 8297 27999 8355 28005
rect 8297 27996 8309 27999
rect 7892 27968 8309 27996
rect 7892 27956 7898 27968
rect 8297 27965 8309 27968
rect 8343 27996 8355 27999
rect 10042 27996 10048 28008
rect 8343 27968 10048 27996
rect 8343 27965 8355 27968
rect 8297 27959 8355 27965
rect 10042 27956 10048 27968
rect 10100 27956 10106 28008
rect 10594 27956 10600 28008
rect 10652 27996 10658 28008
rect 10689 27999 10747 28005
rect 10689 27996 10701 27999
rect 10652 27968 10701 27996
rect 10652 27956 10658 27968
rect 10689 27965 10701 27968
rect 10735 27965 10747 27999
rect 10689 27959 10747 27965
rect 10980 27928 11008 28024
rect 12066 27956 12072 28008
rect 12124 27996 12130 28008
rect 12342 27996 12348 28008
rect 12124 27968 12348 27996
rect 12124 27956 12130 27968
rect 12342 27956 12348 27968
rect 12400 27956 12406 28008
rect 12434 27956 12440 28008
rect 12492 27956 12498 28008
rect 13173 27999 13231 28005
rect 13173 27965 13185 27999
rect 13219 27996 13231 27999
rect 13354 27996 13360 28008
rect 13219 27968 13360 27996
rect 13219 27965 13231 27968
rect 13173 27959 13231 27965
rect 13354 27956 13360 27968
rect 13412 27956 13418 28008
rect 14001 27999 14059 28005
rect 14001 27965 14013 27999
rect 14047 27996 14059 27999
rect 14734 27996 14740 28008
rect 14047 27968 14740 27996
rect 14047 27965 14059 27968
rect 14001 27959 14059 27965
rect 14734 27956 14740 27968
rect 14792 27956 14798 28008
rect 14829 27999 14887 28005
rect 14829 27965 14841 27999
rect 14875 27965 14887 27999
rect 14829 27959 14887 27965
rect 13446 27928 13452 27940
rect 10980 27900 13452 27928
rect 13446 27888 13452 27900
rect 13504 27888 13510 27940
rect 14844 27928 14872 27959
rect 13556 27900 14872 27928
rect 10686 27820 10692 27872
rect 10744 27860 10750 27872
rect 11885 27863 11943 27869
rect 11885 27860 11897 27863
rect 10744 27832 11897 27860
rect 10744 27820 10750 27832
rect 11885 27829 11897 27832
rect 11931 27829 11943 27863
rect 11885 27823 11943 27829
rect 11974 27820 11980 27872
rect 12032 27860 12038 27872
rect 13556 27860 13584 27900
rect 12032 27832 13584 27860
rect 12032 27820 12038 27832
rect 13998 27820 14004 27872
rect 14056 27860 14062 27872
rect 14277 27863 14335 27869
rect 14277 27860 14289 27863
rect 14056 27832 14289 27860
rect 14056 27820 14062 27832
rect 14277 27829 14289 27832
rect 14323 27829 14335 27863
rect 14936 27860 14964 28036
rect 15930 28024 15936 28076
rect 15988 28064 15994 28076
rect 17972 28064 18000 28104
rect 15988 28036 18000 28064
rect 15988 28024 15994 28036
rect 18046 28024 18052 28076
rect 18104 28064 18110 28076
rect 18417 28067 18475 28073
rect 18417 28064 18429 28067
rect 18104 28036 18429 28064
rect 18104 28024 18110 28036
rect 18417 28033 18429 28036
rect 18463 28064 18475 28067
rect 18598 28064 18604 28076
rect 18463 28036 18604 28064
rect 18463 28033 18475 28036
rect 18417 28027 18475 28033
rect 18598 28024 18604 28036
rect 18656 28024 18662 28076
rect 19260 28073 19288 28104
rect 20898 28092 20904 28144
rect 20956 28132 20962 28144
rect 21453 28135 21511 28141
rect 21453 28132 21465 28135
rect 20956 28104 21465 28132
rect 20956 28092 20962 28104
rect 21453 28101 21465 28104
rect 21499 28101 21511 28135
rect 21453 28095 21511 28101
rect 24394 28092 24400 28144
rect 24452 28132 24458 28144
rect 24765 28135 24823 28141
rect 24765 28132 24777 28135
rect 24452 28104 24777 28132
rect 24452 28092 24458 28104
rect 24765 28101 24777 28104
rect 24811 28101 24823 28135
rect 25332 28132 25360 28172
rect 25406 28160 25412 28212
rect 25464 28160 25470 28212
rect 25498 28132 25504 28144
rect 25332 28104 25504 28132
rect 24765 28095 24823 28101
rect 25498 28092 25504 28104
rect 25556 28092 25562 28144
rect 19245 28067 19303 28073
rect 19245 28033 19257 28067
rect 19291 28033 19303 28067
rect 19245 28027 19303 28033
rect 20438 28024 20444 28076
rect 20496 28024 20502 28076
rect 23477 28067 23535 28073
rect 23477 28033 23489 28067
rect 23523 28033 23535 28067
rect 23477 28027 23535 28033
rect 17405 27999 17463 28005
rect 17405 27996 17417 27999
rect 15948 27968 17417 27996
rect 15948 27940 15976 27968
rect 17405 27965 17417 27968
rect 17451 27965 17463 27999
rect 17405 27959 17463 27965
rect 18693 27999 18751 28005
rect 18693 27965 18705 27999
rect 18739 27996 18751 27999
rect 18782 27996 18788 28008
rect 18739 27968 18788 27996
rect 18739 27965 18751 27968
rect 18693 27959 18751 27965
rect 18782 27956 18788 27968
rect 18840 27956 18846 28008
rect 22189 27999 22247 28005
rect 19352 27968 22094 27996
rect 15930 27888 15936 27940
rect 15988 27888 15994 27940
rect 16482 27888 16488 27940
rect 16540 27928 16546 27940
rect 19352 27928 19380 27968
rect 16540 27900 19380 27928
rect 19429 27931 19487 27937
rect 16540 27888 16546 27900
rect 19429 27897 19441 27931
rect 19475 27928 19487 27931
rect 21634 27928 21640 27940
rect 19475 27900 21640 27928
rect 19475 27897 19487 27900
rect 19429 27891 19487 27897
rect 21634 27888 21640 27900
rect 21692 27888 21698 27940
rect 22066 27928 22094 27968
rect 22189 27965 22201 27999
rect 22235 27996 22247 27999
rect 23492 27996 23520 28027
rect 23934 28024 23940 28076
rect 23992 28024 23998 28076
rect 24670 27996 24676 28008
rect 22235 27968 23428 27996
rect 23492 27968 24676 27996
rect 22235 27965 22247 27968
rect 22189 27959 22247 27965
rect 23293 27931 23351 27937
rect 23293 27928 23305 27931
rect 22066 27900 23305 27928
rect 23293 27897 23305 27900
rect 23339 27897 23351 27931
rect 23400 27928 23428 27968
rect 24670 27956 24676 27968
rect 24728 27956 24734 28008
rect 23934 27928 23940 27940
rect 23400 27900 23940 27928
rect 23293 27891 23351 27897
rect 23934 27888 23940 27900
rect 23992 27888 23998 27940
rect 24210 27888 24216 27940
rect 24268 27928 24274 27940
rect 24581 27931 24639 27937
rect 24581 27928 24593 27931
rect 24268 27900 24593 27928
rect 24268 27888 24274 27900
rect 24581 27897 24593 27900
rect 24627 27897 24639 27931
rect 24581 27891 24639 27897
rect 20070 27860 20076 27872
rect 14936 27832 20076 27860
rect 14277 27823 14335 27829
rect 20070 27820 20076 27832
rect 20128 27860 20134 27872
rect 20530 27860 20536 27872
rect 20128 27832 20536 27860
rect 20128 27820 20134 27832
rect 20530 27820 20536 27832
rect 20588 27820 20594 27872
rect 24118 27820 24124 27872
rect 24176 27820 24182 27872
rect 1104 27770 25852 27792
rect 1104 27718 2950 27770
rect 3002 27718 3014 27770
rect 3066 27718 3078 27770
rect 3130 27718 3142 27770
rect 3194 27718 3206 27770
rect 3258 27718 12950 27770
rect 13002 27718 13014 27770
rect 13066 27718 13078 27770
rect 13130 27718 13142 27770
rect 13194 27718 13206 27770
rect 13258 27718 22950 27770
rect 23002 27718 23014 27770
rect 23066 27718 23078 27770
rect 23130 27718 23142 27770
rect 23194 27718 23206 27770
rect 23258 27718 25852 27770
rect 1104 27696 25852 27718
rect 7650 27616 7656 27668
rect 7708 27656 7714 27668
rect 7708 27628 10916 27656
rect 7708 27616 7714 27628
rect 8389 27591 8447 27597
rect 7944 27560 8156 27588
rect 1302 27480 1308 27532
rect 1360 27520 1366 27532
rect 2041 27523 2099 27529
rect 2041 27520 2053 27523
rect 1360 27492 2053 27520
rect 1360 27480 1366 27492
rect 2041 27489 2053 27492
rect 2087 27489 2099 27523
rect 2041 27483 2099 27489
rect 2682 27480 2688 27532
rect 2740 27520 2746 27532
rect 3973 27523 4031 27529
rect 3973 27520 3985 27523
rect 2740 27492 3985 27520
rect 2740 27480 2746 27492
rect 3973 27489 3985 27492
rect 4019 27489 4031 27523
rect 3973 27483 4031 27489
rect 5534 27480 5540 27532
rect 5592 27520 5598 27532
rect 5813 27523 5871 27529
rect 5813 27520 5825 27523
rect 5592 27492 5825 27520
rect 5592 27480 5598 27492
rect 5813 27489 5825 27492
rect 5859 27520 5871 27523
rect 7944 27520 7972 27560
rect 5859 27492 7972 27520
rect 5859 27489 5871 27492
rect 5813 27483 5871 27489
rect 8018 27480 8024 27532
rect 8076 27480 8082 27532
rect 8128 27520 8156 27560
rect 8389 27557 8401 27591
rect 8435 27588 8447 27591
rect 8570 27588 8576 27600
rect 8435 27560 8576 27588
rect 8435 27557 8447 27560
rect 8389 27551 8447 27557
rect 8570 27548 8576 27560
rect 8628 27548 8634 27600
rect 10042 27548 10048 27600
rect 10100 27588 10106 27600
rect 10318 27588 10324 27600
rect 10100 27560 10324 27588
rect 10100 27548 10106 27560
rect 10318 27548 10324 27560
rect 10376 27548 10382 27600
rect 10888 27588 10916 27628
rect 10962 27616 10968 27668
rect 11020 27656 11026 27668
rect 11974 27656 11980 27668
rect 11020 27628 11980 27656
rect 11020 27616 11026 27628
rect 11974 27616 11980 27628
rect 12032 27616 12038 27668
rect 12342 27656 12348 27668
rect 12084 27628 12348 27656
rect 12084 27588 12112 27628
rect 12342 27616 12348 27628
rect 12400 27616 12406 27668
rect 19334 27616 19340 27668
rect 19392 27656 19398 27668
rect 19429 27659 19487 27665
rect 19429 27656 19441 27659
rect 19392 27628 19441 27656
rect 19392 27616 19398 27628
rect 19429 27625 19441 27628
rect 19475 27656 19487 27659
rect 19518 27656 19524 27668
rect 19475 27628 19524 27656
rect 19475 27625 19487 27628
rect 19429 27619 19487 27625
rect 19518 27616 19524 27628
rect 19576 27616 19582 27668
rect 20714 27656 20720 27668
rect 19904 27628 20720 27656
rect 10888 27560 12112 27588
rect 12176 27560 16620 27588
rect 12176 27520 12204 27560
rect 8128 27492 12204 27520
rect 12897 27523 12955 27529
rect 12897 27489 12909 27523
rect 12943 27520 12955 27523
rect 14550 27520 14556 27532
rect 12943 27492 14556 27520
rect 12943 27489 12955 27492
rect 12897 27483 12955 27489
rect 14550 27480 14556 27492
rect 14608 27480 14614 27532
rect 14829 27523 14887 27529
rect 14829 27489 14841 27523
rect 14875 27520 14887 27523
rect 16022 27520 16028 27532
rect 14875 27492 16028 27520
rect 14875 27489 14887 27492
rect 14829 27483 14887 27489
rect 16022 27480 16028 27492
rect 16080 27480 16086 27532
rect 16209 27523 16267 27529
rect 16209 27489 16221 27523
rect 16255 27520 16267 27523
rect 16592 27520 16620 27560
rect 16666 27548 16672 27600
rect 16724 27588 16730 27600
rect 18966 27588 18972 27600
rect 16724 27560 17356 27588
rect 16724 27548 16730 27560
rect 17328 27529 17356 27560
rect 18156 27560 18972 27588
rect 18156 27529 18184 27560
rect 18966 27548 18972 27560
rect 19024 27588 19030 27600
rect 19904 27588 19932 27628
rect 20714 27616 20720 27628
rect 20772 27616 20778 27668
rect 20919 27659 20977 27665
rect 20919 27625 20931 27659
rect 20965 27656 20977 27659
rect 21082 27656 21088 27668
rect 20965 27628 21088 27656
rect 20965 27625 20977 27628
rect 20919 27619 20977 27625
rect 21082 27616 21088 27628
rect 21140 27616 21146 27668
rect 19024 27560 19932 27588
rect 19024 27548 19030 27560
rect 23934 27548 23940 27600
rect 23992 27588 23998 27600
rect 24029 27591 24087 27597
rect 24029 27588 24041 27591
rect 23992 27560 24041 27588
rect 23992 27548 23998 27560
rect 24029 27557 24041 27560
rect 24075 27557 24087 27591
rect 24029 27551 24087 27557
rect 17313 27523 17371 27529
rect 16255 27492 16344 27520
rect 16592 27492 17264 27520
rect 16255 27489 16267 27492
rect 16209 27483 16267 27489
rect 1765 27455 1823 27461
rect 1765 27421 1777 27455
rect 1811 27452 1823 27455
rect 1946 27452 1952 27464
rect 1811 27424 1952 27452
rect 1811 27421 1823 27424
rect 1765 27415 1823 27421
rect 1946 27412 1952 27424
rect 2004 27412 2010 27464
rect 13081 27455 13139 27461
rect 13081 27421 13093 27455
rect 13127 27452 13139 27455
rect 13354 27452 13360 27464
rect 13127 27424 13360 27452
rect 13127 27421 13139 27424
rect 13081 27415 13139 27421
rect 13354 27412 13360 27424
rect 13412 27412 13418 27464
rect 14737 27455 14795 27461
rect 14737 27421 14749 27455
rect 14783 27452 14795 27455
rect 14918 27452 14924 27464
rect 14783 27424 14924 27452
rect 14783 27421 14795 27424
rect 14737 27415 14795 27421
rect 14918 27412 14924 27424
rect 14976 27412 14982 27464
rect 3970 27344 3976 27396
rect 4028 27384 4034 27396
rect 4157 27387 4215 27393
rect 4157 27384 4169 27387
rect 4028 27356 4169 27384
rect 4028 27344 4034 27356
rect 4157 27353 4169 27356
rect 4203 27353 4215 27387
rect 7466 27384 7472 27396
rect 7314 27356 7472 27384
rect 4157 27347 4215 27353
rect 7466 27344 7472 27356
rect 7524 27384 7530 27396
rect 7745 27387 7803 27393
rect 7524 27356 7696 27384
rect 7524 27344 7530 27356
rect 6273 27319 6331 27325
rect 6273 27285 6285 27319
rect 6319 27316 6331 27319
rect 6914 27316 6920 27328
rect 6319 27288 6920 27316
rect 6319 27285 6331 27288
rect 6273 27279 6331 27285
rect 6914 27276 6920 27288
rect 6972 27276 6978 27328
rect 7668 27316 7696 27356
rect 7745 27353 7757 27387
rect 7791 27384 7803 27387
rect 7834 27384 7840 27396
rect 7791 27356 7840 27384
rect 7791 27353 7803 27356
rect 7745 27347 7803 27353
rect 7834 27344 7840 27356
rect 7892 27344 7898 27396
rect 14645 27387 14703 27393
rect 14645 27384 14657 27387
rect 13464 27356 14657 27384
rect 8570 27316 8576 27328
rect 7668 27288 8576 27316
rect 8570 27276 8576 27288
rect 8628 27276 8634 27328
rect 10594 27276 10600 27328
rect 10652 27316 10658 27328
rect 10689 27319 10747 27325
rect 10689 27316 10701 27319
rect 10652 27288 10701 27316
rect 10652 27276 10658 27288
rect 10689 27285 10701 27288
rect 10735 27285 10747 27319
rect 10689 27279 10747 27285
rect 11514 27276 11520 27328
rect 11572 27316 11578 27328
rect 12345 27319 12403 27325
rect 12345 27316 12357 27319
rect 11572 27288 12357 27316
rect 11572 27276 11578 27288
rect 12345 27285 12357 27288
rect 12391 27316 12403 27319
rect 12434 27316 12440 27328
rect 12391 27288 12440 27316
rect 12391 27285 12403 27288
rect 12345 27279 12403 27285
rect 12434 27276 12440 27288
rect 12492 27316 12498 27328
rect 13464 27325 13492 27356
rect 14645 27353 14657 27356
rect 14691 27353 14703 27387
rect 16316 27384 16344 27492
rect 17034 27412 17040 27464
rect 17092 27452 17098 27464
rect 17129 27455 17187 27461
rect 17129 27452 17141 27455
rect 17092 27424 17141 27452
rect 17092 27412 17098 27424
rect 17129 27421 17141 27424
rect 17175 27421 17187 27455
rect 17236 27452 17264 27492
rect 17313 27489 17325 27523
rect 17359 27489 17371 27523
rect 17313 27483 17371 27489
rect 18141 27523 18199 27529
rect 18141 27489 18153 27523
rect 18187 27489 18199 27523
rect 18141 27483 18199 27489
rect 18233 27523 18291 27529
rect 18233 27489 18245 27523
rect 18279 27520 18291 27523
rect 19061 27523 19119 27529
rect 19061 27520 19073 27523
rect 18279 27492 19073 27520
rect 18279 27489 18291 27492
rect 18233 27483 18291 27489
rect 19061 27489 19073 27492
rect 19107 27520 19119 27523
rect 19242 27520 19248 27532
rect 19107 27492 19248 27520
rect 19107 27489 19119 27492
rect 19061 27483 19119 27489
rect 19242 27480 19248 27492
rect 19300 27480 19306 27532
rect 21545 27523 21603 27529
rect 21545 27520 21557 27523
rect 19812 27492 21557 27520
rect 19812 27464 19840 27492
rect 21545 27489 21557 27492
rect 21591 27520 21603 27523
rect 23566 27520 23572 27532
rect 21591 27492 23572 27520
rect 21591 27489 21603 27492
rect 21545 27483 21603 27489
rect 23566 27480 23572 27492
rect 23624 27480 23630 27532
rect 18046 27452 18052 27464
rect 17236 27424 18052 27452
rect 17129 27415 17187 27421
rect 18046 27412 18052 27424
rect 18104 27412 18110 27464
rect 18322 27412 18328 27464
rect 18380 27412 18386 27464
rect 19794 27412 19800 27464
rect 19852 27412 19858 27464
rect 21177 27455 21235 27461
rect 21177 27421 21189 27455
rect 21223 27452 21235 27455
rect 21450 27452 21456 27464
rect 21223 27424 21456 27452
rect 21223 27421 21235 27424
rect 21177 27415 21235 27421
rect 21450 27412 21456 27424
rect 21508 27452 21514 27464
rect 22278 27452 22284 27464
rect 21508 27424 22284 27452
rect 21508 27412 21514 27424
rect 22278 27412 22284 27424
rect 22336 27412 22342 27464
rect 24302 27412 24308 27464
rect 24360 27452 24366 27464
rect 24765 27455 24823 27461
rect 24765 27452 24777 27455
rect 24360 27424 24777 27452
rect 24360 27412 24366 27424
rect 24765 27421 24777 27424
rect 24811 27421 24823 27455
rect 24765 27415 24823 27421
rect 18340 27384 18368 27412
rect 22557 27387 22615 27393
rect 22557 27384 22569 27387
rect 14645 27347 14703 27353
rect 15488 27356 18368 27384
rect 21008 27356 22569 27384
rect 15488 27328 15516 27356
rect 12989 27319 13047 27325
rect 12989 27316 13001 27319
rect 12492 27288 13001 27316
rect 12492 27276 12498 27288
rect 12989 27285 13001 27288
rect 13035 27285 13047 27319
rect 12989 27279 13047 27285
rect 13449 27319 13507 27325
rect 13449 27285 13461 27319
rect 13495 27285 13507 27319
rect 13449 27279 13507 27285
rect 14274 27276 14280 27328
rect 14332 27276 14338 27328
rect 14458 27276 14464 27328
rect 14516 27316 14522 27328
rect 14826 27316 14832 27328
rect 14516 27288 14832 27316
rect 14516 27276 14522 27288
rect 14826 27276 14832 27288
rect 14884 27276 14890 27328
rect 15470 27276 15476 27328
rect 15528 27276 15534 27328
rect 15562 27276 15568 27328
rect 15620 27276 15626 27328
rect 15930 27276 15936 27328
rect 15988 27276 15994 27328
rect 16025 27319 16083 27325
rect 16025 27285 16037 27319
rect 16071 27316 16083 27319
rect 16482 27316 16488 27328
rect 16071 27288 16488 27316
rect 16071 27285 16083 27288
rect 16025 27279 16083 27285
rect 16482 27276 16488 27288
rect 16540 27276 16546 27328
rect 16758 27276 16764 27328
rect 16816 27276 16822 27328
rect 17218 27276 17224 27328
rect 17276 27276 17282 27328
rect 18325 27319 18383 27325
rect 18325 27285 18337 27319
rect 18371 27316 18383 27319
rect 18414 27316 18420 27328
rect 18371 27288 18420 27316
rect 18371 27285 18383 27288
rect 18325 27279 18383 27285
rect 18414 27276 18420 27288
rect 18472 27276 18478 27328
rect 18690 27276 18696 27328
rect 18748 27276 18754 27328
rect 20070 27276 20076 27328
rect 20128 27316 20134 27328
rect 21008 27316 21036 27356
rect 22557 27353 22569 27356
rect 22603 27384 22615 27387
rect 22830 27384 22836 27396
rect 22603 27356 22836 27384
rect 22603 27353 22615 27356
rect 22557 27347 22615 27353
rect 22830 27344 22836 27356
rect 22888 27344 22894 27396
rect 23782 27356 23888 27384
rect 20128 27288 21036 27316
rect 22848 27316 22876 27344
rect 23290 27316 23296 27328
rect 22848 27288 23296 27316
rect 20128 27276 20134 27288
rect 23290 27276 23296 27288
rect 23348 27276 23354 27328
rect 23566 27276 23572 27328
rect 23624 27316 23630 27328
rect 23860 27316 23888 27356
rect 23934 27344 23940 27396
rect 23992 27384 23998 27396
rect 24581 27387 24639 27393
rect 24581 27384 24593 27387
rect 23992 27356 24593 27384
rect 23992 27344 23998 27356
rect 24581 27353 24593 27356
rect 24627 27353 24639 27387
rect 24581 27347 24639 27353
rect 24394 27316 24400 27328
rect 23624 27288 24400 27316
rect 23624 27276 23630 27288
rect 24394 27276 24400 27288
rect 24452 27276 24458 27328
rect 1104 27226 25852 27248
rect 1104 27174 7950 27226
rect 8002 27174 8014 27226
rect 8066 27174 8078 27226
rect 8130 27174 8142 27226
rect 8194 27174 8206 27226
rect 8258 27174 17950 27226
rect 18002 27174 18014 27226
rect 18066 27174 18078 27226
rect 18130 27174 18142 27226
rect 18194 27174 18206 27226
rect 18258 27174 25852 27226
rect 1104 27152 25852 27174
rect 1762 27072 1768 27124
rect 1820 27112 1826 27124
rect 3510 27121 3516 27124
rect 2041 27115 2099 27121
rect 2041 27112 2053 27115
rect 1820 27084 2053 27112
rect 1820 27072 1826 27084
rect 2041 27081 2053 27084
rect 2087 27081 2099 27115
rect 2041 27075 2099 27081
rect 3467 27115 3516 27121
rect 3467 27081 3479 27115
rect 3513 27081 3516 27115
rect 3467 27075 3516 27081
rect 3510 27072 3516 27075
rect 3568 27072 3574 27124
rect 10321 27115 10379 27121
rect 10321 27081 10333 27115
rect 10367 27112 10379 27115
rect 10870 27112 10876 27124
rect 10367 27084 10876 27112
rect 10367 27081 10379 27084
rect 10321 27075 10379 27081
rect 10870 27072 10876 27084
rect 10928 27072 10934 27124
rect 15378 27112 15384 27124
rect 11716 27084 15384 27112
rect 5994 27004 6000 27056
rect 6052 27044 6058 27056
rect 11514 27044 11520 27056
rect 6052 27016 11520 27044
rect 6052 27004 6058 27016
rect 11514 27004 11520 27016
rect 11572 27004 11578 27056
rect 2222 26936 2228 26988
rect 2280 26936 2286 26988
rect 3326 26936 3332 26988
rect 3384 26985 3390 26988
rect 3384 26979 3422 26985
rect 3410 26945 3422 26979
rect 3384 26939 3422 26945
rect 3384 26936 3390 26939
rect 7190 26936 7196 26988
rect 7248 26976 7254 26988
rect 7837 26979 7895 26985
rect 7837 26976 7849 26979
rect 7248 26948 7849 26976
rect 7248 26936 7254 26948
rect 7837 26945 7849 26948
rect 7883 26945 7895 26979
rect 7837 26939 7895 26945
rect 7929 26979 7987 26985
rect 7929 26945 7941 26979
rect 7975 26976 7987 26979
rect 8662 26976 8668 26988
rect 7975 26948 8668 26976
rect 7975 26945 7987 26948
rect 7929 26939 7987 26945
rect 8662 26936 8668 26948
rect 8720 26936 8726 26988
rect 8846 26936 8852 26988
rect 8904 26976 8910 26988
rect 10413 26979 10471 26985
rect 10413 26976 10425 26979
rect 8904 26948 10425 26976
rect 8904 26936 8910 26948
rect 10413 26945 10425 26948
rect 10459 26945 10471 26979
rect 10413 26939 10471 26945
rect 7742 26868 7748 26920
rect 7800 26868 7806 26920
rect 8294 26868 8300 26920
rect 8352 26908 8358 26920
rect 8757 26911 8815 26917
rect 8757 26908 8769 26911
rect 8352 26880 8769 26908
rect 8352 26868 8358 26880
rect 8757 26877 8769 26880
rect 8803 26877 8815 26911
rect 8757 26871 8815 26877
rect 10137 26911 10195 26917
rect 10137 26877 10149 26911
rect 10183 26877 10195 26911
rect 10137 26871 10195 26877
rect 7282 26800 7288 26852
rect 7340 26840 7346 26852
rect 10152 26840 10180 26871
rect 10502 26868 10508 26920
rect 10560 26908 10566 26920
rect 11716 26917 11744 27084
rect 15378 27072 15384 27084
rect 15436 27072 15442 27124
rect 15746 27072 15752 27124
rect 15804 27072 15810 27124
rect 16298 27072 16304 27124
rect 16356 27112 16362 27124
rect 16356 27084 18368 27112
rect 16356 27072 16362 27084
rect 12526 27004 12532 27056
rect 12584 27004 12590 27056
rect 13814 27004 13820 27056
rect 13872 27004 13878 27056
rect 14918 27004 14924 27056
rect 14976 27044 14982 27056
rect 15105 27047 15163 27053
rect 15105 27044 15117 27047
rect 14976 27016 15117 27044
rect 14976 27004 14982 27016
rect 15105 27013 15117 27016
rect 15151 27044 15163 27047
rect 15764 27044 15792 27072
rect 17037 27047 17095 27053
rect 17037 27044 17049 27047
rect 15151 27016 17049 27044
rect 15151 27013 15163 27016
rect 15105 27007 15163 27013
rect 17037 27013 17049 27016
rect 17083 27044 17095 27047
rect 17773 27047 17831 27053
rect 17773 27044 17785 27047
rect 17083 27016 17785 27044
rect 17083 27013 17095 27016
rect 17037 27007 17095 27013
rect 17773 27013 17785 27016
rect 17819 27013 17831 27047
rect 18340 27044 18368 27084
rect 18414 27072 18420 27124
rect 18472 27072 18478 27124
rect 18598 27072 18604 27124
rect 18656 27112 18662 27124
rect 18693 27115 18751 27121
rect 18693 27112 18705 27115
rect 18656 27084 18705 27112
rect 18656 27072 18662 27084
rect 18693 27081 18705 27084
rect 18739 27112 18751 27115
rect 19242 27112 19248 27124
rect 18739 27084 19248 27112
rect 18739 27081 18751 27084
rect 18693 27075 18751 27081
rect 19242 27072 19248 27084
rect 19300 27072 19306 27124
rect 22278 27072 22284 27124
rect 22336 27112 22342 27124
rect 22336 27084 23980 27112
rect 22336 27072 22342 27084
rect 20346 27044 20352 27056
rect 18340 27016 20352 27044
rect 17773 27007 17831 27013
rect 20346 27004 20352 27016
rect 20404 27004 20410 27056
rect 23566 27044 23572 27056
rect 23230 27016 23572 27044
rect 23566 27004 23572 27016
rect 23624 27004 23630 27056
rect 13446 26936 13452 26988
rect 13504 26936 13510 26988
rect 15013 26979 15071 26985
rect 15013 26945 15025 26979
rect 15059 26976 15071 26979
rect 15059 26948 15424 26976
rect 15059 26945 15071 26948
rect 15013 26939 15071 26945
rect 11701 26911 11759 26917
rect 11701 26908 11713 26911
rect 10560 26880 11713 26908
rect 10560 26868 10566 26880
rect 11701 26877 11713 26880
rect 11747 26877 11759 26911
rect 11701 26871 11759 26877
rect 11974 26868 11980 26920
rect 12032 26908 12038 26920
rect 12526 26908 12532 26920
rect 12032 26880 12532 26908
rect 12032 26868 12038 26880
rect 12526 26868 12532 26880
rect 12584 26868 12590 26920
rect 12802 26868 12808 26920
rect 12860 26908 12866 26920
rect 13173 26911 13231 26917
rect 13173 26908 13185 26911
rect 12860 26880 13185 26908
rect 12860 26868 12866 26880
rect 13173 26877 13185 26880
rect 13219 26877 13231 26911
rect 13173 26871 13231 26877
rect 15197 26911 15255 26917
rect 15197 26877 15209 26911
rect 15243 26877 15255 26911
rect 15197 26871 15255 26877
rect 7340 26812 10180 26840
rect 7340 26800 7346 26812
rect 13630 26800 13636 26852
rect 13688 26840 13694 26852
rect 15212 26840 15240 26871
rect 13688 26812 15240 26840
rect 13688 26800 13694 26812
rect 7190 26732 7196 26784
rect 7248 26732 7254 26784
rect 8297 26775 8355 26781
rect 8297 26741 8309 26775
rect 8343 26772 8355 26775
rect 10318 26772 10324 26784
rect 8343 26744 10324 26772
rect 8343 26741 8355 26744
rect 8297 26735 8355 26741
rect 10318 26732 10324 26744
rect 10376 26732 10382 26784
rect 10781 26775 10839 26781
rect 10781 26741 10793 26775
rect 10827 26772 10839 26775
rect 11514 26772 11520 26784
rect 10827 26744 11520 26772
rect 10827 26741 10839 26744
rect 10781 26735 10839 26741
rect 11514 26732 11520 26744
rect 11572 26732 11578 26784
rect 14642 26732 14648 26784
rect 14700 26732 14706 26784
rect 15396 26772 15424 26948
rect 15930 26936 15936 26988
rect 15988 26976 15994 26988
rect 16390 26976 16396 26988
rect 15988 26948 16396 26976
rect 15988 26936 15994 26948
rect 16390 26936 16396 26948
rect 16448 26936 16454 26988
rect 17310 26936 17316 26988
rect 17368 26976 17374 26988
rect 17681 26979 17739 26985
rect 17681 26976 17693 26979
rect 17368 26948 17693 26976
rect 17368 26936 17374 26948
rect 17681 26945 17693 26948
rect 17727 26976 17739 26979
rect 18598 26976 18604 26988
rect 17727 26948 18604 26976
rect 17727 26945 17739 26948
rect 17681 26939 17739 26945
rect 18598 26936 18604 26948
rect 18656 26936 18662 26988
rect 23952 26985 23980 27084
rect 25406 27072 25412 27124
rect 25464 27072 25470 27124
rect 24762 27004 24768 27056
rect 24820 27004 24826 27056
rect 23937 26979 23995 26985
rect 23937 26945 23949 26979
rect 23983 26945 23995 26979
rect 23937 26939 23995 26945
rect 15470 26800 15476 26852
rect 15528 26840 15534 26852
rect 15948 26840 15976 26936
rect 17589 26911 17647 26917
rect 17589 26877 17601 26911
rect 17635 26877 17647 26911
rect 17589 26871 17647 26877
rect 15528 26812 15976 26840
rect 15528 26800 15534 26812
rect 17402 26800 17408 26852
rect 17460 26840 17466 26852
rect 17604 26840 17632 26871
rect 18782 26868 18788 26920
rect 18840 26908 18846 26920
rect 22189 26911 22247 26917
rect 22189 26908 22201 26911
rect 18840 26880 22201 26908
rect 18840 26868 18846 26880
rect 22189 26877 22201 26880
rect 22235 26877 22247 26911
rect 22189 26871 22247 26877
rect 23661 26911 23719 26917
rect 23661 26877 23673 26911
rect 23707 26908 23719 26911
rect 24854 26908 24860 26920
rect 23707 26880 24860 26908
rect 23707 26877 23719 26880
rect 23661 26871 23719 26877
rect 24854 26868 24860 26880
rect 24912 26868 24918 26920
rect 19886 26840 19892 26852
rect 17460 26812 19892 26840
rect 17460 26800 17466 26812
rect 19886 26800 19892 26812
rect 19944 26800 19950 26852
rect 24302 26800 24308 26852
rect 24360 26840 24366 26852
rect 24581 26843 24639 26849
rect 24581 26840 24593 26843
rect 24360 26812 24593 26840
rect 24360 26800 24366 26812
rect 24581 26809 24593 26812
rect 24627 26809 24639 26843
rect 24581 26803 24639 26809
rect 15841 26775 15899 26781
rect 15841 26772 15853 26775
rect 15396 26744 15853 26772
rect 15841 26741 15853 26744
rect 15887 26772 15899 26775
rect 16298 26772 16304 26784
rect 15887 26744 16304 26772
rect 15887 26741 15899 26744
rect 15841 26735 15899 26741
rect 16298 26732 16304 26744
rect 16356 26732 16362 26784
rect 16482 26732 16488 26784
rect 16540 26772 16546 26784
rect 16669 26775 16727 26781
rect 16669 26772 16681 26775
rect 16540 26744 16681 26772
rect 16540 26732 16546 26744
rect 16669 26741 16681 26744
rect 16715 26741 16727 26775
rect 16669 26735 16727 26741
rect 18141 26775 18199 26781
rect 18141 26741 18153 26775
rect 18187 26772 18199 26775
rect 18322 26772 18328 26784
rect 18187 26744 18328 26772
rect 18187 26741 18199 26744
rect 18141 26735 18199 26741
rect 18322 26732 18328 26744
rect 18380 26732 18386 26784
rect 24213 26775 24271 26781
rect 24213 26741 24225 26775
rect 24259 26772 24271 26775
rect 24394 26772 24400 26784
rect 24259 26744 24400 26772
rect 24259 26741 24271 26744
rect 24213 26735 24271 26741
rect 24394 26732 24400 26744
rect 24452 26772 24458 26784
rect 25133 26775 25191 26781
rect 25133 26772 25145 26775
rect 24452 26744 25145 26772
rect 24452 26732 24458 26744
rect 25133 26741 25145 26744
rect 25179 26741 25191 26775
rect 25133 26735 25191 26741
rect 1104 26682 25852 26704
rect 1104 26630 2950 26682
rect 3002 26630 3014 26682
rect 3066 26630 3078 26682
rect 3130 26630 3142 26682
rect 3194 26630 3206 26682
rect 3258 26630 12950 26682
rect 13002 26630 13014 26682
rect 13066 26630 13078 26682
rect 13130 26630 13142 26682
rect 13194 26630 13206 26682
rect 13258 26630 22950 26682
rect 23002 26630 23014 26682
rect 23066 26630 23078 26682
rect 23130 26630 23142 26682
rect 23194 26630 23206 26682
rect 23258 26630 25852 26682
rect 1104 26608 25852 26630
rect 7650 26528 7656 26580
rect 7708 26568 7714 26580
rect 8021 26571 8079 26577
rect 8021 26568 8033 26571
rect 7708 26540 8033 26568
rect 7708 26528 7714 26540
rect 8021 26537 8033 26540
rect 8067 26537 8079 26571
rect 8021 26531 8079 26537
rect 8389 26571 8447 26577
rect 8389 26537 8401 26571
rect 8435 26568 8447 26571
rect 8570 26568 8576 26580
rect 8435 26540 8576 26568
rect 8435 26537 8447 26540
rect 8389 26531 8447 26537
rect 2590 26392 2596 26444
rect 2648 26432 2654 26444
rect 3973 26435 4031 26441
rect 3973 26432 3985 26435
rect 2648 26404 3985 26432
rect 2648 26392 2654 26404
rect 3973 26401 3985 26404
rect 4019 26401 4031 26435
rect 3973 26395 4031 26401
rect 5813 26435 5871 26441
rect 5813 26401 5825 26435
rect 5859 26432 5871 26435
rect 5994 26432 6000 26444
rect 5859 26404 6000 26432
rect 5859 26401 5871 26404
rect 5813 26395 5871 26401
rect 5994 26392 6000 26404
rect 6052 26392 6058 26444
rect 6270 26392 6276 26444
rect 6328 26392 6334 26444
rect 6549 26435 6607 26441
rect 6549 26401 6561 26435
rect 6595 26432 6607 26435
rect 6914 26432 6920 26444
rect 6595 26404 6920 26432
rect 6595 26401 6607 26404
rect 6549 26395 6607 26401
rect 6914 26392 6920 26404
rect 6972 26432 6978 26444
rect 7834 26432 7840 26444
rect 6972 26404 7840 26432
rect 6972 26392 6978 26404
rect 7834 26392 7840 26404
rect 7892 26392 7898 26444
rect 8404 26376 8432 26531
rect 8570 26528 8576 26540
rect 8628 26568 8634 26580
rect 11974 26568 11980 26580
rect 8628 26540 11980 26568
rect 8628 26528 8634 26540
rect 11974 26528 11980 26540
rect 12032 26528 12038 26580
rect 13906 26528 13912 26580
rect 13964 26568 13970 26580
rect 15010 26568 15016 26580
rect 13964 26540 15016 26568
rect 13964 26528 13970 26540
rect 15010 26528 15016 26540
rect 15068 26568 15074 26580
rect 15930 26568 15936 26580
rect 15068 26540 15936 26568
rect 15068 26528 15074 26540
rect 15930 26528 15936 26540
rect 15988 26528 15994 26580
rect 16022 26528 16028 26580
rect 16080 26568 16086 26580
rect 16206 26568 16212 26580
rect 16080 26540 16212 26568
rect 16080 26528 16086 26540
rect 16206 26528 16212 26540
rect 16264 26568 16270 26580
rect 16301 26571 16359 26577
rect 16301 26568 16313 26571
rect 16264 26540 16313 26568
rect 16264 26528 16270 26540
rect 16301 26537 16313 26540
rect 16347 26537 16359 26571
rect 16301 26531 16359 26537
rect 16482 26528 16488 26580
rect 16540 26568 16546 26580
rect 20533 26571 20591 26577
rect 16540 26540 20484 26568
rect 16540 26528 16546 26540
rect 10965 26503 11023 26509
rect 10965 26469 10977 26503
rect 11011 26500 11023 26503
rect 13541 26503 13599 26509
rect 11011 26472 13216 26500
rect 11011 26469 11023 26472
rect 10965 26463 11023 26469
rect 10413 26435 10471 26441
rect 10413 26401 10425 26435
rect 10459 26432 10471 26435
rect 10502 26432 10508 26444
rect 10459 26404 10508 26432
rect 10459 26401 10471 26404
rect 10413 26395 10471 26401
rect 10502 26392 10508 26404
rect 10560 26392 10566 26444
rect 12618 26392 12624 26444
rect 12676 26432 12682 26444
rect 12897 26435 12955 26441
rect 12897 26432 12909 26435
rect 12676 26404 12909 26432
rect 12676 26392 12682 26404
rect 12897 26401 12909 26404
rect 12943 26401 12955 26435
rect 12897 26395 12955 26401
rect 8386 26364 8392 26376
rect 7682 26336 8392 26364
rect 8386 26324 8392 26336
rect 8444 26324 8450 26376
rect 9030 26324 9036 26376
rect 9088 26364 9094 26376
rect 9125 26367 9183 26373
rect 9125 26364 9137 26367
rect 9088 26336 9137 26364
rect 9088 26324 9094 26336
rect 9125 26333 9137 26336
rect 9171 26364 9183 26367
rect 9171 26336 9628 26364
rect 9171 26333 9183 26336
rect 9125 26327 9183 26333
rect 3878 26256 3884 26308
rect 3936 26296 3942 26308
rect 4157 26299 4215 26305
rect 4157 26296 4169 26299
rect 3936 26268 4169 26296
rect 3936 26256 3942 26268
rect 4157 26265 4169 26268
rect 4203 26265 4215 26299
rect 4157 26259 4215 26265
rect 8570 26256 8576 26308
rect 8628 26296 8634 26308
rect 9493 26299 9551 26305
rect 9493 26296 9505 26299
rect 8628 26268 9505 26296
rect 8628 26256 8634 26268
rect 9493 26265 9505 26268
rect 9539 26265 9551 26299
rect 9600 26296 9628 26336
rect 9674 26324 9680 26376
rect 9732 26324 9738 26376
rect 10594 26324 10600 26376
rect 10652 26324 10658 26376
rect 13188 26373 13216 26472
rect 13541 26469 13553 26503
rect 13587 26500 13599 26503
rect 13722 26500 13728 26512
rect 13587 26472 13728 26500
rect 13587 26469 13599 26472
rect 13541 26463 13599 26469
rect 13722 26460 13728 26472
rect 13780 26460 13786 26512
rect 18141 26503 18199 26509
rect 18141 26469 18153 26503
rect 18187 26500 18199 26503
rect 19518 26500 19524 26512
rect 18187 26472 19524 26500
rect 18187 26469 18199 26472
rect 18141 26463 18199 26469
rect 19518 26460 19524 26472
rect 19576 26460 19582 26512
rect 20456 26500 20484 26540
rect 20533 26537 20545 26571
rect 20579 26568 20591 26571
rect 22830 26568 22836 26580
rect 20579 26540 22836 26568
rect 20579 26537 20591 26540
rect 20533 26531 20591 26537
rect 22830 26528 22836 26540
rect 22888 26528 22894 26580
rect 23201 26571 23259 26577
rect 23201 26537 23213 26571
rect 23247 26568 23259 26571
rect 23290 26568 23296 26580
rect 23247 26540 23296 26568
rect 23247 26537 23259 26540
rect 23201 26531 23259 26537
rect 23290 26528 23296 26540
rect 23348 26528 23354 26580
rect 20806 26500 20812 26512
rect 20456 26472 20812 26500
rect 20806 26460 20812 26472
rect 20864 26460 20870 26512
rect 23845 26503 23903 26509
rect 23845 26469 23857 26503
rect 23891 26469 23903 26503
rect 23845 26463 23903 26469
rect 13556 26404 17540 26432
rect 13556 26376 13584 26404
rect 13173 26367 13231 26373
rect 13173 26333 13185 26367
rect 13219 26333 13231 26367
rect 13173 26327 13231 26333
rect 13538 26324 13544 26376
rect 13596 26324 13602 26376
rect 14550 26324 14556 26376
rect 14608 26324 14614 26376
rect 15930 26324 15936 26376
rect 15988 26364 15994 26376
rect 16577 26367 16635 26373
rect 16577 26364 16589 26367
rect 15988 26336 16589 26364
rect 15988 26324 15994 26336
rect 16577 26333 16589 26336
rect 16623 26364 16635 26367
rect 16666 26364 16672 26376
rect 16623 26336 16672 26364
rect 16623 26333 16635 26336
rect 16577 26327 16635 26333
rect 16666 26324 16672 26336
rect 16724 26324 16730 26376
rect 17512 26364 17540 26404
rect 17586 26392 17592 26444
rect 17644 26432 17650 26444
rect 18598 26432 18604 26444
rect 17644 26404 18604 26432
rect 17644 26392 17650 26404
rect 18598 26392 18604 26404
rect 18656 26392 18662 26444
rect 19981 26435 20039 26441
rect 19981 26401 19993 26435
rect 20027 26432 20039 26435
rect 20070 26432 20076 26444
rect 20027 26404 20076 26432
rect 20027 26401 20039 26404
rect 19981 26395 20039 26401
rect 20070 26392 20076 26404
rect 20128 26392 20134 26444
rect 23860 26432 23888 26463
rect 24394 26460 24400 26512
rect 24452 26500 24458 26512
rect 24670 26500 24676 26512
rect 24452 26472 24676 26500
rect 24452 26460 24458 26472
rect 24670 26460 24676 26472
rect 24728 26500 24734 26512
rect 25133 26503 25191 26509
rect 25133 26500 25145 26503
rect 24728 26472 25145 26500
rect 24728 26460 24734 26472
rect 25133 26469 25145 26472
rect 25179 26469 25191 26503
rect 25133 26463 25191 26469
rect 25406 26432 25412 26444
rect 20180 26404 23888 26432
rect 24044 26404 25412 26432
rect 17681 26367 17739 26373
rect 17681 26364 17693 26367
rect 17512 26336 17693 26364
rect 17681 26333 17693 26336
rect 17727 26364 17739 26367
rect 20180 26364 20208 26404
rect 17727 26336 20208 26364
rect 17727 26333 17739 26336
rect 17681 26327 17739 26333
rect 21450 26324 21456 26376
rect 21508 26324 21514 26376
rect 24044 26373 24072 26404
rect 25406 26392 25412 26404
rect 25464 26392 25470 26444
rect 24029 26367 24087 26373
rect 24029 26333 24041 26367
rect 24075 26333 24087 26367
rect 24029 26327 24087 26333
rect 24486 26324 24492 26376
rect 24544 26364 24550 26376
rect 24673 26367 24731 26373
rect 24673 26364 24685 26367
rect 24544 26336 24685 26364
rect 24544 26324 24550 26336
rect 24673 26333 24685 26336
rect 24719 26333 24731 26367
rect 24673 26327 24731 26333
rect 10042 26296 10048 26308
rect 9600 26268 10048 26296
rect 9493 26259 9551 26265
rect 10042 26256 10048 26268
rect 10100 26296 10106 26308
rect 10505 26299 10563 26305
rect 10505 26296 10517 26299
rect 10100 26268 10517 26296
rect 10100 26256 10106 26268
rect 10505 26265 10517 26268
rect 10551 26265 10563 26299
rect 10505 26259 10563 26265
rect 13081 26299 13139 26305
rect 13081 26265 13093 26299
rect 13127 26296 13139 26299
rect 14458 26296 14464 26308
rect 13127 26268 14464 26296
rect 13127 26265 13139 26268
rect 13081 26259 13139 26265
rect 14458 26256 14464 26268
rect 14516 26256 14522 26308
rect 14829 26299 14887 26305
rect 14829 26265 14841 26299
rect 14875 26296 14887 26299
rect 17034 26296 17040 26308
rect 14875 26268 15056 26296
rect 14875 26265 14887 26268
rect 14829 26259 14887 26265
rect 15028 26228 15056 26268
rect 16132 26268 17040 26296
rect 16132 26228 16160 26268
rect 17034 26256 17040 26268
rect 17092 26256 17098 26308
rect 17126 26256 17132 26308
rect 17184 26296 17190 26308
rect 17773 26299 17831 26305
rect 17773 26296 17785 26299
rect 17184 26268 17785 26296
rect 17184 26256 17190 26268
rect 17773 26265 17785 26268
rect 17819 26265 17831 26299
rect 17773 26259 17831 26265
rect 19429 26299 19487 26305
rect 19429 26265 19441 26299
rect 19475 26265 19487 26299
rect 19429 26259 19487 26265
rect 15028 26200 16160 26228
rect 16298 26188 16304 26240
rect 16356 26228 16362 26240
rect 19444 26228 19472 26259
rect 19702 26256 19708 26308
rect 19760 26296 19766 26308
rect 20073 26299 20131 26305
rect 20073 26296 20085 26299
rect 19760 26268 20085 26296
rect 19760 26256 19766 26268
rect 20073 26265 20085 26268
rect 20119 26265 20131 26299
rect 20073 26259 20131 26265
rect 20165 26299 20223 26305
rect 20165 26265 20177 26299
rect 20211 26265 20223 26299
rect 20165 26259 20223 26265
rect 20180 26228 20208 26259
rect 21726 26256 21732 26308
rect 21784 26256 21790 26308
rect 23106 26296 23112 26308
rect 22954 26268 23112 26296
rect 23106 26256 23112 26268
rect 23164 26296 23170 26308
rect 23566 26296 23572 26308
rect 23164 26268 23572 26296
rect 23164 26256 23170 26268
rect 23566 26256 23572 26268
rect 23624 26256 23630 26308
rect 24857 26299 24915 26305
rect 24857 26265 24869 26299
rect 24903 26296 24915 26299
rect 25222 26296 25228 26308
rect 24903 26268 25228 26296
rect 24903 26265 24915 26268
rect 24857 26259 24915 26265
rect 25222 26256 25228 26268
rect 25280 26256 25286 26308
rect 16356 26200 20208 26228
rect 16356 26188 16362 26200
rect 1104 26138 25852 26160
rect 1104 26086 7950 26138
rect 8002 26086 8014 26138
rect 8066 26086 8078 26138
rect 8130 26086 8142 26138
rect 8194 26086 8206 26138
rect 8258 26086 17950 26138
rect 18002 26086 18014 26138
rect 18066 26086 18078 26138
rect 18130 26086 18142 26138
rect 18194 26086 18206 26138
rect 18258 26086 25852 26138
rect 1104 26064 25852 26086
rect 2222 25984 2228 26036
rect 2280 26024 2286 26036
rect 2593 26027 2651 26033
rect 2593 26024 2605 26027
rect 2280 25996 2605 26024
rect 2280 25984 2286 25996
rect 2593 25993 2605 25996
rect 2639 25993 2651 26027
rect 2593 25987 2651 25993
rect 3835 26027 3893 26033
rect 3835 25993 3847 26027
rect 3881 26024 3893 26027
rect 4062 26024 4068 26036
rect 3881 25996 4068 26024
rect 3881 25993 3893 25996
rect 3835 25987 3893 25993
rect 4062 25984 4068 25996
rect 4120 25984 4126 26036
rect 7837 26027 7895 26033
rect 7837 25993 7849 26027
rect 7883 26024 7895 26027
rect 8294 26024 8300 26036
rect 7883 25996 8300 26024
rect 7883 25993 7895 25996
rect 7837 25987 7895 25993
rect 8294 25984 8300 25996
rect 8352 25984 8358 26036
rect 8662 25984 8668 26036
rect 8720 25984 8726 26036
rect 10318 25984 10324 26036
rect 10376 25984 10382 26036
rect 13906 25984 13912 26036
rect 13964 25984 13970 26036
rect 18690 25984 18696 26036
rect 18748 26024 18754 26036
rect 19705 26027 19763 26033
rect 19705 26024 19717 26027
rect 18748 25996 19717 26024
rect 18748 25984 18754 25996
rect 19705 25993 19717 25996
rect 19751 25993 19763 26027
rect 19705 25987 19763 25993
rect 22373 26027 22431 26033
rect 22373 25993 22385 26027
rect 22419 26024 22431 26027
rect 23382 26024 23388 26036
rect 22419 25996 23388 26024
rect 22419 25993 22431 25996
rect 22373 25987 22431 25993
rect 23382 25984 23388 25996
rect 23440 25984 23446 26036
rect 10229 25959 10287 25965
rect 10229 25925 10241 25959
rect 10275 25956 10287 25959
rect 10410 25956 10416 25968
rect 10275 25928 10416 25956
rect 10275 25925 10287 25928
rect 10229 25919 10287 25925
rect 10410 25916 10416 25928
rect 10468 25916 10474 25968
rect 11974 25916 11980 25968
rect 12032 25956 12038 25968
rect 12032 25928 12098 25956
rect 12032 25916 12038 25928
rect 13262 25916 13268 25968
rect 13320 25956 13326 25968
rect 13320 25928 13584 25956
rect 13320 25916 13326 25928
rect 13556 25900 13584 25928
rect 16666 25916 16672 25968
rect 16724 25956 16730 25968
rect 16724 25928 17710 25956
rect 16724 25916 16730 25928
rect 19610 25916 19616 25968
rect 19668 25916 19674 25968
rect 22462 25916 22468 25968
rect 22520 25916 22526 25968
rect 22646 25916 22652 25968
rect 22704 25956 22710 25968
rect 23106 25956 23112 25968
rect 22704 25928 23112 25956
rect 22704 25916 22710 25928
rect 23106 25916 23112 25928
rect 23164 25916 23170 25968
rect 23566 25916 23572 25968
rect 23624 25916 23630 25968
rect 24026 25916 24032 25968
rect 24084 25956 24090 25968
rect 24305 25959 24363 25965
rect 24305 25956 24317 25959
rect 24084 25928 24317 25956
rect 24084 25916 24090 25928
rect 24305 25925 24317 25928
rect 24351 25925 24363 25959
rect 24305 25919 24363 25925
rect 25038 25916 25044 25968
rect 25096 25916 25102 25968
rect 2866 25848 2872 25900
rect 2924 25888 2930 25900
rect 3732 25891 3790 25897
rect 3732 25888 3744 25891
rect 2924 25860 3744 25888
rect 2924 25848 2930 25860
rect 3732 25857 3744 25860
rect 3778 25857 3790 25891
rect 3732 25851 3790 25857
rect 13538 25848 13544 25900
rect 13596 25848 13602 25900
rect 13906 25848 13912 25900
rect 13964 25888 13970 25900
rect 14182 25888 14188 25900
rect 13964 25860 14188 25888
rect 13964 25848 13970 25860
rect 14182 25848 14188 25860
rect 14240 25848 14246 25900
rect 20993 25891 21051 25897
rect 20993 25857 21005 25891
rect 21039 25888 21051 25891
rect 21453 25891 21511 25897
rect 21453 25888 21465 25891
rect 21039 25860 21465 25888
rect 21039 25857 21051 25860
rect 20993 25851 21051 25857
rect 21453 25857 21465 25860
rect 21499 25888 21511 25891
rect 22278 25888 22284 25900
rect 21499 25860 22284 25888
rect 21499 25857 21511 25860
rect 21453 25851 21511 25857
rect 22278 25848 22284 25860
rect 22336 25848 22342 25900
rect 22480 25888 22508 25916
rect 25409 25891 25467 25897
rect 25409 25888 25421 25891
rect 22480 25860 25421 25888
rect 25409 25857 25421 25860
rect 25455 25857 25467 25891
rect 25409 25851 25467 25857
rect 3053 25823 3111 25829
rect 3053 25789 3065 25823
rect 3099 25789 3111 25823
rect 3053 25783 3111 25789
rect 3237 25823 3295 25829
rect 3237 25789 3249 25823
rect 3283 25820 3295 25823
rect 4246 25820 4252 25832
rect 3283 25792 4252 25820
rect 3283 25789 3295 25792
rect 3237 25783 3295 25789
rect 3068 25752 3096 25783
rect 4246 25780 4252 25792
rect 4304 25780 4310 25832
rect 7558 25780 7564 25832
rect 7616 25780 7622 25832
rect 7745 25823 7803 25829
rect 7745 25789 7757 25823
rect 7791 25789 7803 25823
rect 7745 25783 7803 25789
rect 3326 25752 3332 25764
rect 3068 25724 3332 25752
rect 3326 25712 3332 25724
rect 3384 25712 3390 25764
rect 7760 25752 7788 25783
rect 7834 25780 7840 25832
rect 7892 25820 7898 25832
rect 10045 25823 10103 25829
rect 10045 25820 10057 25823
rect 7892 25792 10057 25820
rect 7892 25780 7898 25792
rect 10045 25789 10057 25792
rect 10091 25789 10103 25823
rect 10045 25783 10103 25789
rect 12618 25780 12624 25832
rect 12676 25820 12682 25832
rect 13265 25823 13323 25829
rect 13265 25820 13277 25823
rect 12676 25792 13277 25820
rect 12676 25780 12682 25792
rect 13265 25789 13277 25792
rect 13311 25820 13323 25823
rect 13630 25820 13636 25832
rect 13311 25792 13636 25820
rect 13311 25789 13323 25792
rect 13265 25783 13323 25789
rect 13630 25780 13636 25792
rect 13688 25780 13694 25832
rect 16942 25780 16948 25832
rect 17000 25780 17006 25832
rect 17218 25780 17224 25832
rect 17276 25780 17282 25832
rect 18598 25780 18604 25832
rect 18656 25820 18662 25832
rect 18693 25823 18751 25829
rect 18693 25820 18705 25823
rect 18656 25792 18705 25820
rect 18656 25780 18662 25792
rect 18693 25789 18705 25792
rect 18739 25789 18751 25823
rect 18693 25783 18751 25789
rect 19889 25823 19947 25829
rect 19889 25789 19901 25823
rect 19935 25820 19947 25823
rect 20162 25820 20168 25832
rect 19935 25792 20168 25820
rect 19935 25789 19947 25792
rect 19889 25783 19947 25789
rect 20162 25780 20168 25792
rect 20220 25780 20226 25832
rect 20438 25780 20444 25832
rect 20496 25780 20502 25832
rect 22554 25780 22560 25832
rect 22612 25780 22618 25832
rect 23385 25823 23443 25829
rect 23385 25820 23397 25823
rect 22664 25792 23397 25820
rect 7116 25724 7788 25752
rect 8205 25755 8263 25761
rect 4706 25644 4712 25696
rect 4764 25684 4770 25696
rect 7006 25684 7012 25696
rect 4764 25656 7012 25684
rect 4764 25644 4770 25656
rect 7006 25644 7012 25656
rect 7064 25684 7070 25696
rect 7116 25693 7144 25724
rect 8205 25721 8217 25755
rect 8251 25752 8263 25755
rect 8846 25752 8852 25764
rect 8251 25724 8852 25752
rect 8251 25721 8263 25724
rect 8205 25715 8263 25721
rect 8846 25712 8852 25724
rect 8904 25712 8910 25764
rect 18506 25712 18512 25764
rect 18564 25752 18570 25764
rect 21269 25755 21327 25761
rect 21269 25752 21281 25755
rect 18564 25724 21281 25752
rect 18564 25712 18570 25724
rect 21269 25721 21281 25724
rect 21315 25721 21327 25755
rect 21269 25715 21327 25721
rect 22278 25712 22284 25764
rect 22336 25752 22342 25764
rect 22664 25752 22692 25792
rect 23385 25789 23397 25792
rect 23431 25789 23443 25823
rect 23385 25783 23443 25789
rect 22336 25724 22692 25752
rect 22336 25712 22342 25724
rect 23290 25712 23296 25764
rect 23348 25752 23354 25764
rect 24121 25755 24179 25761
rect 24121 25752 24133 25755
rect 23348 25724 24133 25752
rect 23348 25712 23354 25724
rect 24121 25721 24133 25724
rect 24167 25721 24179 25755
rect 24121 25715 24179 25721
rect 24762 25712 24768 25764
rect 24820 25752 24826 25764
rect 24857 25755 24915 25761
rect 24857 25752 24869 25755
rect 24820 25724 24869 25752
rect 24820 25712 24826 25724
rect 24857 25721 24869 25724
rect 24903 25721 24915 25755
rect 24857 25715 24915 25721
rect 7101 25687 7159 25693
rect 7101 25684 7113 25687
rect 7064 25656 7113 25684
rect 7064 25644 7070 25656
rect 7101 25653 7113 25656
rect 7147 25653 7159 25687
rect 7101 25647 7159 25653
rect 10689 25687 10747 25693
rect 10689 25653 10701 25687
rect 10735 25684 10747 25687
rect 11698 25684 11704 25696
rect 10735 25656 11704 25684
rect 10735 25653 10747 25656
rect 10689 25647 10747 25653
rect 11698 25644 11704 25656
rect 11756 25644 11762 25696
rect 11793 25687 11851 25693
rect 11793 25653 11805 25687
rect 11839 25684 11851 25687
rect 12802 25684 12808 25696
rect 11839 25656 12808 25684
rect 11839 25653 11851 25656
rect 11793 25647 11851 25653
rect 12802 25644 12808 25656
rect 12860 25684 12866 25696
rect 13446 25684 13452 25696
rect 12860 25656 13452 25684
rect 12860 25644 12866 25656
rect 13446 25644 13452 25656
rect 13504 25644 13510 25696
rect 16114 25644 16120 25696
rect 16172 25684 16178 25696
rect 16298 25684 16304 25696
rect 16172 25656 16304 25684
rect 16172 25644 16178 25656
rect 16298 25644 16304 25656
rect 16356 25644 16362 25696
rect 18782 25644 18788 25696
rect 18840 25684 18846 25696
rect 19245 25687 19303 25693
rect 19245 25684 19257 25687
rect 18840 25656 19257 25684
rect 18840 25644 18846 25656
rect 19245 25653 19257 25656
rect 19291 25653 19303 25687
rect 19245 25647 19303 25653
rect 21542 25644 21548 25696
rect 21600 25684 21606 25696
rect 22005 25687 22063 25693
rect 22005 25684 22017 25687
rect 21600 25656 22017 25684
rect 21600 25644 21606 25656
rect 22005 25653 22017 25656
rect 22051 25653 22063 25687
rect 22005 25647 22063 25653
rect 1104 25594 25852 25616
rect 1104 25542 2950 25594
rect 3002 25542 3014 25594
rect 3066 25542 3078 25594
rect 3130 25542 3142 25594
rect 3194 25542 3206 25594
rect 3258 25542 12950 25594
rect 13002 25542 13014 25594
rect 13066 25542 13078 25594
rect 13130 25542 13142 25594
rect 13194 25542 13206 25594
rect 13258 25542 22950 25594
rect 23002 25542 23014 25594
rect 23066 25542 23078 25594
rect 23130 25542 23142 25594
rect 23194 25542 23206 25594
rect 23258 25542 25852 25594
rect 1104 25520 25852 25542
rect 3602 25440 3608 25492
rect 3660 25440 3666 25492
rect 4154 25440 4160 25492
rect 4212 25440 4218 25492
rect 16114 25480 16120 25492
rect 6012 25452 16120 25480
rect 6012 25356 6040 25452
rect 16114 25440 16120 25452
rect 16172 25440 16178 25492
rect 16666 25440 16672 25492
rect 16724 25480 16730 25492
rect 18141 25483 18199 25489
rect 16724 25452 18092 25480
rect 16724 25440 16730 25452
rect 8386 25372 8392 25424
rect 8444 25372 8450 25424
rect 13814 25372 13820 25424
rect 13872 25412 13878 25424
rect 18064 25412 18092 25452
rect 18141 25449 18153 25483
rect 18187 25480 18199 25483
rect 20898 25480 20904 25492
rect 18187 25452 20904 25480
rect 18187 25449 18199 25452
rect 18141 25443 18199 25449
rect 20898 25440 20904 25452
rect 20956 25440 20962 25492
rect 23474 25480 23480 25492
rect 22756 25452 23480 25480
rect 18877 25415 18935 25421
rect 18877 25412 18889 25415
rect 13872 25384 18000 25412
rect 18064 25384 18889 25412
rect 13872 25372 13878 25384
rect 1302 25304 1308 25356
rect 1360 25344 1366 25356
rect 2041 25347 2099 25353
rect 2041 25344 2053 25347
rect 1360 25316 2053 25344
rect 1360 25304 1366 25316
rect 2041 25313 2053 25316
rect 2087 25313 2099 25347
rect 2041 25307 2099 25313
rect 3326 25304 3332 25356
rect 3384 25344 3390 25356
rect 3973 25347 4031 25353
rect 3973 25344 3985 25347
rect 3384 25316 3985 25344
rect 3384 25304 3390 25316
rect 3973 25313 3985 25316
rect 4019 25313 4031 25347
rect 3973 25307 4031 25313
rect 5718 25304 5724 25356
rect 5776 25344 5782 25356
rect 5994 25344 6000 25356
rect 5776 25316 6000 25344
rect 5776 25304 5782 25316
rect 5994 25304 6000 25316
rect 6052 25304 6058 25356
rect 6270 25304 6276 25356
rect 6328 25344 6334 25356
rect 6365 25347 6423 25353
rect 6365 25344 6377 25347
rect 6328 25316 6377 25344
rect 6328 25304 6334 25316
rect 6365 25313 6377 25316
rect 6411 25313 6423 25347
rect 6365 25307 6423 25313
rect 6641 25347 6699 25353
rect 6641 25313 6653 25347
rect 6687 25344 6699 25347
rect 7650 25344 7656 25356
rect 6687 25316 7656 25344
rect 6687 25313 6699 25316
rect 6641 25307 6699 25313
rect 7650 25304 7656 25316
rect 7708 25304 7714 25356
rect 8404 25344 8432 25372
rect 7760 25316 8432 25344
rect 1762 25236 1768 25288
rect 1820 25236 1826 25288
rect 3602 25236 3608 25288
rect 3660 25276 3666 25288
rect 4338 25276 4344 25288
rect 3660 25248 4344 25276
rect 3660 25236 3666 25248
rect 4338 25236 4344 25248
rect 4396 25276 4402 25288
rect 4433 25279 4491 25285
rect 4433 25276 4445 25279
rect 4396 25248 4445 25276
rect 4396 25236 4402 25248
rect 4433 25245 4445 25248
rect 4479 25245 4491 25279
rect 7760 25262 7788 25316
rect 15562 25304 15568 25356
rect 15620 25304 15626 25356
rect 15654 25304 15660 25356
rect 15712 25304 15718 25356
rect 16574 25304 16580 25356
rect 16632 25344 16638 25356
rect 16761 25347 16819 25353
rect 16761 25344 16773 25347
rect 16632 25316 16773 25344
rect 16632 25304 16638 25316
rect 16761 25313 16773 25316
rect 16807 25313 16819 25347
rect 16761 25307 16819 25313
rect 16945 25347 17003 25353
rect 16945 25313 16957 25347
rect 16991 25344 17003 25347
rect 17034 25344 17040 25356
rect 16991 25316 17040 25344
rect 16991 25313 17003 25316
rect 16945 25307 17003 25313
rect 17034 25304 17040 25316
rect 17092 25344 17098 25356
rect 17494 25344 17500 25356
rect 17092 25316 17500 25344
rect 17092 25304 17098 25316
rect 17494 25304 17500 25316
rect 17552 25304 17558 25356
rect 15473 25279 15531 25285
rect 4433 25239 4491 25245
rect 15473 25245 15485 25279
rect 15519 25276 15531 25279
rect 17678 25276 17684 25288
rect 15519 25248 17684 25276
rect 15519 25245 15531 25248
rect 15473 25239 15531 25245
rect 17678 25236 17684 25248
rect 17736 25236 17742 25288
rect 17972 25285 18000 25384
rect 18877 25381 18889 25384
rect 18923 25381 18935 25415
rect 18877 25375 18935 25381
rect 20441 25347 20499 25353
rect 20441 25313 20453 25347
rect 20487 25344 20499 25347
rect 21450 25344 21456 25356
rect 20487 25316 21456 25344
rect 20487 25313 20499 25316
rect 20441 25307 20499 25313
rect 21450 25304 21456 25316
rect 21508 25344 21514 25356
rect 22002 25344 22008 25356
rect 21508 25316 22008 25344
rect 21508 25304 21514 25316
rect 22002 25304 22008 25316
rect 22060 25304 22066 25356
rect 22756 25353 22784 25452
rect 23474 25440 23480 25452
rect 23532 25480 23538 25492
rect 23842 25480 23848 25492
rect 23532 25452 23848 25480
rect 23532 25440 23538 25452
rect 23842 25440 23848 25452
rect 23900 25440 23906 25492
rect 23385 25415 23443 25421
rect 23385 25381 23397 25415
rect 23431 25412 23443 25415
rect 25038 25412 25044 25424
rect 23431 25384 25044 25412
rect 23431 25381 23443 25384
rect 23385 25375 23443 25381
rect 25038 25372 25044 25384
rect 25096 25372 25102 25424
rect 22741 25347 22799 25353
rect 22741 25313 22753 25347
rect 22787 25313 22799 25347
rect 22741 25307 22799 25313
rect 22830 25304 22836 25356
rect 22888 25344 22894 25356
rect 22925 25347 22983 25353
rect 22925 25344 22937 25347
rect 22888 25316 22937 25344
rect 22888 25304 22894 25316
rect 22925 25313 22937 25316
rect 22971 25313 22983 25347
rect 22925 25307 22983 25313
rect 17957 25279 18015 25285
rect 17957 25245 17969 25279
rect 18003 25245 18015 25279
rect 17957 25239 18015 25245
rect 23382 25236 23388 25288
rect 23440 25276 23446 25288
rect 23440 25248 23980 25276
rect 23440 25236 23446 25248
rect 16114 25168 16120 25220
rect 16172 25208 16178 25220
rect 16669 25211 16727 25217
rect 16669 25208 16681 25211
rect 16172 25180 16681 25208
rect 16172 25168 16178 25180
rect 16669 25177 16681 25180
rect 16715 25177 16727 25211
rect 16669 25171 16727 25177
rect 19334 25168 19340 25220
rect 19392 25208 19398 25220
rect 20717 25211 20775 25217
rect 20717 25208 20729 25211
rect 19392 25180 20729 25208
rect 19392 25168 19398 25180
rect 20717 25177 20729 25180
rect 20763 25177 20775 25211
rect 22646 25208 22652 25220
rect 21942 25180 22652 25208
rect 20717 25171 20775 25177
rect 22646 25168 22652 25180
rect 22704 25168 22710 25220
rect 23017 25211 23075 25217
rect 23017 25177 23029 25211
rect 23063 25208 23075 25211
rect 23845 25211 23903 25217
rect 23845 25208 23857 25211
rect 23063 25180 23857 25208
rect 23063 25177 23075 25180
rect 23017 25171 23075 25177
rect 23845 25177 23857 25180
rect 23891 25177 23903 25211
rect 23952 25208 23980 25248
rect 24118 25236 24124 25288
rect 24176 25276 24182 25288
rect 24765 25279 24823 25285
rect 24765 25276 24777 25279
rect 24176 25248 24777 25276
rect 24176 25236 24182 25248
rect 24765 25245 24777 25248
rect 24811 25245 24823 25279
rect 24765 25239 24823 25245
rect 25041 25211 25099 25217
rect 25041 25208 25053 25211
rect 23952 25180 25053 25208
rect 23845 25171 23903 25177
rect 25041 25177 25053 25180
rect 25087 25177 25099 25211
rect 25041 25171 25099 25177
rect 7926 25100 7932 25152
rect 7984 25140 7990 25152
rect 8113 25143 8171 25149
rect 8113 25140 8125 25143
rect 7984 25112 8125 25140
rect 7984 25100 7990 25112
rect 8113 25109 8125 25112
rect 8159 25109 8171 25143
rect 8113 25103 8171 25109
rect 9122 25100 9128 25152
rect 9180 25100 9186 25152
rect 12526 25100 12532 25152
rect 12584 25140 12590 25152
rect 12621 25143 12679 25149
rect 12621 25140 12633 25143
rect 12584 25112 12633 25140
rect 12584 25100 12590 25112
rect 12621 25109 12633 25112
rect 12667 25109 12679 25143
rect 12621 25103 12679 25109
rect 15102 25100 15108 25152
rect 15160 25100 15166 25152
rect 16298 25100 16304 25152
rect 16356 25100 16362 25152
rect 21082 25100 21088 25152
rect 21140 25140 21146 25152
rect 21726 25140 21732 25152
rect 21140 25112 21732 25140
rect 21140 25100 21146 25112
rect 21726 25100 21732 25112
rect 21784 25140 21790 25152
rect 22189 25143 22247 25149
rect 22189 25140 22201 25143
rect 21784 25112 22201 25140
rect 21784 25100 21790 25112
rect 22189 25109 22201 25112
rect 22235 25109 22247 25143
rect 22189 25103 22247 25109
rect 24118 25100 24124 25152
rect 24176 25140 24182 25152
rect 24581 25143 24639 25149
rect 24581 25140 24593 25143
rect 24176 25112 24593 25140
rect 24176 25100 24182 25112
rect 24581 25109 24593 25112
rect 24627 25109 24639 25143
rect 24581 25103 24639 25109
rect 1104 25050 25852 25072
rect 1104 24998 7950 25050
rect 8002 24998 8014 25050
rect 8066 24998 8078 25050
rect 8130 24998 8142 25050
rect 8194 24998 8206 25050
rect 8258 24998 17950 25050
rect 18002 24998 18014 25050
rect 18066 24998 18078 25050
rect 18130 24998 18142 25050
rect 18194 24998 18206 25050
rect 18258 24998 25852 25050
rect 1104 24976 25852 24998
rect 8386 24896 8392 24948
rect 8444 24936 8450 24948
rect 8444 24908 9352 24936
rect 8444 24896 8450 24908
rect 4062 24828 4068 24880
rect 4120 24828 4126 24880
rect 2222 24760 2228 24812
rect 2280 24760 2286 24812
rect 4801 24803 4859 24809
rect 4801 24769 4813 24803
rect 4847 24800 4859 24803
rect 6270 24800 6276 24812
rect 4847 24772 6276 24800
rect 4847 24769 4859 24772
rect 4801 24763 4859 24769
rect 6270 24760 6276 24772
rect 6328 24800 6334 24812
rect 7929 24803 7987 24809
rect 7929 24800 7941 24803
rect 6328 24772 7941 24800
rect 6328 24760 6334 24772
rect 7929 24769 7941 24772
rect 7975 24769 7987 24803
rect 9324 24800 9352 24908
rect 12526 24896 12532 24948
rect 12584 24896 12590 24948
rect 15010 24896 15016 24948
rect 15068 24896 15074 24948
rect 18325 24939 18383 24945
rect 18325 24905 18337 24939
rect 18371 24936 18383 24939
rect 19426 24936 19432 24948
rect 18371 24908 19432 24936
rect 18371 24905 18383 24908
rect 18325 24899 18383 24905
rect 19426 24896 19432 24908
rect 19484 24896 19490 24948
rect 19613 24939 19671 24945
rect 19613 24905 19625 24939
rect 19659 24936 19671 24939
rect 20438 24936 20444 24948
rect 19659 24908 20444 24936
rect 19659 24905 19671 24908
rect 19613 24899 19671 24905
rect 20438 24896 20444 24908
rect 20496 24896 20502 24948
rect 22373 24939 22431 24945
rect 22373 24905 22385 24939
rect 22419 24936 22431 24939
rect 22738 24936 22744 24948
rect 22419 24908 22744 24936
rect 22419 24905 22431 24908
rect 22373 24899 22431 24905
rect 22738 24896 22744 24908
rect 22796 24896 22802 24948
rect 12437 24871 12495 24877
rect 12437 24868 12449 24871
rect 12268 24840 12449 24868
rect 9582 24800 9588 24812
rect 9324 24786 9588 24800
rect 9338 24772 9588 24786
rect 7929 24763 7987 24769
rect 9582 24760 9588 24772
rect 9640 24800 9646 24812
rect 9953 24803 10011 24809
rect 9953 24800 9965 24803
rect 9640 24772 9965 24800
rect 9640 24760 9646 24772
rect 9953 24769 9965 24772
rect 9999 24769 10011 24803
rect 9953 24763 10011 24769
rect 10686 24760 10692 24812
rect 10744 24760 10750 24812
rect 10778 24760 10784 24812
rect 10836 24760 10842 24812
rect 11422 24760 11428 24812
rect 11480 24800 11486 24812
rect 11882 24800 11888 24812
rect 11480 24772 11888 24800
rect 11480 24760 11486 24772
rect 11882 24760 11888 24772
rect 11940 24800 11946 24812
rect 12268 24800 12296 24840
rect 12437 24837 12449 24840
rect 12483 24837 12495 24871
rect 12437 24831 12495 24837
rect 14550 24828 14556 24880
rect 14608 24828 14614 24880
rect 15028 24868 15056 24896
rect 15028 24840 15318 24868
rect 12618 24800 12624 24812
rect 11940 24772 12296 24800
rect 12360 24772 12624 24800
rect 11940 24760 11946 24772
rect 3053 24735 3111 24741
rect 3053 24701 3065 24735
rect 3099 24732 3111 24735
rect 4154 24732 4160 24744
rect 3099 24704 4160 24732
rect 3099 24701 3111 24704
rect 3053 24695 3111 24701
rect 4154 24692 4160 24704
rect 4212 24692 4218 24744
rect 4525 24735 4583 24741
rect 4525 24701 4537 24735
rect 4571 24732 4583 24735
rect 5718 24732 5724 24744
rect 4571 24704 5724 24732
rect 4571 24701 4583 24704
rect 4525 24695 4583 24701
rect 5718 24692 5724 24704
rect 5776 24692 5782 24744
rect 7466 24692 7472 24744
rect 7524 24692 7530 24744
rect 7834 24692 7840 24744
rect 7892 24732 7898 24744
rect 12360 24741 12388 24772
rect 12618 24760 12624 24772
rect 12676 24760 12682 24812
rect 8205 24735 8263 24741
rect 8205 24732 8217 24735
rect 7892 24704 8217 24732
rect 7892 24692 7898 24704
rect 8205 24701 8217 24704
rect 8251 24732 8263 24735
rect 10505 24735 10563 24741
rect 10505 24732 10517 24735
rect 8251 24704 10517 24732
rect 8251 24701 8263 24704
rect 8205 24695 8263 24701
rect 10505 24701 10517 24704
rect 10551 24701 10563 24735
rect 10505 24695 10563 24701
rect 12345 24735 12403 24741
rect 12345 24701 12357 24735
rect 12391 24701 12403 24735
rect 14182 24732 14188 24744
rect 12345 24695 12403 24701
rect 12820 24704 14188 24732
rect 1946 24624 1952 24676
rect 2004 24664 2010 24676
rect 2041 24667 2099 24673
rect 2041 24664 2053 24667
rect 2004 24636 2053 24664
rect 2004 24624 2010 24636
rect 2041 24633 2053 24636
rect 2087 24633 2099 24667
rect 2041 24627 2099 24633
rect 9677 24667 9735 24673
rect 9677 24633 9689 24667
rect 9723 24664 9735 24667
rect 9766 24664 9772 24676
rect 9723 24636 9772 24664
rect 9723 24633 9735 24636
rect 9677 24627 9735 24633
rect 9766 24624 9772 24636
rect 9824 24664 9830 24676
rect 10962 24664 10968 24676
rect 9824 24636 10968 24664
rect 9824 24624 9830 24636
rect 10962 24624 10968 24636
rect 11020 24624 11026 24676
rect 11149 24667 11207 24673
rect 11149 24633 11161 24667
rect 11195 24664 11207 24667
rect 12820 24664 12848 24704
rect 14182 24692 14188 24704
rect 14240 24692 14246 24744
rect 14568 24741 14596 24828
rect 16114 24760 16120 24812
rect 16172 24800 16178 24812
rect 16666 24800 16672 24812
rect 16172 24772 16672 24800
rect 16172 24760 16178 24772
rect 16666 24760 16672 24772
rect 16724 24760 16730 24812
rect 18414 24760 18420 24812
rect 18472 24760 18478 24812
rect 19518 24760 19524 24812
rect 19576 24760 19582 24812
rect 21358 24760 21364 24812
rect 21416 24800 21422 24812
rect 22281 24803 22339 24809
rect 22281 24800 22293 24803
rect 21416 24772 22293 24800
rect 21416 24760 21422 24772
rect 22281 24769 22293 24772
rect 22327 24769 22339 24803
rect 22281 24763 22339 24769
rect 24578 24760 24584 24812
rect 24636 24800 24642 24812
rect 25225 24803 25283 24809
rect 25225 24800 25237 24803
rect 24636 24772 25237 24800
rect 24636 24760 24642 24772
rect 25225 24769 25237 24772
rect 25271 24769 25283 24803
rect 25225 24763 25283 24769
rect 14553 24735 14611 24741
rect 14553 24701 14565 24735
rect 14599 24701 14611 24735
rect 14553 24695 14611 24701
rect 14829 24735 14887 24741
rect 14829 24701 14841 24735
rect 14875 24732 14887 24735
rect 16206 24732 16212 24744
rect 14875 24704 16212 24732
rect 14875 24701 14887 24704
rect 14829 24695 14887 24701
rect 11195 24636 12848 24664
rect 12897 24667 12955 24673
rect 11195 24633 11207 24636
rect 11149 24627 11207 24633
rect 12897 24633 12909 24667
rect 12943 24664 12955 24667
rect 13814 24664 13820 24676
rect 12943 24636 13820 24664
rect 12943 24633 12955 24636
rect 12897 24627 12955 24633
rect 13814 24624 13820 24636
rect 13872 24624 13878 24676
rect 5169 24599 5227 24605
rect 5169 24565 5181 24599
rect 5215 24596 5227 24599
rect 5626 24596 5632 24608
rect 5215 24568 5632 24596
rect 5215 24565 5227 24568
rect 5169 24559 5227 24565
rect 5626 24556 5632 24568
rect 5684 24556 5690 24608
rect 13265 24599 13323 24605
rect 13265 24565 13277 24599
rect 13311 24596 13323 24599
rect 13630 24596 13636 24608
rect 13311 24568 13636 24596
rect 13311 24565 13323 24568
rect 13265 24559 13323 24565
rect 13630 24556 13636 24568
rect 13688 24556 13694 24608
rect 14568 24596 14596 24695
rect 16206 24692 16212 24704
rect 16264 24692 16270 24744
rect 16301 24735 16359 24741
rect 16301 24701 16313 24735
rect 16347 24732 16359 24735
rect 16574 24732 16580 24744
rect 16347 24704 16580 24732
rect 16347 24701 16359 24704
rect 16301 24695 16359 24701
rect 16574 24692 16580 24704
rect 16632 24732 16638 24744
rect 17218 24732 17224 24744
rect 16632 24704 17224 24732
rect 16632 24692 16638 24704
rect 17218 24692 17224 24704
rect 17276 24692 17282 24744
rect 18598 24692 18604 24744
rect 18656 24692 18662 24744
rect 19334 24692 19340 24744
rect 19392 24692 19398 24744
rect 22094 24692 22100 24744
rect 22152 24692 22158 24744
rect 23201 24735 23259 24741
rect 23201 24701 23213 24735
rect 23247 24701 23259 24735
rect 23201 24695 23259 24701
rect 16942 24664 16948 24676
rect 15856 24636 16948 24664
rect 15856 24596 15884 24636
rect 16942 24624 16948 24636
rect 17000 24624 17006 24676
rect 22186 24624 22192 24676
rect 22244 24664 22250 24676
rect 22830 24664 22836 24676
rect 22244 24636 22836 24664
rect 22244 24624 22250 24636
rect 22830 24624 22836 24636
rect 22888 24664 22894 24676
rect 23216 24664 23244 24695
rect 23474 24692 23480 24744
rect 23532 24692 23538 24744
rect 24854 24692 24860 24744
rect 24912 24732 24918 24744
rect 24949 24735 25007 24741
rect 24949 24732 24961 24735
rect 24912 24704 24961 24732
rect 24912 24692 24918 24704
rect 24949 24701 24961 24704
rect 24995 24732 25007 24735
rect 25406 24732 25412 24744
rect 24995 24704 25412 24732
rect 24995 24701 25007 24704
rect 24949 24695 25007 24701
rect 25406 24692 25412 24704
rect 25464 24692 25470 24744
rect 22888 24636 23244 24664
rect 22888 24624 22894 24636
rect 14568 24568 15884 24596
rect 16666 24556 16672 24608
rect 16724 24596 16730 24608
rect 17586 24596 17592 24608
rect 16724 24568 17592 24596
rect 16724 24556 16730 24568
rect 17586 24556 17592 24568
rect 17644 24556 17650 24608
rect 17957 24599 18015 24605
rect 17957 24565 17969 24599
rect 18003 24596 18015 24599
rect 18322 24596 18328 24608
rect 18003 24568 18328 24596
rect 18003 24565 18015 24568
rect 17957 24559 18015 24565
rect 18322 24556 18328 24568
rect 18380 24556 18386 24608
rect 19886 24556 19892 24608
rect 19944 24596 19950 24608
rect 19981 24599 20039 24605
rect 19981 24596 19993 24599
rect 19944 24568 19993 24596
rect 19944 24556 19950 24568
rect 19981 24565 19993 24568
rect 20027 24565 20039 24599
rect 19981 24559 20039 24565
rect 22738 24556 22744 24608
rect 22796 24556 22802 24608
rect 1104 24506 25852 24528
rect 1104 24454 2950 24506
rect 3002 24454 3014 24506
rect 3066 24454 3078 24506
rect 3130 24454 3142 24506
rect 3194 24454 3206 24506
rect 3258 24454 12950 24506
rect 13002 24454 13014 24506
rect 13066 24454 13078 24506
rect 13130 24454 13142 24506
rect 13194 24454 13206 24506
rect 13258 24454 22950 24506
rect 23002 24454 23014 24506
rect 23066 24454 23078 24506
rect 23130 24454 23142 24506
rect 23194 24454 23206 24506
rect 23258 24454 25852 24506
rect 1104 24432 25852 24454
rect 2866 24352 2872 24404
rect 2924 24352 2930 24404
rect 3142 24352 3148 24404
rect 3200 24352 3206 24404
rect 4062 24352 4068 24404
rect 4120 24392 4126 24404
rect 4525 24395 4583 24401
rect 4525 24392 4537 24395
rect 4120 24364 4537 24392
rect 4120 24352 4126 24364
rect 4525 24361 4537 24364
rect 4571 24392 4583 24395
rect 5626 24392 5632 24404
rect 4571 24364 5632 24392
rect 4571 24361 4583 24364
rect 4525 24355 4583 24361
rect 5626 24352 5632 24364
rect 5684 24352 5690 24404
rect 7374 24352 7380 24404
rect 7432 24392 7438 24404
rect 7469 24395 7527 24401
rect 7469 24392 7481 24395
rect 7432 24364 7481 24392
rect 7432 24352 7438 24364
rect 7469 24361 7481 24364
rect 7515 24392 7527 24395
rect 7558 24392 7564 24404
rect 7515 24364 7564 24392
rect 7515 24361 7527 24364
rect 7469 24355 7527 24361
rect 7558 24352 7564 24364
rect 7616 24392 7622 24404
rect 8573 24395 8631 24401
rect 7616 24364 8156 24392
rect 7616 24352 7622 24364
rect 7650 24216 7656 24268
rect 7708 24256 7714 24268
rect 8128 24265 8156 24364
rect 8573 24361 8585 24395
rect 8619 24392 8631 24395
rect 10778 24392 10784 24404
rect 8619 24364 10784 24392
rect 8619 24361 8631 24364
rect 8573 24355 8631 24361
rect 10778 24352 10784 24364
rect 10836 24352 10842 24404
rect 10962 24352 10968 24404
rect 11020 24352 11026 24404
rect 11241 24395 11299 24401
rect 11241 24361 11253 24395
rect 11287 24392 11299 24395
rect 11330 24392 11336 24404
rect 11287 24364 11336 24392
rect 11287 24361 11299 24364
rect 11241 24355 11299 24361
rect 11330 24352 11336 24364
rect 11388 24352 11394 24404
rect 12434 24352 12440 24404
rect 12492 24392 12498 24404
rect 12621 24395 12679 24401
rect 12621 24392 12633 24395
rect 12492 24364 12633 24392
rect 12492 24352 12498 24364
rect 12621 24361 12633 24364
rect 12667 24361 12679 24395
rect 17494 24392 17500 24404
rect 12621 24355 12679 24361
rect 13372 24364 17500 24392
rect 10980 24324 11008 24352
rect 10796 24296 11008 24324
rect 7929 24259 7987 24265
rect 7929 24256 7941 24259
rect 7708 24228 7941 24256
rect 7708 24216 7714 24228
rect 7929 24225 7941 24228
rect 7975 24225 7987 24259
rect 7929 24219 7987 24225
rect 8113 24259 8171 24265
rect 8113 24225 8125 24259
rect 8159 24225 8171 24259
rect 8113 24219 8171 24225
rect 10597 24259 10655 24265
rect 10597 24225 10609 24259
rect 10643 24256 10655 24259
rect 10796 24256 10824 24296
rect 10643 24228 10824 24256
rect 10643 24225 10655 24228
rect 10597 24219 10655 24225
rect 10962 24216 10968 24268
rect 11020 24256 11026 24268
rect 12069 24259 12127 24265
rect 12069 24256 12081 24259
rect 11020 24228 12081 24256
rect 11020 24216 11026 24228
rect 12069 24225 12081 24228
rect 12115 24225 12127 24259
rect 12069 24219 12127 24225
rect 13173 24259 13231 24265
rect 13173 24225 13185 24259
rect 13219 24256 13231 24259
rect 13372 24256 13400 24364
rect 17494 24352 17500 24364
rect 17552 24352 17558 24404
rect 24394 24352 24400 24404
rect 24452 24392 24458 24404
rect 24578 24392 24584 24404
rect 24452 24364 24584 24392
rect 24452 24352 24458 24364
rect 24578 24352 24584 24364
rect 24636 24352 24642 24404
rect 15013 24327 15071 24333
rect 15013 24293 15025 24327
rect 15059 24324 15071 24327
rect 17218 24324 17224 24336
rect 15059 24296 17224 24324
rect 15059 24293 15071 24296
rect 15013 24287 15071 24293
rect 17218 24284 17224 24296
rect 17276 24284 17282 24336
rect 18966 24324 18972 24336
rect 17972 24296 18972 24324
rect 13219 24228 13400 24256
rect 13219 24225 13231 24228
rect 13173 24219 13231 24225
rect 13446 24216 13452 24268
rect 13504 24256 13510 24268
rect 14369 24259 14427 24265
rect 14369 24256 14381 24259
rect 13504 24228 14381 24256
rect 13504 24216 13510 24228
rect 14369 24225 14381 24228
rect 14415 24225 14427 24259
rect 14369 24219 14427 24225
rect 14553 24259 14611 24265
rect 14553 24225 14565 24259
rect 14599 24256 14611 24259
rect 14642 24256 14648 24268
rect 14599 24228 14648 24256
rect 14599 24225 14611 24228
rect 14553 24219 14611 24225
rect 14642 24216 14648 24228
rect 14700 24216 14706 24268
rect 15657 24259 15715 24265
rect 15657 24225 15669 24259
rect 15703 24225 15715 24259
rect 15657 24219 15715 24225
rect 15749 24259 15807 24265
rect 15749 24225 15761 24259
rect 15795 24256 15807 24259
rect 16298 24256 16304 24268
rect 15795 24228 16304 24256
rect 15795 24225 15807 24228
rect 15749 24219 15807 24225
rect 3329 24191 3387 24197
rect 3329 24188 3341 24191
rect 2746 24160 3341 24188
rect 2593 24123 2651 24129
rect 2593 24089 2605 24123
rect 2639 24120 2651 24123
rect 2746 24120 2774 24160
rect 3329 24157 3341 24160
rect 3375 24188 3387 24191
rect 3602 24188 3608 24200
rect 3375 24160 3608 24188
rect 3375 24157 3387 24160
rect 3329 24151 3387 24157
rect 3602 24148 3608 24160
rect 3660 24148 3666 24200
rect 4062 24197 4068 24200
rect 4040 24191 4068 24197
rect 4040 24157 4052 24191
rect 4040 24151 4068 24157
rect 4062 24148 4068 24151
rect 4120 24148 4126 24200
rect 7466 24148 7472 24200
rect 7524 24188 7530 24200
rect 8205 24191 8263 24197
rect 8205 24188 8217 24191
rect 7524 24160 8217 24188
rect 7524 24148 7530 24160
rect 8205 24157 8217 24160
rect 8251 24157 8263 24191
rect 8205 24151 8263 24157
rect 10870 24148 10876 24200
rect 10928 24148 10934 24200
rect 11885 24191 11943 24197
rect 11885 24157 11897 24191
rect 11931 24188 11943 24191
rect 13630 24188 13636 24200
rect 11931 24160 13636 24188
rect 11931 24157 11943 24160
rect 11885 24151 11943 24157
rect 13630 24148 13636 24160
rect 13688 24148 13694 24200
rect 15672 24188 15700 24219
rect 16298 24216 16304 24228
rect 16356 24216 16362 24268
rect 17972 24265 18000 24296
rect 18966 24284 18972 24296
rect 19024 24284 19030 24336
rect 17957 24259 18015 24265
rect 17957 24225 17969 24259
rect 18003 24225 18015 24259
rect 17957 24219 18015 24225
rect 18049 24259 18107 24265
rect 18049 24225 18061 24259
rect 18095 24256 18107 24259
rect 18506 24256 18512 24268
rect 18095 24228 18512 24256
rect 18095 24225 18107 24228
rect 18049 24219 18107 24225
rect 18506 24216 18512 24228
rect 18564 24216 18570 24268
rect 19978 24216 19984 24268
rect 20036 24216 20042 24268
rect 20165 24259 20223 24265
rect 20165 24225 20177 24259
rect 20211 24256 20223 24259
rect 21082 24256 21088 24268
rect 20211 24228 21088 24256
rect 20211 24225 20223 24228
rect 20165 24219 20223 24225
rect 21082 24216 21088 24228
rect 21140 24216 21146 24268
rect 21174 24216 21180 24268
rect 21232 24256 21238 24268
rect 21361 24259 21419 24265
rect 21361 24256 21373 24259
rect 21232 24228 21373 24256
rect 21232 24216 21238 24228
rect 21361 24225 21373 24228
rect 21407 24256 21419 24259
rect 21450 24256 21456 24268
rect 21407 24228 21456 24256
rect 21407 24225 21419 24228
rect 21361 24219 21419 24225
rect 21450 24216 21456 24228
rect 21508 24216 21514 24268
rect 23385 24259 23443 24265
rect 23385 24225 23397 24259
rect 23431 24256 23443 24259
rect 24854 24256 24860 24268
rect 23431 24228 24860 24256
rect 23431 24225 23443 24228
rect 23385 24219 23443 24225
rect 24854 24216 24860 24228
rect 24912 24216 24918 24268
rect 16206 24188 16212 24200
rect 15672 24160 16212 24188
rect 16206 24148 16212 24160
rect 16264 24148 16270 24200
rect 19886 24148 19892 24200
rect 19944 24148 19950 24200
rect 24029 24191 24087 24197
rect 22066 24160 23060 24188
rect 2639 24092 2774 24120
rect 2639 24089 2651 24092
rect 2593 24083 2651 24089
rect 4522 24080 4528 24132
rect 4580 24120 4586 24132
rect 9030 24120 9036 24132
rect 4580 24092 9036 24120
rect 4580 24080 4586 24092
rect 9030 24080 9036 24092
rect 9088 24080 9094 24132
rect 9582 24080 9588 24132
rect 9640 24080 9646 24132
rect 11330 24080 11336 24132
rect 11388 24120 11394 24132
rect 11977 24123 12035 24129
rect 11977 24120 11989 24123
rect 11388 24092 11989 24120
rect 11388 24080 11394 24092
rect 11977 24089 11989 24092
rect 12023 24089 12035 24123
rect 11977 24083 12035 24089
rect 12434 24080 12440 24132
rect 12492 24120 12498 24132
rect 13265 24123 13323 24129
rect 13265 24120 13277 24123
rect 12492 24092 13277 24120
rect 12492 24080 12498 24092
rect 13265 24089 13277 24092
rect 13311 24089 13323 24123
rect 15841 24123 15899 24129
rect 15841 24120 15853 24123
rect 13265 24083 13323 24089
rect 13740 24092 15853 24120
rect 3970 24012 3976 24064
rect 4028 24052 4034 24064
rect 4111 24055 4169 24061
rect 4111 24052 4123 24055
rect 4028 24024 4123 24052
rect 4028 24012 4034 24024
rect 4111 24021 4123 24024
rect 4157 24021 4169 24055
rect 4111 24015 4169 24021
rect 9125 24055 9183 24061
rect 9125 24021 9137 24055
rect 9171 24052 9183 24055
rect 9858 24052 9864 24064
rect 9171 24024 9864 24052
rect 9171 24021 9183 24024
rect 9125 24015 9183 24021
rect 9858 24012 9864 24024
rect 9916 24012 9922 24064
rect 11517 24055 11575 24061
rect 11517 24021 11529 24055
rect 11563 24052 11575 24055
rect 11606 24052 11612 24064
rect 11563 24024 11612 24052
rect 11563 24021 11575 24024
rect 11517 24015 11575 24021
rect 11606 24012 11612 24024
rect 11664 24012 11670 24064
rect 13357 24055 13415 24061
rect 13357 24021 13369 24055
rect 13403 24052 13415 24055
rect 13538 24052 13544 24064
rect 13403 24024 13544 24052
rect 13403 24021 13415 24024
rect 13357 24015 13415 24021
rect 13538 24012 13544 24024
rect 13596 24012 13602 24064
rect 13740 24061 13768 24092
rect 15841 24089 15853 24092
rect 15887 24089 15899 24123
rect 15841 24083 15899 24089
rect 18874 24080 18880 24132
rect 18932 24120 18938 24132
rect 21177 24123 21235 24129
rect 21177 24120 21189 24123
rect 18932 24092 21189 24120
rect 18932 24080 18938 24092
rect 21177 24089 21189 24092
rect 21223 24089 21235 24123
rect 21177 24083 21235 24089
rect 13725 24055 13783 24061
rect 13725 24021 13737 24055
rect 13771 24021 13783 24055
rect 13725 24015 13783 24021
rect 13814 24012 13820 24064
rect 13872 24052 13878 24064
rect 14645 24055 14703 24061
rect 14645 24052 14657 24055
rect 13872 24024 14657 24052
rect 13872 24012 13878 24024
rect 14645 24021 14657 24024
rect 14691 24021 14703 24055
rect 14645 24015 14703 24021
rect 15930 24012 15936 24064
rect 15988 24052 15994 24064
rect 16209 24055 16267 24061
rect 16209 24052 16221 24055
rect 15988 24024 16221 24052
rect 15988 24012 15994 24024
rect 16209 24021 16221 24024
rect 16255 24021 16267 24055
rect 16209 24015 16267 24021
rect 17126 24012 17132 24064
rect 17184 24052 17190 24064
rect 17405 24055 17463 24061
rect 17405 24052 17417 24055
rect 17184 24024 17417 24052
rect 17184 24012 17190 24024
rect 17405 24021 17417 24024
rect 17451 24052 17463 24055
rect 18141 24055 18199 24061
rect 18141 24052 18153 24055
rect 17451 24024 18153 24052
rect 17451 24021 17463 24024
rect 17405 24015 17463 24021
rect 18141 24021 18153 24024
rect 18187 24021 18199 24055
rect 18141 24015 18199 24021
rect 18506 24012 18512 24064
rect 18564 24012 18570 24064
rect 18782 24012 18788 24064
rect 18840 24052 18846 24064
rect 19521 24055 19579 24061
rect 19521 24052 19533 24055
rect 18840 24024 19533 24052
rect 18840 24012 18846 24024
rect 19521 24021 19533 24024
rect 19567 24021 19579 24055
rect 19521 24015 19579 24021
rect 20714 24012 20720 24064
rect 20772 24012 20778 24064
rect 21082 24012 21088 24064
rect 21140 24012 21146 24064
rect 21192 24052 21220 24083
rect 21266 24080 21272 24132
rect 21324 24120 21330 24132
rect 22066 24120 22094 24160
rect 21324 24092 22094 24120
rect 23032 24120 23060 24160
rect 24029 24157 24041 24191
rect 24075 24188 24087 24191
rect 24486 24188 24492 24200
rect 24075 24160 24492 24188
rect 24075 24157 24087 24160
rect 24029 24151 24087 24157
rect 24486 24148 24492 24160
rect 24544 24148 24550 24200
rect 24765 24123 24823 24129
rect 24765 24120 24777 24123
rect 23032 24092 24777 24120
rect 21324 24080 21330 24092
rect 24765 24089 24777 24092
rect 24811 24089 24823 24123
rect 24765 24083 24823 24089
rect 24486 24052 24492 24064
rect 21192 24024 24492 24052
rect 24486 24012 24492 24024
rect 24544 24012 24550 24064
rect 24670 24012 24676 24064
rect 24728 24012 24734 24064
rect 1104 23962 25852 23984
rect 1104 23910 7950 23962
rect 8002 23910 8014 23962
rect 8066 23910 8078 23962
rect 8130 23910 8142 23962
rect 8194 23910 8206 23962
rect 8258 23910 17950 23962
rect 18002 23910 18014 23962
rect 18066 23910 18078 23962
rect 18130 23910 18142 23962
rect 18194 23910 18206 23962
rect 18258 23910 25852 23962
rect 1104 23888 25852 23910
rect 5626 23848 5632 23860
rect 3436 23820 5632 23848
rect 3436 23780 3464 23820
rect 3082 23752 3464 23780
rect 3513 23783 3571 23789
rect 3513 23749 3525 23783
rect 3559 23780 3571 23783
rect 4154 23780 4160 23792
rect 3559 23752 4160 23780
rect 3559 23749 3571 23752
rect 3513 23743 3571 23749
rect 4154 23740 4160 23752
rect 4212 23740 4218 23792
rect 5368 23780 5396 23820
rect 5626 23808 5632 23820
rect 5684 23848 5690 23860
rect 6730 23848 6736 23860
rect 5684 23820 6736 23848
rect 5684 23808 5690 23820
rect 6730 23808 6736 23820
rect 6788 23808 6794 23860
rect 8849 23851 8907 23857
rect 8849 23817 8861 23851
rect 8895 23848 8907 23851
rect 9122 23848 9128 23860
rect 8895 23820 9128 23848
rect 8895 23817 8907 23820
rect 8849 23811 8907 23817
rect 9122 23808 9128 23820
rect 9180 23808 9186 23860
rect 9398 23808 9404 23860
rect 9456 23848 9462 23860
rect 9953 23851 10011 23857
rect 9953 23848 9965 23851
rect 9456 23820 9965 23848
rect 9456 23808 9462 23820
rect 9953 23817 9965 23820
rect 9999 23817 10011 23851
rect 9953 23811 10011 23817
rect 10413 23851 10471 23857
rect 10413 23817 10425 23851
rect 10459 23848 10471 23851
rect 12713 23851 12771 23857
rect 12713 23848 12725 23851
rect 10459 23820 12725 23848
rect 10459 23817 10471 23820
rect 10413 23811 10471 23817
rect 12713 23817 12725 23820
rect 12759 23817 12771 23851
rect 12713 23811 12771 23817
rect 13538 23808 13544 23860
rect 13596 23808 13602 23860
rect 15930 23808 15936 23860
rect 15988 23808 15994 23860
rect 16025 23851 16083 23857
rect 16025 23817 16037 23851
rect 16071 23848 16083 23851
rect 16850 23848 16856 23860
rect 16071 23820 16856 23848
rect 16071 23817 16083 23820
rect 16025 23811 16083 23817
rect 16850 23808 16856 23820
rect 16908 23808 16914 23860
rect 17862 23808 17868 23860
rect 17920 23848 17926 23860
rect 20533 23851 20591 23857
rect 20533 23848 20545 23851
rect 17920 23820 20545 23848
rect 17920 23808 17926 23820
rect 20533 23817 20545 23820
rect 20579 23848 20591 23851
rect 21082 23848 21088 23860
rect 20579 23820 21088 23848
rect 20579 23817 20591 23820
rect 20533 23811 20591 23817
rect 21082 23808 21088 23820
rect 21140 23808 21146 23860
rect 5290 23752 5396 23780
rect 5442 23740 5448 23792
rect 5500 23780 5506 23792
rect 8941 23783 8999 23789
rect 5500 23752 6040 23780
rect 5500 23740 5506 23752
rect 6012 23721 6040 23752
rect 8941 23749 8953 23783
rect 8987 23780 8999 23783
rect 9030 23780 9036 23792
rect 8987 23752 9036 23780
rect 8987 23749 8999 23752
rect 8941 23743 8999 23749
rect 9030 23740 9036 23752
rect 9088 23780 9094 23792
rect 11974 23780 11980 23792
rect 9088 23752 11980 23780
rect 9088 23740 9094 23752
rect 11974 23740 11980 23752
rect 12032 23740 12038 23792
rect 12621 23783 12679 23789
rect 12621 23749 12633 23783
rect 12667 23780 12679 23783
rect 13998 23780 14004 23792
rect 12667 23752 14004 23780
rect 12667 23749 12679 23752
rect 12621 23743 12679 23749
rect 13998 23740 14004 23752
rect 14056 23740 14062 23792
rect 25130 23740 25136 23792
rect 25188 23740 25194 23792
rect 5997 23715 6055 23721
rect 5997 23681 6009 23715
rect 6043 23712 6055 23715
rect 6270 23712 6276 23724
rect 6043 23684 6276 23712
rect 6043 23681 6055 23684
rect 5997 23675 6055 23681
rect 6270 23672 6276 23684
rect 6328 23712 6334 23724
rect 7282 23712 7288 23724
rect 6328 23684 7288 23712
rect 6328 23672 6334 23684
rect 7282 23672 7288 23684
rect 7340 23672 7346 23724
rect 10045 23715 10103 23721
rect 7392 23684 9904 23712
rect 3789 23647 3847 23653
rect 3789 23613 3801 23647
rect 3835 23644 3847 23647
rect 5350 23644 5356 23656
rect 3835 23616 5356 23644
rect 3835 23613 3847 23616
rect 3789 23607 3847 23613
rect 5350 23604 5356 23616
rect 5408 23604 5414 23656
rect 5626 23604 5632 23656
rect 5684 23644 5690 23656
rect 5721 23647 5779 23653
rect 5721 23644 5733 23647
rect 5684 23616 5733 23644
rect 5684 23604 5690 23616
rect 5721 23613 5733 23616
rect 5767 23613 5779 23647
rect 5721 23607 5779 23613
rect 6638 23604 6644 23656
rect 6696 23644 6702 23656
rect 7392 23644 7420 23684
rect 6696 23616 7420 23644
rect 9033 23647 9091 23653
rect 6696 23604 6702 23616
rect 9033 23613 9045 23647
rect 9079 23613 9091 23647
rect 9033 23607 9091 23613
rect 6457 23579 6515 23585
rect 6457 23545 6469 23579
rect 6503 23576 6515 23579
rect 6730 23576 6736 23588
rect 6503 23548 6736 23576
rect 6503 23545 6515 23548
rect 6457 23539 6515 23545
rect 6730 23536 6736 23548
rect 6788 23536 6794 23588
rect 7006 23536 7012 23588
rect 7064 23576 7070 23588
rect 9048 23576 9076 23607
rect 9766 23604 9772 23656
rect 9824 23604 9830 23656
rect 9876 23644 9904 23684
rect 10045 23681 10057 23715
rect 10091 23712 10103 23715
rect 10873 23715 10931 23721
rect 10873 23712 10885 23715
rect 10091 23684 10885 23712
rect 10091 23681 10103 23684
rect 10045 23675 10103 23681
rect 10873 23681 10885 23684
rect 10919 23681 10931 23715
rect 10873 23675 10931 23681
rect 13722 23672 13728 23724
rect 13780 23712 13786 23724
rect 17497 23715 17555 23721
rect 17497 23712 17509 23715
rect 13780 23684 17509 23712
rect 13780 23672 13786 23684
rect 17497 23681 17509 23684
rect 17543 23681 17555 23715
rect 17497 23675 17555 23681
rect 23293 23715 23351 23721
rect 23293 23681 23305 23715
rect 23339 23712 23351 23715
rect 23934 23712 23940 23724
rect 23339 23684 23940 23712
rect 23339 23681 23351 23684
rect 23293 23675 23351 23681
rect 23934 23672 23940 23684
rect 23992 23672 23998 23724
rect 24118 23672 24124 23724
rect 24176 23672 24182 23724
rect 11330 23644 11336 23656
rect 9876 23616 11336 23644
rect 11330 23604 11336 23616
rect 11388 23604 11394 23656
rect 12437 23647 12495 23653
rect 12437 23613 12449 23647
rect 12483 23613 12495 23647
rect 12437 23607 12495 23613
rect 7064 23548 9076 23576
rect 7064 23536 7070 23548
rect 9858 23536 9864 23588
rect 9916 23576 9922 23588
rect 12452 23576 12480 23607
rect 13630 23604 13636 23656
rect 13688 23644 13694 23656
rect 16022 23644 16028 23656
rect 13688 23616 16028 23644
rect 13688 23604 13694 23616
rect 16022 23604 16028 23616
rect 16080 23604 16086 23656
rect 16209 23647 16267 23653
rect 16209 23613 16221 23647
rect 16255 23644 16267 23647
rect 16574 23644 16580 23656
rect 16255 23616 16580 23644
rect 16255 23613 16267 23616
rect 16209 23607 16267 23613
rect 16574 23604 16580 23616
rect 16632 23604 16638 23656
rect 23017 23647 23075 23653
rect 23017 23613 23029 23647
rect 23063 23644 23075 23647
rect 23382 23644 23388 23656
rect 23063 23616 23388 23644
rect 23063 23613 23075 23616
rect 23017 23607 23075 23613
rect 23382 23604 23388 23616
rect 23440 23604 23446 23656
rect 9916 23548 12480 23576
rect 9916 23536 9922 23548
rect 2041 23511 2099 23517
rect 2041 23477 2053 23511
rect 2087 23508 2099 23511
rect 3142 23508 3148 23520
rect 2087 23480 3148 23508
rect 2087 23477 2099 23480
rect 2041 23471 2099 23477
rect 3142 23468 3148 23480
rect 3200 23508 3206 23520
rect 4154 23508 4160 23520
rect 3200 23480 4160 23508
rect 3200 23468 3206 23480
rect 4154 23468 4160 23480
rect 4212 23468 4218 23520
rect 4249 23511 4307 23517
rect 4249 23477 4261 23511
rect 4295 23508 4307 23511
rect 5718 23508 5724 23520
rect 4295 23480 5724 23508
rect 4295 23477 4307 23480
rect 4249 23471 4307 23477
rect 5718 23468 5724 23480
rect 5776 23468 5782 23520
rect 6546 23468 6552 23520
rect 6604 23508 6610 23520
rect 8481 23511 8539 23517
rect 8481 23508 8493 23511
rect 6604 23480 8493 23508
rect 6604 23468 6610 23480
rect 8481 23477 8493 23480
rect 8527 23477 8539 23511
rect 8481 23471 8539 23477
rect 9582 23468 9588 23520
rect 9640 23508 9646 23520
rect 10686 23508 10692 23520
rect 9640 23480 10692 23508
rect 9640 23468 9646 23480
rect 10686 23468 10692 23480
rect 10744 23508 10750 23520
rect 11517 23511 11575 23517
rect 11517 23508 11529 23511
rect 10744 23480 11529 23508
rect 10744 23468 10750 23480
rect 11517 23477 11529 23480
rect 11563 23477 11575 23511
rect 11517 23471 11575 23477
rect 13081 23511 13139 23517
rect 13081 23477 13093 23511
rect 13127 23508 13139 23511
rect 14826 23508 14832 23520
rect 13127 23480 14832 23508
rect 13127 23477 13139 23480
rect 13081 23471 13139 23477
rect 14826 23468 14832 23480
rect 14884 23468 14890 23520
rect 15565 23511 15623 23517
rect 15565 23477 15577 23511
rect 15611 23508 15623 23511
rect 15746 23508 15752 23520
rect 15611 23480 15752 23508
rect 15611 23477 15623 23480
rect 15565 23471 15623 23477
rect 15746 23468 15752 23480
rect 15804 23468 15810 23520
rect 17681 23511 17739 23517
rect 17681 23477 17693 23511
rect 17727 23508 17739 23511
rect 20438 23508 20444 23520
rect 17727 23480 20444 23508
rect 17727 23477 17739 23480
rect 17681 23471 17739 23477
rect 20438 23468 20444 23480
rect 20496 23468 20502 23520
rect 1104 23418 25852 23440
rect 1104 23366 2950 23418
rect 3002 23366 3014 23418
rect 3066 23366 3078 23418
rect 3130 23366 3142 23418
rect 3194 23366 3206 23418
rect 3258 23366 12950 23418
rect 13002 23366 13014 23418
rect 13066 23366 13078 23418
rect 13130 23366 13142 23418
rect 13194 23366 13206 23418
rect 13258 23366 22950 23418
rect 23002 23366 23014 23418
rect 23066 23366 23078 23418
rect 23130 23366 23142 23418
rect 23194 23366 23206 23418
rect 23258 23366 25852 23418
rect 1104 23344 25852 23366
rect 4157 23307 4215 23313
rect 4157 23273 4169 23307
rect 4203 23304 4215 23307
rect 4246 23304 4252 23316
rect 4203 23276 4252 23304
rect 4203 23273 4215 23276
rect 4157 23267 4215 23273
rect 4246 23264 4252 23276
rect 4304 23264 4310 23316
rect 9030 23264 9036 23316
rect 9088 23264 9094 23316
rect 9217 23307 9275 23313
rect 9217 23273 9229 23307
rect 9263 23304 9275 23307
rect 9398 23304 9404 23316
rect 9263 23276 9404 23304
rect 9263 23273 9275 23276
rect 9217 23267 9275 23273
rect 8294 23196 8300 23248
rect 8352 23236 8358 23248
rect 9232 23236 9260 23267
rect 9398 23264 9404 23276
rect 9456 23264 9462 23316
rect 13170 23264 13176 23316
rect 13228 23304 13234 23316
rect 13722 23304 13728 23316
rect 13228 23276 13728 23304
rect 13228 23264 13234 23276
rect 13722 23264 13728 23276
rect 13780 23264 13786 23316
rect 18598 23264 18604 23316
rect 18656 23304 18662 23316
rect 18874 23304 18880 23316
rect 18656 23276 18880 23304
rect 18656 23264 18662 23276
rect 18874 23264 18880 23276
rect 18932 23264 18938 23316
rect 20162 23264 20168 23316
rect 20220 23264 20226 23316
rect 22281 23307 22339 23313
rect 22281 23304 22293 23307
rect 22066 23276 22293 23304
rect 8352 23208 9260 23236
rect 8352 23196 8358 23208
rect 9306 23196 9312 23248
rect 9364 23236 9370 23248
rect 11425 23239 11483 23245
rect 11425 23236 11437 23239
rect 9364 23208 11437 23236
rect 9364 23196 9370 23208
rect 11425 23205 11437 23208
rect 11471 23205 11483 23239
rect 11425 23199 11483 23205
rect 12066 23196 12072 23248
rect 12124 23236 12130 23248
rect 17126 23236 17132 23248
rect 12124 23208 17132 23236
rect 12124 23196 12130 23208
rect 17126 23196 17132 23208
rect 17184 23196 17190 23248
rect 6362 23168 6368 23180
rect 4356 23140 6368 23168
rect 2774 23060 2780 23112
rect 2832 23060 2838 23112
rect 4356 23109 4384 23140
rect 6362 23128 6368 23140
rect 6420 23128 6426 23180
rect 7006 23128 7012 23180
rect 7064 23128 7070 23180
rect 7282 23128 7288 23180
rect 7340 23128 7346 23180
rect 7653 23171 7711 23177
rect 7653 23137 7665 23171
rect 7699 23168 7711 23171
rect 9122 23168 9128 23180
rect 7699 23140 9128 23168
rect 7699 23137 7711 23140
rect 7653 23131 7711 23137
rect 4341 23103 4399 23109
rect 4341 23069 4353 23103
rect 4387 23069 4399 23103
rect 4341 23063 4399 23069
rect 934 22992 940 23044
rect 992 23032 998 23044
rect 1765 23035 1823 23041
rect 1765 23032 1777 23035
rect 992 23004 1777 23032
rect 992 22992 998 23004
rect 1765 23001 1777 23004
rect 1811 23001 1823 23035
rect 6730 23032 6736 23044
rect 6578 23004 6736 23032
rect 1765 22995 1823 23001
rect 6730 22992 6736 23004
rect 6788 23032 6794 23044
rect 7098 23032 7104 23044
rect 6788 23004 7104 23032
rect 6788 22992 6794 23004
rect 7098 22992 7104 23004
rect 7156 23032 7162 23044
rect 7668 23032 7696 23131
rect 9122 23128 9128 23140
rect 9180 23168 9186 23180
rect 9582 23168 9588 23180
rect 9180 23140 9588 23168
rect 9180 23128 9186 23140
rect 9582 23128 9588 23140
rect 9640 23168 9646 23180
rect 9766 23168 9772 23180
rect 9640 23140 9772 23168
rect 9640 23128 9646 23140
rect 9766 23128 9772 23140
rect 9824 23128 9830 23180
rect 10226 23128 10232 23180
rect 10284 23128 10290 23180
rect 11977 23171 12035 23177
rect 11977 23168 11989 23171
rect 10336 23140 11989 23168
rect 8662 23060 8668 23112
rect 8720 23100 8726 23112
rect 10336 23100 10364 23140
rect 11977 23137 11989 23140
rect 12023 23137 12035 23171
rect 12618 23168 12624 23180
rect 11977 23131 12035 23137
rect 12176 23140 12624 23168
rect 8720 23072 10364 23100
rect 11885 23103 11943 23109
rect 8720 23060 8726 23072
rect 11885 23069 11897 23103
rect 11931 23100 11943 23103
rect 12176 23100 12204 23140
rect 12618 23128 12624 23140
rect 12676 23128 12682 23180
rect 13265 23171 13323 23177
rect 13265 23137 13277 23171
rect 13311 23168 13323 23171
rect 13630 23168 13636 23180
rect 13311 23140 13636 23168
rect 13311 23137 13323 23140
rect 13265 23131 13323 23137
rect 13630 23128 13636 23140
rect 13688 23128 13694 23180
rect 15286 23128 15292 23180
rect 15344 23168 15350 23180
rect 17034 23168 17040 23180
rect 15344 23140 17040 23168
rect 15344 23128 15350 23140
rect 17034 23128 17040 23140
rect 17092 23128 17098 23180
rect 17402 23128 17408 23180
rect 17460 23128 17466 23180
rect 18966 23128 18972 23180
rect 19024 23168 19030 23180
rect 21266 23168 21272 23180
rect 19024 23140 21272 23168
rect 19024 23128 19030 23140
rect 21266 23128 21272 23140
rect 21324 23168 21330 23180
rect 21637 23171 21695 23177
rect 21637 23168 21649 23171
rect 21324 23140 21649 23168
rect 21324 23128 21330 23140
rect 21637 23137 21649 23140
rect 21683 23137 21695 23171
rect 21637 23131 21695 23137
rect 12986 23100 12992 23112
rect 11931 23072 12204 23100
rect 12452 23072 12992 23100
rect 11931 23069 11943 23072
rect 11885 23063 11943 23069
rect 7156 23004 7696 23032
rect 9953 23035 10011 23041
rect 7156 22992 7162 23004
rect 9953 23001 9965 23035
rect 9999 23032 10011 23035
rect 10781 23035 10839 23041
rect 10781 23032 10793 23035
rect 9999 23004 10793 23032
rect 9999 23001 10011 23004
rect 9953 22995 10011 23001
rect 10781 23001 10793 23004
rect 10827 23001 10839 23035
rect 10781 22995 10839 23001
rect 11793 23035 11851 23041
rect 11793 23001 11805 23035
rect 11839 23032 11851 23035
rect 12452 23032 12480 23072
rect 12986 23060 12992 23072
rect 13044 23100 13050 23112
rect 15304 23100 15332 23128
rect 13044 23072 15332 23100
rect 13044 23060 13050 23072
rect 16942 23060 16948 23112
rect 17000 23100 17006 23112
rect 17129 23103 17187 23109
rect 17129 23100 17141 23103
rect 17000 23072 17141 23100
rect 17000 23060 17006 23072
rect 17129 23069 17141 23072
rect 17175 23069 17187 23103
rect 17129 23063 17187 23069
rect 21910 23060 21916 23112
rect 21968 23060 21974 23112
rect 11839 23004 12480 23032
rect 11839 23001 11851 23004
rect 11793 22995 11851 23001
rect 12526 22992 12532 23044
rect 12584 23032 12590 23044
rect 13081 23035 13139 23041
rect 13081 23032 13093 23035
rect 12584 23004 13093 23032
rect 12584 22992 12590 23004
rect 13081 23001 13093 23004
rect 13127 23001 13139 23035
rect 19337 23035 19395 23041
rect 19337 23032 19349 23035
rect 18630 23004 19349 23032
rect 13081 22995 13139 23001
rect 19337 23001 19349 23004
rect 19383 23001 19395 23035
rect 22066 23032 22094 23276
rect 22281 23273 22293 23276
rect 22327 23304 22339 23307
rect 22370 23304 22376 23316
rect 22327 23276 22376 23304
rect 22327 23273 22339 23276
rect 22281 23267 22339 23273
rect 22370 23264 22376 23276
rect 22428 23304 22434 23316
rect 24394 23304 24400 23316
rect 22428 23276 24400 23304
rect 22428 23264 22434 23276
rect 24394 23264 24400 23276
rect 24452 23264 24458 23316
rect 23385 23171 23443 23177
rect 23385 23137 23397 23171
rect 23431 23168 23443 23171
rect 24854 23168 24860 23180
rect 23431 23140 24860 23168
rect 23431 23137 23443 23140
rect 23385 23131 23443 23137
rect 24854 23128 24860 23140
rect 24912 23128 24918 23180
rect 25225 23171 25283 23177
rect 25225 23137 25237 23171
rect 25271 23168 25283 23171
rect 25406 23168 25412 23180
rect 25271 23140 25412 23168
rect 25271 23137 25283 23140
rect 25225 23131 25283 23137
rect 25406 23128 25412 23140
rect 25464 23128 25470 23180
rect 24029 23103 24087 23109
rect 24029 23069 24041 23103
rect 24075 23100 24087 23103
rect 24302 23100 24308 23112
rect 24075 23072 24308 23100
rect 24075 23069 24087 23072
rect 24029 23063 24087 23069
rect 24302 23060 24308 23072
rect 24360 23060 24366 23112
rect 24949 23103 25007 23109
rect 24949 23069 24961 23103
rect 24995 23100 25007 23103
rect 25038 23100 25044 23112
rect 24995 23072 25044 23100
rect 24995 23069 25007 23072
rect 24949 23063 25007 23069
rect 25038 23060 25044 23072
rect 25096 23060 25102 23112
rect 21206 23004 22094 23032
rect 19337 22995 19395 23001
rect 5537 22967 5595 22973
rect 5537 22933 5549 22967
rect 5583 22964 5595 22967
rect 5626 22964 5632 22976
rect 5583 22936 5632 22964
rect 5583 22933 5595 22936
rect 5537 22927 5595 22933
rect 5626 22924 5632 22936
rect 5684 22964 5690 22976
rect 6822 22964 6828 22976
rect 5684 22936 6828 22964
rect 5684 22924 5690 22936
rect 6822 22924 6828 22936
rect 6880 22924 6886 22976
rect 8386 22924 8392 22976
rect 8444 22924 8450 22976
rect 9582 22924 9588 22976
rect 9640 22924 9646 22976
rect 10045 22967 10103 22973
rect 10045 22933 10057 22967
rect 10091 22964 10103 22967
rect 11054 22964 11060 22976
rect 10091 22936 11060 22964
rect 10091 22933 10103 22936
rect 10045 22927 10103 22933
rect 11054 22924 11060 22936
rect 11112 22924 11118 22976
rect 12434 22924 12440 22976
rect 12492 22964 12498 22976
rect 12621 22967 12679 22973
rect 12621 22964 12633 22967
rect 12492 22936 12633 22964
rect 12492 22924 12498 22936
rect 12621 22933 12633 22936
rect 12667 22933 12679 22967
rect 12621 22927 12679 22933
rect 12989 22967 13047 22973
rect 12989 22933 13001 22967
rect 13035 22964 13047 22967
rect 13170 22964 13176 22976
rect 13035 22936 13176 22964
rect 13035 22933 13047 22936
rect 12989 22927 13047 22933
rect 13170 22924 13176 22936
rect 13228 22924 13234 22976
rect 13722 22924 13728 22976
rect 13780 22964 13786 22976
rect 15378 22964 15384 22976
rect 13780 22936 15384 22964
rect 13780 22924 13786 22936
rect 15378 22924 15384 22936
rect 15436 22924 15442 22976
rect 19352 22964 19380 22995
rect 21284 22964 21312 23004
rect 19352 22936 21312 22964
rect 24578 22924 24584 22976
rect 24636 22924 24642 22976
rect 25041 22967 25099 22973
rect 25041 22933 25053 22967
rect 25087 22964 25099 22967
rect 25498 22964 25504 22976
rect 25087 22936 25504 22964
rect 25087 22933 25099 22936
rect 25041 22927 25099 22933
rect 25498 22924 25504 22936
rect 25556 22924 25562 22976
rect 1104 22874 25852 22896
rect 1104 22822 7950 22874
rect 8002 22822 8014 22874
rect 8066 22822 8078 22874
rect 8130 22822 8142 22874
rect 8194 22822 8206 22874
rect 8258 22822 17950 22874
rect 18002 22822 18014 22874
rect 18066 22822 18078 22874
rect 18130 22822 18142 22874
rect 18194 22822 18206 22874
rect 18258 22822 25852 22874
rect 1104 22800 25852 22822
rect 1762 22720 1768 22772
rect 1820 22760 1826 22772
rect 1949 22763 2007 22769
rect 1949 22760 1961 22763
rect 1820 22732 1961 22760
rect 1820 22720 1826 22732
rect 1949 22729 1961 22732
rect 1995 22729 2007 22763
rect 1949 22723 2007 22729
rect 2222 22720 2228 22772
rect 2280 22760 2286 22772
rect 2593 22763 2651 22769
rect 2593 22760 2605 22763
rect 2280 22732 2605 22760
rect 2280 22720 2286 22732
rect 2593 22729 2605 22732
rect 2639 22729 2651 22763
rect 2593 22723 2651 22729
rect 3878 22720 3884 22772
rect 3936 22760 3942 22772
rect 4019 22763 4077 22769
rect 4019 22760 4031 22763
rect 3936 22732 4031 22760
rect 3936 22720 3942 22732
rect 4019 22729 4031 22732
rect 4065 22729 4077 22763
rect 8386 22760 8392 22772
rect 4019 22723 4077 22729
rect 8220 22732 8392 22760
rect 7282 22652 7288 22704
rect 7340 22692 7346 22704
rect 8220 22701 8248 22732
rect 8386 22720 8392 22732
rect 8444 22760 8450 22772
rect 10502 22760 10508 22772
rect 8444 22732 10508 22760
rect 8444 22720 8450 22732
rect 10502 22720 10508 22732
rect 10560 22720 10566 22772
rect 10781 22763 10839 22769
rect 10781 22729 10793 22763
rect 10827 22760 10839 22763
rect 11054 22760 11060 22772
rect 10827 22732 11060 22760
rect 10827 22729 10839 22732
rect 10781 22723 10839 22729
rect 11054 22720 11060 22732
rect 11112 22760 11118 22772
rect 12250 22760 12256 22772
rect 11112 22732 12256 22760
rect 11112 22720 11118 22732
rect 12250 22720 12256 22732
rect 12308 22720 12314 22772
rect 12713 22763 12771 22769
rect 12713 22729 12725 22763
rect 12759 22760 12771 22763
rect 12986 22760 12992 22772
rect 12759 22732 12992 22760
rect 12759 22729 12771 22732
rect 12713 22723 12771 22729
rect 12986 22720 12992 22732
rect 13044 22720 13050 22772
rect 13446 22720 13452 22772
rect 13504 22760 13510 22772
rect 13504 22732 13676 22760
rect 13504 22720 13510 22732
rect 7377 22695 7435 22701
rect 7377 22692 7389 22695
rect 7340 22664 7389 22692
rect 7340 22652 7346 22664
rect 7377 22661 7389 22664
rect 7423 22661 7435 22695
rect 7377 22655 7435 22661
rect 8205 22695 8263 22701
rect 8205 22661 8217 22695
rect 8251 22661 8263 22695
rect 8205 22655 8263 22661
rect 9122 22652 9128 22704
rect 9180 22652 9186 22704
rect 9858 22652 9864 22704
rect 9916 22692 9922 22704
rect 10137 22695 10195 22701
rect 10137 22692 10149 22695
rect 9916 22664 10149 22692
rect 9916 22652 9922 22664
rect 10137 22661 10149 22664
rect 10183 22661 10195 22695
rect 10137 22655 10195 22661
rect 10686 22652 10692 22704
rect 10744 22692 10750 22704
rect 10965 22695 11023 22701
rect 10965 22692 10977 22695
rect 10744 22664 10977 22692
rect 10744 22652 10750 22664
rect 10965 22661 10977 22664
rect 11011 22661 11023 22695
rect 10965 22655 11023 22661
rect 12526 22652 12532 22704
rect 12584 22652 12590 22704
rect 12897 22695 12955 22701
rect 12897 22661 12909 22695
rect 12943 22692 12955 22695
rect 13538 22692 13544 22704
rect 12943 22664 13544 22692
rect 12943 22661 12955 22664
rect 12897 22655 12955 22661
rect 13538 22652 13544 22664
rect 13596 22652 13602 22704
rect 13648 22701 13676 22732
rect 14550 22720 14556 22772
rect 14608 22760 14614 22772
rect 15105 22763 15163 22769
rect 15105 22760 15117 22763
rect 14608 22732 15117 22760
rect 14608 22720 14614 22732
rect 15105 22729 15117 22732
rect 15151 22760 15163 22763
rect 15654 22760 15660 22772
rect 15151 22732 15660 22760
rect 15151 22729 15163 22732
rect 15105 22723 15163 22729
rect 15654 22720 15660 22732
rect 15712 22720 15718 22772
rect 15749 22763 15807 22769
rect 15749 22729 15761 22763
rect 15795 22760 15807 22763
rect 21082 22760 21088 22772
rect 15795 22732 21088 22760
rect 15795 22729 15807 22732
rect 15749 22723 15807 22729
rect 21082 22720 21088 22732
rect 21140 22720 21146 22772
rect 21450 22720 21456 22772
rect 21508 22760 21514 22772
rect 22186 22760 22192 22772
rect 21508 22732 22192 22760
rect 21508 22720 21514 22732
rect 22186 22720 22192 22732
rect 22244 22760 22250 22772
rect 22244 22732 23244 22760
rect 22244 22720 22250 22732
rect 13633 22695 13691 22701
rect 13633 22661 13645 22695
rect 13679 22692 13691 22695
rect 13722 22692 13728 22704
rect 13679 22664 13728 22692
rect 13679 22661 13691 22664
rect 13633 22655 13691 22661
rect 13722 22652 13728 22664
rect 13780 22652 13786 22704
rect 16114 22692 16120 22704
rect 14858 22664 16120 22692
rect 16114 22652 16120 22664
rect 16172 22652 16178 22704
rect 16485 22695 16543 22701
rect 16485 22661 16497 22695
rect 16531 22692 16543 22695
rect 17129 22695 17187 22701
rect 17129 22692 17141 22695
rect 16531 22664 17141 22692
rect 16531 22661 16543 22664
rect 16485 22655 16543 22661
rect 17129 22661 17141 22664
rect 17175 22692 17187 22695
rect 17862 22692 17868 22704
rect 17175 22664 17868 22692
rect 17175 22661 17187 22664
rect 17129 22655 17187 22661
rect 17862 22652 17868 22664
rect 17920 22652 17926 22704
rect 21361 22695 21419 22701
rect 21361 22692 21373 22695
rect 20378 22664 21373 22692
rect 21361 22661 21373 22664
rect 21407 22661 21419 22695
rect 21361 22655 21419 22661
rect 2130 22584 2136 22636
rect 2188 22584 2194 22636
rect 2866 22584 2872 22636
rect 2924 22624 2930 22636
rect 3053 22627 3111 22633
rect 3053 22624 3065 22627
rect 2924 22596 3065 22624
rect 2924 22584 2930 22596
rect 3053 22593 3065 22596
rect 3099 22624 3111 22627
rect 3326 22624 3332 22636
rect 3099 22596 3332 22624
rect 3099 22593 3111 22596
rect 3053 22587 3111 22593
rect 3326 22584 3332 22596
rect 3384 22584 3390 22636
rect 3878 22584 3884 22636
rect 3936 22633 3942 22636
rect 3936 22627 3974 22633
rect 3962 22593 3974 22627
rect 3936 22587 3974 22593
rect 3936 22584 3942 22587
rect 5534 22584 5540 22636
rect 5592 22584 5598 22636
rect 5629 22627 5687 22633
rect 5629 22593 5641 22627
rect 5675 22624 5687 22627
rect 7742 22624 7748 22636
rect 5675 22596 7748 22624
rect 5675 22593 5687 22596
rect 5629 22587 5687 22593
rect 7742 22584 7748 22596
rect 7800 22584 7806 22636
rect 10413 22627 10471 22633
rect 10413 22593 10425 22627
rect 10459 22624 10471 22627
rect 10870 22624 10876 22636
rect 10459 22596 10876 22624
rect 10459 22593 10471 22596
rect 10413 22587 10471 22593
rect 10870 22584 10876 22596
rect 10928 22624 10934 22636
rect 11238 22624 11244 22636
rect 10928 22596 11244 22624
rect 10928 22584 10934 22596
rect 11238 22584 11244 22596
rect 11296 22624 11302 22636
rect 13354 22624 13360 22636
rect 11296 22596 13360 22624
rect 11296 22584 11302 22596
rect 13354 22584 13360 22596
rect 13412 22584 13418 22636
rect 15565 22627 15623 22633
rect 15565 22593 15577 22627
rect 15611 22593 15623 22627
rect 15565 22587 15623 22593
rect 17221 22627 17279 22633
rect 17221 22593 17233 22627
rect 17267 22624 17279 22627
rect 18049 22627 18107 22633
rect 18049 22624 18061 22627
rect 17267 22596 18061 22624
rect 17267 22593 17279 22596
rect 17221 22587 17279 22593
rect 18049 22593 18061 22596
rect 18095 22593 18107 22627
rect 21376 22624 21404 22655
rect 21634 22652 21640 22704
rect 21692 22692 21698 22704
rect 23216 22701 23244 22732
rect 24486 22720 24492 22772
rect 24544 22760 24550 22772
rect 25133 22763 25191 22769
rect 25133 22760 25145 22763
rect 24544 22732 25145 22760
rect 24544 22720 24550 22732
rect 25133 22729 25145 22732
rect 25179 22729 25191 22763
rect 25133 22723 25191 22729
rect 22281 22695 22339 22701
rect 22281 22692 22293 22695
rect 21692 22664 22293 22692
rect 21692 22652 21698 22664
rect 22281 22661 22293 22664
rect 22327 22661 22339 22695
rect 22281 22655 22339 22661
rect 23201 22695 23259 22701
rect 23201 22661 23213 22695
rect 23247 22661 23259 22695
rect 23201 22655 23259 22661
rect 22370 22624 22376 22636
rect 21376 22596 22376 22624
rect 18049 22587 18107 22593
rect 3237 22559 3295 22565
rect 3237 22525 3249 22559
rect 3283 22556 3295 22559
rect 4890 22556 4896 22568
rect 3283 22528 4896 22556
rect 3283 22525 3295 22528
rect 3237 22519 3295 22525
rect 4890 22516 4896 22528
rect 4948 22516 4954 22568
rect 5718 22516 5724 22568
rect 5776 22516 5782 22568
rect 8662 22516 8668 22568
rect 8720 22516 8726 22568
rect 12345 22559 12403 22565
rect 12345 22525 12357 22559
rect 12391 22556 12403 22559
rect 12618 22556 12624 22568
rect 12391 22528 12624 22556
rect 12391 22525 12403 22528
rect 12345 22519 12403 22525
rect 12618 22516 12624 22528
rect 12676 22556 12682 22568
rect 13170 22556 13176 22568
rect 12676 22528 13176 22556
rect 12676 22516 12682 22528
rect 13170 22516 13176 22528
rect 13228 22516 13234 22568
rect 15580 22556 15608 22587
rect 22370 22584 22376 22596
rect 22428 22584 22434 22636
rect 22830 22584 22836 22636
rect 22888 22624 22894 22636
rect 22925 22627 22983 22633
rect 22925 22624 22937 22627
rect 22888 22596 22937 22624
rect 22888 22584 22894 22596
rect 22925 22593 22937 22596
rect 22971 22593 22983 22627
rect 24486 22624 24492 22636
rect 24334 22596 24492 22624
rect 22925 22587 22983 22593
rect 24486 22584 24492 22596
rect 24544 22584 24550 22636
rect 25314 22584 25320 22636
rect 25372 22584 25378 22636
rect 14660 22528 15608 22556
rect 17037 22559 17095 22565
rect 11514 22448 11520 22500
rect 11572 22488 11578 22500
rect 11572 22460 13492 22488
rect 11572 22448 11578 22460
rect 4154 22380 4160 22432
rect 4212 22420 4218 22432
rect 5169 22423 5227 22429
rect 5169 22420 5181 22423
rect 4212 22392 5181 22420
rect 4212 22380 4218 22392
rect 5169 22389 5181 22392
rect 5215 22389 5227 22423
rect 13464 22420 13492 22460
rect 14660 22420 14688 22528
rect 17037 22525 17049 22559
rect 17083 22525 17095 22559
rect 17037 22519 17095 22525
rect 17052 22488 17080 22519
rect 17494 22516 17500 22568
rect 17552 22556 17558 22568
rect 19061 22559 19119 22565
rect 19061 22556 19073 22559
rect 17552 22528 19073 22556
rect 17552 22516 17558 22528
rect 19061 22525 19073 22528
rect 19107 22525 19119 22559
rect 19061 22519 19119 22525
rect 20806 22516 20812 22568
rect 20864 22516 20870 22568
rect 21085 22559 21143 22565
rect 21085 22525 21097 22559
rect 21131 22556 21143 22559
rect 21910 22556 21916 22568
rect 21131 22528 21916 22556
rect 21131 22525 21143 22528
rect 21085 22519 21143 22525
rect 18966 22488 18972 22500
rect 17052 22460 18972 22488
rect 18966 22448 18972 22460
rect 19024 22448 19030 22500
rect 13464 22392 14688 22420
rect 17589 22423 17647 22429
rect 5169 22383 5227 22389
rect 17589 22389 17601 22423
rect 17635 22420 17647 22423
rect 18414 22420 18420 22432
rect 17635 22392 18420 22420
rect 17635 22389 17647 22392
rect 17589 22383 17647 22389
rect 18414 22380 18420 22392
rect 18472 22380 18478 22432
rect 18690 22380 18696 22432
rect 18748 22420 18754 22432
rect 21100 22420 21128 22519
rect 21910 22516 21916 22528
rect 21968 22516 21974 22568
rect 21266 22448 21272 22500
rect 21324 22488 21330 22500
rect 21634 22488 21640 22500
rect 21324 22460 21640 22488
rect 21324 22448 21330 22460
rect 21634 22448 21640 22460
rect 21692 22448 21698 22500
rect 18748 22392 21128 22420
rect 22373 22423 22431 22429
rect 18748 22380 18754 22392
rect 22373 22389 22385 22423
rect 22419 22420 22431 22423
rect 23934 22420 23940 22432
rect 22419 22392 23940 22420
rect 22419 22389 22431 22392
rect 22373 22383 22431 22389
rect 23934 22380 23940 22392
rect 23992 22380 23998 22432
rect 24302 22380 24308 22432
rect 24360 22420 24366 22432
rect 24673 22423 24731 22429
rect 24673 22420 24685 22423
rect 24360 22392 24685 22420
rect 24360 22380 24366 22392
rect 24673 22389 24685 22392
rect 24719 22389 24731 22423
rect 24673 22383 24731 22389
rect 1104 22330 25852 22352
rect 1104 22278 2950 22330
rect 3002 22278 3014 22330
rect 3066 22278 3078 22330
rect 3130 22278 3142 22330
rect 3194 22278 3206 22330
rect 3258 22278 12950 22330
rect 13002 22278 13014 22330
rect 13066 22278 13078 22330
rect 13130 22278 13142 22330
rect 13194 22278 13206 22330
rect 13258 22278 22950 22330
rect 23002 22278 23014 22330
rect 23066 22278 23078 22330
rect 23130 22278 23142 22330
rect 23194 22278 23206 22330
rect 23258 22278 25852 22330
rect 1104 22256 25852 22278
rect 5534 22176 5540 22228
rect 5592 22216 5598 22228
rect 6181 22219 6239 22225
rect 6181 22216 6193 22219
rect 5592 22188 6193 22216
rect 5592 22176 5598 22188
rect 6181 22185 6193 22188
rect 6227 22185 6239 22219
rect 6181 22179 6239 22185
rect 12158 22176 12164 22228
rect 12216 22216 12222 22228
rect 12526 22216 12532 22228
rect 12216 22188 12532 22216
rect 12216 22176 12222 22188
rect 12526 22176 12532 22188
rect 12584 22176 12590 22228
rect 13538 22176 13544 22228
rect 13596 22216 13602 22228
rect 15930 22216 15936 22228
rect 13596 22188 15936 22216
rect 13596 22176 13602 22188
rect 15930 22176 15936 22188
rect 15988 22176 15994 22228
rect 17402 22176 17408 22228
rect 17460 22176 17466 22228
rect 19702 22216 19708 22228
rect 19306 22188 19708 22216
rect 3418 22148 3424 22160
rect 2884 22120 3424 22148
rect 2884 22080 2912 22120
rect 3418 22108 3424 22120
rect 3476 22108 3482 22160
rect 5258 22108 5264 22160
rect 5316 22148 5322 22160
rect 5316 22120 8064 22148
rect 5316 22108 5322 22120
rect 2240 22052 2912 22080
rect 2240 22021 2268 22052
rect 6822 22040 6828 22092
rect 6880 22040 6886 22092
rect 8036 22089 8064 22120
rect 12452 22120 14872 22148
rect 8021 22083 8079 22089
rect 8021 22080 8033 22083
rect 7979 22052 8033 22080
rect 8021 22049 8033 22052
rect 8067 22080 8079 22083
rect 8386 22080 8392 22092
rect 8067 22052 8392 22080
rect 8067 22049 8079 22052
rect 8021 22043 8079 22049
rect 8386 22040 8392 22052
rect 8444 22040 8450 22092
rect 11330 22040 11336 22092
rect 11388 22040 11394 22092
rect 11882 22040 11888 22092
rect 11940 22080 11946 22092
rect 12452 22089 12480 22120
rect 12437 22083 12495 22089
rect 12437 22080 12449 22083
rect 11940 22052 12449 22080
rect 11940 22040 11946 22052
rect 12437 22049 12449 22052
rect 12483 22049 12495 22083
rect 12437 22043 12495 22049
rect 12986 22040 12992 22092
rect 13044 22080 13050 22092
rect 13538 22080 13544 22092
rect 13044 22052 13544 22080
rect 13044 22040 13050 22052
rect 13538 22040 13544 22052
rect 13596 22040 13602 22092
rect 14844 22089 14872 22120
rect 17310 22108 17316 22160
rect 17368 22148 17374 22160
rect 19306 22148 19334 22188
rect 19702 22176 19708 22188
rect 19760 22176 19766 22228
rect 22005 22219 22063 22225
rect 22005 22185 22017 22219
rect 22051 22216 22063 22219
rect 22370 22216 22376 22228
rect 22051 22188 22376 22216
rect 22051 22185 22063 22188
rect 22005 22179 22063 22185
rect 22370 22176 22376 22188
rect 22428 22176 22434 22228
rect 25314 22176 25320 22228
rect 25372 22216 25378 22228
rect 25409 22219 25467 22225
rect 25409 22216 25421 22219
rect 25372 22188 25421 22216
rect 25372 22176 25378 22188
rect 25409 22185 25421 22188
rect 25455 22185 25467 22219
rect 25409 22179 25467 22185
rect 22094 22148 22100 22160
rect 17368 22120 19334 22148
rect 19628 22120 22100 22148
rect 17368 22108 17374 22120
rect 14829 22083 14887 22089
rect 14829 22049 14841 22083
rect 14875 22080 14887 22083
rect 15657 22083 15715 22089
rect 14875 22052 14909 22080
rect 14875 22049 14887 22052
rect 14829 22043 14887 22049
rect 15657 22049 15669 22083
rect 15703 22080 15715 22083
rect 16942 22080 16948 22092
rect 15703 22052 16948 22080
rect 15703 22049 15715 22052
rect 15657 22043 15715 22049
rect 16942 22040 16948 22052
rect 17000 22080 17006 22092
rect 18690 22080 18696 22092
rect 17000 22052 18696 22080
rect 17000 22040 17006 22052
rect 18690 22040 18696 22052
rect 18748 22040 18754 22092
rect 19628 22089 19656 22120
rect 22094 22108 22100 22120
rect 22152 22148 22158 22160
rect 24302 22148 24308 22160
rect 22152 22120 24308 22148
rect 22152 22108 22158 22120
rect 24302 22108 24308 22120
rect 24360 22108 24366 22160
rect 24486 22108 24492 22160
rect 24544 22148 24550 22160
rect 24765 22151 24823 22157
rect 24765 22148 24777 22151
rect 24544 22120 24777 22148
rect 24544 22108 24550 22120
rect 24765 22117 24777 22120
rect 24811 22148 24823 22151
rect 24811 22120 24992 22148
rect 24811 22117 24823 22120
rect 24765 22111 24823 22117
rect 19613 22083 19671 22089
rect 19613 22049 19625 22083
rect 19659 22080 19671 22083
rect 21453 22083 21511 22089
rect 19659 22052 19693 22080
rect 19659 22049 19671 22052
rect 19613 22043 19671 22049
rect 21453 22049 21465 22083
rect 21499 22080 21511 22083
rect 22830 22080 22836 22092
rect 21499 22052 22836 22080
rect 21499 22049 21511 22052
rect 21453 22043 21511 22049
rect 22830 22040 22836 22052
rect 22888 22040 22894 22092
rect 23385 22083 23443 22089
rect 23385 22049 23397 22083
rect 23431 22080 23443 22083
rect 24854 22080 24860 22092
rect 23431 22052 24860 22080
rect 23431 22049 23443 22052
rect 23385 22043 23443 22049
rect 24854 22040 24860 22052
rect 24912 22040 24918 22092
rect 24964 22080 24992 22120
rect 25038 22080 25044 22092
rect 24964 22052 25044 22080
rect 25038 22040 25044 22052
rect 25096 22040 25102 22092
rect 2225 22015 2283 22021
rect 2225 21981 2237 22015
rect 2271 21981 2283 22015
rect 2225 21975 2283 21981
rect 2866 21972 2872 22024
rect 2924 21972 2930 22024
rect 6546 21972 6552 22024
rect 6604 21972 6610 22024
rect 7745 22015 7803 22021
rect 7745 21981 7757 22015
rect 7791 22012 7803 22015
rect 9582 22012 9588 22024
rect 7791 21984 9588 22012
rect 7791 21981 7803 21984
rect 7745 21975 7803 21981
rect 9582 21972 9588 21984
rect 9640 21972 9646 22024
rect 13357 22015 13415 22021
rect 13357 21981 13369 22015
rect 13403 22012 13415 22015
rect 14274 22012 14280 22024
rect 13403 21984 14280 22012
rect 13403 21981 13415 21984
rect 13357 21975 13415 21981
rect 14274 21972 14280 21984
rect 14332 21972 14338 22024
rect 14645 22015 14703 22021
rect 14645 21981 14657 22015
rect 14691 22012 14703 22015
rect 19705 22015 19763 22021
rect 14691 21984 15608 22012
rect 14691 21981 14703 21984
rect 14645 21975 14703 21981
rect 10502 21904 10508 21956
rect 10560 21944 10566 21956
rect 11514 21944 11520 21956
rect 10560 21916 11520 21944
rect 10560 21904 10566 21916
rect 11514 21904 11520 21916
rect 11572 21904 11578 21956
rect 12158 21904 12164 21956
rect 12216 21944 12222 21956
rect 12345 21947 12403 21953
rect 12345 21944 12357 21947
rect 12216 21916 12357 21944
rect 12216 21904 12222 21916
rect 12345 21913 12357 21916
rect 12391 21913 12403 21947
rect 12345 21907 12403 21913
rect 1762 21836 1768 21888
rect 1820 21876 1826 21888
rect 2041 21879 2099 21885
rect 2041 21876 2053 21879
rect 1820 21848 2053 21876
rect 1820 21836 1826 21848
rect 2041 21845 2053 21848
rect 2087 21845 2099 21879
rect 2041 21839 2099 21845
rect 2685 21879 2743 21885
rect 2685 21845 2697 21879
rect 2731 21876 2743 21879
rect 2774 21876 2780 21888
rect 2731 21848 2780 21876
rect 2731 21845 2743 21848
rect 2685 21839 2743 21845
rect 2774 21836 2780 21848
rect 2832 21836 2838 21888
rect 6641 21879 6699 21885
rect 6641 21845 6653 21879
rect 6687 21876 6699 21879
rect 7282 21876 7288 21888
rect 6687 21848 7288 21876
rect 6687 21845 6699 21848
rect 6641 21839 6699 21845
rect 7282 21836 7288 21848
rect 7340 21836 7346 21888
rect 7374 21836 7380 21888
rect 7432 21836 7438 21888
rect 7834 21836 7840 21888
rect 7892 21836 7898 21888
rect 9030 21836 9036 21888
rect 9088 21876 9094 21888
rect 11885 21879 11943 21885
rect 11885 21876 11897 21879
rect 9088 21848 11897 21876
rect 9088 21836 9094 21848
rect 11885 21845 11897 21848
rect 11931 21845 11943 21879
rect 11885 21839 11943 21845
rect 12253 21879 12311 21885
rect 12253 21845 12265 21879
rect 12299 21876 12311 21879
rect 12986 21876 12992 21888
rect 12299 21848 12992 21876
rect 12299 21845 12311 21848
rect 12253 21839 12311 21845
rect 12986 21836 12992 21848
rect 13044 21836 13050 21888
rect 13173 21879 13231 21885
rect 13173 21845 13185 21879
rect 13219 21876 13231 21879
rect 13722 21876 13728 21888
rect 13219 21848 13728 21876
rect 13219 21845 13231 21848
rect 13173 21839 13231 21845
rect 13722 21836 13728 21848
rect 13780 21836 13786 21888
rect 13814 21836 13820 21888
rect 13872 21836 13878 21888
rect 14274 21836 14280 21888
rect 14332 21836 14338 21888
rect 14366 21836 14372 21888
rect 14424 21876 14430 21888
rect 14642 21876 14648 21888
rect 14424 21848 14648 21876
rect 14424 21836 14430 21848
rect 14642 21836 14648 21848
rect 14700 21836 14706 21888
rect 14734 21836 14740 21888
rect 14792 21836 14798 21888
rect 15381 21879 15439 21885
rect 15381 21845 15393 21879
rect 15427 21876 15439 21879
rect 15580 21876 15608 21984
rect 19705 21981 19717 22015
rect 19751 22012 19763 22015
rect 20714 22012 20720 22024
rect 19751 21984 20720 22012
rect 19751 21981 19763 21984
rect 19705 21975 19763 21981
rect 20714 21972 20720 21984
rect 20772 21972 20778 22024
rect 24029 22015 24087 22021
rect 24029 21981 24041 22015
rect 24075 22012 24087 22015
rect 24210 22012 24216 22024
rect 24075 21984 24216 22012
rect 24075 21981 24087 21984
rect 24029 21975 24087 21981
rect 24210 21972 24216 21984
rect 24268 21972 24274 22024
rect 15933 21947 15991 21953
rect 15933 21913 15945 21947
rect 15979 21944 15991 21947
rect 16022 21944 16028 21956
rect 15979 21916 16028 21944
rect 15979 21913 15991 21916
rect 15933 21907 15991 21913
rect 16022 21904 16028 21916
rect 16080 21904 16086 21956
rect 16206 21904 16212 21956
rect 16264 21944 16270 21956
rect 16264 21916 16422 21944
rect 16264 21904 16270 21916
rect 17770 21904 17776 21956
rect 17828 21944 17834 21956
rect 17957 21947 18015 21953
rect 17957 21944 17969 21947
rect 17828 21916 17969 21944
rect 17828 21904 17834 21916
rect 17957 21913 17969 21916
rect 18003 21944 18015 21947
rect 20625 21947 20683 21953
rect 20625 21944 20637 21947
rect 18003 21916 20637 21944
rect 18003 21913 18015 21916
rect 17957 21907 18015 21913
rect 20625 21913 20637 21916
rect 20671 21944 20683 21947
rect 21821 21947 21879 21953
rect 21821 21944 21833 21947
rect 20671 21916 21833 21944
rect 20671 21913 20683 21916
rect 20625 21907 20683 21913
rect 21821 21913 21833 21916
rect 21867 21913 21879 21947
rect 22370 21944 22376 21956
rect 21821 21907 21879 21913
rect 22066 21916 22376 21944
rect 17310 21876 17316 21888
rect 15427 21848 17316 21876
rect 15427 21845 15439 21848
rect 15381 21839 15439 21845
rect 17310 21836 17316 21848
rect 17368 21836 17374 21888
rect 19794 21836 19800 21888
rect 19852 21836 19858 21888
rect 20165 21879 20223 21885
rect 20165 21845 20177 21879
rect 20211 21876 20223 21879
rect 22066 21876 22094 21916
rect 22370 21904 22376 21916
rect 22428 21904 22434 21956
rect 20211 21848 22094 21876
rect 20211 21845 20223 21848
rect 20165 21839 20223 21845
rect 1104 21786 25852 21808
rect 1104 21734 7950 21786
rect 8002 21734 8014 21786
rect 8066 21734 8078 21786
rect 8130 21734 8142 21786
rect 8194 21734 8206 21786
rect 8258 21734 17950 21786
rect 18002 21734 18014 21786
rect 18066 21734 18078 21786
rect 18130 21734 18142 21786
rect 18194 21734 18206 21786
rect 18258 21734 25852 21786
rect 1104 21712 25852 21734
rect 2130 21632 2136 21684
rect 2188 21672 2194 21684
rect 2501 21675 2559 21681
rect 2501 21672 2513 21675
rect 2188 21644 2513 21672
rect 2188 21632 2194 21644
rect 2501 21641 2513 21644
rect 2547 21641 2559 21675
rect 2501 21635 2559 21641
rect 6454 21632 6460 21684
rect 6512 21672 6518 21684
rect 6549 21675 6607 21681
rect 6549 21672 6561 21675
rect 6512 21644 6561 21672
rect 6512 21632 6518 21644
rect 6549 21641 6561 21644
rect 6595 21641 6607 21675
rect 6549 21635 6607 21641
rect 6917 21675 6975 21681
rect 6917 21641 6929 21675
rect 6963 21672 6975 21675
rect 7374 21672 7380 21684
rect 6963 21644 7380 21672
rect 6963 21641 6975 21644
rect 6917 21635 6975 21641
rect 7374 21632 7380 21644
rect 7432 21632 7438 21684
rect 7742 21632 7748 21684
rect 7800 21632 7806 21684
rect 8205 21675 8263 21681
rect 8205 21641 8217 21675
rect 8251 21672 8263 21675
rect 9398 21672 9404 21684
rect 8251 21644 9404 21672
rect 8251 21641 8263 21644
rect 8205 21635 8263 21641
rect 9398 21632 9404 21644
rect 9456 21632 9462 21684
rect 10321 21675 10379 21681
rect 10321 21641 10333 21675
rect 10367 21672 10379 21675
rect 11054 21672 11060 21684
rect 10367 21644 11060 21672
rect 10367 21641 10379 21644
rect 10321 21635 10379 21641
rect 11054 21632 11060 21644
rect 11112 21632 11118 21684
rect 11514 21632 11520 21684
rect 11572 21672 11578 21684
rect 11609 21675 11667 21681
rect 11609 21672 11621 21675
rect 11572 21644 11621 21672
rect 11572 21632 11578 21644
rect 11609 21641 11621 21644
rect 11655 21672 11667 21675
rect 15194 21672 15200 21684
rect 11655 21644 15200 21672
rect 11655 21641 11667 21644
rect 11609 21635 11667 21641
rect 15194 21632 15200 21644
rect 15252 21672 15258 21684
rect 17770 21672 17776 21684
rect 15252 21644 17776 21672
rect 15252 21632 15258 21644
rect 17770 21632 17776 21644
rect 17828 21632 17834 21684
rect 18414 21632 18420 21684
rect 18472 21672 18478 21684
rect 18509 21675 18567 21681
rect 18509 21672 18521 21675
rect 18472 21644 18521 21672
rect 18472 21632 18478 21644
rect 18509 21641 18521 21644
rect 18555 21641 18567 21675
rect 18509 21635 18567 21641
rect 19794 21632 19800 21684
rect 19852 21672 19858 21684
rect 22005 21675 22063 21681
rect 22005 21672 22017 21675
rect 19852 21644 22017 21672
rect 19852 21632 19858 21644
rect 22005 21641 22017 21644
rect 22051 21641 22063 21675
rect 22005 21635 22063 21641
rect 25038 21632 25044 21684
rect 25096 21632 25102 21684
rect 6822 21564 6828 21616
rect 6880 21604 6886 21616
rect 6880 21576 8248 21604
rect 6880 21564 6886 21576
rect 3881 21539 3939 21545
rect 3881 21505 3893 21539
rect 3927 21536 3939 21539
rect 4154 21536 4160 21548
rect 3927 21508 4160 21536
rect 3927 21505 3939 21508
rect 3881 21499 3939 21505
rect 4154 21496 4160 21508
rect 4212 21496 4218 21548
rect 4338 21496 4344 21548
rect 4396 21536 4402 21548
rect 4893 21539 4951 21545
rect 4893 21536 4905 21539
rect 4396 21508 4905 21536
rect 4396 21496 4402 21508
rect 4893 21505 4905 21508
rect 4939 21505 4951 21539
rect 4893 21499 4951 21505
rect 7009 21539 7067 21545
rect 7009 21505 7021 21539
rect 7055 21536 7067 21539
rect 7055 21508 8064 21536
rect 7055 21505 7067 21508
rect 7009 21499 7067 21505
rect 2774 21428 2780 21480
rect 2832 21468 2838 21480
rect 2961 21471 3019 21477
rect 2961 21468 2973 21471
rect 2832 21440 2973 21468
rect 2832 21428 2838 21440
rect 2961 21437 2973 21440
rect 3007 21437 3019 21471
rect 2961 21431 3019 21437
rect 3145 21471 3203 21477
rect 3145 21437 3157 21471
rect 3191 21468 3203 21471
rect 3970 21468 3976 21480
rect 3191 21440 3976 21468
rect 3191 21437 3203 21440
rect 3145 21431 3203 21437
rect 2976 21400 3004 21431
rect 3970 21428 3976 21440
rect 4028 21428 4034 21480
rect 7101 21471 7159 21477
rect 7101 21437 7113 21471
rect 7147 21437 7159 21471
rect 7101 21431 7159 21437
rect 4062 21400 4068 21412
rect 2976 21372 4068 21400
rect 4062 21360 4068 21372
rect 4120 21400 4126 21412
rect 4433 21403 4491 21409
rect 4433 21400 4445 21403
rect 4120 21372 4445 21400
rect 4120 21360 4126 21372
rect 4433 21369 4445 21372
rect 4479 21369 4491 21403
rect 4433 21363 4491 21369
rect 6914 21360 6920 21412
rect 6972 21400 6978 21412
rect 7116 21400 7144 21431
rect 6972 21372 7144 21400
rect 6972 21360 6978 21372
rect 3418 21292 3424 21344
rect 3476 21332 3482 21344
rect 3697 21335 3755 21341
rect 3697 21332 3709 21335
rect 3476 21304 3709 21332
rect 3476 21292 3482 21304
rect 3697 21301 3709 21304
rect 3743 21301 3755 21335
rect 3697 21295 3755 21301
rect 4801 21335 4859 21341
rect 4801 21301 4813 21335
rect 4847 21332 4859 21335
rect 5718 21332 5724 21344
rect 4847 21304 5724 21332
rect 4847 21301 4859 21304
rect 4801 21295 4859 21301
rect 5718 21292 5724 21304
rect 5776 21292 5782 21344
rect 8036 21332 8064 21508
rect 8110 21496 8116 21548
rect 8168 21496 8174 21548
rect 8220 21536 8248 21576
rect 9950 21564 9956 21616
rect 10008 21604 10014 21616
rect 11701 21607 11759 21613
rect 11701 21604 11713 21607
rect 10008 21576 11713 21604
rect 10008 21564 10014 21576
rect 11701 21573 11713 21576
rect 11747 21604 11759 21607
rect 12158 21604 12164 21616
rect 11747 21576 12164 21604
rect 11747 21573 11759 21576
rect 11701 21567 11759 21573
rect 12158 21564 12164 21576
rect 12216 21564 12222 21616
rect 12618 21564 12624 21616
rect 12676 21604 12682 21616
rect 12989 21607 13047 21613
rect 12989 21604 13001 21607
rect 12676 21576 13001 21604
rect 12676 21564 12682 21576
rect 12989 21573 13001 21576
rect 13035 21573 13047 21607
rect 12989 21567 13047 21573
rect 15013 21607 15071 21613
rect 15013 21573 15025 21607
rect 15059 21604 15071 21607
rect 19334 21604 19340 21616
rect 15059 21576 19340 21604
rect 15059 21573 15071 21576
rect 15013 21567 15071 21573
rect 13081 21539 13139 21545
rect 8220 21508 8340 21536
rect 8312 21477 8340 21508
rect 13081 21505 13093 21539
rect 13127 21536 13139 21539
rect 13538 21536 13544 21548
rect 13127 21508 13544 21536
rect 13127 21505 13139 21508
rect 13081 21499 13139 21505
rect 13538 21496 13544 21508
rect 13596 21496 13602 21548
rect 14292 21545 14504 21560
rect 14277 21539 14504 21545
rect 14277 21505 14289 21539
rect 14323 21536 14504 21539
rect 15028 21536 15056 21567
rect 19334 21564 19340 21576
rect 19392 21564 19398 21616
rect 19426 21564 19432 21616
rect 19484 21604 19490 21616
rect 19484 21576 19918 21604
rect 19484 21564 19490 21576
rect 21634 21564 21640 21616
rect 21692 21604 21698 21616
rect 22649 21607 22707 21613
rect 22649 21604 22661 21607
rect 21692 21576 22661 21604
rect 21692 21564 21698 21576
rect 22649 21573 22661 21576
rect 22695 21573 22707 21607
rect 24854 21604 24860 21616
rect 23966 21576 24860 21604
rect 22649 21567 22707 21573
rect 24854 21564 24860 21576
rect 24912 21604 24918 21616
rect 25056 21604 25084 21632
rect 24912 21576 25084 21604
rect 24912 21564 24918 21576
rect 14323 21532 15056 21536
rect 14323 21505 14335 21532
rect 14476 21508 15056 21532
rect 14277 21499 14335 21505
rect 15470 21496 15476 21548
rect 15528 21496 15534 21548
rect 18417 21539 18475 21545
rect 18417 21505 18429 21539
rect 18463 21536 18475 21539
rect 18506 21536 18512 21548
rect 18463 21508 18512 21536
rect 18463 21505 18475 21508
rect 18417 21499 18475 21505
rect 18506 21496 18512 21508
rect 18564 21496 18570 21548
rect 21361 21539 21419 21545
rect 21361 21505 21373 21539
rect 21407 21536 21419 21539
rect 22094 21536 22100 21548
rect 21407 21508 22100 21536
rect 21407 21505 21419 21508
rect 21361 21499 21419 21505
rect 22094 21496 22100 21508
rect 22152 21536 22158 21548
rect 22830 21536 22836 21548
rect 22152 21508 22836 21536
rect 22152 21496 22158 21508
rect 22830 21496 22836 21508
rect 22888 21496 22894 21548
rect 8297 21471 8355 21477
rect 8297 21437 8309 21471
rect 8343 21437 8355 21471
rect 8297 21431 8355 21437
rect 9677 21471 9735 21477
rect 9677 21437 9689 21471
rect 9723 21468 9735 21471
rect 10226 21468 10232 21480
rect 9723 21440 10232 21468
rect 9723 21437 9735 21440
rect 9677 21431 9735 21437
rect 10226 21428 10232 21440
rect 10284 21468 10290 21480
rect 10413 21471 10471 21477
rect 10413 21468 10425 21471
rect 10284 21440 10425 21468
rect 10284 21428 10290 21440
rect 10413 21437 10425 21440
rect 10459 21437 10471 21471
rect 10413 21431 10471 21437
rect 10597 21471 10655 21477
rect 10597 21437 10609 21471
rect 10643 21468 10655 21471
rect 12710 21468 12716 21480
rect 10643 21440 12716 21468
rect 10643 21437 10655 21440
rect 10597 21431 10655 21437
rect 8478 21360 8484 21412
rect 8536 21400 8542 21412
rect 9953 21403 10011 21409
rect 9953 21400 9965 21403
rect 8536 21372 9965 21400
rect 8536 21360 8542 21372
rect 9953 21369 9965 21372
rect 9999 21369 10011 21403
rect 10428 21400 10456 21431
rect 12710 21428 12716 21440
rect 12768 21428 12774 21480
rect 12894 21428 12900 21480
rect 12952 21428 12958 21480
rect 14366 21428 14372 21480
rect 14424 21428 14430 21480
rect 14461 21471 14519 21477
rect 14461 21437 14473 21471
rect 14507 21437 14519 21471
rect 14461 21431 14519 21437
rect 11422 21400 11428 21412
rect 10428 21372 11428 21400
rect 9953 21363 10011 21369
rect 11422 21360 11428 21372
rect 11480 21360 11486 21412
rect 13909 21403 13967 21409
rect 13909 21400 13921 21403
rect 13188 21372 13921 21400
rect 9122 21332 9128 21344
rect 8036 21304 9128 21332
rect 9122 21292 9128 21304
rect 9180 21292 9186 21344
rect 12158 21292 12164 21344
rect 12216 21332 12222 21344
rect 13188 21332 13216 21372
rect 13909 21369 13921 21372
rect 13955 21369 13967 21403
rect 13909 21363 13967 21369
rect 13998 21360 14004 21412
rect 14056 21400 14062 21412
rect 14476 21400 14504 21431
rect 14642 21428 14648 21480
rect 14700 21468 14706 21480
rect 15105 21471 15163 21477
rect 15105 21468 15117 21471
rect 14700 21440 15117 21468
rect 14700 21428 14706 21440
rect 15105 21437 15117 21440
rect 15151 21437 15163 21471
rect 15105 21431 15163 21437
rect 18325 21471 18383 21477
rect 18325 21437 18337 21471
rect 18371 21468 18383 21471
rect 20070 21468 20076 21480
rect 18371 21440 20076 21468
rect 18371 21437 18383 21440
rect 18325 21431 18383 21437
rect 20070 21428 20076 21440
rect 20128 21468 20134 21480
rect 21085 21471 21143 21477
rect 21085 21468 21097 21471
rect 20128 21440 21097 21468
rect 20128 21428 20134 21440
rect 21085 21437 21097 21440
rect 21131 21437 21143 21471
rect 21085 21431 21143 21437
rect 24394 21428 24400 21480
rect 24452 21428 24458 21480
rect 24673 21471 24731 21477
rect 24673 21437 24685 21471
rect 24719 21468 24731 21471
rect 25038 21468 25044 21480
rect 24719 21440 25044 21468
rect 24719 21437 24731 21440
rect 24673 21431 24731 21437
rect 14056 21372 14504 21400
rect 15657 21403 15715 21409
rect 14056 21360 14062 21372
rect 15657 21369 15669 21403
rect 15703 21400 15715 21403
rect 17862 21400 17868 21412
rect 15703 21372 17868 21400
rect 15703 21369 15715 21372
rect 15657 21363 15715 21369
rect 17862 21360 17868 21372
rect 17920 21360 17926 21412
rect 19426 21400 19432 21412
rect 18432 21372 19432 21400
rect 12216 21304 13216 21332
rect 13449 21335 13507 21341
rect 12216 21292 12222 21304
rect 13449 21301 13461 21335
rect 13495 21332 13507 21335
rect 14734 21332 14740 21344
rect 13495 21304 14740 21332
rect 13495 21301 13507 21304
rect 13449 21295 13507 21301
rect 14734 21292 14740 21304
rect 14792 21292 14798 21344
rect 16206 21292 16212 21344
rect 16264 21332 16270 21344
rect 17497 21335 17555 21341
rect 17497 21332 17509 21335
rect 16264 21304 17509 21332
rect 16264 21292 16270 21304
rect 17497 21301 17509 21304
rect 17543 21332 17555 21335
rect 18432 21332 18460 21372
rect 19426 21360 19432 21372
rect 19484 21360 19490 21412
rect 17543 21304 18460 21332
rect 17543 21301 17555 21304
rect 17497 21295 17555 21301
rect 18506 21292 18512 21344
rect 18564 21332 18570 21344
rect 18877 21335 18935 21341
rect 18877 21332 18889 21335
rect 18564 21304 18889 21332
rect 18564 21292 18570 21304
rect 18877 21301 18889 21304
rect 18923 21301 18935 21335
rect 18877 21295 18935 21301
rect 19610 21292 19616 21344
rect 19668 21332 19674 21344
rect 20714 21332 20720 21344
rect 19668 21304 20720 21332
rect 19668 21292 19674 21304
rect 20714 21292 20720 21304
rect 20772 21292 20778 21344
rect 22830 21292 22836 21344
rect 22888 21332 22894 21344
rect 24688 21332 24716 21431
rect 25038 21428 25044 21440
rect 25096 21428 25102 21480
rect 22888 21304 24716 21332
rect 22888 21292 22894 21304
rect 1104 21242 25852 21264
rect 1104 21190 2950 21242
rect 3002 21190 3014 21242
rect 3066 21190 3078 21242
rect 3130 21190 3142 21242
rect 3194 21190 3206 21242
rect 3258 21190 12950 21242
rect 13002 21190 13014 21242
rect 13066 21190 13078 21242
rect 13130 21190 13142 21242
rect 13194 21190 13206 21242
rect 13258 21190 22950 21242
rect 23002 21190 23014 21242
rect 23066 21190 23078 21242
rect 23130 21190 23142 21242
rect 23194 21190 23206 21242
rect 23258 21190 25852 21242
rect 1104 21168 25852 21190
rect 2866 21088 2872 21140
rect 2924 21088 2930 21140
rect 7282 21088 7288 21140
rect 7340 21128 7346 21140
rect 7653 21131 7711 21137
rect 7653 21128 7665 21131
rect 7340 21100 7665 21128
rect 7340 21088 7346 21100
rect 7653 21097 7665 21100
rect 7699 21097 7711 21131
rect 7653 21091 7711 21097
rect 8110 21088 8116 21140
rect 8168 21128 8174 21140
rect 10321 21131 10379 21137
rect 10321 21128 10333 21131
rect 8168 21100 10333 21128
rect 8168 21088 8174 21100
rect 10321 21097 10333 21100
rect 10367 21097 10379 21131
rect 10321 21091 10379 21097
rect 11425 21131 11483 21137
rect 11425 21097 11437 21131
rect 11471 21128 11483 21131
rect 12342 21128 12348 21140
rect 11471 21100 12348 21128
rect 11471 21097 11483 21100
rect 11425 21091 11483 21097
rect 12342 21088 12348 21100
rect 12400 21088 12406 21140
rect 12618 21088 12624 21140
rect 12676 21088 12682 21140
rect 12710 21088 12716 21140
rect 12768 21128 12774 21140
rect 13998 21128 14004 21140
rect 12768 21100 14004 21128
rect 12768 21088 12774 21100
rect 13998 21088 14004 21100
rect 14056 21088 14062 21140
rect 16206 21088 16212 21140
rect 16264 21128 16270 21140
rect 16301 21131 16359 21137
rect 16301 21128 16313 21131
rect 16264 21100 16313 21128
rect 16264 21088 16270 21100
rect 16301 21097 16313 21100
rect 16347 21097 16359 21131
rect 16301 21091 16359 21097
rect 19613 21131 19671 21137
rect 19613 21097 19625 21131
rect 19659 21128 19671 21131
rect 24302 21128 24308 21140
rect 19659 21100 24308 21128
rect 19659 21097 19671 21100
rect 19613 21091 19671 21097
rect 24302 21088 24308 21100
rect 24360 21088 24366 21140
rect 7006 21020 7012 21072
rect 7064 21060 7070 21072
rect 7064 21032 8248 21060
rect 7064 21020 7070 21032
rect 3418 20952 3424 21004
rect 3476 20952 3482 21004
rect 5258 20952 5264 21004
rect 5316 20952 5322 21004
rect 5810 20952 5816 21004
rect 5868 20992 5874 21004
rect 6270 20992 6276 21004
rect 5868 20964 6276 20992
rect 5868 20952 5874 20964
rect 6270 20952 6276 20964
rect 6328 20992 6334 21004
rect 8220 21001 8248 21032
rect 11698 21020 11704 21072
rect 11756 21060 11762 21072
rect 11756 21032 12020 21060
rect 11756 21020 11762 21032
rect 8205 20995 8263 21001
rect 6328 20964 8156 20992
rect 6328 20952 6334 20964
rect 3237 20927 3295 20933
rect 3237 20893 3249 20927
rect 3283 20924 3295 20927
rect 3878 20924 3884 20936
rect 3283 20896 3884 20924
rect 3283 20893 3295 20896
rect 3237 20887 3295 20893
rect 3878 20884 3884 20896
rect 3936 20924 3942 20936
rect 4062 20924 4068 20936
rect 3936 20896 4068 20924
rect 3936 20884 3942 20896
rect 4062 20884 4068 20896
rect 4120 20884 4126 20936
rect 4982 20884 4988 20936
rect 5040 20884 5046 20936
rect 6362 20884 6368 20936
rect 6420 20924 6426 20936
rect 7009 20927 7067 20933
rect 7009 20924 7021 20927
rect 6420 20896 7021 20924
rect 6420 20884 6426 20896
rect 7009 20893 7021 20896
rect 7055 20924 7067 20927
rect 7098 20924 7104 20936
rect 7055 20896 7104 20924
rect 7055 20893 7067 20896
rect 7009 20887 7067 20893
rect 7098 20884 7104 20896
rect 7156 20884 7162 20936
rect 8128 20924 8156 20964
rect 8205 20961 8217 20995
rect 8251 20992 8263 20995
rect 10318 20992 10324 21004
rect 8251 20964 10324 20992
rect 8251 20961 8263 20964
rect 8205 20955 8263 20961
rect 10318 20952 10324 20964
rect 10376 20952 10382 21004
rect 10778 20952 10784 21004
rect 10836 20952 10842 21004
rect 11992 21001 12020 21032
rect 22186 21020 22192 21072
rect 22244 21060 22250 21072
rect 22281 21063 22339 21069
rect 22281 21060 22293 21063
rect 22244 21032 22293 21060
rect 22244 21020 22250 21032
rect 22281 21029 22293 21032
rect 22327 21029 22339 21063
rect 22281 21023 22339 21029
rect 23477 21063 23535 21069
rect 23477 21029 23489 21063
rect 23523 21060 23535 21063
rect 24854 21060 24860 21072
rect 23523 21032 24860 21060
rect 23523 21029 23535 21032
rect 23477 21023 23535 21029
rect 10873 20995 10931 21001
rect 10873 20961 10885 20995
rect 10919 20961 10931 20995
rect 10873 20955 10931 20961
rect 11977 20995 12035 21001
rect 11977 20961 11989 20995
rect 12023 20961 12035 20995
rect 11977 20955 12035 20961
rect 10336 20924 10364 20952
rect 10888 20924 10916 20955
rect 13354 20952 13360 21004
rect 13412 20992 13418 21004
rect 14277 20995 14335 21001
rect 14277 20992 14289 20995
rect 13412 20964 14289 20992
rect 13412 20952 13418 20964
rect 14277 20961 14289 20964
rect 14323 20961 14335 20995
rect 14277 20955 14335 20961
rect 14550 20952 14556 21004
rect 14608 20952 14614 21004
rect 18598 20952 18604 21004
rect 18656 20952 18662 21004
rect 18785 20995 18843 21001
rect 18785 20961 18797 20995
rect 18831 20992 18843 20995
rect 19610 20992 19616 21004
rect 18831 20964 19616 20992
rect 18831 20961 18843 20964
rect 18785 20955 18843 20961
rect 19610 20952 19616 20964
rect 19668 20952 19674 21004
rect 20533 20995 20591 21001
rect 20533 20961 20545 20995
rect 20579 20992 20591 20995
rect 22094 20992 22100 21004
rect 20579 20964 22100 20992
rect 20579 20961 20591 20964
rect 20533 20955 20591 20961
rect 22094 20952 22100 20964
rect 22152 20952 22158 21004
rect 8128 20896 9674 20924
rect 10336 20896 10916 20924
rect 7742 20816 7748 20868
rect 7800 20856 7806 20868
rect 8113 20859 8171 20865
rect 8113 20856 8125 20859
rect 7800 20828 8125 20856
rect 7800 20816 7806 20828
rect 8113 20825 8125 20828
rect 8159 20825 8171 20859
rect 9646 20856 9674 20896
rect 13538 20884 13544 20936
rect 13596 20884 13602 20936
rect 18506 20884 18512 20936
rect 18564 20884 18570 20936
rect 19429 20927 19487 20933
rect 19429 20893 19441 20927
rect 19475 20893 19487 20927
rect 19429 20887 19487 20893
rect 10689 20859 10747 20865
rect 9646 20828 10640 20856
rect 8113 20819 8171 20825
rect 4338 20748 4344 20800
rect 4396 20748 4402 20800
rect 6733 20791 6791 20797
rect 6733 20757 6745 20791
rect 6779 20788 6791 20791
rect 6914 20788 6920 20800
rect 6779 20760 6920 20788
rect 6779 20757 6791 20760
rect 6733 20751 6791 20757
rect 6914 20748 6920 20760
rect 6972 20748 6978 20800
rect 7282 20748 7288 20800
rect 7340 20788 7346 20800
rect 8021 20791 8079 20797
rect 8021 20788 8033 20791
rect 7340 20760 8033 20788
rect 7340 20748 7346 20760
rect 8021 20757 8033 20760
rect 8067 20788 8079 20791
rect 8294 20788 8300 20800
rect 8067 20760 8300 20788
rect 8067 20757 8079 20760
rect 8021 20751 8079 20757
rect 8294 20748 8300 20760
rect 8352 20748 8358 20800
rect 8938 20748 8944 20800
rect 8996 20788 9002 20800
rect 9950 20788 9956 20800
rect 8996 20760 9956 20788
rect 8996 20748 9002 20760
rect 9950 20748 9956 20760
rect 10008 20748 10014 20800
rect 10612 20788 10640 20828
rect 10689 20825 10701 20859
rect 10735 20856 10747 20859
rect 11606 20856 11612 20868
rect 10735 20828 11612 20856
rect 10735 20825 10747 20828
rect 10689 20819 10747 20825
rect 11606 20816 11612 20828
rect 11664 20816 11670 20868
rect 12066 20856 12072 20868
rect 11992 20828 12072 20856
rect 11517 20791 11575 20797
rect 11517 20788 11529 20791
rect 10612 20760 11529 20788
rect 11517 20757 11529 20760
rect 11563 20788 11575 20791
rect 11992 20788 12020 20828
rect 12066 20816 12072 20828
rect 12124 20856 12130 20868
rect 12161 20859 12219 20865
rect 12161 20856 12173 20859
rect 12124 20828 12173 20856
rect 12124 20816 12130 20828
rect 12161 20825 12173 20828
rect 12207 20825 12219 20859
rect 16206 20856 16212 20868
rect 15778 20828 16212 20856
rect 12161 20819 12219 20825
rect 16206 20816 16212 20828
rect 16264 20816 16270 20868
rect 17218 20816 17224 20868
rect 17276 20856 17282 20868
rect 19444 20856 19472 20887
rect 21818 20884 21824 20936
rect 21876 20924 21882 20936
rect 23492 20924 23520 21023
rect 24854 21020 24860 21032
rect 24912 21020 24918 21072
rect 21876 20896 23520 20924
rect 21876 20884 21882 20896
rect 17276 20828 19472 20856
rect 17276 20816 17282 20828
rect 20714 20816 20720 20868
rect 20772 20856 20778 20868
rect 20809 20859 20867 20865
rect 20809 20856 20821 20859
rect 20772 20828 20821 20856
rect 20772 20816 20778 20828
rect 20809 20825 20821 20828
rect 20855 20825 20867 20859
rect 20809 20819 20867 20825
rect 21266 20816 21272 20868
rect 21324 20816 21330 20868
rect 22925 20859 22983 20865
rect 22925 20825 22937 20859
rect 22971 20825 22983 20859
rect 22925 20819 22983 20825
rect 23109 20859 23167 20865
rect 23109 20825 23121 20859
rect 23155 20856 23167 20859
rect 23750 20856 23756 20868
rect 23155 20828 23756 20856
rect 23155 20825 23167 20828
rect 23109 20819 23167 20825
rect 11563 20760 12020 20788
rect 12253 20791 12311 20797
rect 11563 20757 11575 20760
rect 11517 20751 11575 20757
rect 12253 20757 12265 20791
rect 12299 20788 12311 20791
rect 12342 20788 12348 20800
rect 12299 20760 12348 20788
rect 12299 20757 12311 20760
rect 12253 20751 12311 20757
rect 12342 20748 12348 20760
rect 12400 20748 12406 20800
rect 16022 20748 16028 20800
rect 16080 20748 16086 20800
rect 16850 20748 16856 20800
rect 16908 20748 16914 20800
rect 17126 20748 17132 20800
rect 17184 20788 17190 20800
rect 18141 20791 18199 20797
rect 18141 20788 18153 20791
rect 17184 20760 18153 20788
rect 17184 20748 17190 20760
rect 18141 20757 18153 20760
rect 18187 20757 18199 20791
rect 18141 20751 18199 20757
rect 20898 20748 20904 20800
rect 20956 20788 20962 20800
rect 22940 20788 22968 20819
rect 23750 20816 23756 20828
rect 23808 20816 23814 20868
rect 20956 20760 22968 20788
rect 20956 20748 20962 20760
rect 1104 20698 25852 20720
rect 1104 20646 7950 20698
rect 8002 20646 8014 20698
rect 8066 20646 8078 20698
rect 8130 20646 8142 20698
rect 8194 20646 8206 20698
rect 8258 20646 17950 20698
rect 18002 20646 18014 20698
rect 18066 20646 18078 20698
rect 18130 20646 18142 20698
rect 18194 20646 18206 20698
rect 18258 20646 25852 20698
rect 1104 20624 25852 20646
rect 4982 20584 4988 20596
rect 3896 20556 4988 20584
rect 1762 20408 1768 20460
rect 1820 20408 1826 20460
rect 3896 20457 3924 20556
rect 4982 20544 4988 20556
rect 5040 20584 5046 20596
rect 5442 20584 5448 20596
rect 5040 20556 5448 20584
rect 5040 20544 5046 20556
rect 5442 20544 5448 20556
rect 5500 20584 5506 20596
rect 5500 20556 8616 20584
rect 5500 20544 5506 20556
rect 4157 20519 4215 20525
rect 4157 20485 4169 20519
rect 4203 20516 4215 20519
rect 4246 20516 4252 20528
rect 4203 20488 4252 20516
rect 4203 20485 4215 20488
rect 4157 20479 4215 20485
rect 4246 20476 4252 20488
rect 4304 20476 4310 20528
rect 3881 20451 3939 20457
rect 3881 20417 3893 20451
rect 3927 20417 3939 20451
rect 5290 20420 6040 20448
rect 3881 20411 3939 20417
rect 1302 20340 1308 20392
rect 1360 20380 1366 20392
rect 2041 20383 2099 20389
rect 2041 20380 2053 20383
rect 1360 20352 2053 20380
rect 1360 20340 1366 20352
rect 2041 20349 2053 20352
rect 2087 20349 2099 20383
rect 2041 20343 2099 20349
rect 5629 20247 5687 20253
rect 5629 20213 5641 20247
rect 5675 20244 5687 20247
rect 5718 20244 5724 20256
rect 5675 20216 5724 20244
rect 5675 20213 5687 20216
rect 5629 20207 5687 20213
rect 5718 20204 5724 20216
rect 5776 20204 5782 20256
rect 6012 20253 6040 20420
rect 7006 20408 7012 20460
rect 7064 20448 7070 20460
rect 7190 20448 7196 20460
rect 7064 20420 7196 20448
rect 7064 20408 7070 20420
rect 7190 20408 7196 20420
rect 7248 20448 7254 20460
rect 8588 20457 8616 20556
rect 10318 20544 10324 20596
rect 10376 20544 10382 20596
rect 12069 20587 12127 20593
rect 12069 20553 12081 20587
rect 12115 20584 12127 20587
rect 12434 20584 12440 20596
rect 12115 20556 12440 20584
rect 12115 20553 12127 20556
rect 12069 20547 12127 20553
rect 12434 20544 12440 20556
rect 12492 20544 12498 20596
rect 14734 20544 14740 20596
rect 14792 20544 14798 20596
rect 14829 20587 14887 20593
rect 14829 20553 14841 20587
rect 14875 20584 14887 20587
rect 15102 20584 15108 20596
rect 14875 20556 15108 20584
rect 14875 20553 14887 20556
rect 14829 20547 14887 20553
rect 15102 20544 15108 20556
rect 15160 20544 15166 20596
rect 16390 20544 16396 20596
rect 16448 20544 16454 20596
rect 16850 20544 16856 20596
rect 16908 20584 16914 20596
rect 17221 20587 17279 20593
rect 17221 20584 17233 20587
rect 16908 20556 17233 20584
rect 16908 20544 16914 20556
rect 17221 20553 17233 20556
rect 17267 20553 17279 20587
rect 20717 20587 20775 20593
rect 20717 20584 20729 20587
rect 17221 20547 17279 20553
rect 19352 20556 20729 20584
rect 9858 20476 9864 20528
rect 9916 20476 9922 20528
rect 11974 20476 11980 20528
rect 12032 20516 12038 20528
rect 13446 20516 13452 20528
rect 12032 20488 13452 20516
rect 12032 20476 12038 20488
rect 13446 20476 13452 20488
rect 13504 20476 13510 20528
rect 16408 20516 16436 20544
rect 17129 20519 17187 20525
rect 17129 20516 17141 20519
rect 16408 20488 17141 20516
rect 17129 20485 17141 20488
rect 17175 20485 17187 20519
rect 18874 20516 18880 20528
rect 17129 20479 17187 20485
rect 18340 20488 18880 20516
rect 7745 20451 7803 20457
rect 7745 20448 7757 20451
rect 7248 20420 7757 20448
rect 7248 20408 7254 20420
rect 7745 20417 7757 20420
rect 7791 20417 7803 20451
rect 7745 20411 7803 20417
rect 8573 20451 8631 20457
rect 8573 20417 8585 20451
rect 8619 20417 8631 20451
rect 8573 20411 8631 20417
rect 12161 20451 12219 20457
rect 12161 20417 12173 20451
rect 12207 20448 12219 20451
rect 13630 20448 13636 20460
rect 12207 20420 13636 20448
rect 12207 20417 12219 20420
rect 12161 20411 12219 20417
rect 13630 20408 13636 20420
rect 13688 20408 13694 20460
rect 15749 20451 15807 20457
rect 15749 20417 15761 20451
rect 15795 20448 15807 20451
rect 16758 20448 16764 20460
rect 15795 20420 16764 20448
rect 15795 20417 15807 20420
rect 15749 20411 15807 20417
rect 16758 20408 16764 20420
rect 16816 20408 16822 20460
rect 7561 20383 7619 20389
rect 7561 20349 7573 20383
rect 7607 20349 7619 20383
rect 7561 20343 7619 20349
rect 7653 20383 7711 20389
rect 7653 20349 7665 20383
rect 7699 20380 7711 20383
rect 8294 20380 8300 20392
rect 7699 20352 8300 20380
rect 7699 20349 7711 20352
rect 7653 20343 7711 20349
rect 7576 20312 7604 20343
rect 8294 20340 8300 20352
rect 8352 20340 8358 20392
rect 8849 20383 8907 20389
rect 8849 20349 8861 20383
rect 8895 20380 8907 20383
rect 9858 20380 9864 20392
rect 8895 20352 9864 20380
rect 8895 20349 8907 20352
rect 8849 20343 8907 20349
rect 9858 20340 9864 20352
rect 9916 20380 9922 20392
rect 10962 20380 10968 20392
rect 9916 20352 10968 20380
rect 9916 20340 9922 20352
rect 10962 20340 10968 20352
rect 11020 20340 11026 20392
rect 11149 20383 11207 20389
rect 11149 20349 11161 20383
rect 11195 20380 11207 20383
rect 11698 20380 11704 20392
rect 11195 20352 11704 20380
rect 11195 20349 11207 20352
rect 11149 20343 11207 20349
rect 11698 20340 11704 20352
rect 11756 20340 11762 20392
rect 12253 20383 12311 20389
rect 12253 20349 12265 20383
rect 12299 20349 12311 20383
rect 12253 20343 12311 20349
rect 15013 20383 15071 20389
rect 15013 20349 15025 20383
rect 15059 20380 15071 20383
rect 16022 20380 16028 20392
rect 15059 20352 16028 20380
rect 15059 20349 15071 20352
rect 15013 20343 15071 20349
rect 7576 20284 7696 20312
rect 5997 20247 6055 20253
rect 5997 20213 6009 20247
rect 6043 20244 6055 20247
rect 6362 20244 6368 20256
rect 6043 20216 6368 20244
rect 6043 20213 6055 20216
rect 5997 20207 6055 20213
rect 6362 20204 6368 20216
rect 6420 20204 6426 20256
rect 7006 20204 7012 20256
rect 7064 20204 7070 20256
rect 7098 20204 7104 20256
rect 7156 20244 7162 20256
rect 7668 20244 7696 20284
rect 7834 20272 7840 20324
rect 7892 20312 7898 20324
rect 8113 20315 8171 20321
rect 8113 20312 8125 20315
rect 7892 20284 8125 20312
rect 7892 20272 7898 20284
rect 8113 20281 8125 20284
rect 8159 20281 8171 20315
rect 8113 20275 8171 20281
rect 10134 20272 10140 20324
rect 10192 20312 10198 20324
rect 10686 20312 10692 20324
rect 10192 20284 10692 20312
rect 10192 20272 10198 20284
rect 10686 20272 10692 20284
rect 10744 20312 10750 20324
rect 12268 20312 12296 20343
rect 16022 20340 16028 20352
rect 16080 20340 16086 20392
rect 17037 20383 17095 20389
rect 17037 20349 17049 20383
rect 17083 20380 17095 20383
rect 18340 20380 18368 20488
rect 18874 20476 18880 20488
rect 18932 20516 18938 20528
rect 18969 20519 19027 20525
rect 18969 20516 18981 20519
rect 18932 20488 18981 20516
rect 18932 20476 18938 20488
rect 18969 20485 18981 20488
rect 19015 20485 19027 20519
rect 19352 20516 19380 20556
rect 20717 20553 20729 20556
rect 20763 20584 20775 20587
rect 21266 20584 21272 20596
rect 20763 20556 21272 20584
rect 20763 20553 20775 20556
rect 20717 20547 20775 20553
rect 21266 20544 21272 20556
rect 21324 20584 21330 20596
rect 21818 20584 21824 20596
rect 21324 20556 21824 20584
rect 21324 20544 21330 20556
rect 21818 20544 21824 20556
rect 21876 20544 21882 20596
rect 22370 20544 22376 20596
rect 22428 20544 22434 20596
rect 22465 20587 22523 20593
rect 22465 20553 22477 20587
rect 22511 20584 22523 20587
rect 22738 20584 22744 20596
rect 22511 20556 22744 20584
rect 22511 20553 22523 20556
rect 22465 20547 22523 20553
rect 22738 20544 22744 20556
rect 22796 20544 22802 20596
rect 23293 20587 23351 20593
rect 23293 20553 23305 20587
rect 23339 20584 23351 20587
rect 24394 20584 24400 20596
rect 23339 20556 24400 20584
rect 23339 20553 23351 20556
rect 23293 20547 23351 20553
rect 19426 20516 19432 20528
rect 19352 20488 19432 20516
rect 18969 20479 19027 20485
rect 19426 20476 19432 20488
rect 19484 20476 19490 20528
rect 18690 20408 18696 20460
rect 18748 20408 18754 20460
rect 17083 20352 18368 20380
rect 20441 20383 20499 20389
rect 17083 20349 17095 20352
rect 17037 20343 17095 20349
rect 20441 20349 20453 20383
rect 20487 20380 20499 20383
rect 20714 20380 20720 20392
rect 20487 20352 20720 20380
rect 20487 20349 20499 20352
rect 20441 20343 20499 20349
rect 20714 20340 20720 20352
rect 20772 20340 20778 20392
rect 22649 20383 22707 20389
rect 22649 20349 22661 20383
rect 22695 20380 22707 20383
rect 23308 20380 23336 20547
rect 24394 20544 24400 20556
rect 24452 20544 24458 20596
rect 24854 20544 24860 20596
rect 24912 20584 24918 20596
rect 25317 20587 25375 20593
rect 25317 20584 25329 20587
rect 24912 20556 25329 20584
rect 24912 20544 24918 20556
rect 25317 20553 25329 20556
rect 25363 20553 25375 20587
rect 25317 20547 25375 20553
rect 24872 20516 24900 20544
rect 24334 20488 24900 20516
rect 25038 20408 25044 20460
rect 25096 20408 25102 20460
rect 22695 20352 23336 20380
rect 22695 20349 22707 20352
rect 22649 20343 22707 20349
rect 24210 20340 24216 20392
rect 24268 20380 24274 20392
rect 24765 20383 24823 20389
rect 24765 20380 24777 20383
rect 24268 20352 24777 20380
rect 24268 20340 24274 20352
rect 24765 20349 24777 20352
rect 24811 20349 24823 20383
rect 24765 20343 24823 20349
rect 10744 20284 12296 20312
rect 10744 20272 10750 20284
rect 20622 20272 20628 20324
rect 20680 20312 20686 20324
rect 22005 20315 22063 20321
rect 22005 20312 22017 20315
rect 20680 20284 22017 20312
rect 20680 20272 20686 20284
rect 22005 20281 22017 20284
rect 22051 20281 22063 20315
rect 22005 20275 22063 20281
rect 10152 20244 10180 20272
rect 7156 20216 10180 20244
rect 7156 20204 7162 20216
rect 10410 20204 10416 20256
rect 10468 20244 10474 20256
rect 11701 20247 11759 20253
rect 11701 20244 11713 20247
rect 10468 20216 11713 20244
rect 10468 20204 10474 20216
rect 11701 20213 11713 20216
rect 11747 20213 11759 20247
rect 11701 20207 11759 20213
rect 14366 20204 14372 20256
rect 14424 20204 14430 20256
rect 15565 20247 15623 20253
rect 15565 20213 15577 20247
rect 15611 20244 15623 20247
rect 15654 20244 15660 20256
rect 15611 20216 15660 20244
rect 15611 20213 15623 20216
rect 15565 20207 15623 20213
rect 15654 20204 15660 20216
rect 15712 20204 15718 20256
rect 17589 20247 17647 20253
rect 17589 20213 17601 20247
rect 17635 20244 17647 20247
rect 18230 20244 18236 20256
rect 17635 20216 18236 20244
rect 17635 20213 17647 20216
rect 17589 20207 17647 20213
rect 18230 20204 18236 20216
rect 18288 20204 18294 20256
rect 1104 20154 25852 20176
rect 1104 20102 2950 20154
rect 3002 20102 3014 20154
rect 3066 20102 3078 20154
rect 3130 20102 3142 20154
rect 3194 20102 3206 20154
rect 3258 20102 12950 20154
rect 13002 20102 13014 20154
rect 13066 20102 13078 20154
rect 13130 20102 13142 20154
rect 13194 20102 13206 20154
rect 13258 20102 22950 20154
rect 23002 20102 23014 20154
rect 23066 20102 23078 20154
rect 23130 20102 23142 20154
rect 23194 20102 23206 20154
rect 23258 20102 25852 20154
rect 1104 20080 25852 20102
rect 5350 20000 5356 20052
rect 5408 20040 5414 20052
rect 5445 20043 5503 20049
rect 5445 20040 5457 20043
rect 5408 20012 5457 20040
rect 5408 20000 5414 20012
rect 5445 20009 5457 20012
rect 5491 20009 5503 20043
rect 5445 20003 5503 20009
rect 6935 20043 6993 20049
rect 6935 20009 6947 20043
rect 6981 20040 6993 20043
rect 7098 20040 7104 20052
rect 6981 20012 7104 20040
rect 6981 20009 6993 20012
rect 6935 20003 6993 20009
rect 7098 20000 7104 20012
rect 7156 20000 7162 20052
rect 8386 20000 8392 20052
rect 8444 20040 8450 20052
rect 8444 20012 8524 20040
rect 8444 20000 8450 20012
rect 6822 19864 6828 19916
rect 6880 19904 6886 19916
rect 7193 19907 7251 19913
rect 7193 19904 7205 19907
rect 6880 19876 7205 19904
rect 6880 19864 6886 19876
rect 7193 19873 7205 19876
rect 7239 19873 7251 19907
rect 7193 19867 7251 19873
rect 7374 19864 7380 19916
rect 7432 19904 7438 19916
rect 8389 19907 8447 19913
rect 8389 19904 8401 19907
rect 7432 19876 8401 19904
rect 7432 19864 7438 19876
rect 8389 19873 8401 19876
rect 8435 19873 8447 19907
rect 8496 19904 8524 20012
rect 9122 20000 9128 20052
rect 9180 20000 9186 20052
rect 9950 20000 9956 20052
rect 10008 20040 10014 20052
rect 10505 20043 10563 20049
rect 10505 20040 10517 20043
rect 10008 20012 10517 20040
rect 10008 20000 10014 20012
rect 10505 20009 10517 20012
rect 10551 20009 10563 20043
rect 12437 20043 12495 20049
rect 12437 20040 12449 20043
rect 10505 20003 10563 20009
rect 11808 20012 12449 20040
rect 11808 19913 11836 20012
rect 12437 20009 12449 20012
rect 12483 20040 12495 20043
rect 12526 20040 12532 20052
rect 12483 20012 12532 20040
rect 12483 20009 12495 20012
rect 12437 20003 12495 20009
rect 12526 20000 12532 20012
rect 12584 20000 12590 20052
rect 24210 20000 24216 20052
rect 24268 20040 24274 20052
rect 24854 20040 24860 20052
rect 24268 20012 24860 20040
rect 24268 20000 24274 20012
rect 24854 20000 24860 20012
rect 24912 20000 24918 20052
rect 16117 19975 16175 19981
rect 16117 19941 16129 19975
rect 16163 19972 16175 19975
rect 19794 19972 19800 19984
rect 16163 19944 19800 19972
rect 16163 19941 16175 19944
rect 16117 19935 16175 19941
rect 19794 19932 19800 19944
rect 19852 19932 19858 19984
rect 9677 19907 9735 19913
rect 9677 19904 9689 19907
rect 8496 19876 9689 19904
rect 8389 19867 8447 19873
rect 9677 19873 9689 19876
rect 9723 19873 9735 19907
rect 9677 19867 9735 19873
rect 11793 19907 11851 19913
rect 11793 19873 11805 19907
rect 11839 19873 11851 19907
rect 11793 19867 11851 19873
rect 11974 19864 11980 19916
rect 12032 19864 12038 19916
rect 18322 19864 18328 19916
rect 18380 19864 18386 19916
rect 18509 19907 18567 19913
rect 18509 19873 18521 19907
rect 18555 19904 18567 19907
rect 20714 19904 20720 19916
rect 18555 19876 20720 19904
rect 18555 19873 18567 19876
rect 18509 19867 18567 19873
rect 20714 19864 20720 19876
rect 20772 19864 20778 19916
rect 23385 19907 23443 19913
rect 23385 19873 23397 19907
rect 23431 19904 23443 19907
rect 25130 19904 25136 19916
rect 23431 19876 25136 19904
rect 23431 19873 23443 19876
rect 23385 19867 23443 19873
rect 25130 19864 25136 19876
rect 25188 19864 25194 19916
rect 2225 19839 2283 19845
rect 2225 19805 2237 19839
rect 2271 19836 2283 19839
rect 3326 19836 3332 19848
rect 2271 19808 3332 19836
rect 2271 19805 2283 19808
rect 2225 19799 2283 19805
rect 3326 19796 3332 19808
rect 3384 19796 3390 19848
rect 8297 19839 8355 19845
rect 8297 19805 8309 19839
rect 8343 19836 8355 19839
rect 8478 19836 8484 19848
rect 8343 19808 8484 19836
rect 8343 19805 8355 19808
rect 8297 19799 8355 19805
rect 8478 19796 8484 19808
rect 8536 19796 8542 19848
rect 9493 19839 9551 19845
rect 9493 19805 9505 19839
rect 9539 19836 9551 19839
rect 10410 19836 10416 19848
rect 9539 19808 10416 19836
rect 9539 19805 9551 19808
rect 9493 19799 9551 19805
rect 10410 19796 10416 19808
rect 10468 19796 10474 19848
rect 11698 19796 11704 19848
rect 11756 19796 11762 19848
rect 14182 19796 14188 19848
rect 14240 19836 14246 19848
rect 15933 19839 15991 19845
rect 15933 19836 15945 19839
rect 14240 19808 15945 19836
rect 14240 19796 14246 19808
rect 15933 19805 15945 19808
rect 15979 19805 15991 19839
rect 15933 19799 15991 19805
rect 16853 19839 16911 19845
rect 16853 19805 16865 19839
rect 16899 19836 16911 19839
rect 17218 19836 17224 19848
rect 16899 19808 17224 19836
rect 16899 19805 16911 19808
rect 16853 19799 16911 19805
rect 17218 19796 17224 19808
rect 17276 19796 17282 19848
rect 18230 19796 18236 19848
rect 18288 19796 18294 19848
rect 19613 19839 19671 19845
rect 19613 19805 19625 19839
rect 19659 19836 19671 19839
rect 20990 19836 20996 19848
rect 19659 19808 20996 19836
rect 19659 19805 19671 19808
rect 19613 19799 19671 19805
rect 20990 19796 20996 19808
rect 21048 19796 21054 19848
rect 21082 19796 21088 19848
rect 21140 19836 21146 19848
rect 21269 19839 21327 19845
rect 21269 19836 21281 19839
rect 21140 19808 21281 19836
rect 21140 19796 21146 19808
rect 21269 19805 21281 19808
rect 21315 19805 21327 19839
rect 21269 19799 21327 19805
rect 24029 19839 24087 19845
rect 24029 19805 24041 19839
rect 24075 19836 24087 19839
rect 24762 19836 24768 19848
rect 24075 19808 24768 19836
rect 24075 19805 24087 19808
rect 24029 19799 24087 19805
rect 24762 19796 24768 19808
rect 24820 19796 24826 19848
rect 6362 19728 6368 19780
rect 6420 19728 6426 19780
rect 7650 19768 7656 19780
rect 7484 19740 7656 19768
rect 7484 19712 7512 19740
rect 7650 19728 7656 19740
rect 7708 19768 7714 19780
rect 8205 19771 8263 19777
rect 8205 19768 8217 19771
rect 7708 19740 8217 19768
rect 7708 19728 7714 19740
rect 8205 19737 8217 19740
rect 8251 19737 8263 19771
rect 8205 19731 8263 19737
rect 10778 19728 10784 19780
rect 10836 19768 10842 19780
rect 13078 19768 13084 19780
rect 10836 19740 13084 19768
rect 10836 19728 10842 19740
rect 13078 19728 13084 19740
rect 13136 19728 13142 19780
rect 20438 19728 20444 19780
rect 20496 19768 20502 19780
rect 22005 19771 22063 19777
rect 22005 19768 22017 19771
rect 20496 19740 22017 19768
rect 20496 19728 20502 19740
rect 22005 19737 22017 19740
rect 22051 19737 22063 19771
rect 22005 19731 22063 19737
rect 22189 19771 22247 19777
rect 22189 19737 22201 19771
rect 22235 19768 22247 19771
rect 22646 19768 22652 19780
rect 22235 19740 22652 19768
rect 22235 19737 22247 19740
rect 22189 19731 22247 19737
rect 22646 19728 22652 19740
rect 22704 19728 22710 19780
rect 1854 19660 1860 19712
rect 1912 19700 1918 19712
rect 2041 19703 2099 19709
rect 2041 19700 2053 19703
rect 1912 19672 2053 19700
rect 1912 19660 1918 19672
rect 2041 19669 2053 19672
rect 2087 19669 2099 19703
rect 2041 19663 2099 19669
rect 6178 19660 6184 19712
rect 6236 19700 6242 19712
rect 6730 19700 6736 19712
rect 6236 19672 6736 19700
rect 6236 19660 6242 19672
rect 6730 19660 6736 19672
rect 6788 19660 6794 19712
rect 7466 19660 7472 19712
rect 7524 19660 7530 19712
rect 7834 19660 7840 19712
rect 7892 19660 7898 19712
rect 9582 19660 9588 19712
rect 9640 19660 9646 19712
rect 10594 19660 10600 19712
rect 10652 19700 10658 19712
rect 11333 19703 11391 19709
rect 11333 19700 11345 19703
rect 10652 19672 11345 19700
rect 10652 19660 10658 19672
rect 11333 19669 11345 19672
rect 11379 19669 11391 19703
rect 11333 19663 11391 19669
rect 17034 19660 17040 19712
rect 17092 19700 17098 19712
rect 17313 19703 17371 19709
rect 17313 19700 17325 19703
rect 17092 19672 17325 19700
rect 17092 19660 17098 19672
rect 17313 19669 17325 19672
rect 17359 19669 17371 19703
rect 17313 19663 17371 19669
rect 17494 19660 17500 19712
rect 17552 19700 17558 19712
rect 17865 19703 17923 19709
rect 17865 19700 17877 19703
rect 17552 19672 17877 19700
rect 17552 19660 17558 19672
rect 17865 19669 17877 19672
rect 17911 19669 17923 19703
rect 17865 19663 17923 19669
rect 19429 19703 19487 19709
rect 19429 19669 19441 19703
rect 19475 19700 19487 19703
rect 19886 19700 19892 19712
rect 19475 19672 19892 19700
rect 19475 19669 19487 19672
rect 19429 19663 19487 19669
rect 19886 19660 19892 19672
rect 19944 19660 19950 19712
rect 21361 19703 21419 19709
rect 21361 19669 21373 19703
rect 21407 19700 21419 19703
rect 21726 19700 21732 19712
rect 21407 19672 21732 19700
rect 21407 19669 21419 19672
rect 21361 19663 21419 19669
rect 21726 19660 21732 19672
rect 21784 19660 21790 19712
rect 1104 19610 25852 19632
rect 1104 19558 7950 19610
rect 8002 19558 8014 19610
rect 8066 19558 8078 19610
rect 8130 19558 8142 19610
rect 8194 19558 8206 19610
rect 8258 19558 17950 19610
rect 18002 19558 18014 19610
rect 18066 19558 18078 19610
rect 18130 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 25852 19610
rect 1104 19536 25852 19558
rect 4890 19456 4896 19508
rect 4948 19456 4954 19508
rect 5718 19456 5724 19508
rect 5776 19496 5782 19508
rect 5776 19468 8800 19496
rect 5776 19456 5782 19468
rect 6362 19388 6368 19440
rect 6420 19428 6426 19440
rect 6917 19431 6975 19437
rect 6917 19428 6929 19431
rect 6420 19400 6929 19428
rect 6420 19388 6426 19400
rect 6917 19397 6929 19400
rect 6963 19428 6975 19431
rect 6963 19400 7958 19428
rect 6963 19397 6975 19400
rect 6917 19391 6975 19397
rect 5077 19363 5135 19369
rect 5077 19329 5089 19363
rect 5123 19360 5135 19363
rect 6454 19360 6460 19372
rect 5123 19332 6460 19360
rect 5123 19329 5135 19332
rect 5077 19323 5135 19329
rect 6454 19320 6460 19332
rect 6512 19320 6518 19372
rect 6822 19320 6828 19372
rect 6880 19360 6886 19372
rect 7193 19363 7251 19369
rect 7193 19360 7205 19363
rect 6880 19332 7205 19360
rect 6880 19320 6886 19332
rect 7193 19329 7205 19332
rect 7239 19329 7251 19363
rect 8772 19360 8800 19468
rect 9398 19456 9404 19508
rect 9456 19496 9462 19508
rect 10413 19499 10471 19505
rect 10413 19496 10425 19499
rect 9456 19468 10425 19496
rect 9456 19456 9462 19468
rect 10413 19465 10425 19468
rect 10459 19465 10471 19499
rect 11882 19496 11888 19508
rect 10413 19459 10471 19465
rect 10796 19468 11888 19496
rect 9217 19431 9275 19437
rect 9217 19397 9229 19431
rect 9263 19428 9275 19431
rect 10796 19428 10824 19468
rect 11882 19456 11888 19468
rect 11940 19456 11946 19508
rect 13078 19456 13084 19508
rect 13136 19456 13142 19508
rect 18141 19499 18199 19505
rect 18141 19465 18153 19499
rect 18187 19496 18199 19499
rect 19242 19496 19248 19508
rect 18187 19468 19248 19496
rect 18187 19465 18199 19468
rect 18141 19459 18199 19465
rect 19242 19456 19248 19468
rect 19300 19456 19306 19508
rect 9263 19400 10824 19428
rect 10873 19431 10931 19437
rect 9263 19397 9275 19400
rect 9217 19391 9275 19397
rect 10873 19397 10885 19431
rect 10919 19428 10931 19431
rect 11606 19428 11612 19440
rect 10919 19400 11612 19428
rect 10919 19397 10931 19400
rect 10873 19391 10931 19397
rect 11606 19388 11612 19400
rect 11664 19388 11670 19440
rect 12710 19388 12716 19440
rect 12768 19428 12774 19440
rect 13906 19428 13912 19440
rect 12768 19400 13912 19428
rect 12768 19388 12774 19400
rect 13906 19388 13912 19400
rect 13964 19388 13970 19440
rect 16945 19431 17003 19437
rect 16945 19397 16957 19431
rect 16991 19428 17003 19431
rect 17313 19431 17371 19437
rect 17313 19428 17325 19431
rect 16991 19400 17325 19428
rect 16991 19397 17003 19400
rect 16945 19391 17003 19397
rect 17313 19397 17325 19400
rect 17359 19428 17371 19431
rect 19150 19428 19156 19440
rect 17359 19400 19156 19428
rect 17359 19397 17371 19400
rect 17313 19391 17371 19397
rect 19150 19388 19156 19400
rect 19208 19388 19214 19440
rect 20533 19431 20591 19437
rect 20533 19397 20545 19431
rect 20579 19428 20591 19431
rect 22094 19428 22100 19440
rect 20579 19400 22100 19428
rect 20579 19397 20591 19400
rect 20533 19391 20591 19397
rect 22094 19388 22100 19400
rect 22152 19388 22158 19440
rect 22557 19431 22615 19437
rect 22557 19397 22569 19431
rect 22603 19428 22615 19431
rect 24854 19428 24860 19440
rect 22603 19400 24860 19428
rect 22603 19397 22615 19400
rect 22557 19391 22615 19397
rect 24854 19388 24860 19400
rect 24912 19388 24918 19440
rect 9674 19360 9680 19372
rect 8772 19332 9680 19360
rect 7193 19323 7251 19329
rect 9674 19320 9680 19332
rect 9732 19320 9738 19372
rect 10781 19363 10839 19369
rect 10781 19329 10793 19363
rect 10827 19360 10839 19363
rect 12434 19360 12440 19372
rect 10827 19332 12440 19360
rect 10827 19329 10839 19332
rect 10781 19323 10839 19329
rect 12434 19320 12440 19332
rect 12492 19320 12498 19372
rect 13449 19363 13507 19369
rect 13449 19329 13461 19363
rect 13495 19360 13507 19363
rect 13495 19332 14228 19360
rect 13495 19329 13507 19332
rect 13449 19323 13507 19329
rect 6914 19252 6920 19304
rect 6972 19292 6978 19304
rect 7469 19295 7527 19301
rect 7469 19292 7481 19295
rect 6972 19264 7481 19292
rect 6972 19252 6978 19264
rect 7469 19261 7481 19264
rect 7515 19261 7527 19295
rect 7469 19255 7527 19261
rect 9585 19295 9643 19301
rect 9585 19261 9597 19295
rect 9631 19292 9643 19295
rect 9950 19292 9956 19304
rect 9631 19264 9956 19292
rect 9631 19261 9643 19264
rect 9585 19255 9643 19261
rect 9950 19252 9956 19264
rect 10008 19252 10014 19304
rect 10318 19252 10324 19304
rect 10376 19292 10382 19304
rect 10965 19295 11023 19301
rect 10965 19292 10977 19295
rect 10376 19264 10977 19292
rect 10376 19252 10382 19264
rect 10965 19261 10977 19264
rect 11011 19261 11023 19295
rect 10965 19255 11023 19261
rect 12805 19295 12863 19301
rect 12805 19261 12817 19295
rect 12851 19292 12863 19295
rect 13538 19292 13544 19304
rect 12851 19264 13544 19292
rect 12851 19261 12863 19264
rect 12805 19255 12863 19261
rect 8754 19184 8760 19236
rect 8812 19224 8818 19236
rect 12820 19224 12848 19255
rect 13538 19252 13544 19264
rect 13596 19252 13602 19304
rect 13633 19295 13691 19301
rect 13633 19261 13645 19295
rect 13679 19261 13691 19295
rect 13633 19255 13691 19261
rect 8812 19196 12848 19224
rect 8812 19184 8818 19196
rect 13354 19184 13360 19236
rect 13412 19224 13418 19236
rect 13648 19224 13676 19255
rect 14200 19233 14228 19332
rect 14826 19320 14832 19372
rect 14884 19360 14890 19372
rect 17957 19363 18015 19369
rect 17957 19360 17969 19363
rect 14884 19332 17969 19360
rect 14884 19320 14890 19332
rect 17957 19329 17969 19332
rect 18003 19329 18015 19363
rect 17957 19323 18015 19329
rect 18782 19320 18788 19372
rect 18840 19320 18846 19372
rect 21453 19363 21511 19369
rect 21453 19329 21465 19363
rect 21499 19360 21511 19363
rect 22278 19360 22284 19372
rect 21499 19332 22284 19360
rect 21499 19329 21511 19332
rect 21453 19323 21511 19329
rect 22278 19320 22284 19332
rect 22336 19320 22342 19372
rect 23382 19320 23388 19372
rect 23440 19320 23446 19372
rect 24397 19363 24455 19369
rect 24397 19329 24409 19363
rect 24443 19360 24455 19363
rect 24486 19360 24492 19372
rect 24443 19332 24492 19360
rect 24443 19329 24455 19332
rect 24397 19323 24455 19329
rect 24486 19320 24492 19332
rect 24544 19320 24550 19372
rect 25222 19320 25228 19372
rect 25280 19320 25286 19372
rect 13412 19196 13676 19224
rect 14185 19227 14243 19233
rect 13412 19184 13418 19196
rect 14185 19193 14197 19227
rect 14231 19224 14243 19227
rect 18506 19224 18512 19236
rect 14231 19196 18512 19224
rect 14231 19193 14243 19196
rect 14185 19187 14243 19193
rect 18506 19184 18512 19196
rect 18564 19184 18570 19236
rect 9858 19116 9864 19168
rect 9916 19156 9922 19168
rect 13372 19156 13400 19184
rect 9916 19128 13400 19156
rect 9916 19116 9922 19128
rect 17402 19116 17408 19168
rect 17460 19116 17466 19168
rect 18601 19159 18659 19165
rect 18601 19125 18613 19159
rect 18647 19156 18659 19159
rect 18782 19156 18788 19168
rect 18647 19128 18788 19156
rect 18647 19125 18659 19128
rect 18601 19119 18659 19125
rect 18782 19116 18788 19128
rect 18840 19116 18846 19168
rect 1104 19066 25852 19088
rect 1104 19014 2950 19066
rect 3002 19014 3014 19066
rect 3066 19014 3078 19066
rect 3130 19014 3142 19066
rect 3194 19014 3206 19066
rect 3258 19014 12950 19066
rect 13002 19014 13014 19066
rect 13066 19014 13078 19066
rect 13130 19014 13142 19066
rect 13194 19014 13206 19066
rect 13258 19014 22950 19066
rect 23002 19014 23014 19066
rect 23066 19014 23078 19066
rect 23130 19014 23142 19066
rect 23194 19014 23206 19066
rect 23258 19014 25852 19066
rect 1104 18992 25852 19014
rect 3970 18912 3976 18964
rect 4028 18912 4034 18964
rect 8294 18912 8300 18964
rect 8352 18952 8358 18964
rect 10689 18955 10747 18961
rect 10689 18952 10701 18955
rect 8352 18924 10701 18952
rect 8352 18912 8358 18924
rect 10689 18921 10701 18924
rect 10735 18921 10747 18955
rect 10689 18915 10747 18921
rect 11422 18912 11428 18964
rect 11480 18952 11486 18964
rect 12437 18955 12495 18961
rect 12437 18952 12449 18955
rect 11480 18924 12449 18952
rect 11480 18912 11486 18924
rect 12437 18921 12449 18924
rect 12483 18952 12495 18955
rect 12618 18952 12624 18964
rect 12483 18924 12624 18952
rect 12483 18921 12495 18924
rect 12437 18915 12495 18921
rect 12618 18912 12624 18924
rect 12676 18952 12682 18964
rect 19058 18952 19064 18964
rect 12676 18924 13216 18952
rect 12676 18912 12682 18924
rect 9766 18844 9772 18896
rect 9824 18884 9830 18896
rect 9950 18884 9956 18896
rect 9824 18856 9956 18884
rect 9824 18844 9830 18856
rect 9950 18844 9956 18856
rect 10008 18844 10014 18896
rect 12066 18844 12072 18896
rect 12124 18884 12130 18896
rect 12713 18887 12771 18893
rect 12713 18884 12725 18887
rect 12124 18856 12725 18884
rect 12124 18844 12130 18856
rect 12713 18853 12725 18856
rect 12759 18853 12771 18887
rect 12713 18847 12771 18853
rect 6914 18776 6920 18828
rect 6972 18816 6978 18828
rect 7926 18816 7932 18828
rect 6972 18788 7932 18816
rect 6972 18776 6978 18788
rect 7926 18776 7932 18788
rect 7984 18776 7990 18828
rect 8297 18819 8355 18825
rect 8297 18785 8309 18819
rect 8343 18816 8355 18819
rect 8662 18816 8668 18828
rect 8343 18788 8668 18816
rect 8343 18785 8355 18788
rect 8297 18779 8355 18785
rect 8662 18776 8668 18788
rect 8720 18776 8726 18828
rect 11333 18819 11391 18825
rect 11333 18785 11345 18819
rect 11379 18816 11391 18819
rect 12802 18816 12808 18828
rect 11379 18788 12808 18816
rect 11379 18785 11391 18788
rect 11333 18779 11391 18785
rect 12544 18760 12572 18788
rect 12802 18776 12808 18788
rect 12860 18776 12866 18828
rect 13188 18825 13216 18924
rect 17328 18924 19064 18952
rect 13998 18884 14004 18896
rect 13372 18856 14004 18884
rect 13372 18825 13400 18856
rect 13998 18844 14004 18856
rect 14056 18844 14062 18896
rect 13173 18819 13231 18825
rect 13173 18785 13185 18819
rect 13219 18785 13231 18819
rect 13173 18779 13231 18785
rect 13357 18819 13415 18825
rect 13357 18785 13369 18819
rect 13403 18785 13415 18819
rect 15654 18816 15660 18828
rect 13357 18779 13415 18785
rect 13464 18788 15660 18816
rect 2225 18751 2283 18757
rect 2225 18717 2237 18751
rect 2271 18748 2283 18751
rect 2774 18748 2780 18760
rect 2271 18720 2780 18748
rect 2271 18717 2283 18720
rect 2225 18711 2283 18717
rect 2774 18708 2780 18720
rect 2832 18708 2838 18760
rect 4154 18708 4160 18760
rect 4212 18708 4218 18760
rect 8570 18708 8576 18760
rect 8628 18708 8634 18760
rect 12526 18708 12532 18760
rect 12584 18708 12590 18760
rect 13081 18751 13139 18757
rect 13081 18717 13093 18751
rect 13127 18748 13139 18751
rect 13464 18748 13492 18788
rect 15654 18776 15660 18788
rect 15712 18776 15718 18828
rect 17328 18825 17356 18924
rect 19058 18912 19064 18924
rect 19116 18912 19122 18964
rect 22554 18912 22560 18964
rect 22612 18952 22618 18964
rect 23198 18952 23204 18964
rect 22612 18924 23204 18952
rect 22612 18912 22618 18924
rect 23198 18912 23204 18924
rect 23256 18952 23262 18964
rect 23581 18955 23639 18961
rect 23581 18952 23593 18955
rect 23256 18924 23593 18952
rect 23256 18912 23262 18924
rect 23581 18921 23593 18924
rect 23627 18921 23639 18955
rect 23581 18915 23639 18921
rect 24210 18912 24216 18964
rect 24268 18912 24274 18964
rect 17865 18887 17923 18893
rect 17865 18853 17877 18887
rect 17911 18884 17923 18887
rect 19978 18884 19984 18896
rect 17911 18856 19984 18884
rect 17911 18853 17923 18856
rect 17865 18847 17923 18853
rect 19978 18844 19984 18856
rect 20036 18844 20042 18896
rect 20165 18887 20223 18893
rect 20165 18853 20177 18887
rect 20211 18884 20223 18887
rect 20530 18884 20536 18896
rect 20211 18856 20536 18884
rect 20211 18853 20223 18856
rect 20165 18847 20223 18853
rect 20530 18844 20536 18856
rect 20588 18844 20594 18896
rect 21729 18887 21787 18893
rect 21729 18884 21741 18887
rect 20732 18856 21741 18884
rect 17313 18819 17371 18825
rect 17313 18785 17325 18819
rect 17359 18785 17371 18819
rect 17313 18779 17371 18785
rect 17405 18819 17463 18825
rect 17405 18785 17417 18819
rect 17451 18816 17463 18819
rect 17586 18816 17592 18828
rect 17451 18788 17592 18816
rect 17451 18785 17463 18788
rect 17405 18779 17463 18785
rect 17586 18776 17592 18788
rect 17644 18816 17650 18828
rect 18141 18819 18199 18825
rect 18141 18816 18153 18819
rect 17644 18788 18153 18816
rect 17644 18776 17650 18788
rect 18141 18785 18153 18788
rect 18187 18785 18199 18819
rect 18141 18779 18199 18785
rect 19610 18776 19616 18828
rect 19668 18776 19674 18828
rect 19705 18819 19763 18825
rect 19705 18785 19717 18819
rect 19751 18816 19763 18819
rect 20438 18816 20444 18828
rect 19751 18788 20444 18816
rect 19751 18785 19763 18788
rect 19705 18779 19763 18785
rect 20438 18776 20444 18788
rect 20496 18816 20502 18828
rect 20732 18816 20760 18856
rect 21729 18853 21741 18856
rect 21775 18853 21787 18887
rect 21729 18847 21787 18853
rect 20496 18788 20760 18816
rect 20901 18819 20959 18825
rect 20496 18776 20502 18788
rect 20901 18785 20913 18819
rect 20947 18816 20959 18819
rect 20947 18788 22140 18816
rect 20947 18785 20959 18788
rect 20901 18779 20959 18785
rect 13127 18720 13492 18748
rect 13127 18717 13139 18720
rect 13081 18711 13139 18717
rect 13538 18708 13544 18760
rect 13596 18748 13602 18760
rect 16853 18751 16911 18757
rect 16853 18748 16865 18751
rect 13596 18720 16865 18748
rect 13596 18708 13602 18720
rect 16853 18717 16865 18720
rect 16899 18748 16911 18751
rect 17497 18751 17555 18757
rect 17497 18748 17509 18751
rect 16899 18720 17509 18748
rect 16899 18717 16911 18720
rect 16853 18711 16911 18717
rect 17497 18717 17509 18720
rect 17543 18717 17555 18751
rect 17497 18711 17555 18717
rect 20993 18751 21051 18757
rect 20993 18717 21005 18751
rect 21039 18748 21051 18751
rect 21542 18748 21548 18760
rect 21039 18720 21548 18748
rect 21039 18717 21051 18720
rect 20993 18711 21051 18717
rect 21542 18708 21548 18720
rect 21600 18708 21606 18760
rect 9766 18680 9772 18692
rect 7866 18652 9772 18680
rect 7944 18624 7972 18652
rect 9766 18640 9772 18652
rect 9824 18640 9830 18692
rect 11057 18683 11115 18689
rect 11057 18649 11069 18683
rect 11103 18680 11115 18683
rect 13722 18680 13728 18692
rect 11103 18652 13728 18680
rect 11103 18649 11115 18652
rect 11057 18643 11115 18649
rect 13556 18624 13584 18652
rect 13722 18640 13728 18652
rect 13780 18640 13786 18692
rect 1762 18572 1768 18624
rect 1820 18612 1826 18624
rect 2041 18615 2099 18621
rect 2041 18612 2053 18615
rect 1820 18584 2053 18612
rect 1820 18572 1826 18584
rect 2041 18581 2053 18584
rect 2087 18581 2099 18615
rect 2041 18575 2099 18581
rect 6825 18615 6883 18621
rect 6825 18581 6837 18615
rect 6871 18612 6883 18615
rect 7650 18612 7656 18624
rect 6871 18584 7656 18612
rect 6871 18581 6883 18584
rect 6825 18575 6883 18581
rect 7650 18572 7656 18584
rect 7708 18572 7714 18624
rect 7926 18572 7932 18624
rect 7984 18572 7990 18624
rect 9214 18572 9220 18624
rect 9272 18572 9278 18624
rect 10134 18572 10140 18624
rect 10192 18612 10198 18624
rect 10321 18615 10379 18621
rect 10321 18612 10333 18615
rect 10192 18584 10333 18612
rect 10192 18572 10198 18584
rect 10321 18581 10333 18584
rect 10367 18612 10379 18615
rect 11149 18615 11207 18621
rect 11149 18612 11161 18615
rect 10367 18584 11161 18612
rect 10367 18581 10379 18584
rect 10321 18575 10379 18581
rect 11149 18581 11161 18584
rect 11195 18612 11207 18615
rect 11790 18612 11796 18624
rect 11195 18584 11796 18612
rect 11195 18581 11207 18584
rect 11149 18575 11207 18581
rect 11790 18572 11796 18584
rect 11848 18572 11854 18624
rect 13538 18572 13544 18624
rect 13596 18572 13602 18624
rect 14182 18572 14188 18624
rect 14240 18612 14246 18624
rect 19061 18615 19119 18621
rect 19061 18612 19073 18615
rect 14240 18584 19073 18612
rect 14240 18572 14246 18584
rect 19061 18581 19073 18584
rect 19107 18612 19119 18615
rect 19797 18615 19855 18621
rect 19797 18612 19809 18615
rect 19107 18584 19809 18612
rect 19107 18581 19119 18584
rect 19061 18575 19119 18581
rect 19797 18581 19809 18584
rect 19843 18581 19855 18615
rect 19797 18575 19855 18581
rect 20346 18572 20352 18624
rect 20404 18612 20410 18624
rect 21085 18615 21143 18621
rect 21085 18612 21097 18615
rect 20404 18584 21097 18612
rect 20404 18572 20410 18584
rect 21085 18581 21097 18584
rect 21131 18581 21143 18615
rect 21085 18575 21143 18581
rect 21450 18572 21456 18624
rect 21508 18572 21514 18624
rect 22112 18621 22140 18788
rect 22830 18776 22836 18828
rect 22888 18816 22894 18828
rect 23845 18819 23903 18825
rect 23845 18816 23857 18819
rect 22888 18788 23857 18816
rect 22888 18776 22894 18788
rect 23845 18785 23857 18788
rect 23891 18785 23903 18819
rect 23845 18779 23903 18785
rect 24302 18708 24308 18760
rect 24360 18748 24366 18760
rect 24765 18751 24823 18757
rect 24765 18748 24777 18751
rect 24360 18720 24777 18748
rect 24360 18708 24366 18720
rect 24765 18717 24777 18720
rect 24811 18717 24823 18751
rect 24765 18711 24823 18717
rect 23138 18652 23244 18680
rect 22097 18615 22155 18621
rect 22097 18581 22109 18615
rect 22143 18612 22155 18615
rect 22554 18612 22560 18624
rect 22143 18584 22560 18612
rect 22143 18581 22155 18584
rect 22097 18575 22155 18581
rect 22554 18572 22560 18584
rect 22612 18572 22618 18624
rect 22738 18572 22744 18624
rect 22796 18612 22802 18624
rect 23216 18612 23244 18652
rect 23658 18640 23664 18692
rect 23716 18680 23722 18692
rect 24581 18683 24639 18689
rect 24581 18680 24593 18683
rect 23716 18652 24593 18680
rect 23716 18640 23722 18652
rect 24581 18649 24593 18652
rect 24627 18649 24639 18683
rect 24581 18643 24639 18649
rect 24210 18612 24216 18624
rect 22796 18584 24216 18612
rect 22796 18572 22802 18584
rect 24210 18572 24216 18584
rect 24268 18572 24274 18624
rect 1104 18522 25852 18544
rect 1104 18470 7950 18522
rect 8002 18470 8014 18522
rect 8066 18470 8078 18522
rect 8130 18470 8142 18522
rect 8194 18470 8206 18522
rect 8258 18470 17950 18522
rect 18002 18470 18014 18522
rect 18066 18470 18078 18522
rect 18130 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 25852 18522
rect 1104 18448 25852 18470
rect 11238 18408 11244 18420
rect 9784 18380 11244 18408
rect 9784 18284 9812 18380
rect 11238 18368 11244 18380
rect 11296 18408 11302 18420
rect 11517 18411 11575 18417
rect 11517 18408 11529 18411
rect 11296 18380 11529 18408
rect 11296 18368 11302 18380
rect 11517 18377 11529 18380
rect 11563 18377 11575 18411
rect 11517 18371 11575 18377
rect 12434 18368 12440 18420
rect 12492 18368 12498 18420
rect 13630 18368 13636 18420
rect 13688 18368 13694 18420
rect 17681 18411 17739 18417
rect 17681 18377 17693 18411
rect 17727 18408 17739 18411
rect 17770 18408 17776 18420
rect 17727 18380 17776 18408
rect 17727 18377 17739 18380
rect 17681 18371 17739 18377
rect 17770 18368 17776 18380
rect 17828 18408 17834 18420
rect 19981 18411 20039 18417
rect 19981 18408 19993 18411
rect 17828 18380 19993 18408
rect 17828 18368 17834 18380
rect 10873 18343 10931 18349
rect 10873 18309 10885 18343
rect 10919 18340 10931 18343
rect 10919 18312 11652 18340
rect 10919 18309 10931 18312
rect 10873 18303 10931 18309
rect 1765 18275 1823 18281
rect 1765 18241 1777 18275
rect 1811 18272 1823 18275
rect 1854 18272 1860 18284
rect 1811 18244 1860 18272
rect 1811 18241 1823 18244
rect 1765 18235 1823 18241
rect 1854 18232 1860 18244
rect 1912 18232 1918 18284
rect 7929 18275 7987 18281
rect 7929 18241 7941 18275
rect 7975 18272 7987 18275
rect 8294 18272 8300 18284
rect 7975 18244 8300 18272
rect 7975 18241 7987 18244
rect 7929 18235 7987 18241
rect 8294 18232 8300 18244
rect 8352 18232 8358 18284
rect 9766 18232 9772 18284
rect 9824 18232 9830 18284
rect 11624 18272 11652 18312
rect 17126 18300 17132 18352
rect 17184 18300 17190 18352
rect 18892 18349 18920 18380
rect 19981 18377 19993 18380
rect 20027 18408 20039 18411
rect 20027 18380 20392 18408
rect 20027 18377 20039 18380
rect 19981 18371 20039 18377
rect 20364 18349 20392 18380
rect 21818 18368 21824 18420
rect 21876 18408 21882 18420
rect 22738 18408 22744 18420
rect 21876 18380 22744 18408
rect 21876 18368 21882 18380
rect 22738 18368 22744 18380
rect 22796 18368 22802 18420
rect 22922 18368 22928 18420
rect 22980 18408 22986 18420
rect 23198 18408 23204 18420
rect 22980 18380 23204 18408
rect 22980 18368 22986 18380
rect 23198 18368 23204 18380
rect 23256 18408 23262 18420
rect 24397 18411 24455 18417
rect 24397 18408 24409 18411
rect 23256 18380 24409 18408
rect 23256 18368 23262 18380
rect 24397 18377 24409 18380
rect 24443 18377 24455 18411
rect 24397 18371 24455 18377
rect 18877 18343 18935 18349
rect 18877 18309 18889 18343
rect 18923 18340 18935 18343
rect 20349 18343 20407 18349
rect 18923 18312 18957 18340
rect 18923 18309 18935 18312
rect 18877 18303 18935 18309
rect 20349 18309 20361 18343
rect 20395 18309 20407 18343
rect 22830 18340 22836 18352
rect 20349 18303 20407 18309
rect 22664 18312 22836 18340
rect 12434 18272 12440 18284
rect 11624 18244 12440 18272
rect 12434 18232 12440 18244
rect 12492 18232 12498 18284
rect 12805 18275 12863 18281
rect 12805 18241 12817 18275
rect 12851 18272 12863 18275
rect 13906 18272 13912 18284
rect 12851 18244 13912 18272
rect 12851 18241 12863 18244
rect 12805 18235 12863 18241
rect 13906 18232 13912 18244
rect 13964 18232 13970 18284
rect 14001 18275 14059 18281
rect 14001 18241 14013 18275
rect 14047 18272 14059 18275
rect 18782 18272 18788 18284
rect 14047 18244 18788 18272
rect 14047 18241 14059 18244
rect 14001 18235 14059 18241
rect 18782 18232 18788 18244
rect 18840 18232 18846 18284
rect 21177 18275 21235 18281
rect 21177 18241 21189 18275
rect 21223 18272 21235 18275
rect 22002 18272 22008 18284
rect 21223 18244 22008 18272
rect 21223 18241 21235 18244
rect 21177 18235 21235 18241
rect 22002 18232 22008 18244
rect 22060 18272 22066 18284
rect 22664 18281 22692 18312
rect 22830 18300 22836 18312
rect 22888 18300 22894 18352
rect 24210 18340 24216 18352
rect 24150 18312 24216 18340
rect 24210 18300 24216 18312
rect 24268 18340 24274 18352
rect 24673 18343 24731 18349
rect 24673 18340 24685 18343
rect 24268 18312 24685 18340
rect 24268 18300 24274 18312
rect 24673 18309 24685 18312
rect 24719 18309 24731 18343
rect 24673 18303 24731 18309
rect 22649 18275 22707 18281
rect 22649 18272 22661 18275
rect 22060 18244 22661 18272
rect 22060 18232 22066 18244
rect 22649 18241 22661 18244
rect 22695 18241 22707 18275
rect 22649 18235 22707 18241
rect 1302 18164 1308 18216
rect 1360 18204 1366 18216
rect 2041 18207 2099 18213
rect 2041 18204 2053 18207
rect 1360 18176 2053 18204
rect 1360 18164 1366 18176
rect 2041 18173 2053 18176
rect 2087 18173 2099 18207
rect 2041 18167 2099 18173
rect 6270 18164 6276 18216
rect 6328 18204 6334 18216
rect 6822 18204 6828 18216
rect 6328 18176 6828 18204
rect 6328 18164 6334 18176
rect 6822 18164 6828 18176
rect 6880 18204 6886 18216
rect 8570 18204 8576 18216
rect 6880 18176 8576 18204
rect 6880 18164 6886 18176
rect 8570 18164 8576 18176
rect 8628 18204 8634 18216
rect 8665 18207 8723 18213
rect 8665 18204 8677 18207
rect 8628 18176 8677 18204
rect 8628 18164 8634 18176
rect 8665 18173 8677 18176
rect 8711 18173 8723 18207
rect 8665 18167 8723 18173
rect 11146 18164 11152 18216
rect 11204 18164 11210 18216
rect 12161 18207 12219 18213
rect 12161 18173 12173 18207
rect 12207 18204 12219 18207
rect 12710 18204 12716 18216
rect 12207 18176 12716 18204
rect 12207 18173 12219 18176
rect 12161 18167 12219 18173
rect 12710 18164 12716 18176
rect 12768 18204 12774 18216
rect 12897 18207 12955 18213
rect 12897 18204 12909 18207
rect 12768 18176 12909 18204
rect 12768 18164 12774 18176
rect 12897 18173 12909 18176
rect 12943 18173 12955 18207
rect 12897 18167 12955 18173
rect 13081 18207 13139 18213
rect 13081 18173 13093 18207
rect 13127 18204 13139 18207
rect 13354 18204 13360 18216
rect 13127 18176 13360 18204
rect 13127 18173 13139 18176
rect 13081 18167 13139 18173
rect 13354 18164 13360 18176
rect 13412 18164 13418 18216
rect 13814 18164 13820 18216
rect 13872 18204 13878 18216
rect 14093 18207 14151 18213
rect 14093 18204 14105 18207
rect 13872 18176 14105 18204
rect 13872 18164 13878 18176
rect 14093 18173 14105 18176
rect 14139 18173 14151 18207
rect 14093 18167 14151 18173
rect 14185 18207 14243 18213
rect 14185 18173 14197 18207
rect 14231 18173 14243 18207
rect 14185 18167 14243 18173
rect 12434 18096 12440 18148
rect 12492 18136 12498 18148
rect 14200 18136 14228 18167
rect 17770 18164 17776 18216
rect 17828 18204 17834 18216
rect 18049 18207 18107 18213
rect 18049 18204 18061 18207
rect 17828 18176 18061 18204
rect 17828 18164 17834 18176
rect 18049 18173 18061 18176
rect 18095 18173 18107 18207
rect 18049 18167 18107 18173
rect 18506 18164 18512 18216
rect 18564 18204 18570 18216
rect 20070 18204 20076 18216
rect 18564 18176 20076 18204
rect 18564 18164 18570 18176
rect 20070 18164 20076 18176
rect 20128 18164 20134 18216
rect 22925 18207 22983 18213
rect 22925 18173 22937 18207
rect 22971 18204 22983 18207
rect 23290 18204 23296 18216
rect 22971 18176 23296 18204
rect 22971 18173 22983 18176
rect 22925 18167 22983 18173
rect 23290 18164 23296 18176
rect 23348 18164 23354 18216
rect 12492 18108 14228 18136
rect 12492 18096 12498 18108
rect 2130 18028 2136 18080
rect 2188 18068 2194 18080
rect 7282 18068 7288 18080
rect 2188 18040 7288 18068
rect 2188 18028 2194 18040
rect 7282 18028 7288 18040
rect 7340 18028 7346 18080
rect 9401 18071 9459 18077
rect 9401 18037 9413 18071
rect 9447 18068 9459 18071
rect 10686 18068 10692 18080
rect 9447 18040 10692 18068
rect 9447 18037 9459 18040
rect 9401 18031 9459 18037
rect 10686 18028 10692 18040
rect 10744 18028 10750 18080
rect 13906 18028 13912 18080
rect 13964 18068 13970 18080
rect 17037 18071 17095 18077
rect 17037 18068 17049 18071
rect 13964 18040 17049 18068
rect 13964 18028 13970 18040
rect 17037 18037 17049 18040
rect 17083 18068 17095 18071
rect 18506 18068 18512 18080
rect 17083 18040 18512 18068
rect 17083 18037 17095 18040
rect 17037 18031 17095 18037
rect 18506 18028 18512 18040
rect 18564 18028 18570 18080
rect 21637 18071 21695 18077
rect 21637 18037 21649 18071
rect 21683 18068 21695 18071
rect 21818 18068 21824 18080
rect 21683 18040 21824 18068
rect 21683 18037 21695 18040
rect 21637 18031 21695 18037
rect 21818 18028 21824 18040
rect 21876 18028 21882 18080
rect 1104 17978 25852 18000
rect 1104 17926 2950 17978
rect 3002 17926 3014 17978
rect 3066 17926 3078 17978
rect 3130 17926 3142 17978
rect 3194 17926 3206 17978
rect 3258 17926 12950 17978
rect 13002 17926 13014 17978
rect 13066 17926 13078 17978
rect 13130 17926 13142 17978
rect 13194 17926 13206 17978
rect 13258 17926 22950 17978
rect 23002 17926 23014 17978
rect 23066 17926 23078 17978
rect 23130 17926 23142 17978
rect 23194 17926 23206 17978
rect 23258 17926 25852 17978
rect 1104 17904 25852 17926
rect 4338 17824 4344 17876
rect 4396 17864 4402 17876
rect 4396 17836 7052 17864
rect 4396 17824 4402 17836
rect 6914 17756 6920 17808
rect 6972 17756 6978 17808
rect 7024 17796 7052 17836
rect 8294 17824 8300 17876
rect 8352 17864 8358 17876
rect 8665 17867 8723 17873
rect 8665 17864 8677 17867
rect 8352 17836 8677 17864
rect 8352 17824 8358 17836
rect 8665 17833 8677 17836
rect 8711 17833 8723 17867
rect 8665 17827 8723 17833
rect 9493 17867 9551 17873
rect 9493 17833 9505 17867
rect 9539 17864 9551 17867
rect 11882 17864 11888 17876
rect 9539 17836 11888 17864
rect 9539 17833 9551 17836
rect 9493 17827 9551 17833
rect 7024 17768 8340 17796
rect 6270 17688 6276 17740
rect 6328 17728 6334 17740
rect 6549 17731 6607 17737
rect 6549 17728 6561 17731
rect 6328 17700 6561 17728
rect 6328 17688 6334 17700
rect 6549 17697 6561 17700
rect 6595 17697 6607 17731
rect 6549 17691 6607 17697
rect 7650 17688 7656 17740
rect 7708 17688 7714 17740
rect 7837 17663 7895 17669
rect 7837 17629 7849 17663
rect 7883 17660 7895 17663
rect 8202 17660 8208 17672
rect 7883 17632 8208 17660
rect 7883 17629 7895 17632
rect 7837 17623 7895 17629
rect 8202 17620 8208 17632
rect 8260 17620 8266 17672
rect 5718 17552 5724 17604
rect 5776 17552 5782 17604
rect 6273 17595 6331 17601
rect 6273 17561 6285 17595
rect 6319 17592 6331 17595
rect 6546 17592 6552 17604
rect 6319 17564 6552 17592
rect 6319 17561 6331 17564
rect 6273 17555 6331 17561
rect 6546 17552 6552 17564
rect 6604 17552 6610 17604
rect 7193 17595 7251 17601
rect 7193 17592 7205 17595
rect 6656 17564 7205 17592
rect 4798 17484 4804 17536
rect 4856 17484 4862 17536
rect 4890 17484 4896 17536
rect 4948 17524 4954 17536
rect 6656 17524 6684 17564
rect 7193 17561 7205 17564
rect 7239 17592 7251 17595
rect 7929 17595 7987 17601
rect 7929 17592 7941 17595
rect 7239 17564 7941 17592
rect 7239 17561 7251 17564
rect 7193 17555 7251 17561
rect 7929 17561 7941 17564
rect 7975 17561 7987 17595
rect 8312 17592 8340 17768
rect 8680 17728 8708 17827
rect 11882 17824 11888 17836
rect 11940 17824 11946 17876
rect 12802 17824 12808 17876
rect 12860 17864 12866 17876
rect 13541 17867 13599 17873
rect 13541 17864 13553 17867
rect 12860 17836 13553 17864
rect 12860 17824 12866 17836
rect 13541 17833 13553 17836
rect 13587 17864 13599 17867
rect 13722 17864 13728 17876
rect 13587 17836 13728 17864
rect 13587 17833 13599 17836
rect 13541 17827 13599 17833
rect 13722 17824 13728 17836
rect 13780 17824 13786 17876
rect 15286 17824 15292 17876
rect 15344 17864 15350 17876
rect 16025 17867 16083 17873
rect 16025 17864 16037 17867
rect 15344 17836 16037 17864
rect 15344 17824 15350 17836
rect 16025 17833 16037 17836
rect 16071 17833 16083 17867
rect 16025 17827 16083 17833
rect 18322 17824 18328 17876
rect 18380 17864 18386 17876
rect 18966 17864 18972 17876
rect 18380 17836 18972 17864
rect 18380 17824 18386 17836
rect 18966 17824 18972 17836
rect 19024 17824 19030 17876
rect 11514 17728 11520 17740
rect 8680 17700 11520 17728
rect 8386 17620 8392 17672
rect 8444 17660 8450 17672
rect 9306 17660 9312 17672
rect 8444 17632 9312 17660
rect 8444 17620 8450 17632
rect 9306 17620 9312 17632
rect 9364 17620 9370 17672
rect 11256 17669 11284 17700
rect 11514 17688 11520 17700
rect 11572 17688 11578 17740
rect 11974 17688 11980 17740
rect 12032 17728 12038 17740
rect 13081 17731 13139 17737
rect 13081 17728 13093 17731
rect 12032 17700 13093 17728
rect 12032 17688 12038 17700
rect 13081 17697 13093 17700
rect 13127 17728 13139 17731
rect 13630 17728 13636 17740
rect 13127 17700 13636 17728
rect 13127 17697 13139 17700
rect 13081 17691 13139 17697
rect 13630 17688 13636 17700
rect 13688 17688 13694 17740
rect 13906 17688 13912 17740
rect 13964 17728 13970 17740
rect 14737 17731 14795 17737
rect 14737 17728 14749 17731
rect 13964 17700 14749 17728
rect 13964 17688 13970 17700
rect 14737 17697 14749 17700
rect 14783 17697 14795 17731
rect 14737 17691 14795 17697
rect 14921 17731 14979 17737
rect 14921 17697 14933 17731
rect 14967 17728 14979 17731
rect 15470 17728 15476 17740
rect 14967 17700 15476 17728
rect 14967 17697 14979 17700
rect 14921 17691 14979 17697
rect 15470 17688 15476 17700
rect 15528 17688 15534 17740
rect 16850 17688 16856 17740
rect 16908 17728 16914 17740
rect 17770 17728 17776 17740
rect 16908 17700 17776 17728
rect 16908 17688 16914 17700
rect 17770 17688 17776 17700
rect 17828 17688 17834 17740
rect 17862 17688 17868 17740
rect 17920 17728 17926 17740
rect 19429 17731 19487 17737
rect 17920 17700 18736 17728
rect 17920 17688 17926 17700
rect 9585 17663 9643 17669
rect 9585 17629 9597 17663
rect 9631 17660 9643 17663
rect 9861 17663 9919 17669
rect 9861 17660 9873 17663
rect 9631 17632 9873 17660
rect 9631 17629 9643 17632
rect 9585 17623 9643 17629
rect 9861 17629 9873 17632
rect 9907 17629 9919 17663
rect 9861 17623 9919 17629
rect 11241 17663 11299 17669
rect 11241 17629 11253 17663
rect 11287 17629 11299 17663
rect 11241 17623 11299 17629
rect 12989 17663 13047 17669
rect 12989 17629 13001 17663
rect 13035 17660 13047 17663
rect 14274 17660 14280 17672
rect 13035 17632 14280 17660
rect 13035 17629 13047 17632
rect 12989 17623 13047 17629
rect 9600 17592 9628 17623
rect 14274 17620 14280 17632
rect 14332 17620 14338 17672
rect 18598 17660 18604 17672
rect 18248 17632 18604 17660
rect 8312 17564 9628 17592
rect 10505 17595 10563 17601
rect 7929 17555 7987 17561
rect 10505 17561 10517 17595
rect 10551 17592 10563 17595
rect 10594 17592 10600 17604
rect 10551 17564 10600 17592
rect 10551 17561 10563 17564
rect 10505 17555 10563 17561
rect 10594 17552 10600 17564
rect 10652 17592 10658 17604
rect 11146 17592 11152 17604
rect 10652 17564 11152 17592
rect 10652 17552 10658 17564
rect 11146 17552 11152 17564
rect 11204 17552 11210 17604
rect 12897 17595 12955 17601
rect 12897 17561 12909 17595
rect 12943 17592 12955 17595
rect 12943 17564 14320 17592
rect 12943 17561 12955 17564
rect 12897 17555 12955 17561
rect 4948 17496 6684 17524
rect 4948 17484 4954 17496
rect 8294 17484 8300 17536
rect 8352 17484 8358 17536
rect 9122 17484 9128 17536
rect 9180 17484 9186 17536
rect 12526 17484 12532 17536
rect 12584 17484 12590 17536
rect 14292 17533 14320 17564
rect 16482 17552 16488 17604
rect 16540 17552 16546 17604
rect 17497 17595 17555 17601
rect 17497 17561 17509 17595
rect 17543 17592 17555 17595
rect 18248 17592 18276 17632
rect 18598 17620 18604 17632
rect 18656 17620 18662 17672
rect 18708 17660 18736 17700
rect 19429 17697 19441 17731
rect 19475 17728 19487 17731
rect 22002 17728 22008 17740
rect 19475 17700 22008 17728
rect 19475 17697 19487 17700
rect 19429 17691 19487 17697
rect 22002 17688 22008 17700
rect 22060 17688 22066 17740
rect 23382 17688 23388 17740
rect 23440 17688 23446 17740
rect 24029 17663 24087 17669
rect 18708 17632 19012 17660
rect 17543 17564 18276 17592
rect 17543 17561 17555 17564
rect 17497 17555 17555 17561
rect 18322 17552 18328 17604
rect 18380 17552 18386 17604
rect 18509 17595 18567 17601
rect 18509 17561 18521 17595
rect 18555 17592 18567 17595
rect 18874 17592 18880 17604
rect 18555 17564 18880 17592
rect 18555 17561 18567 17564
rect 18509 17555 18567 17561
rect 18874 17552 18880 17564
rect 18932 17552 18938 17604
rect 14277 17527 14335 17533
rect 14277 17493 14289 17527
rect 14323 17493 14335 17527
rect 14277 17487 14335 17493
rect 14645 17527 14703 17533
rect 14645 17493 14657 17527
rect 14691 17524 14703 17527
rect 15381 17527 15439 17533
rect 15381 17524 15393 17527
rect 14691 17496 15393 17524
rect 14691 17493 14703 17496
rect 14645 17487 14703 17493
rect 15381 17493 15393 17496
rect 15427 17524 15439 17527
rect 17862 17524 17868 17536
rect 15427 17496 17868 17524
rect 15427 17493 15439 17496
rect 15381 17487 15439 17493
rect 17862 17484 17868 17496
rect 17920 17484 17926 17536
rect 18690 17484 18696 17536
rect 18748 17524 18754 17536
rect 18785 17527 18843 17533
rect 18785 17524 18797 17527
rect 18748 17496 18797 17524
rect 18748 17484 18754 17496
rect 18785 17493 18797 17496
rect 18831 17493 18843 17527
rect 18984 17524 19012 17632
rect 24029 17629 24041 17663
rect 24075 17660 24087 17663
rect 24670 17660 24676 17672
rect 24075 17632 24676 17660
rect 24075 17629 24087 17632
rect 24029 17623 24087 17629
rect 24670 17620 24676 17632
rect 24728 17620 24734 17672
rect 19058 17552 19064 17604
rect 19116 17592 19122 17604
rect 19705 17595 19763 17601
rect 19705 17592 19717 17595
rect 19116 17564 19717 17592
rect 19116 17552 19122 17564
rect 19705 17561 19717 17564
rect 19751 17561 19763 17595
rect 19705 17555 19763 17561
rect 20714 17552 20720 17604
rect 20772 17552 20778 17604
rect 21729 17595 21787 17601
rect 21729 17592 21741 17595
rect 21008 17564 21741 17592
rect 21008 17524 21036 17564
rect 21729 17561 21741 17564
rect 21775 17561 21787 17595
rect 21729 17555 21787 17561
rect 21913 17595 21971 17601
rect 21913 17561 21925 17595
rect 21959 17592 21971 17595
rect 22094 17592 22100 17604
rect 21959 17564 22100 17592
rect 21959 17561 21971 17564
rect 21913 17555 21971 17561
rect 22094 17552 22100 17564
rect 22152 17552 22158 17604
rect 18984 17496 21036 17524
rect 18785 17487 18843 17493
rect 21174 17484 21180 17536
rect 21232 17484 21238 17536
rect 21818 17484 21824 17536
rect 21876 17524 21882 17536
rect 22189 17527 22247 17533
rect 22189 17524 22201 17527
rect 21876 17496 22201 17524
rect 21876 17484 21882 17496
rect 22189 17493 22201 17496
rect 22235 17493 22247 17527
rect 22189 17487 22247 17493
rect 1104 17434 25852 17456
rect 1104 17382 7950 17434
rect 8002 17382 8014 17434
rect 8066 17382 8078 17434
rect 8130 17382 8142 17434
rect 8194 17382 8206 17434
rect 8258 17382 17950 17434
rect 18002 17382 18014 17434
rect 18066 17382 18078 17434
rect 18130 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 25852 17434
rect 1104 17360 25852 17382
rect 4154 17280 4160 17332
rect 4212 17320 4218 17332
rect 5261 17323 5319 17329
rect 5261 17320 5273 17323
rect 4212 17292 5273 17320
rect 4212 17280 4218 17292
rect 5261 17289 5273 17292
rect 5307 17289 5319 17323
rect 5261 17283 5319 17289
rect 5629 17323 5687 17329
rect 5629 17289 5641 17323
rect 5675 17320 5687 17323
rect 7009 17323 7067 17329
rect 7009 17320 7021 17323
rect 5675 17292 7021 17320
rect 5675 17289 5687 17292
rect 5629 17283 5687 17289
rect 7009 17289 7021 17292
rect 7055 17289 7067 17323
rect 7009 17283 7067 17289
rect 7469 17323 7527 17329
rect 7469 17289 7481 17323
rect 7515 17320 7527 17323
rect 7834 17320 7840 17332
rect 7515 17292 7840 17320
rect 7515 17289 7527 17292
rect 7469 17283 7527 17289
rect 7834 17280 7840 17292
rect 7892 17280 7898 17332
rect 9582 17280 9588 17332
rect 9640 17320 9646 17332
rect 10137 17323 10195 17329
rect 10137 17320 10149 17323
rect 9640 17292 10149 17320
rect 9640 17280 9646 17292
rect 10137 17289 10149 17292
rect 10183 17289 10195 17323
rect 11701 17323 11759 17329
rect 11701 17320 11713 17323
rect 10137 17283 10195 17289
rect 10428 17292 11713 17320
rect 5718 17212 5724 17264
rect 5776 17252 5782 17264
rect 9125 17255 9183 17261
rect 5776 17224 5948 17252
rect 5776 17212 5782 17224
rect 4798 17144 4804 17196
rect 4856 17184 4862 17196
rect 5920 17184 5948 17224
rect 9125 17221 9137 17255
rect 9171 17252 9183 17255
rect 10428 17252 10456 17292
rect 11701 17289 11713 17292
rect 11747 17289 11759 17323
rect 11701 17283 11759 17289
rect 12066 17280 12072 17332
rect 12124 17280 12130 17332
rect 12158 17280 12164 17332
rect 12216 17280 12222 17332
rect 12710 17280 12716 17332
rect 12768 17320 12774 17332
rect 13633 17323 13691 17329
rect 12768 17292 13032 17320
rect 12768 17280 12774 17292
rect 9171 17224 10456 17252
rect 10597 17255 10655 17261
rect 9171 17221 9183 17224
rect 9125 17215 9183 17221
rect 10597 17221 10609 17255
rect 10643 17252 10655 17255
rect 10643 17224 12434 17252
rect 10643 17221 10655 17224
rect 10597 17215 10655 17221
rect 6914 17184 6920 17196
rect 4856 17156 5856 17184
rect 5920 17156 6920 17184
rect 4856 17144 4862 17156
rect 5828 17125 5856 17156
rect 6914 17144 6920 17156
rect 6972 17144 6978 17196
rect 7377 17187 7435 17193
rect 7377 17153 7389 17187
rect 7423 17184 7435 17187
rect 8754 17184 8760 17196
rect 7423 17156 8760 17184
rect 7423 17153 7435 17156
rect 7377 17147 7435 17153
rect 8754 17144 8760 17156
rect 8812 17144 8818 17196
rect 9217 17187 9275 17193
rect 9217 17153 9229 17187
rect 9263 17184 9275 17187
rect 10505 17187 10563 17193
rect 9263 17156 10456 17184
rect 9263 17153 9275 17156
rect 9217 17147 9275 17153
rect 5721 17119 5779 17125
rect 5721 17085 5733 17119
rect 5767 17085 5779 17119
rect 5721 17079 5779 17085
rect 5813 17119 5871 17125
rect 5813 17085 5825 17119
rect 5859 17116 5871 17119
rect 6086 17116 6092 17128
rect 5859 17088 6092 17116
rect 5859 17085 5871 17088
rect 5813 17079 5871 17085
rect 5736 17048 5764 17079
rect 6086 17076 6092 17088
rect 6144 17076 6150 17128
rect 6546 17076 6552 17128
rect 6604 17116 6610 17128
rect 7561 17119 7619 17125
rect 7561 17116 7573 17119
rect 6604 17088 7573 17116
rect 6604 17076 6610 17088
rect 7561 17085 7573 17088
rect 7607 17116 7619 17119
rect 9309 17119 9367 17125
rect 7607 17088 9168 17116
rect 7607 17085 7619 17088
rect 7561 17079 7619 17085
rect 8757 17051 8815 17057
rect 8757 17048 8769 17051
rect 5736 17020 8769 17048
rect 8757 17017 8769 17020
rect 8803 17017 8815 17051
rect 9140 17048 9168 17088
rect 9309 17085 9321 17119
rect 9355 17085 9367 17119
rect 9309 17079 9367 17085
rect 9324 17048 9352 17079
rect 9140 17020 9352 17048
rect 8757 17011 8815 17017
rect 4062 16940 4068 16992
rect 4120 16980 4126 16992
rect 9122 16980 9128 16992
rect 4120 16952 9128 16980
rect 4120 16940 4126 16952
rect 9122 16940 9128 16952
rect 9180 16940 9186 16992
rect 10428 16980 10456 17156
rect 10505 17153 10517 17187
rect 10551 17153 10563 17187
rect 12406 17184 12434 17224
rect 12710 17184 12716 17196
rect 12406 17156 12716 17184
rect 10505 17147 10563 17153
rect 10520 17048 10548 17147
rect 12710 17144 12716 17156
rect 12768 17144 12774 17196
rect 10686 17076 10692 17128
rect 10744 17076 10750 17128
rect 11054 17076 11060 17128
rect 11112 17116 11118 17128
rect 13004 17125 13032 17292
rect 13633 17289 13645 17323
rect 13679 17320 13691 17323
rect 13722 17320 13728 17332
rect 13679 17292 13728 17320
rect 13679 17289 13691 17292
rect 13633 17283 13691 17289
rect 13722 17280 13728 17292
rect 13780 17280 13786 17332
rect 15841 17323 15899 17329
rect 15841 17289 15853 17323
rect 15887 17320 15899 17323
rect 16666 17320 16672 17332
rect 15887 17292 16672 17320
rect 15887 17289 15899 17292
rect 15841 17283 15899 17289
rect 16666 17280 16672 17292
rect 16724 17280 16730 17332
rect 19058 17280 19064 17332
rect 19116 17280 19122 17332
rect 19610 17280 19616 17332
rect 19668 17320 19674 17332
rect 19705 17323 19763 17329
rect 19705 17320 19717 17323
rect 19668 17292 19717 17320
rect 19668 17280 19674 17292
rect 19705 17289 19717 17292
rect 19751 17320 19763 17323
rect 19751 17292 22324 17320
rect 19751 17289 19763 17292
rect 19705 17283 19763 17289
rect 14366 17212 14372 17264
rect 14424 17252 14430 17264
rect 14737 17255 14795 17261
rect 14737 17252 14749 17255
rect 14424 17224 14749 17252
rect 14424 17212 14430 17224
rect 14737 17221 14749 17224
rect 14783 17221 14795 17255
rect 14737 17215 14795 17221
rect 20714 17212 20720 17264
rect 20772 17252 20778 17264
rect 21910 17252 21916 17264
rect 20772 17224 21916 17252
rect 20772 17212 20778 17224
rect 21910 17212 21916 17224
rect 21968 17212 21974 17264
rect 22296 17261 22324 17292
rect 23290 17280 23296 17332
rect 23348 17320 23354 17332
rect 23753 17323 23811 17329
rect 23753 17320 23765 17323
rect 23348 17292 23765 17320
rect 23348 17280 23354 17292
rect 23753 17289 23765 17292
rect 23799 17289 23811 17323
rect 23753 17283 23811 17289
rect 24121 17323 24179 17329
rect 24121 17289 24133 17323
rect 24167 17320 24179 17323
rect 24210 17320 24216 17332
rect 24167 17292 24216 17320
rect 24167 17289 24179 17292
rect 24121 17283 24179 17289
rect 22281 17255 22339 17261
rect 22281 17221 22293 17255
rect 22327 17221 22339 17255
rect 24136 17252 24164 17283
rect 24210 17280 24216 17292
rect 24268 17280 24274 17332
rect 23506 17224 24164 17252
rect 22281 17215 22339 17221
rect 13906 17144 13912 17196
rect 13964 17184 13970 17196
rect 15933 17187 15991 17193
rect 15933 17184 15945 17187
rect 13964 17156 15945 17184
rect 13964 17144 13970 17156
rect 15933 17153 15945 17156
rect 15979 17153 15991 17187
rect 15933 17147 15991 17153
rect 18690 17144 18696 17196
rect 18748 17144 18754 17196
rect 12253 17119 12311 17125
rect 12253 17116 12265 17119
rect 11112 17088 12265 17116
rect 11112 17076 11118 17088
rect 12253 17085 12265 17088
rect 12299 17085 12311 17119
rect 12253 17079 12311 17085
rect 12989 17119 13047 17125
rect 12989 17085 13001 17119
rect 13035 17116 13047 17119
rect 13722 17116 13728 17128
rect 13035 17088 13728 17116
rect 13035 17085 13047 17088
rect 12989 17079 13047 17085
rect 13722 17076 13728 17088
rect 13780 17076 13786 17128
rect 13817 17119 13875 17125
rect 13817 17085 13829 17119
rect 13863 17085 13875 17119
rect 13817 17079 13875 17085
rect 15749 17119 15807 17125
rect 15749 17085 15761 17119
rect 15795 17085 15807 17119
rect 15749 17079 15807 17085
rect 13265 17051 13323 17057
rect 13265 17048 13277 17051
rect 10520 17020 13277 17048
rect 13265 17017 13277 17020
rect 13311 17017 13323 17051
rect 13832 17048 13860 17079
rect 13265 17011 13323 17017
rect 13648 17020 13860 17048
rect 15764 17048 15792 17079
rect 16850 17076 16856 17128
rect 16908 17116 16914 17128
rect 17313 17119 17371 17125
rect 17313 17116 17325 17119
rect 16908 17088 17325 17116
rect 16908 17076 16914 17088
rect 17313 17085 17325 17088
rect 17359 17085 17371 17119
rect 17313 17079 17371 17085
rect 17586 17076 17592 17128
rect 17644 17076 17650 17128
rect 18708 17116 18736 17144
rect 19429 17119 19487 17125
rect 19429 17116 19441 17119
rect 18708 17088 19441 17116
rect 19429 17085 19441 17088
rect 19475 17116 19487 17119
rect 20714 17116 20720 17128
rect 19475 17088 20720 17116
rect 19475 17085 19487 17088
rect 19429 17079 19487 17085
rect 20714 17076 20720 17088
rect 20772 17076 20778 17128
rect 21174 17076 21180 17128
rect 21232 17076 21238 17128
rect 21453 17119 21511 17125
rect 21453 17085 21465 17119
rect 21499 17116 21511 17119
rect 21542 17116 21548 17128
rect 21499 17088 21548 17116
rect 21499 17085 21511 17088
rect 21453 17079 21511 17085
rect 21542 17076 21548 17088
rect 21600 17116 21606 17128
rect 22002 17116 22008 17128
rect 21600 17088 22008 17116
rect 21600 17076 21606 17088
rect 22002 17076 22008 17088
rect 22060 17076 22066 17128
rect 16114 17048 16120 17060
rect 15764 17020 16120 17048
rect 11790 16980 11796 16992
rect 10428 16952 11796 16980
rect 11790 16940 11796 16952
rect 11848 16940 11854 16992
rect 12434 16940 12440 16992
rect 12492 16980 12498 16992
rect 13648 16980 13676 17020
rect 16114 17008 16120 17020
rect 16172 17008 16178 17060
rect 16301 17051 16359 17057
rect 16301 17017 16313 17051
rect 16347 17048 16359 17051
rect 16347 17020 17448 17048
rect 16347 17017 16359 17020
rect 16301 17011 16359 17017
rect 12492 16952 13676 16980
rect 12492 16940 12498 16952
rect 14734 16940 14740 16992
rect 14792 16980 14798 16992
rect 14829 16983 14887 16989
rect 14829 16980 14841 16983
rect 14792 16952 14841 16980
rect 14792 16940 14798 16952
rect 14829 16949 14841 16952
rect 14875 16949 14887 16983
rect 17420 16980 17448 17020
rect 18322 16980 18328 16992
rect 17420 16952 18328 16980
rect 14829 16943 14887 16949
rect 18322 16940 18328 16952
rect 18380 16940 18386 16992
rect 1104 16890 25852 16912
rect 1104 16838 2950 16890
rect 3002 16838 3014 16890
rect 3066 16838 3078 16890
rect 3130 16838 3142 16890
rect 3194 16838 3206 16890
rect 3258 16838 12950 16890
rect 13002 16838 13014 16890
rect 13066 16838 13078 16890
rect 13130 16838 13142 16890
rect 13194 16838 13206 16890
rect 13258 16838 22950 16890
rect 23002 16838 23014 16890
rect 23066 16838 23078 16890
rect 23130 16838 23142 16890
rect 23194 16838 23206 16890
rect 23258 16838 25852 16890
rect 1104 16816 25852 16838
rect 5892 16779 5950 16785
rect 5892 16745 5904 16779
rect 5938 16776 5950 16779
rect 6086 16776 6092 16788
rect 5938 16748 6092 16776
rect 5938 16745 5950 16748
rect 5892 16739 5950 16745
rect 6086 16736 6092 16748
rect 6144 16736 6150 16788
rect 6914 16736 6920 16788
rect 6972 16776 6978 16788
rect 7834 16776 7840 16788
rect 6972 16748 7840 16776
rect 6972 16736 6978 16748
rect 2409 16643 2467 16649
rect 2409 16609 2421 16643
rect 2455 16640 2467 16643
rect 2774 16640 2780 16652
rect 2455 16612 2780 16640
rect 2455 16609 2467 16612
rect 2409 16603 2467 16609
rect 2774 16600 2780 16612
rect 2832 16600 2838 16652
rect 5629 16643 5687 16649
rect 5629 16609 5641 16643
rect 5675 16640 5687 16643
rect 6270 16640 6276 16652
rect 5675 16612 6276 16640
rect 5675 16609 5687 16612
rect 5629 16603 5687 16609
rect 6270 16600 6276 16612
rect 6328 16600 6334 16652
rect 2593 16575 2651 16581
rect 2593 16541 2605 16575
rect 2639 16572 2651 16575
rect 4062 16572 4068 16584
rect 2639 16544 4068 16572
rect 2639 16541 2651 16544
rect 2593 16535 2651 16541
rect 4062 16532 4068 16544
rect 4120 16532 4126 16584
rect 7024 16558 7052 16748
rect 7834 16736 7840 16748
rect 7892 16776 7898 16788
rect 7929 16779 7987 16785
rect 7929 16776 7941 16779
rect 7892 16748 7941 16776
rect 7892 16736 7898 16748
rect 7929 16745 7941 16748
rect 7975 16745 7987 16779
rect 7929 16739 7987 16745
rect 11422 16736 11428 16788
rect 11480 16776 11486 16788
rect 14918 16776 14924 16788
rect 11480 16748 14924 16776
rect 11480 16736 11486 16748
rect 14918 16736 14924 16748
rect 14976 16776 14982 16788
rect 15378 16776 15384 16788
rect 14976 16748 15384 16776
rect 14976 16736 14982 16748
rect 15378 16736 15384 16748
rect 15436 16736 15442 16788
rect 16206 16736 16212 16788
rect 16264 16736 16270 16788
rect 18506 16736 18512 16788
rect 18564 16776 18570 16788
rect 18782 16776 18788 16788
rect 18564 16748 18788 16776
rect 18564 16736 18570 16748
rect 18782 16736 18788 16748
rect 18840 16736 18846 16788
rect 21542 16736 21548 16788
rect 21600 16776 21606 16788
rect 21600 16748 23336 16776
rect 21600 16736 21606 16748
rect 9858 16708 9864 16720
rect 8680 16680 9864 16708
rect 7653 16507 7711 16513
rect 7653 16473 7665 16507
rect 7699 16504 7711 16507
rect 8680 16504 8708 16680
rect 9858 16668 9864 16680
rect 9916 16708 9922 16720
rect 9916 16680 10916 16708
rect 9916 16668 9922 16680
rect 9582 16600 9588 16652
rect 9640 16600 9646 16652
rect 9677 16643 9735 16649
rect 9677 16609 9689 16643
rect 9723 16609 9735 16643
rect 9677 16603 9735 16609
rect 8846 16532 8852 16584
rect 8904 16572 8910 16584
rect 9692 16572 9720 16603
rect 10778 16600 10784 16652
rect 10836 16600 10842 16652
rect 10888 16649 10916 16680
rect 11698 16668 11704 16720
rect 11756 16708 11762 16720
rect 15470 16708 15476 16720
rect 11756 16680 12020 16708
rect 11756 16668 11762 16680
rect 10873 16643 10931 16649
rect 10873 16609 10885 16643
rect 10919 16609 10931 16643
rect 11885 16643 11943 16649
rect 11885 16640 11897 16643
rect 10873 16603 10931 16609
rect 10980 16612 11897 16640
rect 8904 16544 9720 16572
rect 8904 16532 8910 16544
rect 10594 16532 10600 16584
rect 10652 16572 10658 16584
rect 10980 16572 11008 16612
rect 11885 16609 11897 16612
rect 11931 16609 11943 16643
rect 11992 16640 12020 16680
rect 13740 16680 15476 16708
rect 12161 16643 12219 16649
rect 12161 16640 12173 16643
rect 11992 16612 12173 16640
rect 11885 16603 11943 16609
rect 12161 16609 12173 16612
rect 12207 16640 12219 16643
rect 13740 16640 13768 16680
rect 15470 16668 15476 16680
rect 15528 16668 15534 16720
rect 14093 16643 14151 16649
rect 14093 16640 14105 16643
rect 12207 16612 13768 16640
rect 13832 16612 14105 16640
rect 12207 16609 12219 16612
rect 12161 16603 12219 16609
rect 13832 16572 13860 16612
rect 14093 16609 14105 16612
rect 14139 16609 14151 16643
rect 14093 16603 14151 16609
rect 19978 16600 19984 16652
rect 20036 16600 20042 16652
rect 20073 16643 20131 16649
rect 20073 16609 20085 16643
rect 20119 16640 20131 16643
rect 21174 16640 21180 16652
rect 20119 16612 21180 16640
rect 20119 16609 20131 16612
rect 20073 16603 20131 16609
rect 21174 16600 21180 16612
rect 21232 16600 21238 16652
rect 22554 16600 22560 16652
rect 22612 16640 22618 16652
rect 23109 16643 23167 16649
rect 23109 16640 23121 16643
rect 22612 16612 23121 16640
rect 22612 16600 22618 16612
rect 23109 16609 23121 16612
rect 23155 16609 23167 16643
rect 23308 16640 23336 16748
rect 24210 16736 24216 16788
rect 24268 16776 24274 16788
rect 24397 16779 24455 16785
rect 24397 16776 24409 16779
rect 24268 16748 24409 16776
rect 24268 16736 24274 16748
rect 24397 16745 24409 16748
rect 24443 16745 24455 16779
rect 24397 16739 24455 16745
rect 23385 16643 23443 16649
rect 23385 16640 23397 16643
rect 23308 16612 23397 16640
rect 23109 16603 23167 16609
rect 23385 16609 23397 16612
rect 23431 16609 23443 16643
rect 23385 16603 23443 16609
rect 10652 16544 11008 16572
rect 13294 16558 13860 16572
rect 13280 16544 13860 16558
rect 10652 16532 10658 16544
rect 9493 16507 9551 16513
rect 7699 16476 8708 16504
rect 9048 16476 9260 16504
rect 7699 16473 7711 16476
rect 7653 16467 7711 16473
rect 7742 16396 7748 16448
rect 7800 16436 7806 16448
rect 9048 16436 9076 16476
rect 7800 16408 9076 16436
rect 7800 16396 7806 16408
rect 9122 16396 9128 16448
rect 9180 16396 9186 16448
rect 9232 16436 9260 16476
rect 9493 16473 9505 16507
rect 9539 16504 9551 16507
rect 10502 16504 10508 16516
rect 9539 16476 10508 16504
rect 9539 16473 9551 16476
rect 9493 16467 9551 16473
rect 10502 16464 10508 16476
rect 10560 16464 10566 16516
rect 10689 16507 10747 16513
rect 10689 16473 10701 16507
rect 10735 16504 10747 16507
rect 11422 16504 11428 16516
rect 10735 16476 11428 16504
rect 10735 16473 10747 16476
rect 10689 16467 10747 16473
rect 11422 16464 11428 16476
rect 11480 16464 11486 16516
rect 10321 16439 10379 16445
rect 10321 16436 10333 16439
rect 9232 16408 10333 16436
rect 10321 16405 10333 16408
rect 10367 16405 10379 16439
rect 10321 16399 10379 16405
rect 11238 16396 11244 16448
rect 11296 16436 11302 16448
rect 13280 16436 13308 16544
rect 15746 16532 15752 16584
rect 15804 16532 15810 16584
rect 19996 16572 20024 16600
rect 20165 16575 20223 16581
rect 20165 16572 20177 16575
rect 19996 16544 20177 16572
rect 20165 16541 20177 16544
rect 20211 16541 20223 16575
rect 20165 16535 20223 16541
rect 22002 16532 22008 16584
rect 22060 16532 22066 16584
rect 11296 16408 13308 16436
rect 11296 16396 11302 16408
rect 13630 16396 13636 16448
rect 13688 16396 13694 16448
rect 15194 16396 15200 16448
rect 15252 16436 15258 16448
rect 15933 16439 15991 16445
rect 15933 16436 15945 16439
rect 15252 16408 15945 16436
rect 15252 16396 15258 16408
rect 15933 16405 15945 16408
rect 15979 16405 15991 16439
rect 15933 16399 15991 16405
rect 20254 16396 20260 16448
rect 20312 16396 20318 16448
rect 20625 16439 20683 16445
rect 20625 16405 20637 16439
rect 20671 16436 20683 16439
rect 21358 16436 21364 16448
rect 20671 16408 21364 16436
rect 20671 16405 20683 16408
rect 20625 16399 20683 16405
rect 21358 16396 21364 16408
rect 21416 16396 21422 16448
rect 21634 16396 21640 16448
rect 21692 16396 21698 16448
rect 21818 16396 21824 16448
rect 21876 16436 21882 16448
rect 23845 16439 23903 16445
rect 23845 16436 23857 16439
rect 21876 16408 23857 16436
rect 21876 16396 21882 16408
rect 23845 16405 23857 16408
rect 23891 16405 23903 16439
rect 23845 16399 23903 16405
rect 1104 16346 25852 16368
rect 1104 16294 7950 16346
rect 8002 16294 8014 16346
rect 8066 16294 8078 16346
rect 8130 16294 8142 16346
rect 8194 16294 8206 16346
rect 8258 16294 17950 16346
rect 18002 16294 18014 16346
rect 18066 16294 18078 16346
rect 18130 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 25852 16346
rect 1104 16272 25852 16294
rect 6454 16192 6460 16244
rect 6512 16232 6518 16244
rect 7561 16235 7619 16241
rect 7561 16232 7573 16235
rect 6512 16204 7573 16232
rect 6512 16192 6518 16204
rect 7561 16201 7573 16204
rect 7607 16201 7619 16235
rect 7561 16195 7619 16201
rect 7929 16235 7987 16241
rect 7929 16201 7941 16235
rect 7975 16232 7987 16235
rect 9122 16232 9128 16244
rect 7975 16204 9128 16232
rect 7975 16201 7987 16204
rect 7929 16195 7987 16201
rect 9122 16192 9128 16204
rect 9180 16192 9186 16244
rect 10781 16235 10839 16241
rect 10781 16201 10793 16235
rect 10827 16232 10839 16235
rect 12526 16232 12532 16244
rect 10827 16204 12532 16232
rect 10827 16201 10839 16204
rect 10781 16195 10839 16201
rect 12526 16192 12532 16204
rect 12584 16192 12590 16244
rect 16942 16192 16948 16244
rect 17000 16232 17006 16244
rect 17770 16232 17776 16244
rect 17000 16204 17776 16232
rect 17000 16192 17006 16204
rect 17770 16192 17776 16204
rect 17828 16192 17834 16244
rect 9214 16164 9220 16176
rect 9140 16136 9220 16164
rect 1762 16056 1768 16108
rect 1820 16056 1826 16108
rect 7834 16056 7840 16108
rect 7892 16096 7898 16108
rect 9140 16105 9168 16136
rect 9214 16124 9220 16136
rect 9272 16124 9278 16176
rect 16206 16124 16212 16176
rect 16264 16124 16270 16176
rect 19242 16124 19248 16176
rect 19300 16164 19306 16176
rect 20533 16167 20591 16173
rect 20533 16164 20545 16167
rect 19300 16136 20545 16164
rect 19300 16124 19306 16136
rect 20533 16133 20545 16136
rect 20579 16133 20591 16167
rect 20533 16127 20591 16133
rect 9125 16099 9183 16105
rect 7892 16068 8156 16096
rect 7892 16056 7898 16068
rect 1302 15988 1308 16040
rect 1360 16028 1366 16040
rect 8128 16037 8156 16068
rect 9125 16065 9137 16099
rect 9171 16065 9183 16099
rect 9398 16096 9404 16108
rect 9125 16059 9183 16065
rect 9232 16068 9404 16096
rect 2041 16031 2099 16037
rect 2041 16028 2053 16031
rect 1360 16000 2053 16028
rect 1360 15988 1366 16000
rect 2041 15997 2053 16000
rect 2087 15997 2099 16031
rect 2041 15991 2099 15997
rect 8021 16031 8079 16037
rect 8021 15997 8033 16031
rect 8067 15997 8079 16031
rect 8021 15991 8079 15997
rect 8113 16031 8171 16037
rect 8113 15997 8125 16031
rect 8159 15997 8171 16031
rect 8113 15991 8171 15997
rect 8036 15960 8064 15991
rect 8478 15988 8484 16040
rect 8536 16028 8542 16040
rect 9232 16037 9260 16068
rect 9398 16056 9404 16068
rect 9456 16056 9462 16108
rect 11698 16056 11704 16108
rect 11756 16096 11762 16108
rect 12802 16096 12808 16108
rect 11756 16068 12808 16096
rect 11756 16056 11762 16068
rect 12802 16056 12808 16068
rect 12860 16056 12866 16108
rect 15197 16099 15255 16105
rect 15197 16065 15209 16099
rect 15243 16065 15255 16099
rect 15197 16059 15255 16065
rect 9217 16031 9275 16037
rect 9217 16028 9229 16031
rect 8536 16000 9229 16028
rect 8536 15988 8542 16000
rect 9217 15997 9229 16000
rect 9263 15997 9275 16031
rect 9217 15991 9275 15997
rect 9306 15988 9312 16040
rect 9364 15988 9370 16040
rect 10870 15988 10876 16040
rect 10928 15988 10934 16040
rect 10965 16031 11023 16037
rect 10965 15997 10977 16031
rect 11011 15997 11023 16031
rect 10965 15991 11023 15997
rect 10413 15963 10471 15969
rect 10413 15960 10425 15963
rect 8036 15932 10425 15960
rect 10413 15929 10425 15932
rect 10459 15929 10471 15963
rect 10980 15960 11008 15991
rect 10413 15923 10471 15929
rect 10888 15932 11008 15960
rect 8754 15852 8760 15904
rect 8812 15852 8818 15904
rect 8846 15852 8852 15904
rect 8904 15892 8910 15904
rect 10888 15892 10916 15932
rect 8904 15864 10916 15892
rect 8904 15852 8910 15864
rect 14826 15852 14832 15904
rect 14884 15852 14890 15904
rect 15212 15892 15240 16059
rect 19794 16056 19800 16108
rect 19852 16096 19858 16108
rect 21269 16099 21327 16105
rect 21269 16096 21281 16099
rect 19852 16068 21281 16096
rect 19852 16056 19858 16068
rect 21269 16065 21281 16068
rect 21315 16065 21327 16099
rect 21269 16059 21327 16065
rect 23385 16099 23443 16105
rect 23385 16065 23397 16099
rect 23431 16096 23443 16099
rect 23658 16096 23664 16108
rect 23431 16068 23664 16096
rect 23431 16065 23443 16068
rect 23385 16059 23443 16065
rect 23658 16056 23664 16068
rect 23716 16056 23722 16108
rect 23934 16056 23940 16108
rect 23992 16056 23998 16108
rect 24854 16096 24860 16108
rect 24044 16068 24860 16096
rect 15286 15988 15292 16040
rect 15344 15988 15350 16040
rect 15470 15988 15476 16040
rect 15528 15988 15534 16040
rect 19518 15988 19524 16040
rect 19576 15988 19582 16040
rect 21453 16031 21511 16037
rect 21453 15997 21465 16031
rect 21499 16028 21511 16031
rect 23017 16031 23075 16037
rect 21499 16000 22094 16028
rect 21499 15997 21511 16000
rect 21453 15991 21511 15997
rect 16022 15920 16028 15972
rect 16080 15920 16086 15972
rect 16574 15920 16580 15972
rect 16632 15960 16638 15972
rect 17773 15963 17831 15969
rect 17773 15960 17785 15963
rect 16632 15932 17785 15960
rect 16632 15920 16638 15932
rect 17773 15929 17785 15932
rect 17819 15929 17831 15963
rect 17773 15923 17831 15929
rect 20717 15963 20775 15969
rect 20717 15929 20729 15963
rect 20763 15960 20775 15963
rect 22066 15960 22094 16000
rect 23017 15997 23029 16031
rect 23063 16028 23075 16031
rect 24044 16028 24072 16068
rect 24854 16056 24860 16068
rect 24912 16056 24918 16108
rect 23063 16000 24072 16028
rect 23063 15997 23075 16000
rect 23017 15991 23075 15997
rect 24762 15988 24768 16040
rect 24820 15988 24826 16040
rect 23934 15960 23940 15972
rect 20763 15932 21496 15960
rect 22066 15932 23940 15960
rect 20763 15929 20775 15932
rect 20717 15923 20775 15929
rect 16666 15892 16672 15904
rect 15212 15864 16672 15892
rect 16666 15852 16672 15864
rect 16724 15892 16730 15904
rect 16761 15895 16819 15901
rect 16761 15892 16773 15895
rect 16724 15864 16773 15892
rect 16724 15852 16730 15864
rect 16761 15861 16773 15864
rect 16807 15892 16819 15895
rect 19426 15892 19432 15904
rect 16807 15864 19432 15892
rect 16807 15861 16819 15864
rect 16761 15855 16819 15861
rect 19426 15852 19432 15864
rect 19484 15852 19490 15904
rect 19794 15852 19800 15904
rect 19852 15892 19858 15904
rect 19981 15895 20039 15901
rect 19981 15892 19993 15895
rect 19852 15864 19993 15892
rect 19852 15852 19858 15864
rect 19981 15861 19993 15864
rect 20027 15861 20039 15895
rect 21468 15892 21496 15932
rect 23934 15920 23940 15932
rect 23992 15920 23998 15972
rect 23658 15892 23664 15904
rect 21468 15864 23664 15892
rect 19981 15855 20039 15861
rect 23658 15852 23664 15864
rect 23716 15852 23722 15904
rect 1104 15802 25852 15824
rect 1104 15750 2950 15802
rect 3002 15750 3014 15802
rect 3066 15750 3078 15802
rect 3130 15750 3142 15802
rect 3194 15750 3206 15802
rect 3258 15750 12950 15802
rect 13002 15750 13014 15802
rect 13066 15750 13078 15802
rect 13130 15750 13142 15802
rect 13194 15750 13206 15802
rect 13258 15750 22950 15802
rect 23002 15750 23014 15802
rect 23066 15750 23078 15802
rect 23130 15750 23142 15802
rect 23194 15750 23206 15802
rect 23258 15750 25852 15802
rect 1104 15728 25852 15750
rect 6181 15691 6239 15697
rect 6181 15657 6193 15691
rect 6227 15688 6239 15691
rect 6546 15688 6552 15700
rect 6227 15660 6552 15688
rect 6227 15657 6239 15660
rect 6181 15651 6239 15657
rect 6546 15648 6552 15660
rect 6604 15648 6610 15700
rect 7282 15648 7288 15700
rect 7340 15688 7346 15700
rect 9306 15688 9312 15700
rect 7340 15660 9312 15688
rect 7340 15648 7346 15660
rect 9306 15648 9312 15660
rect 9364 15688 9370 15700
rect 10502 15688 10508 15700
rect 9364 15660 10508 15688
rect 9364 15648 9370 15660
rect 10502 15648 10508 15660
rect 10560 15688 10566 15700
rect 11054 15688 11060 15700
rect 10560 15660 11060 15688
rect 10560 15648 10566 15660
rect 11054 15648 11060 15660
rect 11112 15648 11118 15700
rect 11882 15648 11888 15700
rect 11940 15688 11946 15700
rect 11977 15691 12035 15697
rect 11977 15688 11989 15691
rect 11940 15660 11989 15688
rect 11940 15648 11946 15660
rect 11977 15657 11989 15660
rect 12023 15657 12035 15691
rect 11977 15651 12035 15657
rect 12802 15648 12808 15700
rect 12860 15648 12866 15700
rect 17586 15648 17592 15700
rect 17644 15688 17650 15700
rect 17681 15691 17739 15697
rect 17681 15688 17693 15691
rect 17644 15660 17693 15688
rect 17644 15648 17650 15660
rect 17681 15657 17693 15660
rect 17727 15657 17739 15691
rect 21085 15691 21143 15697
rect 21085 15688 21097 15691
rect 17681 15651 17739 15657
rect 19352 15660 21097 15688
rect 7926 15580 7932 15632
rect 7984 15620 7990 15632
rect 8297 15623 8355 15629
rect 8297 15620 8309 15623
rect 7984 15592 8309 15620
rect 7984 15580 7990 15592
rect 8297 15589 8309 15592
rect 8343 15589 8355 15623
rect 8297 15583 8355 15589
rect 10229 15555 10287 15561
rect 10229 15521 10241 15555
rect 10275 15552 10287 15555
rect 10594 15552 10600 15564
rect 10275 15524 10600 15552
rect 10275 15521 10287 15524
rect 10229 15515 10287 15521
rect 10594 15512 10600 15524
rect 10652 15512 10658 15564
rect 11238 15512 11244 15564
rect 11296 15552 11302 15564
rect 12437 15555 12495 15561
rect 12437 15552 12449 15555
rect 11296 15524 12449 15552
rect 11296 15512 11302 15524
rect 12437 15521 12449 15524
rect 12483 15521 12495 15555
rect 12437 15515 12495 15521
rect 15933 15555 15991 15561
rect 15933 15521 15945 15555
rect 15979 15552 15991 15555
rect 16850 15552 16856 15564
rect 15979 15524 16856 15552
rect 15979 15521 15991 15524
rect 15933 15515 15991 15521
rect 16850 15512 16856 15524
rect 16908 15512 16914 15564
rect 17696 15552 17724 15651
rect 18233 15555 18291 15561
rect 18233 15552 18245 15555
rect 17696 15524 18245 15552
rect 18233 15521 18245 15524
rect 18279 15521 18291 15555
rect 18233 15515 18291 15521
rect 18322 15512 18328 15564
rect 18380 15552 18386 15564
rect 18417 15555 18475 15561
rect 18417 15552 18429 15555
rect 18380 15524 18429 15552
rect 18380 15512 18386 15524
rect 18417 15521 18429 15524
rect 18463 15521 18475 15555
rect 18417 15515 18475 15521
rect 7929 15487 7987 15493
rect 7929 15453 7941 15487
rect 7975 15453 7987 15487
rect 7929 15447 7987 15453
rect 6914 15376 6920 15428
rect 6972 15376 6978 15428
rect 7374 15376 7380 15428
rect 7432 15416 7438 15428
rect 7653 15419 7711 15425
rect 7653 15416 7665 15419
rect 7432 15388 7665 15416
rect 7432 15376 7438 15388
rect 7653 15385 7665 15388
rect 7699 15385 7711 15419
rect 7653 15379 7711 15385
rect 6270 15308 6276 15360
rect 6328 15348 6334 15360
rect 6822 15348 6828 15360
rect 6328 15320 6828 15348
rect 6328 15308 6334 15320
rect 6822 15308 6828 15320
rect 6880 15348 6886 15360
rect 7944 15348 7972 15447
rect 14458 15444 14464 15496
rect 14516 15484 14522 15496
rect 14829 15487 14887 15493
rect 14829 15484 14841 15487
rect 14516 15456 14841 15484
rect 14516 15444 14522 15456
rect 14829 15453 14841 15456
rect 14875 15453 14887 15487
rect 14829 15447 14887 15453
rect 17770 15444 17776 15496
rect 17828 15484 17834 15496
rect 19352 15484 19380 15660
rect 21085 15657 21097 15660
rect 21131 15657 21143 15691
rect 21085 15651 21143 15657
rect 19613 15555 19671 15561
rect 19613 15521 19625 15555
rect 19659 15552 19671 15555
rect 19978 15552 19984 15564
rect 19659 15524 19984 15552
rect 19659 15521 19671 15524
rect 19613 15515 19671 15521
rect 19978 15512 19984 15524
rect 20036 15512 20042 15564
rect 20254 15512 20260 15564
rect 20312 15552 20318 15564
rect 20625 15555 20683 15561
rect 20625 15552 20637 15555
rect 20312 15524 20637 15552
rect 20312 15512 20318 15524
rect 20625 15521 20637 15524
rect 20671 15521 20683 15555
rect 20625 15515 20683 15521
rect 21637 15555 21695 15561
rect 21637 15521 21649 15555
rect 21683 15552 21695 15555
rect 23290 15552 23296 15564
rect 21683 15524 23296 15552
rect 21683 15521 21695 15524
rect 21637 15515 21695 15521
rect 23290 15512 23296 15524
rect 23348 15512 23354 15564
rect 23845 15555 23903 15561
rect 23845 15521 23857 15555
rect 23891 15552 23903 15555
rect 24854 15552 24860 15564
rect 23891 15524 24860 15552
rect 23891 15521 23903 15524
rect 23845 15515 23903 15521
rect 24854 15512 24860 15524
rect 24912 15512 24918 15564
rect 19705 15487 19763 15493
rect 19705 15484 19717 15487
rect 17828 15456 19717 15484
rect 17828 15444 17834 15456
rect 19705 15453 19717 15456
rect 19751 15453 19763 15487
rect 19705 15447 19763 15453
rect 19996 15456 20208 15484
rect 9674 15376 9680 15428
rect 9732 15416 9738 15428
rect 10505 15419 10563 15425
rect 10505 15416 10517 15419
rect 9732 15388 10517 15416
rect 9732 15376 9738 15388
rect 10505 15385 10517 15388
rect 10551 15385 10563 15419
rect 10505 15379 10563 15385
rect 11238 15376 11244 15428
rect 11296 15376 11302 15428
rect 16114 15376 16120 15428
rect 16172 15416 16178 15428
rect 16209 15419 16267 15425
rect 16209 15416 16221 15419
rect 16172 15388 16221 15416
rect 16172 15376 16178 15388
rect 16209 15385 16221 15388
rect 16255 15385 16267 15419
rect 16209 15379 16267 15385
rect 16666 15376 16672 15428
rect 16724 15376 16730 15428
rect 17862 15376 17868 15428
rect 17920 15416 17926 15428
rect 19794 15416 19800 15428
rect 17920 15388 19800 15416
rect 17920 15376 17926 15388
rect 19794 15376 19800 15388
rect 19852 15376 19858 15428
rect 6880 15320 7972 15348
rect 14369 15351 14427 15357
rect 6880 15308 6886 15320
rect 14369 15317 14381 15351
rect 14415 15348 14427 15351
rect 14642 15348 14648 15360
rect 14415 15320 14648 15348
rect 14415 15317 14427 15320
rect 14369 15311 14427 15317
rect 14642 15308 14648 15320
rect 14700 15308 14706 15360
rect 18506 15308 18512 15360
rect 18564 15308 18570 15360
rect 18877 15351 18935 15357
rect 18877 15317 18889 15351
rect 18923 15348 18935 15351
rect 19996 15348 20024 15456
rect 20180 15416 20208 15456
rect 20530 15444 20536 15496
rect 20588 15484 20594 15496
rect 21729 15487 21787 15493
rect 21729 15484 21741 15487
rect 20588 15456 21741 15484
rect 20588 15444 20594 15456
rect 21729 15453 21741 15456
rect 21775 15453 21787 15487
rect 21729 15447 21787 15453
rect 21818 15444 21824 15496
rect 21876 15444 21882 15496
rect 22646 15444 22652 15496
rect 22704 15444 22710 15496
rect 22002 15416 22008 15428
rect 20180 15388 22008 15416
rect 22002 15376 22008 15388
rect 22060 15376 22066 15428
rect 18923 15320 20024 15348
rect 20165 15351 20223 15357
rect 18923 15317 18935 15320
rect 18877 15311 18935 15317
rect 20165 15317 20177 15351
rect 20211 15348 20223 15351
rect 20990 15348 20996 15360
rect 20211 15320 20996 15348
rect 20211 15317 20223 15320
rect 20165 15311 20223 15317
rect 20990 15308 20996 15320
rect 21048 15308 21054 15360
rect 22189 15351 22247 15357
rect 22189 15317 22201 15351
rect 22235 15348 22247 15351
rect 23290 15348 23296 15360
rect 22235 15320 23296 15348
rect 22235 15317 22247 15320
rect 22189 15311 22247 15317
rect 23290 15308 23296 15320
rect 23348 15308 23354 15360
rect 1104 15258 25852 15280
rect 1104 15206 7950 15258
rect 8002 15206 8014 15258
rect 8066 15206 8078 15258
rect 8130 15206 8142 15258
rect 8194 15206 8206 15258
rect 8258 15206 17950 15258
rect 18002 15206 18014 15258
rect 18066 15206 18078 15258
rect 18130 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 25852 15258
rect 1104 15184 25852 15206
rect 10870 15104 10876 15156
rect 10928 15144 10934 15156
rect 13081 15147 13139 15153
rect 13081 15144 13093 15147
rect 10928 15116 13093 15144
rect 10928 15104 10934 15116
rect 13081 15113 13093 15116
rect 13127 15113 13139 15147
rect 13081 15107 13139 15113
rect 13449 15147 13507 15153
rect 13449 15113 13461 15147
rect 13495 15144 13507 15147
rect 14826 15144 14832 15156
rect 13495 15116 14832 15144
rect 13495 15113 13507 15116
rect 13449 15107 13507 15113
rect 14826 15104 14832 15116
rect 14884 15104 14890 15156
rect 15286 15104 15292 15156
rect 15344 15144 15350 15156
rect 16206 15144 16212 15156
rect 15344 15116 16212 15144
rect 15344 15104 15350 15116
rect 16206 15104 16212 15116
rect 16264 15144 16270 15156
rect 16264 15116 16988 15144
rect 16264 15104 16270 15116
rect 10965 15079 11023 15085
rect 10965 15076 10977 15079
rect 9890 15048 10977 15076
rect 10965 15045 10977 15048
rect 11011 15076 11023 15079
rect 11238 15076 11244 15088
rect 11011 15048 11244 15076
rect 11011 15045 11023 15048
rect 10965 15039 11023 15045
rect 11238 15036 11244 15048
rect 11296 15036 11302 15088
rect 12250 15036 12256 15088
rect 12308 15036 12314 15088
rect 12529 15079 12587 15085
rect 12529 15045 12541 15079
rect 12575 15076 12587 15079
rect 12802 15076 12808 15088
rect 12575 15048 12808 15076
rect 12575 15045 12587 15048
rect 12529 15039 12587 15045
rect 12802 15036 12808 15048
rect 12860 15036 12866 15088
rect 15930 15036 15936 15088
rect 15988 15076 15994 15088
rect 16117 15079 16175 15085
rect 16117 15076 16129 15079
rect 15988 15048 16129 15076
rect 15988 15036 15994 15048
rect 16117 15045 16129 15048
rect 16163 15076 16175 15079
rect 16669 15079 16727 15085
rect 16669 15076 16681 15079
rect 16163 15048 16681 15076
rect 16163 15045 16175 15048
rect 16117 15039 16175 15045
rect 16669 15045 16681 15048
rect 16715 15045 16727 15079
rect 16960 15076 16988 15116
rect 18506 15104 18512 15156
rect 18564 15104 18570 15156
rect 19518 15104 19524 15156
rect 19576 15104 19582 15156
rect 19889 15147 19947 15153
rect 19889 15113 19901 15147
rect 19935 15144 19947 15147
rect 20346 15144 20352 15156
rect 19935 15116 20352 15144
rect 19935 15113 19947 15116
rect 19889 15107 19947 15113
rect 20346 15104 20352 15116
rect 20404 15104 20410 15156
rect 24578 15144 24584 15156
rect 21468 15116 24584 15144
rect 19429 15079 19487 15085
rect 19429 15076 19441 15079
rect 16960 15048 19441 15076
rect 16669 15039 16727 15045
rect 19429 15045 19441 15048
rect 19475 15045 19487 15079
rect 19429 15039 19487 15045
rect 12268 15008 12296 15036
rect 12434 15008 12440 15020
rect 12268 14980 12440 15008
rect 12434 14968 12440 14980
rect 12492 14968 12498 15020
rect 13541 15011 13599 15017
rect 13541 14977 13553 15011
rect 13587 15008 13599 15011
rect 14918 15008 14924 15020
rect 13587 14980 14924 15008
rect 13587 14977 13599 14980
rect 13541 14971 13599 14977
rect 14918 14968 14924 14980
rect 14976 14968 14982 15020
rect 15102 14968 15108 15020
rect 15160 15008 15166 15020
rect 17405 15011 17463 15017
rect 17405 15008 17417 15011
rect 15160 14980 17417 15008
rect 15160 14968 15166 14980
rect 17405 14977 17417 14980
rect 17451 14977 17463 15011
rect 17405 14971 17463 14977
rect 20533 15011 20591 15017
rect 20533 14977 20545 15011
rect 20579 15008 20591 15011
rect 20622 15008 20628 15020
rect 20579 14980 20628 15008
rect 20579 14977 20591 14980
rect 20533 14971 20591 14977
rect 20622 14968 20628 14980
rect 20680 14968 20686 15020
rect 21468 15017 21496 15116
rect 24578 15104 24584 15116
rect 24636 15104 24642 15156
rect 23293 15079 23351 15085
rect 23293 15045 23305 15079
rect 23339 15076 23351 15079
rect 24854 15076 24860 15088
rect 23339 15048 24860 15076
rect 23339 15045 23351 15048
rect 23293 15039 23351 15045
rect 24854 15036 24860 15048
rect 24912 15036 24918 15088
rect 21453 15011 21511 15017
rect 21453 14977 21465 15011
rect 21499 14977 21511 15011
rect 21453 14971 21511 14977
rect 22094 14968 22100 15020
rect 22152 14968 22158 15020
rect 23750 14968 23756 15020
rect 23808 15008 23814 15020
rect 23937 15011 23995 15017
rect 23937 15008 23949 15011
rect 23808 14980 23949 15008
rect 23808 14968 23814 14980
rect 23937 14977 23949 14980
rect 23983 14977 23995 15011
rect 23937 14971 23995 14977
rect 9858 14900 9864 14952
rect 9916 14940 9922 14952
rect 10321 14943 10379 14949
rect 10321 14940 10333 14943
rect 9916 14912 10333 14940
rect 9916 14900 9922 14912
rect 10321 14909 10333 14912
rect 10367 14940 10379 14943
rect 10367 14912 10548 14940
rect 10367 14909 10379 14912
rect 10321 14903 10379 14909
rect 10520 14872 10548 14912
rect 10594 14900 10600 14952
rect 10652 14940 10658 14952
rect 12250 14940 12256 14952
rect 10652 14912 12256 14940
rect 10652 14900 10658 14912
rect 12250 14900 12256 14912
rect 12308 14900 12314 14952
rect 13630 14900 13636 14952
rect 13688 14900 13694 14952
rect 17126 14900 17132 14952
rect 17184 14900 17190 14952
rect 17313 14943 17371 14949
rect 17313 14909 17325 14943
rect 17359 14940 17371 14943
rect 18049 14943 18107 14949
rect 18049 14940 18061 14943
rect 17359 14912 18061 14940
rect 17359 14909 17371 14912
rect 17313 14903 17371 14909
rect 18049 14909 18061 14912
rect 18095 14909 18107 14943
rect 18049 14903 18107 14909
rect 19337 14943 19395 14949
rect 19337 14909 19349 14943
rect 19383 14909 19395 14943
rect 22830 14940 22836 14952
rect 19337 14903 19395 14909
rect 22066 14912 22836 14940
rect 10520 14844 11008 14872
rect 8846 14764 8852 14816
rect 8904 14764 8910 14816
rect 10980 14804 11008 14844
rect 11054 14832 11060 14884
rect 11112 14872 11118 14884
rect 12345 14875 12403 14881
rect 12345 14872 12357 14875
rect 11112 14844 12357 14872
rect 11112 14832 11118 14844
rect 12345 14841 12357 14844
rect 12391 14841 12403 14875
rect 12345 14835 12403 14841
rect 13648 14804 13676 14900
rect 16301 14875 16359 14881
rect 16301 14841 16313 14875
rect 16347 14872 16359 14875
rect 16390 14872 16396 14884
rect 16347 14844 16396 14872
rect 16347 14841 16359 14844
rect 16301 14835 16359 14841
rect 16390 14832 16396 14844
rect 16448 14832 16454 14884
rect 16482 14832 16488 14884
rect 16540 14872 16546 14884
rect 17328 14872 17356 14903
rect 16540 14844 17356 14872
rect 17773 14875 17831 14881
rect 16540 14832 16546 14844
rect 17773 14841 17785 14875
rect 17819 14872 17831 14875
rect 18414 14872 18420 14884
rect 17819 14844 18420 14872
rect 17819 14841 17831 14844
rect 17773 14835 17831 14841
rect 18414 14832 18420 14844
rect 18472 14832 18478 14884
rect 19352 14872 19380 14903
rect 22066 14872 22094 14912
rect 22830 14900 22836 14912
rect 22888 14900 22894 14952
rect 24670 14900 24676 14952
rect 24728 14900 24734 14952
rect 19352 14844 22094 14872
rect 10980 14776 13676 14804
rect 15930 14764 15936 14816
rect 15988 14804 15994 14816
rect 16500 14804 16528 14832
rect 15988 14776 16528 14804
rect 15988 14764 15994 14776
rect 20346 14764 20352 14816
rect 20404 14764 20410 14816
rect 21266 14764 21272 14816
rect 21324 14764 21330 14816
rect 1104 14714 25852 14736
rect 1104 14662 2950 14714
rect 3002 14662 3014 14714
rect 3066 14662 3078 14714
rect 3130 14662 3142 14714
rect 3194 14662 3206 14714
rect 3258 14662 12950 14714
rect 13002 14662 13014 14714
rect 13066 14662 13078 14714
rect 13130 14662 13142 14714
rect 13194 14662 13206 14714
rect 13258 14662 22950 14714
rect 23002 14662 23014 14714
rect 23066 14662 23078 14714
rect 23130 14662 23142 14714
rect 23194 14662 23206 14714
rect 23258 14662 25852 14714
rect 1104 14640 25852 14662
rect 9217 14603 9275 14609
rect 9217 14569 9229 14603
rect 9263 14600 9275 14603
rect 9582 14600 9588 14612
rect 9263 14572 9588 14600
rect 9263 14569 9275 14572
rect 9217 14563 9275 14569
rect 9582 14560 9588 14572
rect 9640 14560 9646 14612
rect 10502 14560 10508 14612
rect 10560 14600 10566 14612
rect 11330 14600 11336 14612
rect 10560 14572 11336 14600
rect 10560 14560 10566 14572
rect 11330 14560 11336 14572
rect 11388 14560 11394 14612
rect 11606 14560 11612 14612
rect 11664 14600 11670 14612
rect 12805 14603 12863 14609
rect 12805 14600 12817 14603
rect 11664 14572 12817 14600
rect 11664 14560 11670 14572
rect 12805 14569 12817 14572
rect 12851 14569 12863 14603
rect 12805 14563 12863 14569
rect 15013 14603 15071 14609
rect 15013 14569 15025 14603
rect 15059 14600 15071 14603
rect 16114 14600 16120 14612
rect 15059 14572 16120 14600
rect 15059 14569 15071 14572
rect 15013 14563 15071 14569
rect 16114 14560 16120 14572
rect 16172 14560 16178 14612
rect 18046 14560 18052 14612
rect 18104 14600 18110 14612
rect 18785 14603 18843 14609
rect 18785 14600 18797 14603
rect 18104 14572 18797 14600
rect 18104 14560 18110 14572
rect 18785 14569 18797 14572
rect 18831 14600 18843 14603
rect 19150 14600 19156 14612
rect 18831 14572 19156 14600
rect 18831 14569 18843 14572
rect 18785 14563 18843 14569
rect 19150 14560 19156 14572
rect 19208 14560 19214 14612
rect 15102 14532 15108 14544
rect 13280 14504 15108 14532
rect 8297 14467 8355 14473
rect 8297 14433 8309 14467
rect 8343 14464 8355 14467
rect 8846 14464 8852 14476
rect 8343 14436 8852 14464
rect 8343 14433 8355 14436
rect 8297 14427 8355 14433
rect 8846 14424 8852 14436
rect 8904 14424 8910 14476
rect 9030 14424 9036 14476
rect 9088 14464 9094 14476
rect 9677 14467 9735 14473
rect 9677 14464 9689 14467
rect 9088 14436 9689 14464
rect 9088 14424 9094 14436
rect 9677 14433 9689 14436
rect 9723 14433 9735 14467
rect 9677 14427 9735 14433
rect 9858 14424 9864 14476
rect 9916 14424 9922 14476
rect 10962 14424 10968 14476
rect 11020 14464 11026 14476
rect 11977 14467 12035 14473
rect 11977 14464 11989 14467
rect 11020 14436 11989 14464
rect 11020 14424 11026 14436
rect 11977 14433 11989 14436
rect 12023 14464 12035 14467
rect 12023 14436 12434 14464
rect 12023 14433 12035 14436
rect 11977 14427 12035 14433
rect 6914 14356 6920 14408
rect 6972 14396 6978 14408
rect 7190 14396 7196 14408
rect 6972 14368 7196 14396
rect 6972 14356 6978 14368
rect 7190 14356 7196 14368
rect 7248 14356 7254 14408
rect 8570 14356 8576 14408
rect 8628 14356 8634 14408
rect 12250 14356 12256 14408
rect 12308 14356 12314 14408
rect 11238 14288 11244 14340
rect 11296 14288 11302 14340
rect 12406 14328 12434 14436
rect 13170 14424 13176 14476
rect 13228 14464 13234 14476
rect 13280 14473 13308 14504
rect 15102 14492 15108 14504
rect 15160 14492 15166 14544
rect 13265 14467 13323 14473
rect 13265 14464 13277 14467
rect 13228 14436 13277 14464
rect 13228 14424 13234 14436
rect 13265 14433 13277 14436
rect 13311 14433 13323 14467
rect 13265 14427 13323 14433
rect 13354 14424 13360 14476
rect 13412 14424 13418 14476
rect 19794 14464 19800 14476
rect 15212 14436 19800 14464
rect 13998 14328 14004 14340
rect 12406 14300 14004 14328
rect 13998 14288 14004 14300
rect 14056 14328 14062 14340
rect 15102 14328 15108 14340
rect 14056 14300 15108 14328
rect 14056 14288 14062 14300
rect 15102 14288 15108 14300
rect 15160 14288 15166 14340
rect 6825 14263 6883 14269
rect 6825 14229 6837 14263
rect 6871 14260 6883 14263
rect 6914 14260 6920 14272
rect 6871 14232 6920 14260
rect 6871 14229 6883 14232
rect 6825 14223 6883 14229
rect 6914 14220 6920 14232
rect 6972 14220 6978 14272
rect 9030 14220 9036 14272
rect 9088 14260 9094 14272
rect 9585 14263 9643 14269
rect 9585 14260 9597 14263
rect 9088 14232 9597 14260
rect 9088 14220 9094 14232
rect 9585 14229 9597 14232
rect 9631 14229 9643 14263
rect 9585 14223 9643 14229
rect 13078 14220 13084 14272
rect 13136 14260 13142 14272
rect 13173 14263 13231 14269
rect 13173 14260 13185 14263
rect 13136 14232 13185 14260
rect 13136 14220 13142 14232
rect 13173 14229 13185 14232
rect 13219 14260 13231 14263
rect 14734 14260 14740 14272
rect 13219 14232 14740 14260
rect 13219 14229 13231 14232
rect 13173 14223 13231 14229
rect 14734 14220 14740 14232
rect 14792 14260 14798 14272
rect 15212 14260 15240 14436
rect 19794 14424 19800 14436
rect 19852 14424 19858 14476
rect 16761 14399 16819 14405
rect 16761 14365 16773 14399
rect 16807 14396 16819 14399
rect 16850 14396 16856 14408
rect 16807 14368 16856 14396
rect 16807 14365 16819 14368
rect 16761 14359 16819 14365
rect 16850 14356 16856 14368
rect 16908 14356 16914 14408
rect 17494 14356 17500 14408
rect 17552 14356 17558 14408
rect 18046 14356 18052 14408
rect 18104 14356 18110 14408
rect 21450 14356 21456 14408
rect 21508 14396 21514 14408
rect 23109 14399 23167 14405
rect 23109 14396 23121 14399
rect 21508 14368 23121 14396
rect 21508 14356 21514 14368
rect 23109 14365 23121 14368
rect 23155 14365 23167 14399
rect 23109 14359 23167 14365
rect 16054 14300 16436 14328
rect 14792 14232 15240 14260
rect 16408 14260 16436 14300
rect 16482 14288 16488 14340
rect 16540 14288 16546 14340
rect 18233 14331 18291 14337
rect 18233 14297 18245 14331
rect 18279 14328 18291 14331
rect 18966 14328 18972 14340
rect 18279 14300 18972 14328
rect 18279 14297 18291 14300
rect 18233 14291 18291 14297
rect 18966 14288 18972 14300
rect 19024 14288 19030 14340
rect 21726 14288 21732 14340
rect 21784 14328 21790 14340
rect 22922 14328 22928 14340
rect 21784 14300 22928 14328
rect 21784 14288 21790 14300
rect 22922 14288 22928 14300
rect 22980 14288 22986 14340
rect 16574 14260 16580 14272
rect 16408 14232 16580 14260
rect 14792 14220 14798 14232
rect 16574 14220 16580 14232
rect 16632 14220 16638 14272
rect 17310 14220 17316 14272
rect 17368 14220 17374 14272
rect 17586 14220 17592 14272
rect 17644 14260 17650 14272
rect 18509 14263 18567 14269
rect 18509 14260 18521 14263
rect 17644 14232 18521 14260
rect 17644 14220 17650 14232
rect 18509 14229 18521 14232
rect 18555 14260 18567 14263
rect 18877 14263 18935 14269
rect 18877 14260 18889 14263
rect 18555 14232 18889 14260
rect 18555 14229 18567 14232
rect 18509 14223 18567 14229
rect 18877 14229 18889 14232
rect 18923 14229 18935 14263
rect 18877 14223 18935 14229
rect 22554 14220 22560 14272
rect 22612 14260 22618 14272
rect 23293 14263 23351 14269
rect 23293 14260 23305 14263
rect 22612 14232 23305 14260
rect 22612 14220 22618 14232
rect 23293 14229 23305 14232
rect 23339 14229 23351 14263
rect 23293 14223 23351 14229
rect 1104 14170 25852 14192
rect 1104 14118 7950 14170
rect 8002 14118 8014 14170
rect 8066 14118 8078 14170
rect 8130 14118 8142 14170
rect 8194 14118 8206 14170
rect 8258 14118 17950 14170
rect 18002 14118 18014 14170
rect 18066 14118 18078 14170
rect 18130 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 25852 14170
rect 1104 14096 25852 14118
rect 7190 14016 7196 14068
rect 7248 14056 7254 14068
rect 8478 14056 8484 14068
rect 7248 14028 8484 14056
rect 7248 14016 7254 14028
rect 8478 14016 8484 14028
rect 8536 14016 8542 14068
rect 10778 14016 10784 14068
rect 10836 14056 10842 14068
rect 10836 14028 12434 14056
rect 10836 14016 10842 14028
rect 10873 13991 10931 13997
rect 10873 13957 10885 13991
rect 10919 13988 10931 13991
rect 10962 13988 10968 14000
rect 10919 13960 10968 13988
rect 10919 13957 10931 13960
rect 10873 13951 10931 13957
rect 10962 13948 10968 13960
rect 11020 13948 11026 14000
rect 11238 13948 11244 14000
rect 11296 13948 11302 14000
rect 12406 13988 12434 14028
rect 12710 14016 12716 14068
rect 12768 14016 12774 14068
rect 13078 14016 13084 14068
rect 13136 14016 13142 14068
rect 13170 14016 13176 14068
rect 13228 14016 13234 14068
rect 14645 14059 14703 14065
rect 14645 14025 14657 14059
rect 14691 14056 14703 14059
rect 17034 14056 17040 14068
rect 14691 14028 17040 14056
rect 14691 14025 14703 14028
rect 14645 14019 14703 14025
rect 17034 14016 17040 14028
rect 17092 14016 17098 14068
rect 18598 14016 18604 14068
rect 18656 14016 18662 14068
rect 20990 14016 20996 14068
rect 21048 14016 21054 14068
rect 21453 14059 21511 14065
rect 21453 14025 21465 14059
rect 21499 14056 21511 14059
rect 21910 14056 21916 14068
rect 21499 14028 21916 14056
rect 21499 14025 21511 14028
rect 21453 14019 21511 14025
rect 21910 14016 21916 14028
rect 21968 14016 21974 14068
rect 22189 14059 22247 14065
rect 22189 14025 22201 14059
rect 22235 14056 22247 14059
rect 22738 14056 22744 14068
rect 22235 14028 22744 14056
rect 22235 14025 22247 14028
rect 22189 14019 22247 14025
rect 22738 14016 22744 14028
rect 22796 14016 22802 14068
rect 14277 13991 14335 13997
rect 14277 13988 14289 13991
rect 12406 13960 14289 13988
rect 14277 13957 14289 13960
rect 14323 13957 14335 13991
rect 14277 13951 14335 13957
rect 15289 13991 15347 13997
rect 15289 13957 15301 13991
rect 15335 13988 15347 13991
rect 16022 13988 16028 14000
rect 15335 13960 16028 13988
rect 15335 13957 15347 13960
rect 15289 13951 15347 13957
rect 16022 13948 16028 13960
rect 16080 13948 16086 14000
rect 16298 13948 16304 14000
rect 16356 13988 16362 14000
rect 16574 13988 16580 14000
rect 16356 13960 16580 13988
rect 16356 13948 16362 13960
rect 16574 13948 16580 13960
rect 16632 13988 16638 14000
rect 17586 13988 17592 14000
rect 16632 13960 17592 13988
rect 16632 13948 16638 13960
rect 17586 13948 17592 13960
rect 17644 13948 17650 14000
rect 19702 13948 19708 14000
rect 19760 13988 19766 14000
rect 19889 13991 19947 13997
rect 19889 13988 19901 13991
rect 19760 13960 19901 13988
rect 19760 13948 19766 13960
rect 19889 13957 19901 13960
rect 19935 13988 19947 13991
rect 20349 13991 20407 13997
rect 20349 13988 20361 13991
rect 19935 13960 20361 13988
rect 19935 13957 19947 13960
rect 19889 13951 19947 13957
rect 20349 13957 20361 13960
rect 20395 13957 20407 13991
rect 20349 13951 20407 13957
rect 21085 13991 21143 13997
rect 21085 13957 21097 13991
rect 21131 13988 21143 13991
rect 22830 13988 22836 14000
rect 21131 13960 22836 13988
rect 21131 13957 21143 13960
rect 21085 13951 21143 13957
rect 22830 13948 22836 13960
rect 22888 13948 22894 14000
rect 25130 13948 25136 14000
rect 25188 13948 25194 14000
rect 2774 13880 2780 13932
rect 2832 13880 2838 13932
rect 11256 13920 11284 13948
rect 12345 13923 12403 13929
rect 12345 13920 12357 13923
rect 10258 13892 12357 13920
rect 12345 13889 12357 13892
rect 12391 13889 12403 13923
rect 12345 13883 12403 13889
rect 14185 13923 14243 13929
rect 14185 13889 14197 13923
rect 14231 13920 14243 13923
rect 20073 13923 20131 13929
rect 14231 13892 15884 13920
rect 14231 13889 14243 13892
rect 14185 13883 14243 13889
rect 1762 13812 1768 13864
rect 1820 13812 1826 13864
rect 6822 13812 6828 13864
rect 6880 13852 6886 13864
rect 8570 13852 8576 13864
rect 6880 13824 8576 13852
rect 6880 13812 6886 13824
rect 8570 13812 8576 13824
rect 8628 13852 8634 13864
rect 8849 13855 8907 13861
rect 8849 13852 8861 13855
rect 8628 13824 8861 13852
rect 8628 13812 8634 13824
rect 8849 13821 8861 13824
rect 8895 13821 8907 13855
rect 9125 13855 9183 13861
rect 9125 13852 9137 13855
rect 8849 13815 8907 13821
rect 8956 13824 9137 13852
rect 6914 13744 6920 13796
rect 6972 13784 6978 13796
rect 7834 13784 7840 13796
rect 6972 13756 7840 13784
rect 6972 13744 6978 13756
rect 7834 13744 7840 13756
rect 7892 13784 7898 13796
rect 8956 13784 8984 13824
rect 9125 13821 9137 13824
rect 9171 13821 9183 13855
rect 9125 13815 9183 13821
rect 12158 13812 12164 13864
rect 12216 13852 12222 13864
rect 13170 13852 13176 13864
rect 12216 13824 13176 13852
rect 12216 13812 12222 13824
rect 13170 13812 13176 13824
rect 13228 13812 13234 13864
rect 13265 13855 13323 13861
rect 13265 13821 13277 13855
rect 13311 13821 13323 13855
rect 13265 13815 13323 13821
rect 14093 13855 14151 13861
rect 14093 13821 14105 13855
rect 14139 13821 14151 13855
rect 14093 13815 14151 13821
rect 15473 13855 15531 13861
rect 15473 13821 15485 13855
rect 15519 13852 15531 13855
rect 15746 13852 15752 13864
rect 15519 13824 15752 13852
rect 15519 13821 15531 13824
rect 15473 13815 15531 13821
rect 7892 13756 8984 13784
rect 7892 13744 7898 13756
rect 12526 13744 12532 13796
rect 12584 13784 12590 13796
rect 13280 13784 13308 13815
rect 12584 13756 13308 13784
rect 14108 13784 14136 13815
rect 15746 13812 15752 13824
rect 15804 13812 15810 13864
rect 15856 13861 15884 13892
rect 20073 13889 20085 13923
rect 20119 13920 20131 13923
rect 21818 13920 21824 13932
rect 20119 13892 21824 13920
rect 20119 13889 20131 13892
rect 20073 13883 20131 13889
rect 21818 13880 21824 13892
rect 21876 13880 21882 13932
rect 22002 13880 22008 13932
rect 22060 13880 22066 13932
rect 22649 13923 22707 13929
rect 22649 13889 22661 13923
rect 22695 13889 22707 13923
rect 22649 13883 22707 13889
rect 15841 13855 15899 13861
rect 15841 13821 15853 13855
rect 15887 13852 15899 13855
rect 15930 13852 15936 13864
rect 15887 13824 15936 13852
rect 15887 13821 15899 13824
rect 15841 13815 15899 13821
rect 15930 13812 15936 13824
rect 15988 13812 15994 13864
rect 16850 13812 16856 13864
rect 16908 13812 16914 13864
rect 17126 13812 17132 13864
rect 17184 13812 17190 13864
rect 19058 13812 19064 13864
rect 19116 13812 19122 13864
rect 20809 13855 20867 13861
rect 20809 13821 20821 13855
rect 20855 13821 20867 13855
rect 20809 13815 20867 13821
rect 14458 13784 14464 13796
rect 14108 13756 14464 13784
rect 12584 13744 12590 13756
rect 14458 13744 14464 13756
rect 14516 13744 14522 13796
rect 20824 13784 20852 13815
rect 21358 13812 21364 13864
rect 21416 13852 21422 13864
rect 22664 13852 22692 13883
rect 22922 13880 22928 13932
rect 22980 13920 22986 13932
rect 23937 13923 23995 13929
rect 23937 13920 23949 13923
rect 22980 13892 23949 13920
rect 22980 13880 22986 13892
rect 23937 13889 23949 13892
rect 23983 13889 23995 13923
rect 23937 13883 23995 13889
rect 23382 13852 23388 13864
rect 21416 13824 22692 13852
rect 22848 13824 23388 13852
rect 21416 13812 21422 13824
rect 20898 13784 20904 13796
rect 20824 13756 20904 13784
rect 20898 13744 20904 13756
rect 20956 13744 20962 13796
rect 22848 13793 22876 13824
rect 23382 13812 23388 13824
rect 23440 13812 23446 13864
rect 22833 13787 22891 13793
rect 22833 13753 22845 13787
rect 22879 13753 22891 13787
rect 22833 13747 22891 13753
rect 16022 13676 16028 13728
rect 16080 13716 16086 13728
rect 17862 13716 17868 13728
rect 16080 13688 17868 13716
rect 16080 13676 16086 13688
rect 17862 13676 17868 13688
rect 17920 13676 17926 13728
rect 21358 13676 21364 13728
rect 21416 13716 21422 13728
rect 21726 13716 21732 13728
rect 21416 13688 21732 13716
rect 21416 13676 21422 13688
rect 21726 13676 21732 13688
rect 21784 13716 21790 13728
rect 23109 13719 23167 13725
rect 23109 13716 23121 13719
rect 21784 13688 23121 13716
rect 21784 13676 21790 13688
rect 23109 13685 23121 13688
rect 23155 13685 23167 13719
rect 23109 13679 23167 13685
rect 1104 13626 25852 13648
rect 1104 13574 2950 13626
rect 3002 13574 3014 13626
rect 3066 13574 3078 13626
rect 3130 13574 3142 13626
rect 3194 13574 3206 13626
rect 3258 13574 12950 13626
rect 13002 13574 13014 13626
rect 13066 13574 13078 13626
rect 13130 13574 13142 13626
rect 13194 13574 13206 13626
rect 13258 13574 22950 13626
rect 23002 13574 23014 13626
rect 23066 13574 23078 13626
rect 23130 13574 23142 13626
rect 23194 13574 23206 13626
rect 23258 13574 25852 13626
rect 1104 13552 25852 13574
rect 8478 13472 8484 13524
rect 8536 13512 8542 13524
rect 8941 13515 8999 13521
rect 8941 13512 8953 13515
rect 8536 13484 8953 13512
rect 8536 13472 8542 13484
rect 8941 13481 8953 13484
rect 8987 13481 8999 13515
rect 8941 13475 8999 13481
rect 12434 13472 12440 13524
rect 12492 13512 12498 13524
rect 13538 13512 13544 13524
rect 12492 13484 13544 13512
rect 12492 13472 12498 13484
rect 13538 13472 13544 13484
rect 13596 13512 13602 13524
rect 13817 13515 13875 13521
rect 13817 13512 13829 13515
rect 13596 13484 13829 13512
rect 13596 13472 13602 13484
rect 13817 13481 13829 13484
rect 13863 13481 13875 13515
rect 13817 13475 13875 13481
rect 14182 13472 14188 13524
rect 14240 13512 14246 13524
rect 14734 13512 14740 13524
rect 14240 13484 14740 13512
rect 14240 13472 14246 13484
rect 14734 13472 14740 13484
rect 14792 13472 14798 13524
rect 15473 13515 15531 13521
rect 15473 13481 15485 13515
rect 15519 13512 15531 13515
rect 15562 13512 15568 13524
rect 15519 13484 15568 13512
rect 15519 13481 15531 13484
rect 15473 13475 15531 13481
rect 12805 13447 12863 13453
rect 12805 13413 12817 13447
rect 12851 13444 12863 13447
rect 14550 13444 14556 13456
rect 12851 13416 14556 13444
rect 12851 13413 12863 13416
rect 12805 13407 12863 13413
rect 14550 13404 14556 13416
rect 14608 13404 14614 13456
rect 7098 13336 7104 13388
rect 7156 13376 7162 13388
rect 7650 13376 7656 13388
rect 7156 13348 7656 13376
rect 7156 13336 7162 13348
rect 7650 13336 7656 13348
rect 7708 13336 7714 13388
rect 12253 13379 12311 13385
rect 12253 13345 12265 13379
rect 12299 13376 12311 13379
rect 12434 13376 12440 13388
rect 12299 13348 12440 13376
rect 12299 13345 12311 13348
rect 12253 13339 12311 13345
rect 12434 13336 12440 13348
rect 12492 13336 12498 13388
rect 13173 13379 13231 13385
rect 13173 13345 13185 13379
rect 13219 13376 13231 13379
rect 14090 13376 14096 13388
rect 13219 13348 14096 13376
rect 13219 13345 13231 13348
rect 13173 13339 13231 13345
rect 6822 13268 6828 13320
rect 6880 13268 6886 13320
rect 8478 13240 8484 13252
rect 8326 13212 8484 13240
rect 8478 13200 8484 13212
rect 8536 13200 8542 13252
rect 9030 13200 9036 13252
rect 9088 13240 9094 13252
rect 12437 13243 12495 13249
rect 12437 13240 12449 13243
rect 9088 13212 12449 13240
rect 9088 13200 9094 13212
rect 12437 13209 12449 13212
rect 12483 13209 12495 13243
rect 12437 13203 12495 13209
rect 8570 13132 8576 13184
rect 8628 13132 8634 13184
rect 12345 13175 12403 13181
rect 12345 13141 12357 13175
rect 12391 13172 12403 13175
rect 13188 13172 13216 13339
rect 14090 13336 14096 13348
rect 14148 13336 14154 13388
rect 14921 13311 14979 13317
rect 14921 13277 14933 13311
rect 14967 13308 14979 13311
rect 15488 13308 15516 13475
rect 15562 13472 15568 13484
rect 15620 13472 15626 13524
rect 18877 13515 18935 13521
rect 18877 13481 18889 13515
rect 18923 13512 18935 13515
rect 21082 13512 21088 13524
rect 18923 13484 21088 13512
rect 18923 13481 18935 13484
rect 18877 13475 18935 13481
rect 21082 13472 21088 13484
rect 21140 13472 21146 13524
rect 18598 13444 18604 13456
rect 18340 13416 18604 13444
rect 18340 13385 18368 13416
rect 18598 13404 18604 13416
rect 18656 13404 18662 13456
rect 19334 13404 19340 13456
rect 19392 13404 19398 13456
rect 19889 13447 19947 13453
rect 19889 13413 19901 13447
rect 19935 13444 19947 13447
rect 21174 13444 21180 13456
rect 19935 13416 21180 13444
rect 19935 13413 19947 13416
rect 19889 13407 19947 13413
rect 21174 13404 21180 13416
rect 21232 13404 21238 13456
rect 18325 13379 18383 13385
rect 18325 13345 18337 13379
rect 18371 13345 18383 13379
rect 18325 13339 18383 13345
rect 18414 13336 18420 13388
rect 18472 13336 18478 13388
rect 21542 13336 21548 13388
rect 21600 13376 21606 13388
rect 22557 13379 22615 13385
rect 22557 13376 22569 13379
rect 21600 13348 22569 13376
rect 21600 13336 21606 13348
rect 22557 13345 22569 13348
rect 22603 13345 22615 13379
rect 22557 13339 22615 13345
rect 22830 13336 22836 13388
rect 22888 13376 22894 13388
rect 23017 13379 23075 13385
rect 23017 13376 23029 13379
rect 22888 13348 23029 13376
rect 22888 13336 22894 13348
rect 23017 13345 23029 13348
rect 23063 13345 23075 13379
rect 23017 13339 23075 13345
rect 14967 13280 15516 13308
rect 18509 13311 18567 13317
rect 14967 13277 14979 13280
rect 14921 13271 14979 13277
rect 18509 13277 18521 13311
rect 18555 13308 18567 13311
rect 19058 13308 19064 13320
rect 18555 13280 19064 13308
rect 18555 13277 18567 13280
rect 18509 13271 18567 13277
rect 19058 13268 19064 13280
rect 19116 13268 19122 13320
rect 19610 13268 19616 13320
rect 19668 13308 19674 13320
rect 19705 13311 19763 13317
rect 19705 13308 19717 13311
rect 19668 13280 19717 13308
rect 19668 13268 19674 13280
rect 19705 13277 19717 13280
rect 19751 13308 19763 13311
rect 20165 13311 20223 13317
rect 20165 13308 20177 13311
rect 19751 13280 20177 13308
rect 19751 13277 19763 13280
rect 19705 13271 19763 13277
rect 20165 13277 20177 13280
rect 20211 13277 20223 13311
rect 20165 13271 20223 13277
rect 17497 13243 17555 13249
rect 17497 13209 17509 13243
rect 17543 13240 17555 13243
rect 19334 13240 19340 13252
rect 17543 13212 19340 13240
rect 17543 13209 17555 13212
rect 17497 13203 17555 13209
rect 19334 13200 19340 13212
rect 19392 13200 19398 13252
rect 12391 13144 13216 13172
rect 12391 13141 12403 13144
rect 12345 13135 12403 13141
rect 15010 13132 15016 13184
rect 15068 13132 15074 13184
rect 16853 13175 16911 13181
rect 16853 13141 16865 13175
rect 16899 13172 16911 13175
rect 17218 13172 17224 13184
rect 16899 13144 17224 13172
rect 16899 13141 16911 13144
rect 16853 13135 16911 13141
rect 17218 13132 17224 13144
rect 17276 13132 17282 13184
rect 17589 13175 17647 13181
rect 17589 13141 17601 13175
rect 17635 13172 17647 13175
rect 18506 13172 18512 13184
rect 17635 13144 18512 13172
rect 17635 13141 17647 13144
rect 17589 13135 17647 13141
rect 18506 13132 18512 13144
rect 18564 13132 18570 13184
rect 20809 13175 20867 13181
rect 20809 13141 20821 13175
rect 20855 13172 20867 13175
rect 20898 13172 20904 13184
rect 20855 13144 20904 13172
rect 20855 13141 20867 13144
rect 20809 13135 20867 13141
rect 20898 13132 20904 13144
rect 20956 13132 20962 13184
rect 21192 13172 21220 13294
rect 23290 13268 23296 13320
rect 23348 13308 23354 13320
rect 23661 13311 23719 13317
rect 23661 13308 23673 13311
rect 23348 13280 23673 13308
rect 23348 13268 23354 13280
rect 23661 13277 23673 13280
rect 23707 13277 23719 13311
rect 23661 13271 23719 13277
rect 22281 13243 22339 13249
rect 22281 13209 22293 13243
rect 22327 13209 22339 13243
rect 22281 13203 22339 13209
rect 21358 13172 21364 13184
rect 21192 13144 21364 13172
rect 21358 13132 21364 13144
rect 21416 13132 21422 13184
rect 21634 13132 21640 13184
rect 21692 13172 21698 13184
rect 22296 13172 22324 13203
rect 21692 13144 22324 13172
rect 21692 13132 21698 13144
rect 23842 13132 23848 13184
rect 23900 13132 23906 13184
rect 1104 13082 25852 13104
rect 1104 13030 7950 13082
rect 8002 13030 8014 13082
rect 8066 13030 8078 13082
rect 8130 13030 8142 13082
rect 8194 13030 8206 13082
rect 8258 13030 17950 13082
rect 18002 13030 18014 13082
rect 18066 13030 18078 13082
rect 18130 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 25852 13082
rect 1104 13008 25852 13030
rect 8294 12928 8300 12980
rect 8352 12968 8358 12980
rect 9125 12971 9183 12977
rect 9125 12968 9137 12971
rect 8352 12940 9137 12968
rect 8352 12928 8358 12940
rect 9125 12937 9137 12940
rect 9171 12937 9183 12971
rect 9125 12931 9183 12937
rect 11790 12928 11796 12980
rect 11848 12928 11854 12980
rect 12802 12928 12808 12980
rect 12860 12968 12866 12980
rect 13173 12971 13231 12977
rect 13173 12968 13185 12971
rect 12860 12940 13185 12968
rect 12860 12928 12866 12940
rect 13173 12937 13185 12940
rect 13219 12968 13231 12971
rect 13446 12968 13452 12980
rect 13219 12940 13452 12968
rect 13219 12937 13231 12940
rect 13173 12931 13231 12937
rect 13446 12928 13452 12940
rect 13504 12928 13510 12980
rect 16850 12968 16856 12980
rect 14200 12940 16856 12968
rect 7558 12860 7564 12912
rect 7616 12900 7622 12912
rect 8478 12900 8484 12912
rect 7616 12872 8484 12900
rect 7616 12860 7622 12872
rect 8478 12860 8484 12872
rect 8536 12900 8542 12912
rect 9582 12900 9588 12912
rect 8536 12872 9588 12900
rect 8536 12860 8542 12872
rect 9582 12860 9588 12872
rect 9640 12860 9646 12912
rect 12253 12903 12311 12909
rect 12253 12869 12265 12903
rect 12299 12900 12311 12903
rect 13998 12900 14004 12912
rect 12299 12872 14004 12900
rect 12299 12869 12311 12872
rect 12253 12863 12311 12869
rect 13998 12860 14004 12872
rect 14056 12860 14062 12912
rect 7282 12792 7288 12844
rect 7340 12832 7346 12844
rect 9217 12835 9275 12841
rect 9217 12832 9229 12835
rect 7340 12804 9229 12832
rect 7340 12792 7346 12804
rect 9217 12801 9229 12804
rect 9263 12801 9275 12835
rect 9217 12795 9275 12801
rect 12161 12835 12219 12841
rect 12161 12801 12173 12835
rect 12207 12832 12219 12835
rect 13446 12832 13452 12844
rect 12207 12804 13452 12832
rect 12207 12801 12219 12804
rect 12161 12795 12219 12801
rect 13446 12792 13452 12804
rect 13504 12792 13510 12844
rect 13538 12792 13544 12844
rect 13596 12792 13602 12844
rect 14200 12841 14228 12940
rect 16850 12928 16856 12940
rect 16908 12928 16914 12980
rect 17034 12928 17040 12980
rect 17092 12968 17098 12980
rect 17129 12971 17187 12977
rect 17129 12968 17141 12971
rect 17092 12940 17141 12968
rect 17092 12928 17098 12940
rect 17129 12937 17141 12940
rect 17175 12937 17187 12971
rect 17129 12931 17187 12937
rect 17218 12928 17224 12980
rect 17276 12928 17282 12980
rect 21358 12968 21364 12980
rect 20824 12940 21364 12968
rect 14458 12860 14464 12912
rect 14516 12860 14522 12912
rect 16298 12900 16304 12912
rect 15686 12886 16304 12900
rect 15672 12872 16304 12886
rect 14185 12835 14243 12841
rect 14185 12801 14197 12835
rect 14231 12801 14243 12835
rect 14185 12795 14243 12801
rect 15672 12776 15700 12872
rect 16298 12860 16304 12872
rect 16356 12860 16362 12912
rect 19061 12903 19119 12909
rect 19061 12900 19073 12903
rect 18340 12872 19073 12900
rect 18340 12841 18368 12872
rect 19061 12869 19073 12872
rect 19107 12869 19119 12903
rect 20824 12900 20852 12940
rect 21358 12928 21364 12940
rect 21416 12928 21422 12980
rect 20746 12872 20852 12900
rect 19061 12863 19119 12869
rect 20898 12860 20904 12912
rect 20956 12900 20962 12912
rect 21177 12903 21235 12909
rect 21177 12900 21189 12903
rect 20956 12872 21189 12900
rect 20956 12860 20962 12872
rect 21177 12869 21189 12872
rect 21223 12869 21235 12903
rect 21177 12863 21235 12869
rect 23293 12903 23351 12909
rect 23293 12869 23305 12903
rect 23339 12900 23351 12903
rect 24854 12900 24860 12912
rect 23339 12872 24860 12900
rect 23339 12869 23351 12872
rect 23293 12863 23351 12869
rect 24854 12860 24860 12872
rect 24912 12860 24918 12912
rect 18325 12835 18383 12841
rect 18325 12832 18337 12835
rect 15764 12804 18337 12832
rect 8570 12724 8576 12776
rect 8628 12764 8634 12776
rect 8846 12764 8852 12776
rect 8628 12736 8852 12764
rect 8628 12724 8634 12736
rect 8846 12724 8852 12736
rect 8904 12764 8910 12776
rect 8941 12767 8999 12773
rect 8941 12764 8953 12767
rect 8904 12736 8953 12764
rect 8904 12724 8910 12736
rect 8941 12733 8953 12736
rect 8987 12733 8999 12767
rect 8941 12727 8999 12733
rect 11330 12724 11336 12776
rect 11388 12764 11394 12776
rect 12345 12767 12403 12773
rect 12345 12764 12357 12767
rect 11388 12736 12357 12764
rect 11388 12724 11394 12736
rect 12345 12733 12357 12736
rect 12391 12733 12403 12767
rect 12345 12727 12403 12733
rect 14090 12724 14096 12776
rect 14148 12764 14154 12776
rect 14148 12736 15608 12764
rect 14148 12724 14154 12736
rect 15580 12696 15608 12736
rect 15654 12724 15660 12776
rect 15712 12724 15718 12776
rect 15764 12696 15792 12804
rect 18325 12801 18337 12804
rect 18371 12801 18383 12835
rect 18325 12795 18383 12801
rect 18414 12792 18420 12844
rect 18472 12792 18478 12844
rect 22094 12792 22100 12844
rect 22152 12792 22158 12844
rect 23934 12792 23940 12844
rect 23992 12792 23998 12844
rect 15933 12767 15991 12773
rect 15933 12733 15945 12767
rect 15979 12764 15991 12767
rect 16482 12764 16488 12776
rect 15979 12736 16488 12764
rect 15979 12733 15991 12736
rect 15933 12727 15991 12733
rect 16482 12724 16488 12736
rect 16540 12764 16546 12776
rect 16945 12767 17003 12773
rect 16945 12764 16957 12767
rect 16540 12736 16957 12764
rect 16540 12724 16546 12736
rect 16945 12733 16957 12736
rect 16991 12733 17003 12767
rect 16945 12727 17003 12733
rect 18233 12767 18291 12773
rect 18233 12733 18245 12767
rect 18279 12764 18291 12767
rect 19426 12764 19432 12776
rect 18279 12736 19432 12764
rect 18279 12733 18291 12736
rect 18233 12727 18291 12733
rect 19426 12724 19432 12736
rect 19484 12764 19490 12776
rect 19705 12767 19763 12773
rect 19705 12764 19717 12767
rect 19484 12736 19717 12764
rect 19484 12724 19490 12736
rect 19705 12733 19717 12736
rect 19751 12733 19763 12767
rect 19705 12727 19763 12733
rect 21450 12724 21456 12776
rect 21508 12724 21514 12776
rect 24762 12724 24768 12776
rect 24820 12724 24826 12776
rect 15580 12668 15792 12696
rect 18785 12699 18843 12705
rect 18785 12665 18797 12699
rect 18831 12696 18843 12699
rect 18831 12668 19748 12696
rect 18831 12665 18843 12668
rect 18785 12659 18843 12665
rect 19720 12640 19748 12668
rect 9585 12631 9643 12637
rect 9585 12597 9597 12631
rect 9631 12628 9643 12631
rect 10962 12628 10968 12640
rect 9631 12600 10968 12628
rect 9631 12597 9643 12600
rect 9585 12591 9643 12597
rect 10962 12588 10968 12600
rect 11020 12588 11026 12640
rect 13633 12631 13691 12637
rect 13633 12597 13645 12631
rect 13679 12628 13691 12631
rect 14274 12628 14280 12640
rect 13679 12600 14280 12628
rect 13679 12597 13691 12600
rect 13633 12591 13691 12597
rect 14274 12588 14280 12600
rect 14332 12588 14338 12640
rect 17589 12631 17647 12637
rect 17589 12597 17601 12631
rect 17635 12628 17647 12631
rect 19518 12628 19524 12640
rect 17635 12600 19524 12628
rect 17635 12597 17647 12600
rect 17589 12591 17647 12597
rect 19518 12588 19524 12600
rect 19576 12588 19582 12640
rect 19702 12588 19708 12640
rect 19760 12588 19766 12640
rect 1104 12538 25852 12560
rect 1104 12486 2950 12538
rect 3002 12486 3014 12538
rect 3066 12486 3078 12538
rect 3130 12486 3142 12538
rect 3194 12486 3206 12538
rect 3258 12486 12950 12538
rect 13002 12486 13014 12538
rect 13066 12486 13078 12538
rect 13130 12486 13142 12538
rect 13194 12486 13206 12538
rect 13258 12486 22950 12538
rect 23002 12486 23014 12538
rect 23066 12486 23078 12538
rect 23130 12486 23142 12538
rect 23194 12486 23206 12538
rect 23258 12486 25852 12538
rect 1104 12464 25852 12486
rect 11057 12427 11115 12433
rect 11057 12393 11069 12427
rect 11103 12424 11115 12427
rect 12434 12424 12440 12436
rect 11103 12396 12440 12424
rect 11103 12393 11115 12396
rect 11057 12387 11115 12393
rect 12434 12384 12440 12396
rect 12492 12384 12498 12436
rect 13446 12384 13452 12436
rect 13504 12424 13510 12436
rect 14277 12427 14335 12433
rect 14277 12424 14289 12427
rect 13504 12396 14289 12424
rect 13504 12384 13510 12396
rect 14277 12393 14289 12396
rect 14323 12393 14335 12427
rect 14277 12387 14335 12393
rect 14458 12384 14464 12436
rect 14516 12424 14522 12436
rect 15562 12424 15568 12436
rect 14516 12396 15568 12424
rect 14516 12384 14522 12396
rect 15562 12384 15568 12396
rect 15620 12424 15626 12436
rect 15620 12396 16344 12424
rect 15620 12384 15626 12396
rect 3326 12316 3332 12368
rect 3384 12356 3390 12368
rect 6730 12356 6736 12368
rect 3384 12328 6736 12356
rect 3384 12316 3390 12328
rect 6730 12316 6736 12328
rect 6788 12316 6794 12368
rect 10962 12316 10968 12368
rect 11020 12356 11026 12368
rect 11020 12328 16252 12356
rect 11020 12316 11026 12328
rect 9309 12291 9367 12297
rect 9309 12257 9321 12291
rect 9355 12288 9367 12291
rect 11238 12288 11244 12300
rect 9355 12260 11244 12288
rect 9355 12257 9367 12260
rect 9309 12251 9367 12257
rect 11238 12248 11244 12260
rect 11296 12248 11302 12300
rect 14921 12291 14979 12297
rect 14921 12257 14933 12291
rect 14967 12288 14979 12291
rect 15102 12288 15108 12300
rect 14967 12260 15108 12288
rect 14967 12257 14979 12260
rect 14921 12251 14979 12257
rect 15102 12248 15108 12260
rect 15160 12248 15166 12300
rect 12802 12180 12808 12232
rect 12860 12180 12866 12232
rect 14645 12223 14703 12229
rect 14645 12189 14657 12223
rect 14691 12220 14703 12223
rect 15194 12220 15200 12232
rect 14691 12192 15200 12220
rect 14691 12189 14703 12192
rect 14645 12183 14703 12189
rect 15194 12180 15200 12192
rect 15252 12180 15258 12232
rect 15378 12180 15384 12232
rect 15436 12220 15442 12232
rect 16224 12229 16252 12328
rect 15565 12223 15623 12229
rect 15565 12220 15577 12223
rect 15436 12192 15577 12220
rect 15436 12180 15442 12192
rect 15565 12189 15577 12192
rect 15611 12189 15623 12223
rect 15565 12183 15623 12189
rect 16209 12223 16267 12229
rect 16209 12189 16221 12223
rect 16255 12189 16267 12223
rect 16316 12220 16344 12396
rect 17126 12384 17132 12436
rect 17184 12384 17190 12436
rect 20993 12427 21051 12433
rect 17604 12396 20852 12424
rect 16393 12359 16451 12365
rect 16393 12325 16405 12359
rect 16439 12356 16451 12359
rect 17604 12356 17632 12396
rect 16439 12328 17632 12356
rect 16439 12325 16451 12328
rect 16393 12319 16451 12325
rect 19978 12316 19984 12368
rect 20036 12316 20042 12368
rect 16850 12248 16856 12300
rect 16908 12288 16914 12300
rect 18877 12291 18935 12297
rect 18877 12288 18889 12291
rect 16908 12260 18889 12288
rect 16908 12248 16914 12260
rect 18877 12257 18889 12260
rect 18923 12257 18935 12291
rect 18877 12251 18935 12257
rect 19521 12223 19579 12229
rect 16316 12206 17526 12220
rect 16316 12192 17540 12206
rect 16209 12183 16267 12189
rect 8846 12112 8852 12164
rect 8904 12152 8910 12164
rect 9585 12155 9643 12161
rect 9585 12152 9597 12155
rect 8904 12124 9597 12152
rect 8904 12112 8910 12124
rect 9585 12121 9597 12124
rect 9631 12121 9643 12155
rect 9585 12115 9643 12121
rect 9674 12112 9680 12164
rect 9732 12152 9738 12164
rect 9732 12124 10074 12152
rect 9732 12112 9738 12124
rect 9968 12084 9996 12124
rect 12618 12112 12624 12164
rect 12676 12152 12682 12164
rect 13446 12152 13452 12164
rect 12676 12124 13452 12152
rect 12676 12112 12682 12124
rect 13446 12112 13452 12124
rect 13504 12152 13510 12164
rect 13541 12155 13599 12161
rect 13541 12152 13553 12155
rect 13504 12124 13553 12152
rect 13504 12112 13510 12124
rect 13541 12121 13553 12124
rect 13587 12121 13599 12155
rect 13541 12115 13599 12121
rect 13725 12155 13783 12161
rect 13725 12121 13737 12155
rect 13771 12152 13783 12155
rect 14182 12152 14188 12164
rect 13771 12124 14188 12152
rect 13771 12121 13783 12124
rect 13725 12115 13783 12121
rect 14182 12112 14188 12124
rect 14240 12112 14246 12164
rect 15580 12152 15608 12183
rect 16669 12155 16727 12161
rect 16669 12152 16681 12155
rect 15580 12124 16681 12152
rect 16669 12121 16681 12124
rect 16715 12121 16727 12155
rect 16669 12115 16727 12121
rect 11333 12087 11391 12093
rect 11333 12084 11345 12087
rect 9968 12056 11345 12084
rect 11333 12053 11345 12056
rect 11379 12084 11391 12087
rect 11974 12084 11980 12096
rect 11379 12056 11980 12084
rect 11379 12053 11391 12056
rect 11333 12047 11391 12053
rect 11974 12044 11980 12056
rect 12032 12044 12038 12096
rect 12710 12044 12716 12096
rect 12768 12084 12774 12096
rect 12897 12087 12955 12093
rect 12897 12084 12909 12087
rect 12768 12056 12909 12084
rect 12768 12044 12774 12056
rect 12897 12053 12909 12056
rect 12943 12053 12955 12087
rect 12897 12047 12955 12053
rect 14734 12044 14740 12096
rect 14792 12044 14798 12096
rect 15654 12044 15660 12096
rect 15712 12044 15718 12096
rect 17512 12084 17540 12192
rect 19521 12189 19533 12223
rect 19567 12220 19579 12223
rect 19996 12220 20024 12316
rect 20824 12229 20852 12396
rect 20993 12393 21005 12427
rect 21039 12424 21051 12427
rect 22094 12424 22100 12436
rect 21039 12396 22100 12424
rect 21039 12393 21051 12396
rect 20993 12387 21051 12393
rect 22094 12384 22100 12396
rect 22152 12384 22158 12436
rect 19567 12192 20024 12220
rect 20809 12223 20867 12229
rect 19567 12189 19579 12192
rect 19521 12183 19579 12189
rect 20809 12189 20821 12223
rect 20855 12189 20867 12223
rect 20809 12183 20867 12189
rect 22646 12180 22652 12232
rect 22704 12180 22710 12232
rect 22738 12180 22744 12232
rect 22796 12220 22802 12232
rect 24765 12223 24823 12229
rect 24765 12220 24777 12223
rect 22796 12192 24777 12220
rect 22796 12180 22802 12192
rect 24765 12189 24777 12192
rect 24811 12189 24823 12223
rect 24765 12183 24823 12189
rect 18601 12155 18659 12161
rect 18170 12124 18552 12152
rect 18248 12084 18276 12124
rect 17512 12056 18276 12084
rect 18524 12084 18552 12124
rect 18601 12121 18613 12155
rect 18647 12152 18659 12155
rect 19242 12152 19248 12164
rect 18647 12124 19248 12152
rect 18647 12121 18659 12124
rect 18601 12115 18659 12121
rect 19242 12112 19248 12124
rect 19300 12112 19306 12164
rect 23845 12155 23903 12161
rect 23845 12121 23857 12155
rect 23891 12152 23903 12155
rect 24946 12152 24952 12164
rect 23891 12124 24952 12152
rect 23891 12121 23903 12124
rect 23845 12115 23903 12121
rect 24946 12112 24952 12124
rect 25004 12112 25010 12164
rect 19058 12084 19064 12096
rect 18524 12056 19064 12084
rect 19058 12044 19064 12056
rect 19116 12044 19122 12096
rect 19426 12044 19432 12096
rect 19484 12084 19490 12096
rect 19613 12087 19671 12093
rect 19613 12084 19625 12087
rect 19484 12056 19625 12084
rect 19484 12044 19490 12056
rect 19613 12053 19625 12056
rect 19659 12053 19671 12087
rect 19613 12047 19671 12053
rect 21358 12044 21364 12096
rect 21416 12084 21422 12096
rect 21545 12087 21603 12093
rect 21545 12084 21557 12087
rect 21416 12056 21557 12084
rect 21416 12044 21422 12056
rect 21545 12053 21557 12056
rect 21591 12053 21603 12087
rect 21545 12047 21603 12053
rect 24578 12044 24584 12096
rect 24636 12044 24642 12096
rect 1104 11994 25852 12016
rect 1104 11942 7950 11994
rect 8002 11942 8014 11994
rect 8066 11942 8078 11994
rect 8130 11942 8142 11994
rect 8194 11942 8206 11994
rect 8258 11942 17950 11994
rect 18002 11942 18014 11994
rect 18066 11942 18078 11994
rect 18130 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 25852 11994
rect 1104 11920 25852 11942
rect 13814 11880 13820 11892
rect 13280 11852 13820 11880
rect 11974 11772 11980 11824
rect 12032 11812 12038 11824
rect 13280 11812 13308 11852
rect 13814 11840 13820 11852
rect 13872 11880 13878 11892
rect 13872 11852 14320 11880
rect 13872 11840 13878 11852
rect 14292 11812 14320 11852
rect 14366 11840 14372 11892
rect 14424 11840 14430 11892
rect 14918 11840 14924 11892
rect 14976 11840 14982 11892
rect 15378 11840 15384 11892
rect 15436 11880 15442 11892
rect 18414 11880 18420 11892
rect 15436 11852 18420 11880
rect 15436 11840 15442 11852
rect 18414 11840 18420 11852
rect 18472 11840 18478 11892
rect 19797 11883 19855 11889
rect 19797 11849 19809 11883
rect 19843 11849 19855 11883
rect 19797 11843 19855 11849
rect 14458 11812 14464 11824
rect 12032 11784 13386 11812
rect 14292 11784 14464 11812
rect 12032 11772 12038 11784
rect 14458 11772 14464 11784
rect 14516 11772 14522 11824
rect 15289 11815 15347 11821
rect 15289 11781 15301 11815
rect 15335 11812 15347 11815
rect 17310 11812 17316 11824
rect 15335 11784 17316 11812
rect 15335 11781 15347 11784
rect 15289 11775 15347 11781
rect 17310 11772 17316 11784
rect 17368 11772 17374 11824
rect 19334 11772 19340 11824
rect 19392 11812 19398 11824
rect 19812 11812 19840 11843
rect 22646 11840 22652 11892
rect 22704 11840 22710 11892
rect 19392 11784 19748 11812
rect 19812 11784 23244 11812
rect 19392 11772 19398 11784
rect 19610 11704 19616 11756
rect 19668 11704 19674 11756
rect 19720 11744 19748 11784
rect 20349 11747 20407 11753
rect 20349 11744 20361 11747
rect 19720 11716 20361 11744
rect 20349 11713 20361 11716
rect 20395 11744 20407 11747
rect 20809 11747 20867 11753
rect 20809 11744 20821 11747
rect 20395 11716 20821 11744
rect 20395 11713 20407 11716
rect 20349 11707 20407 11713
rect 20809 11713 20821 11716
rect 20855 11713 20867 11747
rect 20809 11707 20867 11713
rect 22462 11704 22468 11756
rect 22520 11704 22526 11756
rect 23216 11753 23244 11784
rect 23201 11747 23259 11753
rect 23201 11713 23213 11747
rect 23247 11713 23259 11747
rect 23201 11707 23259 11713
rect 23658 11704 23664 11756
rect 23716 11744 23722 11756
rect 23937 11747 23995 11753
rect 23937 11744 23949 11747
rect 23716 11716 23949 11744
rect 23716 11704 23722 11716
rect 23937 11713 23949 11716
rect 23983 11713 23995 11747
rect 23937 11707 23995 11713
rect 11238 11636 11244 11688
rect 11296 11676 11302 11688
rect 12250 11676 12256 11688
rect 11296 11648 12256 11676
rect 11296 11636 11302 11648
rect 12250 11636 12256 11648
rect 12308 11676 12314 11688
rect 12621 11679 12679 11685
rect 12621 11676 12633 11679
rect 12308 11648 12633 11676
rect 12308 11636 12314 11648
rect 12621 11645 12633 11648
rect 12667 11645 12679 11679
rect 12621 11639 12679 11645
rect 12897 11679 12955 11685
rect 12897 11645 12909 11679
rect 12943 11676 12955 11679
rect 13354 11676 13360 11688
rect 12943 11648 13360 11676
rect 12943 11645 12955 11648
rect 12897 11639 12955 11645
rect 13354 11636 13360 11648
rect 13412 11636 13418 11688
rect 15378 11636 15384 11688
rect 15436 11636 15442 11688
rect 15470 11636 15476 11688
rect 15528 11636 15534 11688
rect 15562 11636 15568 11688
rect 15620 11676 15626 11688
rect 16117 11679 16175 11685
rect 16117 11676 16129 11679
rect 15620 11648 16129 11676
rect 15620 11636 15626 11648
rect 16117 11645 16129 11648
rect 16163 11645 16175 11679
rect 16117 11639 16175 11645
rect 24670 11636 24676 11688
rect 24728 11636 24734 11688
rect 15838 11568 15844 11620
rect 15896 11608 15902 11620
rect 19978 11608 19984 11620
rect 15896 11580 19984 11608
rect 15896 11568 15902 11580
rect 19978 11568 19984 11580
rect 20036 11608 20042 11620
rect 20346 11608 20352 11620
rect 20036 11580 20352 11608
rect 20036 11568 20042 11580
rect 20346 11568 20352 11580
rect 20404 11568 20410 11620
rect 20533 11611 20591 11617
rect 20533 11577 20545 11611
rect 20579 11608 20591 11611
rect 23474 11608 23480 11620
rect 20579 11580 23480 11608
rect 20579 11577 20591 11580
rect 20533 11571 20591 11577
rect 23474 11568 23480 11580
rect 23532 11568 23538 11620
rect 19058 11500 19064 11552
rect 19116 11500 19122 11552
rect 23385 11543 23443 11549
rect 23385 11509 23397 11543
rect 23431 11540 23443 11543
rect 23934 11540 23940 11552
rect 23431 11512 23940 11540
rect 23431 11509 23443 11512
rect 23385 11503 23443 11509
rect 23934 11500 23940 11512
rect 23992 11500 23998 11552
rect 1104 11450 25852 11472
rect 1104 11398 2950 11450
rect 3002 11398 3014 11450
rect 3066 11398 3078 11450
rect 3130 11398 3142 11450
rect 3194 11398 3206 11450
rect 3258 11398 12950 11450
rect 13002 11398 13014 11450
rect 13066 11398 13078 11450
rect 13130 11398 13142 11450
rect 13194 11398 13206 11450
rect 13258 11398 22950 11450
rect 23002 11398 23014 11450
rect 23066 11398 23078 11450
rect 23130 11398 23142 11450
rect 23194 11398 23206 11450
rect 23258 11398 25852 11450
rect 1104 11376 25852 11398
rect 11974 11296 11980 11348
rect 12032 11336 12038 11348
rect 13265 11339 13323 11345
rect 13265 11336 13277 11339
rect 12032 11308 13277 11336
rect 12032 11296 12038 11308
rect 13265 11305 13277 11308
rect 13311 11305 13323 11339
rect 13265 11299 13323 11305
rect 13998 11296 14004 11348
rect 14056 11336 14062 11348
rect 15473 11339 15531 11345
rect 15473 11336 15485 11339
rect 14056 11308 15485 11336
rect 14056 11296 14062 11308
rect 15473 11305 15485 11308
rect 15519 11305 15531 11339
rect 15473 11299 15531 11305
rect 18325 11339 18383 11345
rect 18325 11305 18337 11339
rect 18371 11336 18383 11339
rect 22462 11336 22468 11348
rect 18371 11308 22468 11336
rect 18371 11305 18383 11308
rect 18325 11299 18383 11305
rect 22462 11296 22468 11308
rect 22520 11296 22526 11348
rect 13446 11228 13452 11280
rect 13504 11268 13510 11280
rect 13817 11271 13875 11277
rect 13817 11268 13829 11271
rect 13504 11240 13829 11268
rect 13504 11228 13510 11240
rect 13817 11237 13829 11240
rect 13863 11237 13875 11271
rect 13817 11231 13875 11237
rect 15013 11271 15071 11277
rect 15013 11237 15025 11271
rect 15059 11268 15071 11271
rect 20165 11271 20223 11277
rect 15059 11240 16574 11268
rect 15059 11237 15071 11240
rect 15013 11231 15071 11237
rect 11238 11160 11244 11212
rect 11296 11160 11302 11212
rect 11517 11203 11575 11209
rect 11517 11169 11529 11203
rect 11563 11200 11575 11203
rect 12526 11200 12532 11212
rect 11563 11172 12532 11200
rect 11563 11169 11575 11172
rect 11517 11163 11575 11169
rect 12526 11160 12532 11172
rect 12584 11160 12590 11212
rect 12989 11203 13047 11209
rect 12989 11169 13001 11203
rect 13035 11200 13047 11203
rect 13354 11200 13360 11212
rect 13035 11172 13360 11200
rect 13035 11169 13047 11172
rect 12989 11163 13047 11169
rect 13354 11160 13360 11172
rect 13412 11200 13418 11212
rect 14369 11203 14427 11209
rect 14369 11200 14381 11203
rect 13412 11172 14381 11200
rect 13412 11160 13418 11172
rect 14369 11169 14381 11172
rect 14415 11169 14427 11203
rect 14369 11163 14427 11169
rect 14550 11160 14556 11212
rect 14608 11160 14614 11212
rect 15102 11160 15108 11212
rect 15160 11200 15166 11212
rect 16025 11203 16083 11209
rect 16025 11200 16037 11203
rect 15160 11172 16037 11200
rect 15160 11160 15166 11172
rect 16025 11169 16037 11172
rect 16071 11169 16083 11203
rect 16025 11163 16083 11169
rect 14645 11135 14703 11141
rect 14645 11101 14657 11135
rect 14691 11132 14703 11135
rect 15562 11132 15568 11144
rect 14691 11104 15568 11132
rect 14691 11101 14703 11104
rect 14645 11095 14703 11101
rect 15562 11092 15568 11104
rect 15620 11092 15626 11144
rect 15838 11092 15844 11144
rect 15896 11092 15902 11144
rect 16546 11132 16574 11240
rect 20165 11237 20177 11271
rect 20211 11268 20223 11271
rect 22002 11268 22008 11280
rect 20211 11240 22008 11268
rect 20211 11237 20223 11240
rect 20165 11231 20223 11237
rect 22002 11228 22008 11240
rect 22060 11228 22066 11280
rect 22830 11228 22836 11280
rect 22888 11268 22894 11280
rect 22925 11271 22983 11277
rect 22925 11268 22937 11271
rect 22888 11240 22937 11268
rect 22888 11228 22894 11240
rect 22925 11237 22937 11240
rect 22971 11237 22983 11271
rect 22925 11231 22983 11237
rect 19242 11160 19248 11212
rect 19300 11200 19306 11212
rect 19521 11203 19579 11209
rect 19521 11200 19533 11203
rect 19300 11172 19533 11200
rect 19300 11160 19306 11172
rect 19521 11169 19533 11172
rect 19567 11169 19579 11203
rect 19521 11163 19579 11169
rect 19702 11160 19708 11212
rect 19760 11160 19766 11212
rect 22554 11160 22560 11212
rect 22612 11200 22618 11212
rect 22612 11172 24808 11200
rect 22612 11160 22618 11172
rect 18141 11135 18199 11141
rect 18141 11132 18153 11135
rect 16546 11104 18153 11132
rect 18141 11101 18153 11104
rect 18187 11101 18199 11135
rect 18141 11095 18199 11101
rect 21910 11092 21916 11144
rect 21968 11132 21974 11144
rect 22741 11135 22799 11141
rect 22741 11132 22753 11135
rect 21968 11104 22753 11132
rect 21968 11092 21974 11104
rect 22741 11101 22753 11104
rect 22787 11101 22799 11135
rect 22741 11095 22799 11101
rect 23382 11092 23388 11144
rect 23440 11132 23446 11144
rect 24780 11141 24808 11172
rect 23845 11135 23903 11141
rect 23845 11132 23857 11135
rect 23440 11104 23857 11132
rect 23440 11092 23446 11104
rect 23845 11101 23857 11104
rect 23891 11101 23903 11135
rect 23845 11095 23903 11101
rect 24765 11135 24823 11141
rect 24765 11101 24777 11135
rect 24811 11101 24823 11135
rect 24765 11095 24823 11101
rect 11974 11024 11980 11076
rect 12032 11024 12038 11076
rect 19797 11067 19855 11073
rect 19797 11033 19809 11067
rect 19843 11064 19855 11067
rect 20625 11067 20683 11073
rect 20625 11064 20637 11067
rect 19843 11036 20637 11064
rect 19843 11033 19855 11036
rect 19797 11027 19855 11033
rect 20625 11033 20637 11036
rect 20671 11033 20683 11067
rect 20625 11027 20683 11033
rect 24210 11024 24216 11076
rect 24268 11064 24274 11076
rect 24581 11067 24639 11073
rect 24581 11064 24593 11067
rect 24268 11036 24593 11064
rect 24268 11024 24274 11036
rect 24581 11033 24593 11036
rect 24627 11033 24639 11067
rect 24581 11027 24639 11033
rect 15933 10999 15991 11005
rect 15933 10965 15945 10999
rect 15979 10996 15991 10999
rect 16022 10996 16028 11008
rect 15979 10968 16028 10996
rect 15979 10965 15991 10968
rect 15933 10959 15991 10965
rect 16022 10956 16028 10968
rect 16080 10956 16086 11008
rect 24026 10956 24032 11008
rect 24084 10956 24090 11008
rect 1104 10906 25852 10928
rect 1104 10854 7950 10906
rect 8002 10854 8014 10906
rect 8066 10854 8078 10906
rect 8130 10854 8142 10906
rect 8194 10854 8206 10906
rect 8258 10854 17950 10906
rect 18002 10854 18014 10906
rect 18066 10854 18078 10906
rect 18130 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 25852 10906
rect 1104 10832 25852 10854
rect 13814 10752 13820 10804
rect 13872 10792 13878 10804
rect 14461 10795 14519 10801
rect 14461 10792 14473 10795
rect 13872 10764 14473 10792
rect 13872 10752 13878 10764
rect 14461 10761 14473 10764
rect 14507 10761 14519 10795
rect 14461 10755 14519 10761
rect 15838 10752 15844 10804
rect 15896 10792 15902 10804
rect 16206 10792 16212 10804
rect 15896 10764 16212 10792
rect 15896 10752 15902 10764
rect 16206 10752 16212 10764
rect 16264 10752 16270 10804
rect 18049 10795 18107 10801
rect 18049 10761 18061 10795
rect 18095 10792 18107 10795
rect 19242 10792 19248 10804
rect 18095 10764 19248 10792
rect 18095 10761 18107 10764
rect 18049 10755 18107 10761
rect 19242 10752 19248 10764
rect 19300 10752 19306 10804
rect 19518 10684 19524 10736
rect 19576 10684 19582 10736
rect 18432 10588 18460 10642
rect 21082 10616 21088 10668
rect 21140 10616 21146 10668
rect 23934 10616 23940 10668
rect 23992 10616 23998 10668
rect 19058 10588 19064 10600
rect 18432 10560 19064 10588
rect 19058 10548 19064 10560
rect 19116 10588 19122 10600
rect 19797 10591 19855 10597
rect 19116 10560 19748 10588
rect 19116 10548 19122 10560
rect 19720 10520 19748 10560
rect 19797 10557 19809 10591
rect 19843 10588 19855 10591
rect 21450 10588 21456 10600
rect 19843 10560 21456 10588
rect 19843 10557 19855 10560
rect 19797 10551 19855 10557
rect 21450 10548 21456 10560
rect 21508 10548 21514 10600
rect 24762 10548 24768 10600
rect 24820 10548 24826 10600
rect 20165 10523 20223 10529
rect 20165 10520 20177 10523
rect 19720 10492 20177 10520
rect 20165 10489 20177 10492
rect 20211 10520 20223 10523
rect 21358 10520 21364 10532
rect 20211 10492 21364 10520
rect 20211 10489 20223 10492
rect 20165 10483 20223 10489
rect 21358 10480 21364 10492
rect 21416 10480 21422 10532
rect 15381 10455 15439 10461
rect 15381 10421 15393 10455
rect 15427 10452 15439 10455
rect 16022 10452 16028 10464
rect 15427 10424 16028 10452
rect 15427 10421 15439 10424
rect 15381 10415 15439 10421
rect 16022 10412 16028 10424
rect 16080 10412 16086 10464
rect 21269 10455 21327 10461
rect 21269 10421 21281 10455
rect 21315 10452 21327 10455
rect 24302 10452 24308 10464
rect 21315 10424 24308 10452
rect 21315 10421 21327 10424
rect 21269 10415 21327 10421
rect 24302 10412 24308 10424
rect 24360 10412 24366 10464
rect 1104 10362 25852 10384
rect 1104 10310 2950 10362
rect 3002 10310 3014 10362
rect 3066 10310 3078 10362
rect 3130 10310 3142 10362
rect 3194 10310 3206 10362
rect 3258 10310 12950 10362
rect 13002 10310 13014 10362
rect 13066 10310 13078 10362
rect 13130 10310 13142 10362
rect 13194 10310 13206 10362
rect 13258 10310 22950 10362
rect 23002 10310 23014 10362
rect 23066 10310 23078 10362
rect 23130 10310 23142 10362
rect 23194 10310 23206 10362
rect 23258 10310 25852 10362
rect 1104 10288 25852 10310
rect 23385 10115 23443 10121
rect 23385 10081 23397 10115
rect 23431 10112 23443 10115
rect 24854 10112 24860 10124
rect 23431 10084 24860 10112
rect 23431 10081 23443 10084
rect 23385 10075 23443 10081
rect 24854 10072 24860 10084
rect 24912 10072 24918 10124
rect 9398 10004 9404 10056
rect 9456 10044 9462 10056
rect 11609 10047 11667 10053
rect 11609 10044 11621 10047
rect 9456 10016 11621 10044
rect 9456 10004 9462 10016
rect 11609 10013 11621 10016
rect 11655 10013 11667 10047
rect 11609 10007 11667 10013
rect 17037 10047 17095 10053
rect 17037 10013 17049 10047
rect 17083 10044 17095 10047
rect 19886 10044 19892 10056
rect 17083 10016 19892 10044
rect 17083 10013 17095 10016
rect 17037 10007 17095 10013
rect 19886 10004 19892 10016
rect 19944 10004 19950 10056
rect 24029 10047 24087 10053
rect 24029 10013 24041 10047
rect 24075 10044 24087 10047
rect 24578 10044 24584 10056
rect 24075 10016 24584 10044
rect 24075 10013 24087 10016
rect 24029 10007 24087 10013
rect 24578 10004 24584 10016
rect 24636 10004 24642 10056
rect 24765 10047 24823 10053
rect 24765 10013 24777 10047
rect 24811 10013 24823 10047
rect 24765 10007 24823 10013
rect 11793 9979 11851 9985
rect 11793 9945 11805 9979
rect 11839 9976 11851 9979
rect 12342 9976 12348 9988
rect 11839 9948 12348 9976
rect 11839 9945 11851 9948
rect 11793 9939 11851 9945
rect 12342 9936 12348 9948
rect 12400 9936 12406 9988
rect 16482 9936 16488 9988
rect 16540 9976 16546 9988
rect 16853 9979 16911 9985
rect 16853 9976 16865 9979
rect 16540 9948 16865 9976
rect 16540 9936 16546 9948
rect 16853 9945 16865 9948
rect 16899 9945 16911 9979
rect 16853 9939 16911 9945
rect 23842 9936 23848 9988
rect 23900 9976 23906 9988
rect 24780 9976 24808 10007
rect 23900 9948 24808 9976
rect 23900 9936 23906 9948
rect 24118 9868 24124 9920
rect 24176 9908 24182 9920
rect 24581 9911 24639 9917
rect 24581 9908 24593 9911
rect 24176 9880 24593 9908
rect 24176 9868 24182 9880
rect 24581 9877 24593 9880
rect 24627 9877 24639 9911
rect 24581 9871 24639 9877
rect 1104 9818 25852 9840
rect 1104 9766 7950 9818
rect 8002 9766 8014 9818
rect 8066 9766 8078 9818
rect 8130 9766 8142 9818
rect 8194 9766 8206 9818
rect 8258 9766 17950 9818
rect 18002 9766 18014 9818
rect 18066 9766 18078 9818
rect 18130 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 25852 9818
rect 1104 9744 25852 9766
rect 2866 9596 2872 9648
rect 2924 9636 2930 9648
rect 5626 9636 5632 9648
rect 2924 9608 5632 9636
rect 2924 9596 2930 9608
rect 5626 9596 5632 9608
rect 5684 9596 5690 9648
rect 5718 9596 5724 9648
rect 5776 9636 5782 9648
rect 6825 9639 6883 9645
rect 6825 9636 6837 9639
rect 5776 9608 6837 9636
rect 5776 9596 5782 9608
rect 6825 9605 6837 9608
rect 6871 9605 6883 9639
rect 6825 9599 6883 9605
rect 13538 9596 13544 9648
rect 13596 9636 13602 9648
rect 14369 9639 14427 9645
rect 14369 9636 14381 9639
rect 13596 9608 14381 9636
rect 13596 9596 13602 9608
rect 14369 9605 14381 9608
rect 14415 9605 14427 9639
rect 14369 9599 14427 9605
rect 5997 9571 6055 9577
rect 5997 9537 6009 9571
rect 6043 9568 6055 9571
rect 6917 9571 6975 9577
rect 6917 9568 6929 9571
rect 6043 9540 6929 9568
rect 6043 9537 6055 9540
rect 5997 9531 6055 9537
rect 6917 9537 6929 9540
rect 6963 9537 6975 9571
rect 6917 9531 6975 9537
rect 22002 9528 22008 9580
rect 22060 9528 22066 9580
rect 23934 9528 23940 9580
rect 23992 9528 23998 9580
rect 6733 9503 6791 9509
rect 6733 9469 6745 9503
rect 6779 9469 6791 9503
rect 6733 9463 6791 9469
rect 6748 9432 6776 9463
rect 24762 9460 24768 9512
rect 24820 9460 24826 9512
rect 7098 9432 7104 9444
rect 6748 9404 7104 9432
rect 7098 9392 7104 9404
rect 7156 9392 7162 9444
rect 7282 9392 7288 9444
rect 7340 9392 7346 9444
rect 14553 9435 14611 9441
rect 14553 9401 14565 9435
rect 14599 9432 14611 9435
rect 15194 9432 15200 9444
rect 14599 9404 15200 9432
rect 14599 9401 14611 9404
rect 14553 9395 14611 9401
rect 15194 9392 15200 9404
rect 15252 9392 15258 9444
rect 22189 9367 22247 9373
rect 22189 9333 22201 9367
rect 22235 9364 22247 9367
rect 24486 9364 24492 9376
rect 22235 9336 24492 9364
rect 22235 9333 22247 9336
rect 22189 9327 22247 9333
rect 24486 9324 24492 9336
rect 24544 9324 24550 9376
rect 1104 9274 25852 9296
rect 1104 9222 2950 9274
rect 3002 9222 3014 9274
rect 3066 9222 3078 9274
rect 3130 9222 3142 9274
rect 3194 9222 3206 9274
rect 3258 9222 12950 9274
rect 13002 9222 13014 9274
rect 13066 9222 13078 9274
rect 13130 9222 13142 9274
rect 13194 9222 13206 9274
rect 13258 9222 22950 9274
rect 23002 9222 23014 9274
rect 23066 9222 23078 9274
rect 23130 9222 23142 9274
rect 23194 9222 23206 9274
rect 23258 9222 25852 9274
rect 1104 9200 25852 9222
rect 15930 8916 15936 8968
rect 15988 8956 15994 8968
rect 16117 8959 16175 8965
rect 16117 8956 16129 8959
rect 15988 8928 16129 8956
rect 15988 8916 15994 8928
rect 16117 8925 16129 8928
rect 16163 8925 16175 8959
rect 16117 8919 16175 8925
rect 18509 8959 18567 8965
rect 18509 8925 18521 8959
rect 18555 8956 18567 8959
rect 18598 8956 18604 8968
rect 18555 8928 18604 8956
rect 18555 8925 18567 8928
rect 18509 8919 18567 8925
rect 18598 8916 18604 8928
rect 18656 8916 18662 8968
rect 22830 8916 22836 8968
rect 22888 8956 22894 8968
rect 23109 8959 23167 8965
rect 23109 8956 23121 8959
rect 22888 8928 23121 8956
rect 22888 8916 22894 8928
rect 23109 8925 23121 8928
rect 23155 8925 23167 8959
rect 23109 8919 23167 8925
rect 24854 8916 24860 8968
rect 24912 8956 24918 8968
rect 25038 8956 25044 8968
rect 24912 8928 25044 8956
rect 24912 8916 24918 8928
rect 25038 8916 25044 8928
rect 25096 8956 25102 8968
rect 25317 8959 25375 8965
rect 25317 8956 25329 8959
rect 25096 8928 25329 8956
rect 25096 8916 25102 8928
rect 25317 8925 25329 8928
rect 25363 8925 25375 8959
rect 25317 8919 25375 8925
rect 16301 8891 16359 8897
rect 16301 8857 16313 8891
rect 16347 8888 16359 8891
rect 17770 8888 17776 8900
rect 16347 8860 17776 8888
rect 16347 8857 16359 8860
rect 16301 8851 16359 8857
rect 17770 8848 17776 8860
rect 17828 8848 17834 8900
rect 18693 8891 18751 8897
rect 18693 8857 18705 8891
rect 18739 8888 18751 8891
rect 20714 8888 20720 8900
rect 18739 8860 20720 8888
rect 18739 8857 18751 8860
rect 18693 8851 18751 8857
rect 20714 8848 20720 8860
rect 20772 8848 20778 8900
rect 22738 8848 22744 8900
rect 22796 8888 22802 8900
rect 23753 8891 23811 8897
rect 23753 8888 23765 8891
rect 22796 8860 23765 8888
rect 22796 8848 22802 8860
rect 23753 8857 23765 8860
rect 23799 8857 23811 8891
rect 23753 8851 23811 8857
rect 23937 8891 23995 8897
rect 23937 8857 23949 8891
rect 23983 8888 23995 8891
rect 25498 8888 25504 8900
rect 23983 8860 25504 8888
rect 23983 8857 23995 8860
rect 23937 8851 23995 8857
rect 25240 8832 25268 8860
rect 25498 8848 25504 8860
rect 25556 8848 25562 8900
rect 23290 8780 23296 8832
rect 23348 8780 23354 8832
rect 24670 8780 24676 8832
rect 24728 8780 24734 8832
rect 25222 8780 25228 8832
rect 25280 8780 25286 8832
rect 1104 8730 25852 8752
rect 1104 8678 7950 8730
rect 8002 8678 8014 8730
rect 8066 8678 8078 8730
rect 8130 8678 8142 8730
rect 8194 8678 8206 8730
rect 8258 8678 17950 8730
rect 18002 8678 18014 8730
rect 18066 8678 18078 8730
rect 18130 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 25852 8730
rect 1104 8656 25852 8678
rect 6822 8616 6828 8628
rect 3896 8588 6828 8616
rect 3896 8489 3924 8588
rect 6822 8576 6828 8588
rect 6880 8576 6886 8628
rect 5905 8551 5963 8557
rect 5905 8517 5917 8551
rect 5951 8548 5963 8551
rect 12618 8548 12624 8560
rect 5951 8520 12624 8548
rect 5951 8517 5963 8520
rect 5905 8511 5963 8517
rect 12618 8508 12624 8520
rect 12676 8508 12682 8560
rect 24670 8548 24676 8560
rect 23492 8520 24676 8548
rect 3881 8483 3939 8489
rect 3881 8449 3893 8483
rect 3927 8449 3939 8483
rect 6365 8483 6423 8489
rect 6365 8480 6377 8483
rect 5290 8452 6377 8480
rect 3881 8443 3939 8449
rect 6365 8449 6377 8452
rect 6411 8480 6423 8483
rect 7558 8480 7564 8492
rect 6411 8452 7564 8480
rect 6411 8449 6423 8452
rect 6365 8443 6423 8449
rect 7558 8440 7564 8452
rect 7616 8440 7622 8492
rect 23492 8489 23520 8520
rect 24670 8508 24676 8520
rect 24728 8508 24734 8560
rect 25130 8508 25136 8560
rect 25188 8508 25194 8560
rect 23477 8483 23535 8489
rect 23477 8449 23489 8483
rect 23523 8449 23535 8483
rect 23477 8443 23535 8449
rect 24026 8440 24032 8492
rect 24084 8440 24090 8492
rect 2774 8372 2780 8424
rect 2832 8412 2838 8424
rect 4157 8415 4215 8421
rect 4157 8412 4169 8415
rect 2832 8384 4169 8412
rect 2832 8372 2838 8384
rect 4157 8381 4169 8384
rect 4203 8381 4215 8415
rect 4157 8375 4215 8381
rect 23017 8415 23075 8421
rect 23017 8381 23029 8415
rect 23063 8412 23075 8415
rect 24578 8412 24584 8424
rect 23063 8384 24584 8412
rect 23063 8381 23075 8384
rect 23017 8375 23075 8381
rect 24578 8372 24584 8384
rect 24636 8372 24642 8424
rect 1104 8186 25852 8208
rect 1104 8134 2950 8186
rect 3002 8134 3014 8186
rect 3066 8134 3078 8186
rect 3130 8134 3142 8186
rect 3194 8134 3206 8186
rect 3258 8134 12950 8186
rect 13002 8134 13014 8186
rect 13066 8134 13078 8186
rect 13130 8134 13142 8186
rect 13194 8134 13206 8186
rect 13258 8134 22950 8186
rect 23002 8134 23014 8186
rect 23066 8134 23078 8186
rect 23130 8134 23142 8186
rect 23194 8134 23206 8186
rect 23258 8134 25852 8186
rect 1104 8112 25852 8134
rect 23385 7939 23443 7945
rect 23385 7905 23397 7939
rect 23431 7936 23443 7939
rect 24946 7936 24952 7948
rect 23431 7908 24952 7936
rect 23431 7905 23443 7908
rect 23385 7899 23443 7905
rect 24946 7896 24952 7908
rect 25004 7896 25010 7948
rect 18693 7871 18751 7877
rect 18693 7837 18705 7871
rect 18739 7868 18751 7871
rect 18782 7868 18788 7880
rect 18739 7840 18788 7868
rect 18739 7837 18751 7840
rect 18693 7831 18751 7837
rect 18782 7828 18788 7840
rect 18840 7828 18846 7880
rect 20349 7871 20407 7877
rect 20349 7837 20361 7871
rect 20395 7868 20407 7871
rect 21266 7868 21272 7880
rect 20395 7840 21272 7868
rect 20395 7837 20407 7840
rect 20349 7831 20407 7837
rect 21266 7828 21272 7840
rect 21324 7828 21330 7880
rect 24029 7871 24087 7877
rect 24029 7837 24041 7871
rect 24075 7868 24087 7871
rect 24210 7868 24216 7880
rect 24075 7840 24216 7868
rect 24075 7837 24087 7840
rect 24029 7831 24087 7837
rect 24210 7828 24216 7840
rect 24268 7828 24274 7880
rect 24302 7828 24308 7880
rect 24360 7868 24366 7880
rect 24857 7871 24915 7877
rect 24857 7868 24869 7871
rect 24360 7840 24869 7868
rect 24360 7828 24366 7840
rect 24857 7837 24869 7840
rect 24903 7837 24915 7871
rect 24857 7831 24915 7837
rect 18877 7803 18935 7809
rect 18877 7769 18889 7803
rect 18923 7800 18935 7803
rect 20254 7800 20260 7812
rect 18923 7772 20260 7800
rect 18923 7769 18935 7772
rect 18877 7763 18935 7769
rect 20254 7760 20260 7772
rect 20312 7760 20318 7812
rect 20533 7803 20591 7809
rect 20533 7769 20545 7803
rect 20579 7800 20591 7803
rect 21082 7800 21088 7812
rect 20579 7772 21088 7800
rect 20579 7769 20591 7772
rect 20533 7763 20591 7769
rect 21082 7760 21088 7772
rect 21140 7760 21146 7812
rect 24670 7692 24676 7744
rect 24728 7692 24734 7744
rect 1104 7642 25852 7664
rect 1104 7590 7950 7642
rect 8002 7590 8014 7642
rect 8066 7590 8078 7642
rect 8130 7590 8142 7642
rect 8194 7590 8206 7642
rect 8258 7590 17950 7642
rect 18002 7590 18014 7642
rect 18066 7590 18078 7642
rect 18130 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 25852 7642
rect 1104 7568 25852 7590
rect 22738 7460 22744 7472
rect 21468 7432 22744 7460
rect 21468 7401 21496 7432
rect 22738 7420 22744 7432
rect 22796 7420 22802 7472
rect 21453 7395 21511 7401
rect 21453 7361 21465 7395
rect 21499 7361 21511 7395
rect 21453 7355 21511 7361
rect 21542 7352 21548 7404
rect 21600 7392 21606 7404
rect 22097 7395 22155 7401
rect 22097 7392 22109 7395
rect 21600 7364 22109 7392
rect 21600 7352 21606 7364
rect 22097 7361 22109 7364
rect 22143 7361 22155 7395
rect 22097 7355 22155 7361
rect 24118 7352 24124 7404
rect 24176 7352 24182 7404
rect 20990 7284 20996 7336
rect 21048 7284 21054 7336
rect 22462 7284 22468 7336
rect 22520 7324 22526 7336
rect 22557 7327 22615 7333
rect 22557 7324 22569 7327
rect 22520 7296 22569 7324
rect 22520 7284 22526 7296
rect 22557 7293 22569 7296
rect 22603 7293 22615 7327
rect 22557 7287 22615 7293
rect 24762 7284 24768 7336
rect 24820 7284 24826 7336
rect 1104 7098 25852 7120
rect 1104 7046 2950 7098
rect 3002 7046 3014 7098
rect 3066 7046 3078 7098
rect 3130 7046 3142 7098
rect 3194 7046 3206 7098
rect 3258 7046 12950 7098
rect 13002 7046 13014 7098
rect 13066 7046 13078 7098
rect 13130 7046 13142 7098
rect 13194 7046 13206 7098
rect 13258 7046 22950 7098
rect 23002 7046 23014 7098
rect 23066 7046 23078 7098
rect 23130 7046 23142 7098
rect 23194 7046 23206 7098
rect 23258 7046 25852 7098
rect 1104 7024 25852 7046
rect 23385 6851 23443 6857
rect 23385 6817 23397 6851
rect 23431 6848 23443 6851
rect 24854 6848 24860 6860
rect 23431 6820 24860 6848
rect 23431 6817 23443 6820
rect 23385 6811 23443 6817
rect 24854 6808 24860 6820
rect 24912 6808 24918 6860
rect 15286 6740 15292 6792
rect 15344 6780 15350 6792
rect 18233 6783 18291 6789
rect 18233 6780 18245 6783
rect 15344 6752 18245 6780
rect 15344 6740 15350 6752
rect 18233 6749 18245 6752
rect 18279 6749 18291 6783
rect 18233 6743 18291 6749
rect 19429 6783 19487 6789
rect 19429 6749 19441 6783
rect 19475 6780 19487 6783
rect 19794 6780 19800 6792
rect 19475 6752 19800 6780
rect 19475 6749 19487 6752
rect 19429 6743 19487 6749
rect 19794 6740 19800 6752
rect 19852 6740 19858 6792
rect 20809 6783 20867 6789
rect 20809 6749 20821 6783
rect 20855 6749 20867 6783
rect 20809 6743 20867 6749
rect 24029 6783 24087 6789
rect 24029 6749 24041 6783
rect 24075 6749 24087 6783
rect 24029 6743 24087 6749
rect 3418 6672 3424 6724
rect 3476 6712 3482 6724
rect 7006 6712 7012 6724
rect 3476 6684 7012 6712
rect 3476 6672 3482 6684
rect 7006 6672 7012 6684
rect 7064 6672 7070 6724
rect 18417 6715 18475 6721
rect 18417 6681 18429 6715
rect 18463 6712 18475 6715
rect 19702 6712 19708 6724
rect 18463 6684 19708 6712
rect 18463 6681 18475 6684
rect 18417 6675 18475 6681
rect 19702 6672 19708 6684
rect 19760 6672 19766 6724
rect 3142 6604 3148 6656
rect 3200 6644 3206 6656
rect 6270 6644 6276 6656
rect 3200 6616 6276 6644
rect 3200 6604 3206 6616
rect 6270 6604 6276 6616
rect 6328 6604 6334 6656
rect 19613 6647 19671 6653
rect 19613 6613 19625 6647
rect 19659 6644 19671 6647
rect 20824 6644 20852 6743
rect 22002 6672 22008 6724
rect 22060 6672 22066 6724
rect 24044 6712 24072 6743
rect 24486 6740 24492 6792
rect 24544 6780 24550 6792
rect 24765 6783 24823 6789
rect 24765 6780 24777 6783
rect 24544 6752 24777 6780
rect 24544 6740 24550 6752
rect 24765 6749 24777 6752
rect 24811 6749 24823 6783
rect 24765 6743 24823 6749
rect 24044 6684 24624 6712
rect 24596 6653 24624 6684
rect 19659 6616 20852 6644
rect 24581 6647 24639 6653
rect 19659 6613 19671 6616
rect 19613 6607 19671 6613
rect 24581 6613 24593 6647
rect 24627 6613 24639 6647
rect 24581 6607 24639 6613
rect 1104 6554 25852 6576
rect 1104 6502 7950 6554
rect 8002 6502 8014 6554
rect 8066 6502 8078 6554
rect 8130 6502 8142 6554
rect 8194 6502 8206 6554
rect 8258 6502 17950 6554
rect 18002 6502 18014 6554
rect 18066 6502 18078 6554
rect 18130 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 25852 6554
rect 1104 6480 25852 6502
rect 19521 6443 19579 6449
rect 19521 6409 19533 6443
rect 19567 6440 19579 6443
rect 21542 6440 21548 6452
rect 19567 6412 21548 6440
rect 19567 6409 19579 6412
rect 19521 6403 19579 6409
rect 21542 6400 21548 6412
rect 21600 6400 21606 6452
rect 11974 6332 11980 6384
rect 12032 6372 12038 6384
rect 21269 6375 21327 6381
rect 12032 6344 20116 6372
rect 12032 6332 12038 6344
rect 17310 6264 17316 6316
rect 17368 6304 17374 6316
rect 20088 6313 20116 6344
rect 21269 6341 21281 6375
rect 21315 6372 21327 6375
rect 23382 6372 23388 6384
rect 21315 6344 23388 6372
rect 21315 6341 21327 6344
rect 21269 6335 21327 6341
rect 23382 6332 23388 6344
rect 23440 6332 23446 6384
rect 19429 6307 19487 6313
rect 19429 6304 19441 6307
rect 17368 6276 19441 6304
rect 17368 6264 17374 6276
rect 19429 6273 19441 6276
rect 19475 6273 19487 6307
rect 19429 6267 19487 6273
rect 20073 6307 20131 6313
rect 20073 6273 20085 6307
rect 20119 6273 20131 6307
rect 20073 6267 20131 6273
rect 20162 6264 20168 6316
rect 20220 6304 20226 6316
rect 22097 6307 22155 6313
rect 22097 6304 22109 6307
rect 20220 6276 22109 6304
rect 20220 6264 20226 6276
rect 22097 6273 22109 6276
rect 22143 6273 22155 6307
rect 22097 6267 22155 6273
rect 23290 6264 23296 6316
rect 23348 6304 23354 6316
rect 23937 6307 23995 6313
rect 23937 6304 23949 6307
rect 23348 6276 23949 6304
rect 23348 6264 23354 6276
rect 23937 6273 23949 6276
rect 23983 6273 23995 6307
rect 23937 6267 23995 6273
rect 22557 6239 22615 6245
rect 22557 6236 22569 6239
rect 22112 6208 22569 6236
rect 22112 6180 22140 6208
rect 22557 6205 22569 6208
rect 22603 6205 22615 6239
rect 22557 6199 22615 6205
rect 24762 6196 24768 6248
rect 24820 6196 24826 6248
rect 22094 6128 22100 6180
rect 22152 6128 22158 6180
rect 16206 6060 16212 6112
rect 16264 6100 16270 6112
rect 23934 6100 23940 6112
rect 16264 6072 23940 6100
rect 16264 6060 16270 6072
rect 23934 6060 23940 6072
rect 23992 6060 23998 6112
rect 1104 6010 25852 6032
rect 1104 5958 2950 6010
rect 3002 5958 3014 6010
rect 3066 5958 3078 6010
rect 3130 5958 3142 6010
rect 3194 5958 3206 6010
rect 3258 5958 12950 6010
rect 13002 5958 13014 6010
rect 13066 5958 13078 6010
rect 13130 5958 13142 6010
rect 13194 5958 13206 6010
rect 13258 5958 22950 6010
rect 23002 5958 23014 6010
rect 23066 5958 23078 6010
rect 23130 5958 23142 6010
rect 23194 5958 23206 6010
rect 23258 5958 25852 6010
rect 1104 5936 25852 5958
rect 20162 5856 20168 5908
rect 20220 5856 20226 5908
rect 20254 5788 20260 5840
rect 20312 5828 20318 5840
rect 20312 5800 22600 5828
rect 20312 5788 20318 5800
rect 10870 5720 10876 5772
rect 10928 5760 10934 5772
rect 15838 5760 15844 5772
rect 10928 5732 15844 5760
rect 10928 5720 10934 5732
rect 15838 5720 15844 5732
rect 15896 5720 15902 5772
rect 18874 5720 18880 5772
rect 18932 5760 18938 5772
rect 19334 5760 19340 5772
rect 18932 5732 19340 5760
rect 18932 5720 18938 5732
rect 19334 5720 19340 5732
rect 19392 5720 19398 5772
rect 20622 5720 20628 5772
rect 20680 5760 20686 5772
rect 21177 5763 21235 5769
rect 21177 5760 21189 5763
rect 20680 5732 21189 5760
rect 20680 5720 20686 5732
rect 21177 5729 21189 5732
rect 21223 5729 21235 5763
rect 21177 5723 21235 5729
rect 19978 5652 19984 5704
rect 20036 5652 20042 5704
rect 20714 5652 20720 5704
rect 20772 5652 20778 5704
rect 22572 5701 22600 5800
rect 23017 5763 23075 5769
rect 23017 5729 23029 5763
rect 23063 5729 23075 5763
rect 23017 5723 23075 5729
rect 22557 5695 22615 5701
rect 22557 5661 22569 5695
rect 22603 5661 22615 5695
rect 22557 5655 22615 5661
rect 21910 5584 21916 5636
rect 21968 5624 21974 5636
rect 23032 5624 23060 5723
rect 21968 5596 23060 5624
rect 21968 5584 21974 5596
rect 7558 5516 7564 5568
rect 7616 5556 7622 5568
rect 13906 5556 13912 5568
rect 7616 5528 13912 5556
rect 7616 5516 7622 5528
rect 13906 5516 13912 5528
rect 13964 5516 13970 5568
rect 1104 5466 25852 5488
rect 1104 5414 7950 5466
rect 8002 5414 8014 5466
rect 8066 5414 8078 5466
rect 8130 5414 8142 5466
rect 8194 5414 8206 5466
rect 8258 5414 17950 5466
rect 18002 5414 18014 5466
rect 18066 5414 18078 5466
rect 18130 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 25852 5466
rect 1104 5392 25852 5414
rect 15746 5312 15752 5364
rect 15804 5352 15810 5364
rect 16850 5352 16856 5364
rect 15804 5324 16856 5352
rect 15804 5312 15810 5324
rect 16850 5312 16856 5324
rect 16908 5312 16914 5364
rect 16206 5244 16212 5296
rect 16264 5244 16270 5296
rect 19794 5284 19800 5296
rect 19168 5256 19800 5284
rect 16022 5176 16028 5228
rect 16080 5176 16086 5228
rect 19168 5225 19196 5256
rect 19794 5244 19800 5256
rect 19852 5244 19858 5296
rect 19153 5219 19211 5225
rect 19153 5185 19165 5219
rect 19199 5185 19211 5219
rect 19153 5179 19211 5185
rect 19426 5176 19432 5228
rect 19484 5216 19490 5228
rect 19613 5219 19671 5225
rect 19613 5216 19625 5219
rect 19484 5188 19625 5216
rect 19484 5176 19490 5188
rect 19613 5185 19625 5188
rect 19659 5185 19671 5219
rect 19613 5179 19671 5185
rect 19702 5176 19708 5228
rect 19760 5216 19766 5228
rect 22005 5219 22063 5225
rect 22005 5216 22017 5219
rect 19760 5188 22017 5216
rect 19760 5176 19766 5188
rect 22005 5185 22017 5188
rect 22051 5185 22063 5219
rect 22005 5179 22063 5185
rect 24121 5219 24179 5225
rect 24121 5185 24133 5219
rect 24167 5216 24179 5219
rect 24670 5216 24676 5228
rect 24167 5188 24676 5216
rect 24167 5185 24179 5188
rect 24121 5179 24179 5185
rect 24670 5176 24676 5188
rect 24728 5176 24734 5228
rect 18693 5151 18751 5157
rect 18693 5117 18705 5151
rect 18739 5117 18751 5151
rect 18693 5111 18751 5117
rect 18708 5080 18736 5111
rect 19518 5108 19524 5160
rect 19576 5148 19582 5160
rect 20073 5151 20131 5157
rect 20073 5148 20085 5151
rect 19576 5120 20085 5148
rect 19576 5108 19582 5120
rect 20073 5117 20085 5120
rect 20119 5117 20131 5151
rect 20073 5111 20131 5117
rect 22278 5108 22284 5160
rect 22336 5148 22342 5160
rect 22465 5151 22523 5157
rect 22465 5148 22477 5151
rect 22336 5120 22477 5148
rect 22336 5108 22342 5120
rect 22465 5117 22477 5120
rect 22511 5117 22523 5151
rect 22465 5111 22523 5117
rect 24762 5108 24768 5160
rect 24820 5108 24826 5160
rect 20530 5080 20536 5092
rect 18708 5052 20536 5080
rect 20530 5040 20536 5052
rect 20588 5040 20594 5092
rect 16942 4972 16948 5024
rect 17000 5012 17006 5024
rect 18690 5012 18696 5024
rect 17000 4984 18696 5012
rect 17000 4972 17006 4984
rect 18690 4972 18696 4984
rect 18748 4972 18754 5024
rect 1104 4922 25852 4944
rect 1104 4870 2950 4922
rect 3002 4870 3014 4922
rect 3066 4870 3078 4922
rect 3130 4870 3142 4922
rect 3194 4870 3206 4922
rect 3258 4870 12950 4922
rect 13002 4870 13014 4922
rect 13066 4870 13078 4922
rect 13130 4870 13142 4922
rect 13194 4870 13206 4922
rect 13258 4870 22950 4922
rect 23002 4870 23014 4922
rect 23066 4870 23078 4922
rect 23130 4870 23142 4922
rect 23194 4870 23206 4922
rect 23258 4870 25852 4922
rect 1104 4848 25852 4870
rect 3234 4768 3240 4820
rect 3292 4808 3298 4820
rect 6362 4808 6368 4820
rect 3292 4780 6368 4808
rect 3292 4768 3298 4780
rect 6362 4768 6368 4780
rect 6420 4768 6426 4820
rect 25314 4768 25320 4820
rect 25372 4768 25378 4820
rect 5166 4700 5172 4752
rect 5224 4740 5230 4752
rect 10318 4740 10324 4752
rect 5224 4712 10324 4740
rect 5224 4700 5230 4712
rect 10318 4700 10324 4712
rect 10376 4700 10382 4752
rect 19886 4632 19892 4684
rect 19944 4632 19950 4684
rect 21726 4632 21732 4684
rect 21784 4632 21790 4684
rect 16390 4564 16396 4616
rect 16448 4604 16454 4616
rect 17405 4607 17463 4613
rect 17405 4604 17417 4607
rect 16448 4576 17417 4604
rect 16448 4564 16454 4576
rect 17405 4573 17417 4576
rect 17451 4573 17463 4607
rect 17405 4567 17463 4573
rect 19334 4564 19340 4616
rect 19392 4604 19398 4616
rect 19429 4607 19487 4613
rect 19429 4604 19441 4607
rect 19392 4576 19441 4604
rect 19392 4564 19398 4576
rect 19429 4573 19441 4576
rect 19475 4573 19487 4607
rect 19429 4567 19487 4573
rect 21174 4564 21180 4616
rect 21232 4604 21238 4616
rect 21269 4607 21327 4613
rect 21269 4604 21281 4607
rect 21232 4576 21281 4604
rect 21232 4564 21238 4576
rect 21269 4573 21281 4576
rect 21315 4573 21327 4607
rect 21269 4567 21327 4573
rect 18322 4496 18328 4548
rect 18380 4496 18386 4548
rect 1394 4428 1400 4480
rect 1452 4428 1458 4480
rect 1104 4378 25852 4400
rect 1104 4326 7950 4378
rect 8002 4326 8014 4378
rect 8066 4326 8078 4378
rect 8130 4326 8142 4378
rect 8194 4326 8206 4378
rect 8258 4326 17950 4378
rect 18002 4326 18014 4378
rect 18066 4326 18078 4378
rect 18130 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 25852 4378
rect 1104 4304 25852 4326
rect 8386 4224 8392 4276
rect 8444 4264 8450 4276
rect 10042 4264 10048 4276
rect 8444 4236 10048 4264
rect 8444 4224 8450 4236
rect 10042 4224 10048 4236
rect 10100 4224 10106 4276
rect 5074 4156 5080 4208
rect 5132 4196 5138 4208
rect 8938 4196 8944 4208
rect 5132 4168 8944 4196
rect 5132 4156 5138 4168
rect 8938 4156 8944 4168
rect 8996 4156 9002 4208
rect 13722 4156 13728 4208
rect 13780 4196 13786 4208
rect 14642 4196 14648 4208
rect 13780 4168 14648 4196
rect 13780 4156 13786 4168
rect 14642 4156 14648 4168
rect 14700 4156 14706 4208
rect 21818 4156 21824 4208
rect 21876 4196 21882 4208
rect 21876 4168 22140 4196
rect 21876 4156 21882 4168
rect 1118 4088 1124 4140
rect 1176 4128 1182 4140
rect 1394 4128 1400 4140
rect 1176 4100 1400 4128
rect 1176 4088 1182 4100
rect 1394 4088 1400 4100
rect 1452 4128 1458 4140
rect 1581 4131 1639 4137
rect 1581 4128 1593 4131
rect 1452 4100 1593 4128
rect 1452 4088 1458 4100
rect 1581 4097 1593 4100
rect 1627 4097 1639 4131
rect 1581 4091 1639 4097
rect 8113 4131 8171 4137
rect 8113 4097 8125 4131
rect 8159 4128 8171 4131
rect 8159 4100 8524 4128
rect 8159 4097 8171 4100
rect 8113 4091 8171 4097
rect 1765 3995 1823 4001
rect 1765 3961 1777 3995
rect 1811 3992 1823 3995
rect 5718 3992 5724 4004
rect 1811 3964 5724 3992
rect 1811 3961 1823 3964
rect 1765 3955 1823 3961
rect 5718 3952 5724 3964
rect 5776 3952 5782 4004
rect 7834 3952 7840 4004
rect 7892 3992 7898 4004
rect 7929 3995 7987 4001
rect 7929 3992 7941 3995
rect 7892 3964 7941 3992
rect 7892 3952 7898 3964
rect 7929 3961 7941 3964
rect 7975 3961 7987 3995
rect 7929 3955 7987 3961
rect 2225 3927 2283 3933
rect 2225 3893 2237 3927
rect 2271 3924 2283 3927
rect 2682 3924 2688 3936
rect 2271 3896 2688 3924
rect 2271 3893 2283 3896
rect 2225 3887 2283 3893
rect 2682 3884 2688 3896
rect 2740 3884 2746 3936
rect 2866 3884 2872 3936
rect 2924 3884 2930 3936
rect 3237 3927 3295 3933
rect 3237 3893 3249 3927
rect 3283 3924 3295 3927
rect 3326 3924 3332 3936
rect 3283 3896 3332 3924
rect 3283 3893 3295 3896
rect 3237 3887 3295 3893
rect 3326 3884 3332 3896
rect 3384 3884 3390 3936
rect 5534 3884 5540 3936
rect 5592 3884 5598 3936
rect 8496 3933 8524 4100
rect 9214 4088 9220 4140
rect 9272 4128 9278 4140
rect 9309 4131 9367 4137
rect 9309 4128 9321 4131
rect 9272 4100 9321 4128
rect 9272 4088 9278 4100
rect 9309 4097 9321 4100
rect 9355 4128 9367 4131
rect 9861 4131 9919 4137
rect 9861 4128 9873 4131
rect 9355 4100 9873 4128
rect 9355 4097 9367 4100
rect 9309 4091 9367 4097
rect 9861 4097 9873 4100
rect 9907 4097 9919 4131
rect 9861 4091 9919 4097
rect 12710 4088 12716 4140
rect 12768 4128 12774 4140
rect 12989 4131 13047 4137
rect 12989 4128 13001 4131
rect 12768 4100 13001 4128
rect 12768 4088 12774 4100
rect 12989 4097 13001 4100
rect 13035 4097 13047 4131
rect 12989 4091 13047 4097
rect 15194 4088 15200 4140
rect 15252 4128 15258 4140
rect 16853 4131 16911 4137
rect 16853 4128 16865 4131
rect 15252 4100 16865 4128
rect 15252 4088 15258 4100
rect 16853 4097 16865 4100
rect 16899 4097 16911 4131
rect 16853 4091 16911 4097
rect 18598 4088 18604 4140
rect 18656 4128 18662 4140
rect 22112 4137 22140 4168
rect 18693 4131 18751 4137
rect 18693 4128 18705 4131
rect 18656 4100 18705 4128
rect 18656 4088 18662 4100
rect 18693 4097 18705 4100
rect 18739 4097 18751 4131
rect 18693 4091 18751 4097
rect 22097 4131 22155 4137
rect 22097 4097 22109 4131
rect 22143 4097 22155 4131
rect 22097 4091 22155 4097
rect 23474 4088 23480 4140
rect 23532 4128 23538 4140
rect 23845 4131 23903 4137
rect 23845 4128 23857 4131
rect 23532 4100 23857 4128
rect 23532 4088 23538 4100
rect 23845 4097 23857 4100
rect 23891 4097 23903 4131
rect 23845 4091 23903 4097
rect 12802 4020 12808 4072
rect 12860 4060 12866 4072
rect 13449 4063 13507 4069
rect 13449 4060 13461 4063
rect 12860 4032 13461 4060
rect 12860 4020 12866 4032
rect 13449 4029 13461 4032
rect 13495 4029 13507 4063
rect 13449 4023 13507 4029
rect 16206 4020 16212 4072
rect 16264 4060 16270 4072
rect 17313 4063 17371 4069
rect 17313 4060 17325 4063
rect 16264 4032 17325 4060
rect 16264 4020 16270 4032
rect 17313 4029 17325 4032
rect 17359 4029 17371 4063
rect 17313 4023 17371 4029
rect 18414 4020 18420 4072
rect 18472 4060 18478 4072
rect 19153 4063 19211 4069
rect 19153 4060 19165 4063
rect 18472 4032 19165 4060
rect 18472 4020 18478 4032
rect 19153 4029 19165 4032
rect 19199 4029 19211 4063
rect 19153 4023 19211 4029
rect 20254 4020 20260 4072
rect 20312 4060 20318 4072
rect 22465 4063 22523 4069
rect 22465 4060 22477 4063
rect 20312 4032 22477 4060
rect 20312 4020 20318 4032
rect 22465 4029 22477 4032
rect 22511 4029 22523 4063
rect 22465 4023 22523 4029
rect 24305 4063 24363 4069
rect 24305 4029 24317 4063
rect 24351 4029 24363 4063
rect 24305 4023 24363 4029
rect 9493 3995 9551 4001
rect 9493 3961 9505 3995
rect 9539 3992 9551 3995
rect 12066 3992 12072 4004
rect 9539 3964 12072 3992
rect 9539 3961 9551 3964
rect 9493 3955 9551 3961
rect 12066 3952 12072 3964
rect 12124 3952 12130 4004
rect 21358 3952 21364 4004
rect 21416 3992 21422 4004
rect 24320 3992 24348 4023
rect 21416 3964 24348 3992
rect 21416 3952 21422 3964
rect 8481 3927 8539 3933
rect 8481 3893 8493 3927
rect 8527 3924 8539 3927
rect 8754 3924 8760 3936
rect 8527 3896 8760 3924
rect 8527 3893 8539 3896
rect 8481 3887 8539 3893
rect 8754 3884 8760 3896
rect 8812 3884 8818 3936
rect 10962 3884 10968 3936
rect 11020 3924 11026 3936
rect 11241 3927 11299 3933
rect 11241 3924 11253 3927
rect 11020 3896 11253 3924
rect 11020 3884 11026 3896
rect 11241 3893 11253 3896
rect 11287 3893 11299 3927
rect 11241 3887 11299 3893
rect 11790 3884 11796 3936
rect 11848 3924 11854 3936
rect 12621 3927 12679 3933
rect 12621 3924 12633 3927
rect 11848 3896 12633 3924
rect 11848 3884 11854 3896
rect 12621 3893 12633 3896
rect 12667 3893 12679 3927
rect 12621 3887 12679 3893
rect 20990 3884 20996 3936
rect 21048 3924 21054 3936
rect 25314 3924 25320 3936
rect 21048 3896 25320 3924
rect 21048 3884 21054 3896
rect 25314 3884 25320 3896
rect 25372 3884 25378 3936
rect 1104 3834 25852 3856
rect 1104 3782 2950 3834
rect 3002 3782 3014 3834
rect 3066 3782 3078 3834
rect 3130 3782 3142 3834
rect 3194 3782 3206 3834
rect 3258 3782 12950 3834
rect 13002 3782 13014 3834
rect 13066 3782 13078 3834
rect 13130 3782 13142 3834
rect 13194 3782 13206 3834
rect 13258 3782 22950 3834
rect 23002 3782 23014 3834
rect 23066 3782 23078 3834
rect 23130 3782 23142 3834
rect 23194 3782 23206 3834
rect 23258 3782 25852 3834
rect 1104 3760 25852 3782
rect 2501 3723 2559 3729
rect 2501 3689 2513 3723
rect 2547 3720 2559 3723
rect 2774 3720 2780 3732
rect 2547 3692 2780 3720
rect 2547 3689 2559 3692
rect 2501 3683 2559 3689
rect 2774 3680 2780 3692
rect 2832 3680 2838 3732
rect 3237 3723 3295 3729
rect 3237 3689 3249 3723
rect 3283 3720 3295 3723
rect 3418 3720 3424 3732
rect 3283 3692 3424 3720
rect 3283 3689 3295 3692
rect 3237 3683 3295 3689
rect 3418 3680 3424 3692
rect 3476 3680 3482 3732
rect 5074 3680 5080 3732
rect 5132 3680 5138 3732
rect 6549 3723 6607 3729
rect 6549 3689 6561 3723
rect 6595 3720 6607 3723
rect 6638 3720 6644 3732
rect 6595 3692 6644 3720
rect 6595 3689 6607 3692
rect 6549 3683 6607 3689
rect 6638 3680 6644 3692
rect 6696 3680 6702 3732
rect 7653 3723 7711 3729
rect 7653 3689 7665 3723
rect 7699 3720 7711 3723
rect 7742 3720 7748 3732
rect 7699 3692 7748 3720
rect 7699 3689 7711 3692
rect 7653 3683 7711 3689
rect 7742 3680 7748 3692
rect 7800 3680 7806 3732
rect 8386 3680 8392 3732
rect 8444 3680 8450 3732
rect 11517 3723 11575 3729
rect 11517 3689 11529 3723
rect 11563 3720 11575 3723
rect 13630 3720 13636 3732
rect 11563 3692 13636 3720
rect 11563 3689 11575 3692
rect 11517 3683 11575 3689
rect 13630 3680 13636 3692
rect 13688 3680 13694 3732
rect 25222 3680 25228 3732
rect 25280 3680 25286 3732
rect 1857 3655 1915 3661
rect 1857 3621 1869 3655
rect 1903 3652 1915 3655
rect 4890 3652 4896 3664
rect 1903 3624 4896 3652
rect 1903 3621 1915 3624
rect 1857 3615 1915 3621
rect 4890 3612 4896 3624
rect 4948 3612 4954 3664
rect 5813 3655 5871 3661
rect 5813 3621 5825 3655
rect 5859 3652 5871 3655
rect 16022 3652 16028 3664
rect 5859 3624 16028 3652
rect 5859 3621 5871 3624
rect 5813 3615 5871 3621
rect 16022 3612 16028 3624
rect 16080 3612 16086 3664
rect 19794 3612 19800 3664
rect 19852 3652 19858 3664
rect 19852 3624 22094 3652
rect 19852 3612 19858 3624
rect 10321 3587 10379 3593
rect 10321 3553 10333 3587
rect 10367 3584 10379 3587
rect 10367 3556 13952 3584
rect 10367 3553 10379 3556
rect 10321 3547 10379 3553
rect 2317 3519 2375 3525
rect 2317 3485 2329 3519
rect 2363 3516 2375 3519
rect 2774 3516 2780 3528
rect 2363 3488 2780 3516
rect 2363 3485 2375 3488
rect 2317 3479 2375 3485
rect 2774 3476 2780 3488
rect 2832 3476 2838 3528
rect 2866 3476 2872 3528
rect 2924 3516 2930 3528
rect 3053 3519 3111 3525
rect 3053 3516 3065 3519
rect 2924 3488 3065 3516
rect 2924 3476 2930 3488
rect 3053 3485 3065 3488
rect 3099 3485 3111 3519
rect 4893 3519 4951 3525
rect 4893 3516 4905 3519
rect 3053 3479 3111 3485
rect 4816 3488 4905 3516
rect 1486 3408 1492 3460
rect 1544 3448 1550 3460
rect 1673 3451 1731 3457
rect 1673 3448 1685 3451
rect 1544 3420 1685 3448
rect 1544 3408 1550 3420
rect 1673 3417 1685 3420
rect 1719 3417 1731 3451
rect 1673 3411 1731 3417
rect 4816 3392 4844 3488
rect 4893 3485 4905 3488
rect 4939 3485 4951 3519
rect 4893 3479 4951 3485
rect 5534 3476 5540 3528
rect 5592 3516 5598 3528
rect 5629 3519 5687 3525
rect 5629 3516 5641 3519
rect 5592 3488 5641 3516
rect 5592 3476 5598 3488
rect 5629 3485 5641 3488
rect 5675 3485 5687 3519
rect 5629 3479 5687 3485
rect 6270 3476 6276 3528
rect 6328 3516 6334 3528
rect 6365 3519 6423 3525
rect 6365 3516 6377 3519
rect 6328 3488 6377 3516
rect 6328 3476 6334 3488
rect 6365 3485 6377 3488
rect 6411 3516 6423 3519
rect 6917 3519 6975 3525
rect 6917 3516 6929 3519
rect 6411 3488 6929 3516
rect 6411 3485 6423 3488
rect 6365 3479 6423 3485
rect 6917 3485 6929 3488
rect 6963 3485 6975 3519
rect 7469 3519 7527 3525
rect 7469 3516 7481 3519
rect 6917 3479 6975 3485
rect 7392 3488 7481 3516
rect 7392 3392 7420 3488
rect 7469 3485 7481 3488
rect 7515 3485 7527 3519
rect 7469 3479 7527 3485
rect 7834 3476 7840 3528
rect 7892 3516 7898 3528
rect 8205 3519 8263 3525
rect 8205 3516 8217 3519
rect 7892 3488 8217 3516
rect 7892 3476 7898 3488
rect 8205 3485 8217 3488
rect 8251 3485 8263 3519
rect 8205 3479 8263 3485
rect 9582 3476 9588 3528
rect 9640 3476 9646 3528
rect 9950 3476 9956 3528
rect 10008 3516 10014 3528
rect 10045 3519 10103 3525
rect 10045 3516 10057 3519
rect 10008 3488 10057 3516
rect 10008 3476 10014 3488
rect 10045 3485 10057 3488
rect 10091 3485 10103 3519
rect 10045 3479 10103 3485
rect 10686 3476 10692 3528
rect 10744 3516 10750 3528
rect 11333 3519 11391 3525
rect 11333 3516 11345 3519
rect 10744 3488 11345 3516
rect 10744 3476 10750 3488
rect 11333 3485 11345 3488
rect 11379 3516 11391 3519
rect 11885 3519 11943 3525
rect 11885 3516 11897 3519
rect 11379 3488 11897 3516
rect 11379 3485 11391 3488
rect 11333 3479 11391 3485
rect 11885 3485 11897 3488
rect 11931 3485 11943 3519
rect 11885 3479 11943 3485
rect 13722 3476 13728 3528
rect 13780 3476 13786 3528
rect 12526 3408 12532 3460
rect 12584 3408 12590 3460
rect 13924 3448 13952 3556
rect 13998 3544 14004 3596
rect 14056 3584 14062 3596
rect 14737 3587 14795 3593
rect 14737 3584 14749 3587
rect 14056 3556 14749 3584
rect 14056 3544 14062 3556
rect 14737 3553 14749 3556
rect 14783 3553 14795 3587
rect 14737 3547 14795 3553
rect 15470 3544 15476 3596
rect 15528 3584 15534 3596
rect 16577 3587 16635 3593
rect 16577 3584 16589 3587
rect 15528 3556 16589 3584
rect 15528 3544 15534 3556
rect 16577 3553 16589 3556
rect 16623 3553 16635 3587
rect 16577 3547 16635 3553
rect 17678 3544 17684 3596
rect 17736 3584 17742 3596
rect 19889 3587 19947 3593
rect 19889 3584 19901 3587
rect 17736 3556 19901 3584
rect 17736 3544 17742 3556
rect 19889 3553 19901 3556
rect 19935 3553 19947 3587
rect 19889 3547 19947 3553
rect 21729 3587 21787 3593
rect 21729 3553 21741 3587
rect 21775 3553 21787 3587
rect 22066 3584 22094 3624
rect 23477 3587 23535 3593
rect 23477 3584 23489 3587
rect 22066 3556 23489 3584
rect 21729 3547 21787 3553
rect 23477 3553 23489 3556
rect 23523 3553 23535 3587
rect 23477 3547 23535 3553
rect 14274 3476 14280 3528
rect 14332 3476 14338 3528
rect 15010 3476 15016 3528
rect 15068 3516 15074 3528
rect 16117 3519 16175 3525
rect 16117 3516 16129 3519
rect 15068 3488 16129 3516
rect 15068 3476 15074 3488
rect 16117 3485 16129 3488
rect 16163 3485 16175 3519
rect 16117 3479 16175 3485
rect 17770 3476 17776 3528
rect 17828 3516 17834 3528
rect 19429 3519 19487 3525
rect 19429 3516 19441 3519
rect 17828 3488 19441 3516
rect 17828 3476 17834 3488
rect 19429 3485 19441 3488
rect 19475 3485 19487 3519
rect 19429 3479 19487 3485
rect 21082 3476 21088 3528
rect 21140 3516 21146 3528
rect 21269 3519 21327 3525
rect 21269 3516 21281 3519
rect 21140 3488 21281 3516
rect 21140 3476 21146 3488
rect 21269 3485 21281 3488
rect 21315 3485 21327 3519
rect 21269 3479 21327 3485
rect 14734 3448 14740 3460
rect 13924 3420 14740 3448
rect 14734 3408 14740 3420
rect 14792 3408 14798 3460
rect 19150 3408 19156 3460
rect 19208 3448 19214 3460
rect 21744 3448 21772 3547
rect 23201 3519 23259 3525
rect 23201 3516 23213 3519
rect 19208 3420 21772 3448
rect 22066 3488 23213 3516
rect 19208 3408 19214 3420
rect 3694 3340 3700 3392
rect 3752 3380 3758 3392
rect 3881 3383 3939 3389
rect 3881 3380 3893 3383
rect 3752 3352 3893 3380
rect 3752 3340 3758 3352
rect 3881 3349 3893 3352
rect 3927 3349 3939 3383
rect 3881 3343 3939 3349
rect 3970 3340 3976 3392
rect 4028 3380 4034 3392
rect 4157 3383 4215 3389
rect 4157 3380 4169 3383
rect 4028 3352 4169 3380
rect 4028 3340 4034 3352
rect 4157 3349 4169 3352
rect 4203 3349 4215 3383
rect 4157 3343 4215 3349
rect 4430 3340 4436 3392
rect 4488 3340 4494 3392
rect 4617 3383 4675 3389
rect 4617 3349 4629 3383
rect 4663 3380 4675 3383
rect 4798 3380 4804 3392
rect 4663 3352 4804 3380
rect 4663 3349 4675 3352
rect 4617 3343 4675 3349
rect 4798 3340 4804 3352
rect 4856 3340 4862 3392
rect 7193 3383 7251 3389
rect 7193 3349 7205 3383
rect 7239 3380 7251 3383
rect 7374 3380 7380 3392
rect 7239 3352 7380 3380
rect 7239 3349 7251 3352
rect 7193 3343 7251 3349
rect 7374 3340 7380 3352
rect 7432 3340 7438 3392
rect 9401 3383 9459 3389
rect 9401 3349 9413 3383
rect 9447 3380 9459 3383
rect 11882 3380 11888 3392
rect 9447 3352 11888 3380
rect 9447 3349 9459 3352
rect 9401 3343 9459 3349
rect 11882 3340 11888 3352
rect 11940 3340 11946 3392
rect 21450 3340 21456 3392
rect 21508 3380 21514 3392
rect 22066 3380 22094 3488
rect 23201 3485 23213 3488
rect 23247 3516 23259 3519
rect 23842 3516 23848 3528
rect 23247 3488 23848 3516
rect 23247 3485 23259 3488
rect 23201 3479 23259 3485
rect 23842 3476 23848 3488
rect 23900 3516 23906 3528
rect 24397 3519 24455 3525
rect 24397 3516 24409 3519
rect 23900 3488 24409 3516
rect 23900 3476 23906 3488
rect 24397 3485 24409 3488
rect 24443 3485 24455 3519
rect 24397 3479 24455 3485
rect 24765 3519 24823 3525
rect 24765 3485 24777 3519
rect 24811 3516 24823 3519
rect 25038 3516 25044 3528
rect 24811 3488 25044 3516
rect 24811 3485 24823 3488
rect 24765 3479 24823 3485
rect 25038 3476 25044 3488
rect 25096 3476 25102 3528
rect 21508 3352 22094 3380
rect 21508 3340 21514 3352
rect 1104 3290 25852 3312
rect 1104 3238 7950 3290
rect 8002 3238 8014 3290
rect 8066 3238 8078 3290
rect 8130 3238 8142 3290
rect 8194 3238 8206 3290
rect 8258 3238 17950 3290
rect 18002 3238 18014 3290
rect 18066 3238 18078 3290
rect 18130 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 25852 3290
rect 1104 3216 25852 3238
rect 2130 3136 2136 3188
rect 2188 3136 2194 3188
rect 4433 3179 4491 3185
rect 4433 3145 4445 3179
rect 4479 3145 4491 3179
rect 4433 3139 4491 3145
rect 5077 3179 5135 3185
rect 5077 3145 5089 3179
rect 5123 3176 5135 3179
rect 5166 3176 5172 3188
rect 5123 3148 5172 3176
rect 5123 3145 5135 3148
rect 5077 3139 5135 3145
rect 4448 3108 4476 3139
rect 5166 3136 5172 3148
rect 5224 3136 5230 3188
rect 5902 3136 5908 3188
rect 5960 3136 5966 3188
rect 23842 3136 23848 3188
rect 23900 3136 23906 3188
rect 10410 3108 10416 3120
rect 4448 3080 10416 3108
rect 10410 3068 10416 3080
rect 10468 3068 10474 3120
rect 1854 3000 1860 3052
rect 1912 3040 1918 3052
rect 1949 3043 2007 3049
rect 1949 3040 1961 3043
rect 1912 3012 1961 3040
rect 1912 3000 1918 3012
rect 1949 3009 1961 3012
rect 1995 3009 2007 3043
rect 1949 3003 2007 3009
rect 2869 3043 2927 3049
rect 2869 3009 2881 3043
rect 2915 3040 2927 3043
rect 3326 3040 3332 3052
rect 2915 3012 3332 3040
rect 2915 3009 2927 3012
rect 2869 3003 2927 3009
rect 3326 3000 3332 3012
rect 3384 3000 3390 3052
rect 3694 3000 3700 3052
rect 3752 3040 3758 3052
rect 3789 3043 3847 3049
rect 3789 3040 3801 3043
rect 3752 3012 3801 3040
rect 3752 3000 3758 3012
rect 3789 3009 3801 3012
rect 3835 3009 3847 3043
rect 3789 3003 3847 3009
rect 4249 3043 4307 3049
rect 4249 3009 4261 3043
rect 4295 3040 4307 3043
rect 4430 3040 4436 3052
rect 4295 3012 4436 3040
rect 4295 3009 4307 3012
rect 4249 3003 4307 3009
rect 4430 3000 4436 3012
rect 4488 3000 4494 3052
rect 5166 3000 5172 3052
rect 5224 3040 5230 3052
rect 5261 3043 5319 3049
rect 5261 3040 5273 3043
rect 5224 3012 5273 3040
rect 5224 3000 5230 3012
rect 5261 3009 5273 3012
rect 5307 3009 5319 3043
rect 5261 3003 5319 3009
rect 5813 3043 5871 3049
rect 5813 3009 5825 3043
rect 5859 3040 5871 3043
rect 5902 3040 5908 3052
rect 5859 3012 5908 3040
rect 5859 3009 5871 3012
rect 5813 3003 5871 3009
rect 5902 3000 5908 3012
rect 5960 3040 5966 3052
rect 6365 3043 6423 3049
rect 6365 3040 6377 3043
rect 5960 3012 6377 3040
rect 5960 3000 5966 3012
rect 6365 3009 6377 3012
rect 6411 3009 6423 3043
rect 6365 3003 6423 3009
rect 7377 3043 7435 3049
rect 7377 3009 7389 3043
rect 7423 3040 7435 3043
rect 7558 3040 7564 3052
rect 7423 3012 7564 3040
rect 7423 3009 7435 3012
rect 7377 3003 7435 3009
rect 7558 3000 7564 3012
rect 7616 3000 7622 3052
rect 8846 3000 8852 3052
rect 8904 3000 8910 3052
rect 10318 3000 10324 3052
rect 10376 3040 10382 3052
rect 10962 3040 10968 3052
rect 10376 3012 10968 3040
rect 10376 3000 10382 3012
rect 10962 3000 10968 3012
rect 11020 3040 11026 3052
rect 11149 3043 11207 3049
rect 11149 3040 11161 3043
rect 11020 3012 11161 3040
rect 11020 3000 11026 3012
rect 11149 3009 11161 3012
rect 11195 3009 11207 3043
rect 11149 3003 11207 3009
rect 12250 3000 12256 3052
rect 12308 3000 12314 3052
rect 14182 3000 14188 3052
rect 14240 3000 14246 3052
rect 16209 3043 16267 3049
rect 16209 3009 16221 3043
rect 16255 3040 16267 3043
rect 16482 3040 16488 3052
rect 16255 3012 16488 3040
rect 16255 3009 16267 3012
rect 16209 3003 16267 3009
rect 16482 3000 16488 3012
rect 16540 3000 16546 3052
rect 16850 3000 16856 3052
rect 16908 3000 16914 3052
rect 18690 3000 18696 3052
rect 18748 3000 18754 3052
rect 22002 3000 22008 3052
rect 22060 3040 22066 3052
rect 22830 3040 22836 3052
rect 22060 3012 22836 3040
rect 22060 3000 22066 3012
rect 22830 3000 22836 3012
rect 22888 3000 22894 3052
rect 25317 3043 25375 3049
rect 25317 3009 25329 3043
rect 25363 3009 25375 3043
rect 25317 3003 25375 3009
rect 3053 2975 3111 2981
rect 3053 2941 3065 2975
rect 3099 2972 3111 2975
rect 4706 2972 4712 2984
rect 3099 2944 4712 2972
rect 3099 2941 3111 2944
rect 3053 2935 3111 2941
rect 4706 2932 4712 2944
rect 4764 2932 4770 2984
rect 7101 2975 7159 2981
rect 7101 2972 7113 2975
rect 7024 2944 7113 2972
rect 3605 2907 3663 2913
rect 3605 2873 3617 2907
rect 3651 2904 3663 2907
rect 4614 2904 4620 2916
rect 3651 2876 4620 2904
rect 3651 2873 3663 2876
rect 3605 2867 3663 2873
rect 4614 2864 4620 2876
rect 4672 2864 4678 2916
rect 7024 2848 7052 2944
rect 7101 2941 7113 2944
rect 7147 2941 7159 2975
rect 7101 2935 7159 2941
rect 8478 2932 8484 2984
rect 8536 2972 8542 2984
rect 8573 2975 8631 2981
rect 8573 2972 8585 2975
rect 8536 2944 8585 2972
rect 8536 2932 8542 2944
rect 8573 2941 8585 2944
rect 8619 2941 8631 2975
rect 8573 2935 8631 2941
rect 10870 2932 10876 2984
rect 10928 2932 10934 2984
rect 11790 2932 11796 2984
rect 11848 2972 11854 2984
rect 12529 2975 12587 2981
rect 12529 2972 12541 2975
rect 11848 2944 12541 2972
rect 11848 2932 11854 2944
rect 12529 2941 12541 2944
rect 12575 2941 12587 2975
rect 12529 2935 12587 2941
rect 13630 2932 13636 2984
rect 13688 2932 13694 2984
rect 14734 2932 14740 2984
rect 14792 2972 14798 2984
rect 15013 2975 15071 2981
rect 15013 2972 15025 2975
rect 14792 2944 15025 2972
rect 14792 2932 14798 2944
rect 15013 2941 15025 2944
rect 15059 2941 15071 2975
rect 15013 2935 15071 2941
rect 15838 2932 15844 2984
rect 15896 2972 15902 2984
rect 17313 2975 17371 2981
rect 17313 2972 17325 2975
rect 15896 2944 17325 2972
rect 15896 2932 15902 2944
rect 17313 2941 17325 2944
rect 17359 2941 17371 2975
rect 17313 2935 17371 2941
rect 19153 2975 19211 2981
rect 19153 2941 19165 2975
rect 19199 2941 19211 2975
rect 19153 2935 19211 2941
rect 16574 2864 16580 2916
rect 16632 2904 16638 2916
rect 19168 2904 19196 2935
rect 20530 2932 20536 2984
rect 20588 2972 20594 2984
rect 23934 2972 23940 2984
rect 20588 2944 23940 2972
rect 20588 2932 20594 2944
rect 23934 2932 23940 2944
rect 23992 2932 23998 2984
rect 16632 2876 19196 2904
rect 16632 2864 16638 2876
rect 19978 2864 19984 2916
rect 20036 2904 20042 2916
rect 21726 2904 21732 2916
rect 20036 2876 21732 2904
rect 20036 2864 20042 2876
rect 21726 2864 21732 2876
rect 21784 2864 21790 2916
rect 23566 2864 23572 2916
rect 23624 2904 23630 2916
rect 25332 2904 25360 3003
rect 25406 2904 25412 2916
rect 23624 2876 25412 2904
rect 23624 2864 23630 2876
rect 25406 2864 25412 2876
rect 25464 2864 25470 2916
rect 1486 2796 1492 2848
rect 1544 2796 1550 2848
rect 1673 2839 1731 2845
rect 1673 2805 1685 2839
rect 1719 2836 1731 2839
rect 1854 2836 1860 2848
rect 1719 2808 1860 2836
rect 1719 2805 1731 2808
rect 1673 2799 1731 2805
rect 1854 2796 1860 2808
rect 1912 2796 1918 2848
rect 6825 2839 6883 2845
rect 6825 2805 6837 2839
rect 6871 2836 6883 2839
rect 7006 2836 7012 2848
rect 6871 2808 7012 2836
rect 6871 2805 6883 2808
rect 6825 2799 6883 2805
rect 7006 2796 7012 2808
rect 7064 2796 7070 2848
rect 7834 2796 7840 2848
rect 7892 2836 7898 2848
rect 8205 2839 8263 2845
rect 8205 2836 8217 2839
rect 7892 2808 8217 2836
rect 7892 2796 7898 2808
rect 8205 2805 8217 2808
rect 8251 2805 8263 2839
rect 8205 2799 8263 2805
rect 9582 2796 9588 2848
rect 9640 2836 9646 2848
rect 9677 2839 9735 2845
rect 9677 2836 9689 2839
rect 9640 2808 9689 2836
rect 9640 2796 9646 2808
rect 9677 2805 9689 2808
rect 9723 2805 9735 2839
rect 9677 2799 9735 2805
rect 9950 2796 9956 2848
rect 10008 2796 10014 2848
rect 17310 2796 17316 2848
rect 17368 2836 17374 2848
rect 18322 2836 18328 2848
rect 17368 2808 18328 2836
rect 17368 2796 17374 2808
rect 18322 2796 18328 2808
rect 18380 2796 18386 2848
rect 18782 2796 18788 2848
rect 18840 2836 18846 2848
rect 19886 2836 19892 2848
rect 18840 2808 19892 2836
rect 18840 2796 18846 2808
rect 19886 2796 19892 2808
rect 19944 2796 19950 2848
rect 20990 2796 20996 2848
rect 21048 2836 21054 2848
rect 22278 2836 22284 2848
rect 21048 2808 22284 2836
rect 21048 2796 21054 2808
rect 22278 2796 22284 2808
rect 22336 2796 22342 2848
rect 1104 2746 25852 2768
rect 1104 2694 2950 2746
rect 3002 2694 3014 2746
rect 3066 2694 3078 2746
rect 3130 2694 3142 2746
rect 3194 2694 3206 2746
rect 3258 2694 12950 2746
rect 13002 2694 13014 2746
rect 13066 2694 13078 2746
rect 13130 2694 13142 2746
rect 13194 2694 13206 2746
rect 13258 2694 22950 2746
rect 23002 2694 23014 2746
rect 23066 2694 23078 2746
rect 23130 2694 23142 2746
rect 23194 2694 23206 2746
rect 23258 2694 25852 2746
rect 1104 2672 25852 2694
rect 10778 2632 10784 2644
rect 4448 2604 10784 2632
rect 2041 2567 2099 2573
rect 2041 2533 2053 2567
rect 2087 2564 2099 2567
rect 2087 2536 4384 2564
rect 2087 2533 2099 2536
rect 2041 2527 2099 2533
rect 2590 2456 2596 2508
rect 2648 2496 2654 2508
rect 3421 2499 3479 2505
rect 3421 2496 3433 2499
rect 2648 2468 3433 2496
rect 2648 2456 2654 2468
rect 3421 2465 3433 2468
rect 3467 2496 3479 2499
rect 3970 2496 3976 2508
rect 3467 2468 3976 2496
rect 3467 2465 3479 2468
rect 3421 2459 3479 2465
rect 3970 2456 3976 2468
rect 4028 2456 4034 2508
rect 1581 2431 1639 2437
rect 1581 2397 1593 2431
rect 1627 2428 1639 2431
rect 1857 2431 1915 2437
rect 1857 2428 1869 2431
rect 1627 2400 1869 2428
rect 1627 2397 1639 2400
rect 1581 2391 1639 2397
rect 1857 2397 1869 2400
rect 1903 2428 1915 2431
rect 2222 2428 2228 2440
rect 1903 2400 2228 2428
rect 1903 2397 1915 2400
rect 1857 2391 1915 2397
rect 2222 2388 2228 2400
rect 2280 2388 2286 2440
rect 3142 2388 3148 2440
rect 3200 2388 3206 2440
rect 4157 2431 4215 2437
rect 4157 2428 4169 2431
rect 4080 2400 4169 2428
rect 4080 2304 4108 2400
rect 4157 2397 4169 2400
rect 4203 2397 4215 2431
rect 4356 2428 4384 2536
rect 4448 2505 4476 2604
rect 10778 2592 10784 2604
rect 10836 2592 10842 2644
rect 11885 2635 11943 2641
rect 11885 2601 11897 2635
rect 11931 2632 11943 2635
rect 15378 2632 15384 2644
rect 11931 2604 15384 2632
rect 11931 2601 11943 2604
rect 11885 2595 11943 2601
rect 15378 2592 15384 2604
rect 15436 2592 15442 2644
rect 24673 2635 24731 2641
rect 24673 2601 24685 2635
rect 24719 2632 24731 2635
rect 24946 2632 24952 2644
rect 24719 2604 24952 2632
rect 24719 2601 24731 2604
rect 24673 2595 24731 2601
rect 24946 2592 24952 2604
rect 25004 2592 25010 2644
rect 25406 2592 25412 2644
rect 25464 2592 25470 2644
rect 5813 2567 5871 2573
rect 5813 2533 5825 2567
rect 5859 2564 5871 2567
rect 7285 2567 7343 2573
rect 5859 2536 7144 2564
rect 5859 2533 5871 2536
rect 5813 2527 5871 2533
rect 4433 2499 4491 2505
rect 4433 2465 4445 2499
rect 4479 2465 4491 2499
rect 6914 2496 6920 2508
rect 4433 2459 4491 2465
rect 4540 2468 6920 2496
rect 4540 2428 4568 2468
rect 6914 2456 6920 2468
rect 6972 2456 6978 2508
rect 4356 2400 4568 2428
rect 5997 2431 6055 2437
rect 4157 2391 4215 2397
rect 5997 2397 6009 2431
rect 6043 2428 6055 2431
rect 7116 2428 7144 2536
rect 7285 2533 7297 2567
rect 7331 2564 7343 2567
rect 9490 2564 9496 2576
rect 7331 2536 9496 2564
rect 7331 2533 7343 2536
rect 7285 2527 7343 2533
rect 9490 2524 9496 2536
rect 9548 2524 9554 2576
rect 11606 2564 11612 2576
rect 9600 2536 11612 2564
rect 9600 2496 9628 2536
rect 11606 2524 11612 2536
rect 11664 2524 11670 2576
rect 18966 2524 18972 2576
rect 19024 2564 19030 2576
rect 19024 2536 22048 2564
rect 19024 2524 19030 2536
rect 7300 2468 9628 2496
rect 10689 2499 10747 2505
rect 7300 2428 7328 2468
rect 10689 2465 10701 2499
rect 10735 2496 10747 2499
rect 12158 2496 12164 2508
rect 10735 2468 12164 2496
rect 10735 2465 10747 2468
rect 10689 2459 10747 2465
rect 12158 2456 12164 2468
rect 12216 2456 12222 2508
rect 14093 2499 14151 2505
rect 14093 2496 14105 2499
rect 12268 2468 14105 2496
rect 6043 2400 6500 2428
rect 7116 2400 7328 2428
rect 6043 2397 6055 2400
rect 5997 2391 6055 2397
rect 3881 2295 3939 2301
rect 3881 2261 3893 2295
rect 3927 2292 3939 2295
rect 4062 2292 4068 2304
rect 3927 2264 4068 2292
rect 3927 2261 3939 2264
rect 3881 2255 3939 2261
rect 4062 2252 4068 2264
rect 4120 2252 4126 2304
rect 5166 2252 5172 2304
rect 5224 2292 5230 2304
rect 6472 2301 6500 2400
rect 8294 2388 8300 2440
rect 8352 2388 8358 2440
rect 8573 2431 8631 2437
rect 8573 2397 8585 2431
rect 8619 2428 8631 2431
rect 8619 2400 9076 2428
rect 8619 2397 8631 2400
rect 8573 2391 8631 2397
rect 6733 2363 6791 2369
rect 6733 2329 6745 2363
rect 6779 2360 6791 2363
rect 7101 2363 7159 2369
rect 7101 2360 7113 2363
rect 6779 2332 7113 2360
rect 6779 2329 6791 2332
rect 6733 2323 6791 2329
rect 7101 2329 7113 2332
rect 7147 2360 7159 2363
rect 7742 2360 7748 2372
rect 7147 2332 7748 2360
rect 7147 2329 7159 2332
rect 7101 2323 7159 2329
rect 7742 2320 7748 2332
rect 7800 2320 7806 2372
rect 5353 2295 5411 2301
rect 5353 2292 5365 2295
rect 5224 2264 5365 2292
rect 5224 2252 5230 2264
rect 5353 2261 5365 2264
rect 5399 2261 5411 2295
rect 5353 2255 5411 2261
rect 6457 2295 6515 2301
rect 6457 2261 6469 2295
rect 6503 2292 6515 2295
rect 6638 2292 6644 2304
rect 6503 2264 6644 2292
rect 6503 2261 6515 2264
rect 6457 2255 6515 2261
rect 6638 2252 6644 2264
rect 6696 2252 6702 2304
rect 6914 2252 6920 2304
rect 6972 2292 6978 2304
rect 7650 2292 7656 2304
rect 6972 2264 7656 2292
rect 6972 2252 6978 2264
rect 7650 2252 7656 2264
rect 7708 2252 7714 2304
rect 8478 2252 8484 2304
rect 8536 2292 8542 2304
rect 8941 2295 8999 2301
rect 8941 2292 8953 2295
rect 8536 2264 8953 2292
rect 8536 2252 8542 2264
rect 8941 2261 8953 2264
rect 8987 2261 8999 2295
rect 9048 2292 9076 2400
rect 11054 2388 11060 2440
rect 11112 2388 11118 2440
rect 11422 2388 11428 2440
rect 11480 2428 11486 2440
rect 11701 2431 11759 2437
rect 11701 2428 11713 2431
rect 11480 2400 11713 2428
rect 11480 2388 11486 2400
rect 11701 2397 11713 2400
rect 11747 2428 11759 2431
rect 12268 2428 12296 2468
rect 14093 2465 14105 2468
rect 14139 2465 14151 2499
rect 14093 2459 14151 2465
rect 15102 2456 15108 2508
rect 15160 2496 15166 2508
rect 17313 2499 17371 2505
rect 17313 2496 17325 2499
rect 15160 2468 17325 2496
rect 15160 2456 15166 2468
rect 17313 2465 17325 2468
rect 17359 2465 17371 2499
rect 19889 2499 19947 2505
rect 19889 2496 19901 2499
rect 17313 2459 17371 2465
rect 17972 2468 19901 2496
rect 11747 2400 12296 2428
rect 11747 2397 11759 2400
rect 11701 2391 11759 2397
rect 12342 2388 12348 2440
rect 12400 2388 12406 2440
rect 15654 2388 15660 2440
rect 15712 2388 15718 2440
rect 15746 2388 15752 2440
rect 15804 2428 15810 2440
rect 16853 2431 16911 2437
rect 16853 2428 16865 2431
rect 15804 2400 16865 2428
rect 15804 2388 15810 2400
rect 16853 2397 16865 2400
rect 16899 2397 16911 2431
rect 16853 2391 16911 2397
rect 16942 2388 16948 2440
rect 17000 2428 17006 2440
rect 17972 2428 18000 2468
rect 19889 2465 19901 2468
rect 19935 2465 19947 2499
rect 19889 2459 19947 2465
rect 22020 2437 22048 2536
rect 22465 2499 22523 2505
rect 22465 2465 22477 2499
rect 22511 2465 22523 2499
rect 22465 2459 22523 2465
rect 19429 2431 19487 2437
rect 19429 2428 19441 2431
rect 17000 2400 18000 2428
rect 18064 2400 19441 2428
rect 17000 2388 17006 2400
rect 13262 2320 13268 2372
rect 13320 2320 13326 2372
rect 14366 2320 14372 2372
rect 14424 2360 14430 2372
rect 14645 2363 14703 2369
rect 14645 2360 14657 2363
rect 14424 2332 14657 2360
rect 14424 2320 14430 2332
rect 14645 2329 14657 2332
rect 14691 2329 14703 2363
rect 14645 2323 14703 2329
rect 17402 2320 17408 2372
rect 17460 2360 17466 2372
rect 18064 2360 18092 2400
rect 19429 2397 19441 2400
rect 19475 2397 19487 2431
rect 19429 2391 19487 2397
rect 22005 2431 22063 2437
rect 22005 2397 22017 2431
rect 22051 2397 22063 2431
rect 22005 2391 22063 2397
rect 17460 2332 18092 2360
rect 17460 2320 17466 2332
rect 18506 2320 18512 2372
rect 18564 2360 18570 2372
rect 22480 2360 22508 2459
rect 24302 2388 24308 2440
rect 24360 2428 24366 2440
rect 24857 2431 24915 2437
rect 24857 2428 24869 2431
rect 24360 2400 24869 2428
rect 24360 2388 24366 2400
rect 24857 2397 24869 2400
rect 24903 2428 24915 2431
rect 25133 2431 25191 2437
rect 25133 2428 25145 2431
rect 24903 2400 25145 2428
rect 24903 2397 24915 2400
rect 24857 2391 24915 2397
rect 25133 2397 25145 2400
rect 25179 2397 25191 2431
rect 25133 2391 25191 2397
rect 18564 2332 22508 2360
rect 18564 2320 18570 2332
rect 9217 2295 9275 2301
rect 9217 2292 9229 2295
rect 9048 2264 9229 2292
rect 8941 2255 8999 2261
rect 9217 2261 9229 2264
rect 9263 2292 9275 2295
rect 10962 2292 10968 2304
rect 9263 2264 10968 2292
rect 9263 2261 9275 2264
rect 9217 2255 9275 2261
rect 10962 2252 10968 2264
rect 11020 2252 11026 2304
rect 1104 2202 25852 2224
rect 1104 2150 7950 2202
rect 8002 2150 8014 2202
rect 8066 2150 8078 2202
rect 8130 2150 8142 2202
rect 8194 2150 8206 2202
rect 8258 2150 17950 2202
rect 18002 2150 18014 2202
rect 18066 2150 18078 2202
rect 18130 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 25852 2202
rect 1104 2128 25852 2150
rect 3142 2048 3148 2100
rect 3200 2088 3206 2100
rect 9030 2088 9036 2100
rect 3200 2060 9036 2088
rect 3200 2048 3206 2060
rect 9030 2048 9036 2060
rect 9088 2048 9094 2100
rect 8294 1980 8300 2032
rect 8352 2020 8358 2032
rect 15930 2020 15936 2032
rect 8352 1992 15936 2020
rect 8352 1980 8358 1992
rect 15930 1980 15936 1992
rect 15988 1980 15994 2032
<< via1 >>
rect 7950 54374 8002 54426
rect 8014 54374 8066 54426
rect 8078 54374 8130 54426
rect 8142 54374 8194 54426
rect 8206 54374 8258 54426
rect 17950 54374 18002 54426
rect 18014 54374 18066 54426
rect 18078 54374 18130 54426
rect 18142 54374 18194 54426
rect 18206 54374 18258 54426
rect 13820 54315 13872 54324
rect 13820 54281 13829 54315
rect 13829 54281 13863 54315
rect 13863 54281 13872 54315
rect 13820 54272 13872 54281
rect 14556 54272 14608 54324
rect 19340 54272 19392 54324
rect 5908 54136 5960 54188
rect 8484 54204 8536 54256
rect 10876 54247 10928 54256
rect 10876 54213 10885 54247
rect 10885 54213 10919 54247
rect 10919 54213 10928 54247
rect 10876 54204 10928 54213
rect 5356 54068 5408 54120
rect 7196 54068 7248 54120
rect 9404 54068 9456 54120
rect 9864 54179 9916 54188
rect 9864 54145 9873 54179
rect 9873 54145 9907 54179
rect 9907 54145 9916 54179
rect 9864 54136 9916 54145
rect 12072 54179 12124 54188
rect 12072 54145 12081 54179
rect 12081 54145 12115 54179
rect 12115 54145 12124 54179
rect 12072 54136 12124 54145
rect 14924 54204 14976 54256
rect 16028 54204 16080 54256
rect 16672 54204 16724 54256
rect 15292 54136 15344 54188
rect 15844 54136 15896 54188
rect 17500 54204 17552 54256
rect 18420 54247 18472 54256
rect 18420 54213 18429 54247
rect 18429 54213 18463 54247
rect 18463 54213 18472 54247
rect 18420 54204 18472 54213
rect 17132 54136 17184 54188
rect 11888 54068 11940 54120
rect 11980 54068 12032 54120
rect 18604 54136 18656 54188
rect 19340 54136 19392 54188
rect 20076 54204 20128 54256
rect 20720 54204 20772 54256
rect 22652 54204 22704 54256
rect 21180 54136 21232 54188
rect 21824 54136 21876 54188
rect 23940 54179 23992 54188
rect 23940 54145 23949 54179
rect 23949 54145 23983 54179
rect 23983 54145 23992 54179
rect 23940 54136 23992 54145
rect 24124 54068 24176 54120
rect 15660 54043 15712 54052
rect 15660 54009 15669 54043
rect 15669 54009 15703 54043
rect 15703 54009 15712 54043
rect 15660 54000 15712 54009
rect 18604 54043 18656 54052
rect 18604 54009 18613 54043
rect 18613 54009 18647 54043
rect 18647 54009 18656 54043
rect 18604 54000 18656 54009
rect 21732 54000 21784 54052
rect 15108 53932 15160 53984
rect 16488 53932 16540 53984
rect 16948 53932 17000 53984
rect 17776 53932 17828 53984
rect 19616 53975 19668 53984
rect 19616 53941 19625 53975
rect 19625 53941 19659 53975
rect 19659 53941 19668 53975
rect 19616 53932 19668 53941
rect 20536 53932 20588 53984
rect 21180 53932 21232 53984
rect 22008 53975 22060 53984
rect 22008 53941 22017 53975
rect 22017 53941 22051 53975
rect 22051 53941 22060 53975
rect 22008 53932 22060 53941
rect 2950 53830 3002 53882
rect 3014 53830 3066 53882
rect 3078 53830 3130 53882
rect 3142 53830 3194 53882
rect 3206 53830 3258 53882
rect 12950 53830 13002 53882
rect 13014 53830 13066 53882
rect 13078 53830 13130 53882
rect 13142 53830 13194 53882
rect 13206 53830 13258 53882
rect 22950 53830 23002 53882
rect 23014 53830 23066 53882
rect 23078 53830 23130 53882
rect 23142 53830 23194 53882
rect 23206 53830 23258 53882
rect 14924 53728 14976 53780
rect 15568 53728 15620 53780
rect 20444 53728 20496 53780
rect 4620 53592 4672 53644
rect 7564 53592 7616 53644
rect 8300 53635 8352 53644
rect 8300 53601 8309 53635
rect 8309 53601 8343 53635
rect 8343 53601 8352 53635
rect 8300 53592 8352 53601
rect 10508 53635 10560 53644
rect 10508 53601 10517 53635
rect 10517 53601 10551 53635
rect 10551 53601 10560 53635
rect 10508 53592 10560 53601
rect 11612 53592 11664 53644
rect 25596 53660 25648 53712
rect 23296 53592 23348 53644
rect 6184 53524 6236 53576
rect 6644 53567 6696 53576
rect 6644 53533 6653 53567
rect 6653 53533 6687 53567
rect 6687 53533 6696 53567
rect 6644 53524 6696 53533
rect 7380 53567 7432 53576
rect 7380 53533 7389 53567
rect 7389 53533 7423 53567
rect 7423 53533 7432 53567
rect 7380 53524 7432 53533
rect 9036 53524 9088 53576
rect 9680 53524 9732 53576
rect 11060 53567 11112 53576
rect 11060 53533 11069 53567
rect 11069 53533 11103 53567
rect 11103 53533 11112 53567
rect 11060 53524 11112 53533
rect 11888 53567 11940 53576
rect 11888 53533 11897 53567
rect 11897 53533 11931 53567
rect 11931 53533 11940 53567
rect 11888 53524 11940 53533
rect 13820 53524 13872 53576
rect 14188 53524 14240 53576
rect 15568 53524 15620 53576
rect 16396 53524 16448 53576
rect 16764 53524 16816 53576
rect 17868 53524 17920 53576
rect 18328 53524 18380 53576
rect 18972 53524 19024 53576
rect 20444 53524 20496 53576
rect 20812 53524 20864 53576
rect 21548 53524 21600 53576
rect 24032 53567 24084 53576
rect 24032 53533 24041 53567
rect 24041 53533 24075 53567
rect 24075 53533 24084 53567
rect 24032 53524 24084 53533
rect 3792 53431 3844 53440
rect 3792 53397 3801 53431
rect 3801 53397 3835 53431
rect 3835 53397 3844 53431
rect 3792 53388 3844 53397
rect 13636 53388 13688 53440
rect 15752 53388 15804 53440
rect 15936 53431 15988 53440
rect 15936 53397 15945 53431
rect 15945 53397 15979 53431
rect 15979 53397 15988 53431
rect 15936 53388 15988 53397
rect 17040 53388 17092 53440
rect 17408 53431 17460 53440
rect 17408 53397 17417 53431
rect 17417 53397 17451 53431
rect 17451 53397 17460 53431
rect 17408 53388 17460 53397
rect 18512 53388 18564 53440
rect 18696 53431 18748 53440
rect 18696 53397 18705 53431
rect 18705 53397 18739 53431
rect 18739 53397 18748 53431
rect 18696 53388 18748 53397
rect 19524 53431 19576 53440
rect 19524 53397 19533 53431
rect 19533 53397 19567 53431
rect 19567 53397 19576 53431
rect 19524 53388 19576 53397
rect 21272 53388 21324 53440
rect 21456 53431 21508 53440
rect 21456 53397 21465 53431
rect 21465 53397 21499 53431
rect 21499 53397 21508 53431
rect 21456 53388 21508 53397
rect 21548 53388 21600 53440
rect 24492 53388 24544 53440
rect 25320 53388 25372 53440
rect 7950 53286 8002 53338
rect 8014 53286 8066 53338
rect 8078 53286 8130 53338
rect 8142 53286 8194 53338
rect 8206 53286 8258 53338
rect 17950 53286 18002 53338
rect 18014 53286 18066 53338
rect 18078 53286 18130 53338
rect 18142 53286 18194 53338
rect 18206 53286 18258 53338
rect 2780 53184 2832 53236
rect 15844 53184 15896 53236
rect 16396 53227 16448 53236
rect 16396 53193 16405 53227
rect 16405 53193 16439 53227
rect 16439 53193 16448 53227
rect 16396 53184 16448 53193
rect 16672 53227 16724 53236
rect 16672 53193 16681 53227
rect 16681 53193 16715 53227
rect 16715 53193 16724 53227
rect 16672 53184 16724 53193
rect 16764 53184 16816 53236
rect 17868 53227 17920 53236
rect 17868 53193 17877 53227
rect 17877 53193 17911 53227
rect 17911 53193 17920 53227
rect 17868 53184 17920 53193
rect 18328 53184 18380 53236
rect 19340 53227 19392 53236
rect 19340 53193 19349 53227
rect 19349 53193 19383 53227
rect 19383 53193 19392 53227
rect 19340 53184 19392 53193
rect 20720 53227 20772 53236
rect 20720 53193 20729 53227
rect 20729 53193 20763 53227
rect 20763 53193 20772 53227
rect 20720 53184 20772 53193
rect 20812 53184 20864 53236
rect 21640 53184 21692 53236
rect 6368 53116 6420 53168
rect 12716 53116 12768 53168
rect 18420 53116 18472 53168
rect 5816 53091 5868 53100
rect 5816 53057 5825 53091
rect 5825 53057 5859 53091
rect 5859 53057 5868 53091
rect 5816 53048 5868 53057
rect 6736 53048 6788 53100
rect 9128 53091 9180 53100
rect 9128 53057 9137 53091
rect 9137 53057 9171 53091
rect 9171 53057 9180 53091
rect 9128 53048 9180 53057
rect 9404 53048 9456 53100
rect 10692 53048 10744 53100
rect 13452 53048 13504 53100
rect 19708 53048 19760 53100
rect 21916 53048 21968 53100
rect 22284 53048 22336 53100
rect 24952 53048 25004 53100
rect 4252 52980 4304 53032
rect 5724 52980 5776 53032
rect 8668 53023 8720 53032
rect 8668 52989 8677 53023
rect 8677 52989 8711 53023
rect 8711 52989 8720 53023
rect 8668 52980 8720 52989
rect 10140 52980 10192 53032
rect 11244 52980 11296 53032
rect 24860 53023 24912 53032
rect 24860 52989 24869 53023
rect 24869 52989 24903 53023
rect 24903 52989 24912 53023
rect 24860 52980 24912 52989
rect 4068 52844 4120 52896
rect 6000 52844 6052 52896
rect 12808 52844 12860 52896
rect 14372 52887 14424 52896
rect 14372 52853 14381 52887
rect 14381 52853 14415 52887
rect 14415 52853 14424 52887
rect 14372 52844 14424 52853
rect 19800 52887 19852 52896
rect 19800 52853 19809 52887
rect 19809 52853 19843 52887
rect 19843 52853 19852 52887
rect 19800 52844 19852 52853
rect 22192 52887 22244 52896
rect 22192 52853 22201 52887
rect 22201 52853 22235 52887
rect 22235 52853 22244 52887
rect 22192 52844 22244 52853
rect 22744 52887 22796 52896
rect 22744 52853 22753 52887
rect 22753 52853 22787 52887
rect 22787 52853 22796 52887
rect 22744 52844 22796 52853
rect 23480 52844 23532 52896
rect 25228 52844 25280 52896
rect 2950 52742 3002 52794
rect 3014 52742 3066 52794
rect 3078 52742 3130 52794
rect 3142 52742 3194 52794
rect 3206 52742 3258 52794
rect 12950 52742 13002 52794
rect 13014 52742 13066 52794
rect 13078 52742 13130 52794
rect 13142 52742 13194 52794
rect 13206 52742 13258 52794
rect 22950 52742 23002 52794
rect 23014 52742 23066 52794
rect 23078 52742 23130 52794
rect 23142 52742 23194 52794
rect 23206 52742 23258 52794
rect 940 52640 992 52692
rect 4344 52640 4396 52692
rect 12072 52640 12124 52692
rect 13452 52640 13504 52692
rect 21824 52683 21876 52692
rect 21824 52649 21833 52683
rect 21833 52649 21867 52683
rect 21867 52649 21876 52683
rect 21824 52640 21876 52649
rect 23940 52683 23992 52692
rect 23940 52649 23949 52683
rect 23949 52649 23983 52683
rect 23983 52649 23992 52683
rect 23940 52640 23992 52649
rect 1216 52572 1268 52624
rect 3792 52572 3844 52624
rect 3332 52504 3384 52556
rect 13360 52572 13412 52624
rect 24768 52572 24820 52624
rect 25964 52572 26016 52624
rect 4436 52504 4488 52556
rect 6092 52547 6144 52556
rect 6092 52513 6101 52547
rect 6101 52513 6135 52547
rect 6135 52513 6144 52547
rect 6092 52504 6144 52513
rect 6460 52504 6512 52556
rect 6920 52504 6972 52556
rect 7840 52547 7892 52556
rect 7840 52513 7849 52547
rect 7849 52513 7883 52547
rect 7883 52513 7892 52547
rect 7840 52504 7892 52513
rect 9772 52504 9824 52556
rect 4528 52436 4580 52488
rect 6552 52479 6604 52488
rect 6552 52445 6561 52479
rect 6561 52445 6595 52479
rect 6595 52445 6604 52479
rect 6552 52436 6604 52445
rect 9496 52436 9548 52488
rect 9588 52436 9640 52488
rect 11796 52479 11848 52488
rect 11796 52445 11805 52479
rect 11805 52445 11839 52479
rect 11839 52445 11848 52479
rect 11796 52436 11848 52445
rect 12348 52436 12400 52488
rect 13452 52479 13504 52488
rect 13452 52445 13461 52479
rect 13461 52445 13495 52479
rect 13495 52445 13504 52479
rect 13452 52436 13504 52445
rect 23480 52436 23532 52488
rect 24216 52436 24268 52488
rect 25228 52436 25280 52488
rect 12716 52368 12768 52420
rect 23296 52343 23348 52352
rect 23296 52309 23305 52343
rect 23305 52309 23339 52343
rect 23339 52309 23348 52343
rect 23296 52300 23348 52309
rect 24584 52343 24636 52352
rect 24584 52309 24593 52343
rect 24593 52309 24627 52343
rect 24627 52309 24636 52343
rect 24584 52300 24636 52309
rect 7950 52198 8002 52250
rect 8014 52198 8066 52250
rect 8078 52198 8130 52250
rect 8142 52198 8194 52250
rect 8206 52198 8258 52250
rect 17950 52198 18002 52250
rect 18014 52198 18066 52250
rect 18078 52198 18130 52250
rect 18142 52198 18194 52250
rect 18206 52198 18258 52250
rect 11888 52139 11940 52148
rect 11888 52105 11897 52139
rect 11897 52105 11931 52139
rect 11931 52105 11940 52139
rect 11888 52096 11940 52105
rect 12348 52139 12400 52148
rect 12348 52105 12357 52139
rect 12357 52105 12391 52139
rect 12391 52105 12400 52139
rect 12348 52096 12400 52105
rect 23480 52139 23532 52148
rect 23480 52105 23489 52139
rect 23489 52105 23523 52139
rect 23523 52105 23532 52139
rect 23480 52096 23532 52105
rect 24584 52096 24636 52148
rect 4988 52071 5040 52080
rect 4988 52037 4997 52071
rect 4997 52037 5031 52071
rect 5031 52037 5040 52071
rect 4988 52028 5040 52037
rect 5356 51960 5408 52012
rect 7196 52028 7248 52080
rect 7012 52003 7064 52012
rect 7012 51969 7021 52003
rect 7021 51969 7055 52003
rect 7055 51969 7064 52003
rect 7012 51960 7064 51969
rect 10140 51960 10192 52012
rect 11612 51960 11664 52012
rect 24400 51960 24452 52012
rect 24676 51960 24728 52012
rect 25228 52003 25280 52012
rect 25228 51969 25237 52003
rect 25237 51969 25271 52003
rect 25271 51969 25280 52003
rect 25228 51960 25280 51969
rect 3516 51935 3568 51944
rect 3516 51901 3525 51935
rect 3525 51901 3559 51935
rect 3559 51901 3568 51935
rect 3516 51892 3568 51901
rect 7104 51892 7156 51944
rect 9680 51935 9732 51944
rect 9680 51901 9689 51935
rect 9689 51901 9723 51935
rect 9723 51901 9732 51935
rect 9680 51892 9732 51901
rect 24400 51799 24452 51808
rect 24400 51765 24409 51799
rect 24409 51765 24443 51799
rect 24443 51765 24452 51799
rect 24400 51756 24452 51765
rect 25688 51756 25740 51808
rect 2950 51654 3002 51706
rect 3014 51654 3066 51706
rect 3078 51654 3130 51706
rect 3142 51654 3194 51706
rect 3206 51654 3258 51706
rect 12950 51654 13002 51706
rect 13014 51654 13066 51706
rect 13078 51654 13130 51706
rect 13142 51654 13194 51706
rect 13206 51654 13258 51706
rect 22950 51654 23002 51706
rect 23014 51654 23066 51706
rect 23078 51654 23130 51706
rect 23142 51654 23194 51706
rect 23206 51654 23258 51706
rect 5908 51595 5960 51604
rect 5908 51561 5917 51595
rect 5917 51561 5951 51595
rect 5951 51561 5960 51595
rect 5908 51552 5960 51561
rect 24676 51595 24728 51604
rect 24676 51561 24685 51595
rect 24685 51561 24719 51595
rect 24719 51561 24728 51595
rect 24676 51552 24728 51561
rect 2412 51459 2464 51468
rect 2412 51425 2421 51459
rect 2421 51425 2455 51459
rect 2455 51425 2464 51459
rect 2412 51416 2464 51425
rect 4160 51459 4212 51468
rect 4160 51425 4169 51459
rect 4169 51425 4203 51459
rect 4203 51425 4212 51459
rect 4160 51416 4212 51425
rect 6920 51459 6972 51468
rect 6920 51425 6929 51459
rect 6929 51425 6963 51459
rect 6963 51425 6972 51459
rect 6920 51416 6972 51425
rect 6000 51348 6052 51400
rect 7104 51348 7156 51400
rect 7748 51391 7800 51400
rect 7748 51357 7757 51391
rect 7757 51357 7791 51391
rect 7791 51357 7800 51391
rect 7748 51348 7800 51357
rect 24768 51484 24820 51536
rect 25320 51391 25372 51400
rect 25320 51357 25329 51391
rect 25329 51357 25363 51391
rect 25363 51357 25372 51391
rect 25320 51348 25372 51357
rect 6736 51280 6788 51332
rect 20996 51212 21048 51264
rect 22744 51212 22796 51264
rect 23848 51255 23900 51264
rect 23848 51221 23857 51255
rect 23857 51221 23891 51255
rect 23891 51221 23900 51255
rect 23848 51212 23900 51221
rect 25596 51212 25648 51264
rect 7950 51110 8002 51162
rect 8014 51110 8066 51162
rect 8078 51110 8130 51162
rect 8142 51110 8194 51162
rect 8206 51110 8258 51162
rect 17950 51110 18002 51162
rect 18014 51110 18066 51162
rect 18078 51110 18130 51162
rect 18142 51110 18194 51162
rect 18206 51110 18258 51162
rect 9864 51051 9916 51060
rect 9864 51017 9873 51051
rect 9873 51017 9907 51051
rect 9907 51017 9916 51051
rect 9864 51008 9916 51017
rect 10692 51051 10744 51060
rect 10692 51017 10701 51051
rect 10701 51017 10735 51051
rect 10735 51017 10744 51051
rect 10692 51008 10744 51017
rect 2872 50940 2924 50992
rect 6736 50983 6788 50992
rect 6736 50949 6745 50983
rect 6745 50949 6779 50983
rect 6779 50949 6788 50983
rect 6736 50940 6788 50949
rect 1124 50804 1176 50856
rect 4160 50915 4212 50924
rect 4160 50881 4169 50915
rect 4169 50881 4203 50915
rect 4203 50881 4212 50915
rect 4160 50872 4212 50881
rect 8300 50872 8352 50924
rect 8576 50872 8628 50924
rect 9956 50872 10008 50924
rect 25320 50915 25372 50924
rect 25320 50881 25329 50915
rect 25329 50881 25363 50915
rect 25363 50881 25372 50915
rect 25320 50872 25372 50881
rect 6920 50736 6972 50788
rect 25136 50711 25188 50720
rect 25136 50677 25145 50711
rect 25145 50677 25179 50711
rect 25179 50677 25188 50711
rect 25136 50668 25188 50677
rect 2950 50566 3002 50618
rect 3014 50566 3066 50618
rect 3078 50566 3130 50618
rect 3142 50566 3194 50618
rect 3206 50566 3258 50618
rect 12950 50566 13002 50618
rect 13014 50566 13066 50618
rect 13078 50566 13130 50618
rect 13142 50566 13194 50618
rect 13206 50566 13258 50618
rect 22950 50566 23002 50618
rect 23014 50566 23066 50618
rect 23078 50566 23130 50618
rect 23142 50566 23194 50618
rect 23206 50566 23258 50618
rect 1124 50396 1176 50448
rect 9404 50439 9456 50448
rect 9404 50405 9413 50439
rect 9413 50405 9447 50439
rect 9447 50405 9456 50439
rect 9404 50396 9456 50405
rect 2044 50328 2096 50380
rect 4344 50371 4396 50380
rect 4344 50337 4353 50371
rect 4353 50337 4387 50371
rect 4387 50337 4396 50371
rect 4344 50328 4396 50337
rect 3976 50260 4028 50312
rect 8668 50260 8720 50312
rect 25320 50303 25372 50312
rect 25320 50269 25329 50303
rect 25329 50269 25363 50303
rect 25363 50269 25372 50303
rect 25320 50260 25372 50269
rect 7748 50192 7800 50244
rect 23388 50124 23440 50176
rect 7950 50022 8002 50074
rect 8014 50022 8066 50074
rect 8078 50022 8130 50074
rect 8142 50022 8194 50074
rect 8206 50022 8258 50074
rect 17950 50022 18002 50074
rect 18014 50022 18066 50074
rect 18078 50022 18130 50074
rect 18142 50022 18194 50074
rect 18206 50022 18258 50074
rect 7012 49920 7064 49972
rect 7380 49920 7432 49972
rect 21364 49920 21416 49972
rect 1676 49852 1728 49904
rect 7656 49852 7708 49904
rect 9588 49895 9640 49904
rect 9588 49861 9597 49895
rect 9597 49861 9631 49895
rect 9631 49861 9640 49895
rect 9588 49852 9640 49861
rect 3700 49784 3752 49836
rect 6552 49827 6604 49836
rect 6552 49793 6561 49827
rect 6561 49793 6595 49827
rect 6595 49793 6604 49827
rect 6552 49784 6604 49793
rect 7380 49784 7432 49836
rect 24768 49827 24820 49836
rect 24768 49793 24777 49827
rect 24777 49793 24811 49827
rect 24811 49793 24820 49827
rect 24768 49784 24820 49793
rect 2950 49478 3002 49530
rect 3014 49478 3066 49530
rect 3078 49478 3130 49530
rect 3142 49478 3194 49530
rect 3206 49478 3258 49530
rect 12950 49478 13002 49530
rect 13014 49478 13066 49530
rect 13078 49478 13130 49530
rect 13142 49478 13194 49530
rect 13206 49478 13258 49530
rect 22950 49478 23002 49530
rect 23014 49478 23066 49530
rect 23078 49478 23130 49530
rect 23142 49478 23194 49530
rect 23206 49478 23258 49530
rect 1308 49240 1360 49292
rect 9404 49240 9456 49292
rect 3332 49172 3384 49224
rect 10048 49172 10100 49224
rect 25320 49215 25372 49224
rect 25320 49181 25329 49215
rect 25329 49181 25363 49215
rect 25363 49181 25372 49215
rect 25320 49172 25372 49181
rect 4068 49104 4120 49156
rect 9036 49104 9088 49156
rect 19892 49036 19944 49088
rect 7950 48934 8002 48986
rect 8014 48934 8066 48986
rect 8078 48934 8130 48986
rect 8142 48934 8194 48986
rect 8206 48934 8258 48986
rect 17950 48934 18002 48986
rect 18014 48934 18066 48986
rect 18078 48934 18130 48986
rect 18142 48934 18194 48986
rect 18206 48934 18258 48986
rect 11796 48832 11848 48884
rect 11704 48739 11756 48748
rect 11704 48705 11713 48739
rect 11713 48705 11747 48739
rect 11747 48705 11756 48739
rect 11704 48696 11756 48705
rect 24768 48739 24820 48748
rect 24768 48705 24777 48739
rect 24777 48705 24811 48739
rect 24811 48705 24820 48739
rect 24768 48696 24820 48705
rect 21640 48492 21692 48544
rect 2950 48390 3002 48442
rect 3014 48390 3066 48442
rect 3078 48390 3130 48442
rect 3142 48390 3194 48442
rect 3206 48390 3258 48442
rect 12950 48390 13002 48442
rect 13014 48390 13066 48442
rect 13078 48390 13130 48442
rect 13142 48390 13194 48442
rect 13206 48390 13258 48442
rect 22950 48390 23002 48442
rect 23014 48390 23066 48442
rect 23078 48390 23130 48442
rect 23142 48390 23194 48442
rect 23206 48390 23258 48442
rect 20720 48220 20772 48272
rect 25504 48084 25556 48136
rect 1308 48016 1360 48068
rect 4068 47948 4120 48000
rect 24860 47948 24912 48000
rect 7950 47846 8002 47898
rect 8014 47846 8066 47898
rect 8078 47846 8130 47898
rect 8142 47846 8194 47898
rect 8206 47846 8258 47898
rect 17950 47846 18002 47898
rect 18014 47846 18066 47898
rect 18078 47846 18130 47898
rect 18142 47846 18194 47898
rect 18206 47846 18258 47898
rect 23848 47744 23900 47796
rect 24400 47744 24452 47796
rect 24032 47676 24084 47728
rect 24860 47608 24912 47660
rect 25872 47472 25924 47524
rect 16120 47404 16172 47456
rect 25504 47447 25556 47456
rect 25504 47413 25513 47447
rect 25513 47413 25547 47447
rect 25547 47413 25556 47447
rect 25504 47404 25556 47413
rect 2950 47302 3002 47354
rect 3014 47302 3066 47354
rect 3078 47302 3130 47354
rect 3142 47302 3194 47354
rect 3206 47302 3258 47354
rect 12950 47302 13002 47354
rect 13014 47302 13066 47354
rect 13078 47302 13130 47354
rect 13142 47302 13194 47354
rect 13206 47302 13258 47354
rect 22950 47302 23002 47354
rect 23014 47302 23066 47354
rect 23078 47302 23130 47354
rect 23142 47302 23194 47354
rect 23206 47302 23258 47354
rect 6828 47200 6880 47252
rect 11612 47200 11664 47252
rect 13820 47200 13872 47252
rect 14832 47200 14884 47252
rect 14556 47064 14608 47116
rect 16488 47064 16540 47116
rect 10968 46996 11020 47048
rect 11520 47039 11572 47048
rect 11520 47005 11529 47039
rect 11529 47005 11563 47039
rect 11563 47005 11572 47039
rect 11520 46996 11572 47005
rect 16856 47039 16908 47048
rect 16856 47005 16865 47039
rect 16865 47005 16899 47039
rect 16899 47005 16908 47039
rect 16856 46996 16908 47005
rect 17776 47107 17828 47116
rect 17776 47073 17785 47107
rect 17785 47073 17819 47107
rect 17819 47073 17828 47107
rect 17776 47064 17828 47073
rect 23296 47200 23348 47252
rect 24952 47132 25004 47184
rect 18972 46996 19024 47048
rect 16120 46928 16172 46980
rect 16580 46971 16632 46980
rect 16580 46937 16589 46971
rect 16589 46937 16623 46971
rect 16623 46937 16632 46971
rect 16580 46928 16632 46937
rect 24952 46928 25004 46980
rect 17316 46903 17368 46912
rect 17316 46869 17325 46903
rect 17325 46869 17359 46903
rect 17359 46869 17368 46903
rect 17316 46860 17368 46869
rect 7950 46758 8002 46810
rect 8014 46758 8066 46810
rect 8078 46758 8130 46810
rect 8142 46758 8194 46810
rect 8206 46758 8258 46810
rect 17950 46758 18002 46810
rect 18014 46758 18066 46810
rect 18078 46758 18130 46810
rect 18142 46758 18194 46810
rect 18206 46758 18258 46810
rect 7104 46699 7156 46708
rect 7104 46665 7113 46699
rect 7113 46665 7147 46699
rect 7147 46665 7156 46699
rect 7104 46656 7156 46665
rect 13820 46656 13872 46708
rect 16120 46656 16172 46708
rect 17408 46656 17460 46708
rect 18696 46656 18748 46708
rect 19616 46656 19668 46708
rect 20536 46699 20588 46708
rect 20536 46665 20545 46699
rect 20545 46665 20579 46699
rect 20579 46665 20588 46699
rect 20536 46656 20588 46665
rect 16028 46588 16080 46640
rect 18604 46588 18656 46640
rect 7288 46563 7340 46572
rect 7288 46529 7297 46563
rect 7297 46529 7331 46563
rect 7331 46529 7340 46563
rect 7288 46520 7340 46529
rect 16580 46520 16632 46572
rect 15476 46495 15528 46504
rect 15476 46461 15485 46495
rect 15485 46461 15519 46495
rect 15519 46461 15528 46495
rect 15476 46452 15528 46461
rect 16856 46452 16908 46504
rect 17776 46520 17828 46572
rect 18512 46520 18564 46572
rect 23848 46520 23900 46572
rect 24676 46520 24728 46572
rect 18604 46495 18656 46504
rect 18604 46461 18613 46495
rect 18613 46461 18647 46495
rect 18647 46461 18656 46495
rect 18604 46452 18656 46461
rect 26056 46452 26108 46504
rect 24860 46384 24912 46436
rect 17132 46316 17184 46368
rect 18328 46316 18380 46368
rect 23296 46359 23348 46368
rect 23296 46325 23305 46359
rect 23305 46325 23339 46359
rect 23339 46325 23348 46359
rect 23296 46316 23348 46325
rect 23848 46359 23900 46368
rect 23848 46325 23857 46359
rect 23857 46325 23891 46359
rect 23891 46325 23900 46359
rect 23848 46316 23900 46325
rect 2950 46214 3002 46266
rect 3014 46214 3066 46266
rect 3078 46214 3130 46266
rect 3142 46214 3194 46266
rect 3206 46214 3258 46266
rect 12950 46214 13002 46266
rect 13014 46214 13066 46266
rect 13078 46214 13130 46266
rect 13142 46214 13194 46266
rect 13206 46214 13258 46266
rect 22950 46214 23002 46266
rect 23014 46214 23066 46266
rect 23078 46214 23130 46266
rect 23142 46214 23194 46266
rect 23206 46214 23258 46266
rect 16580 46112 16632 46164
rect 18420 46112 18472 46164
rect 18696 46112 18748 46164
rect 25044 46112 25096 46164
rect 15844 45976 15896 46028
rect 16120 45976 16172 46028
rect 1216 45908 1268 45960
rect 9864 45908 9916 45960
rect 16856 45976 16908 46028
rect 19800 45976 19852 46028
rect 22284 46044 22336 46096
rect 24584 46044 24636 46096
rect 21548 45976 21600 46028
rect 20904 45908 20956 45960
rect 24860 45976 24912 46028
rect 24216 45908 24268 45960
rect 17592 45840 17644 45892
rect 18604 45840 18656 45892
rect 19616 45840 19668 45892
rect 20260 45840 20312 45892
rect 20536 45840 20588 45892
rect 24676 45840 24728 45892
rect 20076 45772 20128 45824
rect 24124 45772 24176 45824
rect 7950 45670 8002 45722
rect 8014 45670 8066 45722
rect 8078 45670 8130 45722
rect 8142 45670 8194 45722
rect 8206 45670 8258 45722
rect 17950 45670 18002 45722
rect 18014 45670 18066 45722
rect 18078 45670 18130 45722
rect 18142 45670 18194 45722
rect 18206 45670 18258 45722
rect 1216 45568 1268 45620
rect 6644 45500 6696 45552
rect 11980 45500 12032 45552
rect 14832 45543 14884 45552
rect 14832 45509 14841 45543
rect 14841 45509 14875 45543
rect 14875 45509 14884 45543
rect 14832 45500 14884 45509
rect 22008 45500 22060 45552
rect 7104 45228 7156 45280
rect 8392 45475 8444 45484
rect 8392 45441 8401 45475
rect 8401 45441 8435 45475
rect 8435 45441 8444 45475
rect 8392 45432 8444 45441
rect 9772 45475 9824 45484
rect 9772 45441 9781 45475
rect 9781 45441 9815 45475
rect 9815 45441 9824 45475
rect 9772 45432 9824 45441
rect 12256 45432 12308 45484
rect 13728 45432 13780 45484
rect 15476 45432 15528 45484
rect 17224 45432 17276 45484
rect 19524 45432 19576 45484
rect 22652 45475 22704 45484
rect 22652 45441 22661 45475
rect 22661 45441 22695 45475
rect 22695 45441 22704 45475
rect 22652 45432 22704 45441
rect 24124 45475 24176 45484
rect 24124 45441 24133 45475
rect 24133 45441 24167 45475
rect 24167 45441 24176 45475
rect 24124 45432 24176 45441
rect 13544 45364 13596 45416
rect 8576 45339 8628 45348
rect 8576 45305 8585 45339
rect 8585 45305 8619 45339
rect 8619 45305 8628 45339
rect 8576 45296 8628 45305
rect 9956 45339 10008 45348
rect 9956 45305 9965 45339
rect 9965 45305 9999 45339
rect 9999 45305 10008 45339
rect 9956 45296 10008 45305
rect 19432 45364 19484 45416
rect 20812 45364 20864 45416
rect 24768 45407 24820 45416
rect 24768 45373 24777 45407
rect 24777 45373 24811 45407
rect 24811 45373 24820 45407
rect 24768 45364 24820 45373
rect 8300 45228 8352 45280
rect 12256 45271 12308 45280
rect 12256 45237 12265 45271
rect 12265 45237 12299 45271
rect 12299 45237 12308 45271
rect 12256 45228 12308 45237
rect 12716 45228 12768 45280
rect 15292 45228 15344 45280
rect 15844 45228 15896 45280
rect 16856 45271 16908 45280
rect 16856 45237 16865 45271
rect 16865 45237 16899 45271
rect 16899 45237 16908 45271
rect 16856 45228 16908 45237
rect 18512 45228 18564 45280
rect 18604 45228 18656 45280
rect 19064 45228 19116 45280
rect 19524 45228 19576 45280
rect 19708 45271 19760 45280
rect 19708 45237 19717 45271
rect 19717 45237 19751 45271
rect 19751 45237 19760 45271
rect 19708 45228 19760 45237
rect 2950 45126 3002 45178
rect 3014 45126 3066 45178
rect 3078 45126 3130 45178
rect 3142 45126 3194 45178
rect 3206 45126 3258 45178
rect 12950 45126 13002 45178
rect 13014 45126 13066 45178
rect 13078 45126 13130 45178
rect 13142 45126 13194 45178
rect 13206 45126 13258 45178
rect 22950 45126 23002 45178
rect 23014 45126 23066 45178
rect 23078 45126 23130 45178
rect 23142 45126 23194 45178
rect 23206 45126 23258 45178
rect 10140 45067 10192 45076
rect 10140 45033 10149 45067
rect 10149 45033 10183 45067
rect 10183 45033 10192 45067
rect 10140 45024 10192 45033
rect 15844 45024 15896 45076
rect 5816 44956 5868 45008
rect 7472 44820 7524 44872
rect 10692 44863 10744 44872
rect 10692 44829 10701 44863
rect 10701 44829 10735 44863
rect 10735 44829 10744 44863
rect 10692 44820 10744 44829
rect 14280 44863 14332 44872
rect 14280 44829 14289 44863
rect 14289 44829 14323 44863
rect 14323 44829 14332 44863
rect 14280 44820 14332 44829
rect 8760 44684 8812 44736
rect 9680 44727 9732 44736
rect 9680 44693 9689 44727
rect 9689 44693 9723 44727
rect 9723 44693 9732 44727
rect 11244 44752 11296 44804
rect 9680 44684 9732 44693
rect 12348 44684 12400 44736
rect 14096 44752 14148 44804
rect 14556 44795 14608 44804
rect 14556 44761 14565 44795
rect 14565 44761 14599 44795
rect 14599 44761 14608 44795
rect 14556 44752 14608 44761
rect 15292 44752 15344 44804
rect 13728 44684 13780 44736
rect 16028 44727 16080 44736
rect 16028 44693 16037 44727
rect 16037 44693 16071 44727
rect 16071 44693 16080 44727
rect 16028 44684 16080 44693
rect 22744 44956 22796 45008
rect 21916 44931 21968 44940
rect 21916 44897 21925 44931
rect 21925 44897 21959 44931
rect 21959 44897 21968 44931
rect 21916 44888 21968 44897
rect 24124 44888 24176 44940
rect 21180 44863 21232 44872
rect 21180 44829 21189 44863
rect 21189 44829 21223 44863
rect 21223 44829 21232 44863
rect 21180 44820 21232 44829
rect 22652 44820 22704 44872
rect 24492 44820 24544 44872
rect 25320 44863 25372 44872
rect 25320 44829 25329 44863
rect 25329 44829 25363 44863
rect 25363 44829 25372 44863
rect 25320 44820 25372 44829
rect 17224 44684 17276 44736
rect 17500 44684 17552 44736
rect 19340 44684 19392 44736
rect 20904 44795 20956 44804
rect 20904 44761 20913 44795
rect 20913 44761 20947 44795
rect 20947 44761 20956 44795
rect 20904 44752 20956 44761
rect 21088 44684 21140 44736
rect 21456 44684 21508 44736
rect 22468 44684 22520 44736
rect 22836 44727 22888 44736
rect 22836 44693 22845 44727
rect 22845 44693 22879 44727
rect 22879 44693 22888 44727
rect 22836 44684 22888 44693
rect 23572 44684 23624 44736
rect 7950 44582 8002 44634
rect 8014 44582 8066 44634
rect 8078 44582 8130 44634
rect 8142 44582 8194 44634
rect 8206 44582 8258 44634
rect 17950 44582 18002 44634
rect 18014 44582 18066 44634
rect 18078 44582 18130 44634
rect 18142 44582 18194 44634
rect 18206 44582 18258 44634
rect 7196 44523 7248 44532
rect 7196 44489 7205 44523
rect 7205 44489 7239 44523
rect 7239 44489 7248 44523
rect 7196 44480 7248 44489
rect 7748 44480 7800 44532
rect 9036 44523 9088 44532
rect 9036 44489 9045 44523
rect 9045 44489 9079 44523
rect 9079 44489 9088 44523
rect 9036 44480 9088 44489
rect 9220 44480 9272 44532
rect 7748 44344 7800 44396
rect 8484 44455 8536 44464
rect 8484 44421 8493 44455
rect 8493 44421 8527 44455
rect 8527 44421 8536 44455
rect 8484 44412 8536 44421
rect 10048 44480 10100 44532
rect 11704 44523 11756 44532
rect 11704 44489 11713 44523
rect 11713 44489 11747 44523
rect 11747 44489 11756 44523
rect 11704 44480 11756 44489
rect 13636 44480 13688 44532
rect 11060 44412 11112 44464
rect 6736 44276 6788 44328
rect 8300 44276 8352 44328
rect 8760 44344 8812 44396
rect 9404 44387 9456 44396
rect 9404 44353 9413 44387
rect 9413 44353 9447 44387
rect 9447 44353 9456 44387
rect 9404 44344 9456 44353
rect 12624 44344 12676 44396
rect 11336 44276 11388 44328
rect 12164 44319 12216 44328
rect 12164 44285 12173 44319
rect 12173 44285 12207 44319
rect 12207 44285 12216 44319
rect 12164 44276 12216 44285
rect 12348 44319 12400 44328
rect 12348 44285 12357 44319
rect 12357 44285 12391 44319
rect 12391 44285 12400 44319
rect 12348 44276 12400 44285
rect 11244 44140 11296 44192
rect 11888 44140 11940 44192
rect 15936 44276 15988 44328
rect 17040 44480 17092 44532
rect 18512 44480 18564 44532
rect 24216 44480 24268 44532
rect 19616 44412 19668 44464
rect 21088 44412 21140 44464
rect 18052 44344 18104 44396
rect 25964 44344 26016 44396
rect 19432 44319 19484 44328
rect 19432 44285 19441 44319
rect 19441 44285 19475 44319
rect 19475 44285 19484 44319
rect 19432 44276 19484 44285
rect 21456 44319 21508 44328
rect 21456 44285 21465 44319
rect 21465 44285 21499 44319
rect 21499 44285 21508 44319
rect 21456 44276 21508 44285
rect 22100 44276 22152 44328
rect 23756 44319 23808 44328
rect 23756 44285 23765 44319
rect 23765 44285 23799 44319
rect 23799 44285 23808 44319
rect 23756 44276 23808 44285
rect 25504 44276 25556 44328
rect 14556 44208 14608 44260
rect 15384 44208 15436 44260
rect 20812 44208 20864 44260
rect 14188 44140 14240 44192
rect 19064 44140 19116 44192
rect 21088 44140 21140 44192
rect 2950 44038 3002 44090
rect 3014 44038 3066 44090
rect 3078 44038 3130 44090
rect 3142 44038 3194 44090
rect 3206 44038 3258 44090
rect 12950 44038 13002 44090
rect 13014 44038 13066 44090
rect 13078 44038 13130 44090
rect 13142 44038 13194 44090
rect 13206 44038 13258 44090
rect 22950 44038 23002 44090
rect 23014 44038 23066 44090
rect 23078 44038 23130 44090
rect 23142 44038 23194 44090
rect 23206 44038 23258 44090
rect 9128 43936 9180 43988
rect 20904 43936 20956 43988
rect 22100 43936 22152 43988
rect 24216 43936 24268 43988
rect 24768 43936 24820 43988
rect 6184 43868 6236 43920
rect 7840 43868 7892 43920
rect 9496 43868 9548 43920
rect 1308 43732 1360 43784
rect 14924 43800 14976 43852
rect 15476 43800 15528 43852
rect 18604 43800 18656 43852
rect 23756 43843 23808 43852
rect 23756 43809 23765 43843
rect 23765 43809 23799 43843
rect 23799 43809 23808 43843
rect 23756 43800 23808 43809
rect 25044 43800 25096 43852
rect 10508 43732 10560 43784
rect 10692 43732 10744 43784
rect 11796 43775 11848 43784
rect 11796 43741 11805 43775
rect 11805 43741 11839 43775
rect 11839 43741 11848 43775
rect 11796 43732 11848 43741
rect 19432 43775 19484 43784
rect 19432 43741 19441 43775
rect 19441 43741 19475 43775
rect 19475 43741 19484 43775
rect 19432 43732 19484 43741
rect 20812 43732 20864 43784
rect 21088 43732 21140 43784
rect 22008 43732 22060 43784
rect 24768 43775 24820 43784
rect 24768 43741 24777 43775
rect 24777 43741 24811 43775
rect 24811 43741 24820 43775
rect 24768 43732 24820 43741
rect 1768 43639 1820 43648
rect 1768 43605 1777 43639
rect 1777 43605 1811 43639
rect 1811 43605 1820 43639
rect 1768 43596 1820 43605
rect 11704 43664 11756 43716
rect 12348 43664 12400 43716
rect 15844 43664 15896 43716
rect 17500 43664 17552 43716
rect 18052 43664 18104 43716
rect 19984 43664 20036 43716
rect 23756 43664 23808 43716
rect 9128 43596 9180 43648
rect 10784 43596 10836 43648
rect 13636 43596 13688 43648
rect 13728 43596 13780 43648
rect 17592 43639 17644 43648
rect 17592 43605 17601 43639
rect 17601 43605 17635 43639
rect 17635 43605 17644 43639
rect 17592 43596 17644 43605
rect 25504 43639 25556 43648
rect 25504 43605 25513 43639
rect 25513 43605 25547 43639
rect 25547 43605 25556 43639
rect 25504 43596 25556 43605
rect 7950 43494 8002 43546
rect 8014 43494 8066 43546
rect 8078 43494 8130 43546
rect 8142 43494 8194 43546
rect 8206 43494 8258 43546
rect 17950 43494 18002 43546
rect 18014 43494 18066 43546
rect 18078 43494 18130 43546
rect 18142 43494 18194 43546
rect 18206 43494 18258 43546
rect 1768 43392 1820 43444
rect 6552 43392 6604 43444
rect 8668 43435 8720 43444
rect 8668 43401 8677 43435
rect 8677 43401 8711 43435
rect 8711 43401 8720 43435
rect 8668 43392 8720 43401
rect 12164 43392 12216 43444
rect 17132 43392 17184 43444
rect 10048 43324 10100 43376
rect 10784 43367 10836 43376
rect 10784 43333 10793 43367
rect 10793 43333 10827 43367
rect 10827 43333 10836 43367
rect 10784 43324 10836 43333
rect 19892 43392 19944 43444
rect 22008 43392 22060 43444
rect 22284 43367 22336 43376
rect 22284 43333 22293 43367
rect 22293 43333 22327 43367
rect 22327 43333 22336 43367
rect 22284 43324 22336 43333
rect 22560 43324 22612 43376
rect 23756 43435 23808 43444
rect 23756 43401 23765 43435
rect 23765 43401 23799 43435
rect 23799 43401 23808 43435
rect 23756 43392 23808 43401
rect 24400 43392 24452 43444
rect 23664 43324 23716 43376
rect 24216 43367 24268 43376
rect 24216 43333 24225 43367
rect 24225 43333 24259 43367
rect 24259 43333 24268 43367
rect 24216 43324 24268 43333
rect 4988 43256 5040 43308
rect 5172 43256 5224 43308
rect 10692 43256 10744 43308
rect 15660 43256 15712 43308
rect 25412 43256 25464 43308
rect 10784 43188 10836 43240
rect 11060 43188 11112 43240
rect 11888 43120 11940 43172
rect 14096 43120 14148 43172
rect 22008 43231 22060 43240
rect 22008 43197 22017 43231
rect 22017 43197 22051 43231
rect 22051 43197 22060 43231
rect 22008 43188 22060 43197
rect 8484 43052 8536 43104
rect 16672 43052 16724 43104
rect 25228 43052 25280 43104
rect 2950 42950 3002 43002
rect 3014 42950 3066 43002
rect 3078 42950 3130 43002
rect 3142 42950 3194 43002
rect 3206 42950 3258 43002
rect 12950 42950 13002 43002
rect 13014 42950 13066 43002
rect 13078 42950 13130 43002
rect 13142 42950 13194 43002
rect 13206 42950 13258 43002
rect 22950 42950 23002 43002
rect 23014 42950 23066 43002
rect 23078 42950 23130 43002
rect 23142 42950 23194 43002
rect 23206 42950 23258 43002
rect 12716 42848 12768 42900
rect 17408 42848 17460 42900
rect 15844 42780 15896 42832
rect 16856 42780 16908 42832
rect 4160 42755 4212 42764
rect 4160 42721 4169 42755
rect 4169 42721 4203 42755
rect 4203 42721 4212 42755
rect 4160 42712 4212 42721
rect 6368 42712 6420 42764
rect 8300 42755 8352 42764
rect 8300 42721 8309 42755
rect 8309 42721 8343 42755
rect 8343 42721 8352 42755
rect 8300 42712 8352 42721
rect 9220 42712 9272 42764
rect 12532 42755 12584 42764
rect 12532 42721 12541 42755
rect 12541 42721 12575 42755
rect 12575 42721 12584 42755
rect 12532 42712 12584 42721
rect 14280 42755 14332 42764
rect 14280 42721 14289 42755
rect 14289 42721 14323 42755
rect 14323 42721 14332 42755
rect 14280 42712 14332 42721
rect 25136 42780 25188 42832
rect 25412 42780 25464 42832
rect 7564 42644 7616 42696
rect 6460 42619 6512 42628
rect 6460 42585 6469 42619
rect 6469 42585 6503 42619
rect 6503 42585 6512 42619
rect 6460 42576 6512 42585
rect 8484 42687 8536 42696
rect 8484 42653 8493 42687
rect 8493 42653 8527 42687
rect 8527 42653 8536 42687
rect 8484 42644 8536 42653
rect 9036 42644 9088 42696
rect 9680 42644 9732 42696
rect 11244 42644 11296 42696
rect 11796 42644 11848 42696
rect 18328 42644 18380 42696
rect 21180 42687 21232 42696
rect 21180 42653 21189 42687
rect 21189 42653 21223 42687
rect 21223 42653 21232 42687
rect 21180 42644 21232 42653
rect 22008 42644 22060 42696
rect 22284 42687 22336 42696
rect 22284 42653 22293 42687
rect 22293 42653 22327 42687
rect 22327 42653 22336 42687
rect 22284 42644 22336 42653
rect 23664 42644 23716 42696
rect 9496 42576 9548 42628
rect 10968 42576 11020 42628
rect 6828 42508 6880 42560
rect 7380 42508 7432 42560
rect 7656 42508 7708 42560
rect 9864 42508 9916 42560
rect 11060 42508 11112 42560
rect 13728 42576 13780 42628
rect 15016 42576 15068 42628
rect 20904 42619 20956 42628
rect 20904 42585 20913 42619
rect 20913 42585 20947 42619
rect 20947 42585 20956 42619
rect 20904 42576 20956 42585
rect 12072 42508 12124 42560
rect 12440 42551 12492 42560
rect 12440 42517 12449 42551
rect 12449 42517 12483 42551
rect 12483 42517 12492 42551
rect 12440 42508 12492 42517
rect 15568 42508 15620 42560
rect 16304 42551 16356 42560
rect 16304 42517 16313 42551
rect 16313 42517 16347 42551
rect 16347 42517 16356 42551
rect 16304 42508 16356 42517
rect 17684 42508 17736 42560
rect 17868 42551 17920 42560
rect 17868 42517 17877 42551
rect 17877 42517 17911 42551
rect 17911 42517 17920 42551
rect 17868 42508 17920 42517
rect 19340 42508 19392 42560
rect 20536 42508 20588 42560
rect 20812 42508 20864 42560
rect 22560 42619 22612 42628
rect 22560 42585 22569 42619
rect 22569 42585 22603 42619
rect 22603 42585 22612 42619
rect 22560 42576 22612 42585
rect 21272 42508 21324 42560
rect 24492 42508 24544 42560
rect 24584 42551 24636 42560
rect 24584 42517 24593 42551
rect 24593 42517 24627 42551
rect 24627 42517 24636 42551
rect 24584 42508 24636 42517
rect 24860 42508 24912 42560
rect 25504 42551 25556 42560
rect 25504 42517 25513 42551
rect 25513 42517 25547 42551
rect 25547 42517 25556 42551
rect 25504 42508 25556 42517
rect 7950 42406 8002 42458
rect 8014 42406 8066 42458
rect 8078 42406 8130 42458
rect 8142 42406 8194 42458
rect 8206 42406 8258 42458
rect 17950 42406 18002 42458
rect 18014 42406 18066 42458
rect 18078 42406 18130 42458
rect 18142 42406 18194 42458
rect 18206 42406 18258 42458
rect 6920 42304 6972 42356
rect 7380 42304 7432 42356
rect 3700 42279 3752 42288
rect 3700 42245 3709 42279
rect 3709 42245 3743 42279
rect 3743 42245 3752 42279
rect 3700 42236 3752 42245
rect 9404 42304 9456 42356
rect 10048 42304 10100 42356
rect 10968 42304 11020 42356
rect 11520 42304 11572 42356
rect 12440 42304 12492 42356
rect 16764 42304 16816 42356
rect 19432 42304 19484 42356
rect 22836 42304 22888 42356
rect 4344 42168 4396 42220
rect 8576 42236 8628 42288
rect 12348 42236 12400 42288
rect 13728 42236 13780 42288
rect 15016 42236 15068 42288
rect 16304 42236 16356 42288
rect 13820 42168 13872 42220
rect 15476 42168 15528 42220
rect 18420 42236 18472 42288
rect 21180 42236 21232 42288
rect 22744 42236 22796 42288
rect 23848 42304 23900 42356
rect 24492 42236 24544 42288
rect 24676 42236 24728 42288
rect 19248 42168 19300 42220
rect 8484 42100 8536 42152
rect 11152 42100 11204 42152
rect 15568 42100 15620 42152
rect 19156 42100 19208 42152
rect 11520 42032 11572 42084
rect 21088 42168 21140 42220
rect 22376 42211 22428 42220
rect 22376 42177 22385 42211
rect 22385 42177 22419 42211
rect 22419 42177 22428 42211
rect 22376 42168 22428 42177
rect 23664 42168 23716 42220
rect 22192 42143 22244 42152
rect 22192 42109 22201 42143
rect 22201 42109 22235 42143
rect 22235 42109 22244 42143
rect 22192 42100 22244 42109
rect 22560 42100 22612 42152
rect 25044 42143 25096 42152
rect 25044 42109 25053 42143
rect 25053 42109 25087 42143
rect 25087 42109 25096 42143
rect 25044 42100 25096 42109
rect 20536 42032 20588 42084
rect 4344 42007 4396 42016
rect 4344 41973 4353 42007
rect 4353 41973 4387 42007
rect 4387 41973 4396 42007
rect 4344 41964 4396 41973
rect 8668 41964 8720 42016
rect 11428 41964 11480 42016
rect 14556 41964 14608 42016
rect 19616 42007 19668 42016
rect 19616 41973 19625 42007
rect 19625 41973 19659 42007
rect 19659 41973 19668 42007
rect 19616 41964 19668 41973
rect 21088 41964 21140 42016
rect 25136 41964 25188 42016
rect 2950 41862 3002 41914
rect 3014 41862 3066 41914
rect 3078 41862 3130 41914
rect 3142 41862 3194 41914
rect 3206 41862 3258 41914
rect 12950 41862 13002 41914
rect 13014 41862 13066 41914
rect 13078 41862 13130 41914
rect 13142 41862 13194 41914
rect 13206 41862 13258 41914
rect 22950 41862 23002 41914
rect 23014 41862 23066 41914
rect 23078 41862 23130 41914
rect 23142 41862 23194 41914
rect 23206 41862 23258 41914
rect 4436 41803 4488 41812
rect 4436 41769 4445 41803
rect 4445 41769 4479 41803
rect 4479 41769 4488 41803
rect 4436 41760 4488 41769
rect 5356 41803 5408 41812
rect 5356 41769 5365 41803
rect 5365 41769 5399 41803
rect 5399 41769 5408 41803
rect 5356 41760 5408 41769
rect 7288 41760 7340 41812
rect 16212 41760 16264 41812
rect 8484 41667 8536 41676
rect 8484 41633 8493 41667
rect 8493 41633 8527 41667
rect 8527 41633 8536 41667
rect 8484 41624 8536 41633
rect 11244 41667 11296 41676
rect 11244 41633 11253 41667
rect 11253 41633 11287 41667
rect 11287 41633 11296 41667
rect 11244 41624 11296 41633
rect 11520 41667 11572 41676
rect 11520 41633 11529 41667
rect 11529 41633 11563 41667
rect 11563 41633 11572 41667
rect 11520 41624 11572 41633
rect 15476 41624 15528 41676
rect 17500 41760 17552 41812
rect 19248 41760 19300 41812
rect 21272 41760 21324 41812
rect 23572 41760 23624 41812
rect 19064 41692 19116 41744
rect 19340 41692 19392 41744
rect 6644 41556 6696 41608
rect 8300 41556 8352 41608
rect 13268 41556 13320 41608
rect 13728 41556 13780 41608
rect 18420 41624 18472 41676
rect 19708 41624 19760 41676
rect 23204 41692 23256 41744
rect 24400 41692 24452 41744
rect 20812 41667 20864 41676
rect 20812 41633 20821 41667
rect 20821 41633 20855 41667
rect 20855 41633 20864 41667
rect 20812 41624 20864 41633
rect 20996 41667 21048 41676
rect 20996 41633 21005 41667
rect 21005 41633 21039 41667
rect 21039 41633 21048 41667
rect 20996 41624 21048 41633
rect 22100 41667 22152 41676
rect 22100 41633 22109 41667
rect 22109 41633 22143 41667
rect 22143 41633 22152 41667
rect 22100 41624 22152 41633
rect 23388 41624 23440 41676
rect 23664 41624 23716 41676
rect 21088 41556 21140 41608
rect 21916 41556 21968 41608
rect 23756 41599 23808 41608
rect 23756 41565 23765 41599
rect 23765 41565 23799 41599
rect 23799 41565 23808 41599
rect 23756 41556 23808 41565
rect 24768 41556 24820 41608
rect 1676 41531 1728 41540
rect 1676 41497 1685 41531
rect 1685 41497 1719 41531
rect 1719 41497 1728 41531
rect 1676 41488 1728 41497
rect 3608 41420 3660 41472
rect 6276 41420 6328 41472
rect 9588 41420 9640 41472
rect 12532 41420 12584 41472
rect 13268 41463 13320 41472
rect 13268 41429 13277 41463
rect 13277 41429 13311 41463
rect 13311 41429 13320 41463
rect 13268 41420 13320 41429
rect 19432 41463 19484 41472
rect 19432 41429 19441 41463
rect 19441 41429 19475 41463
rect 19475 41429 19484 41463
rect 19432 41420 19484 41429
rect 19524 41420 19576 41472
rect 21180 41420 21232 41472
rect 22652 41420 22704 41472
rect 23480 41420 23532 41472
rect 24952 41420 25004 41472
rect 7950 41318 8002 41370
rect 8014 41318 8066 41370
rect 8078 41318 8130 41370
rect 8142 41318 8194 41370
rect 8206 41318 8258 41370
rect 17950 41318 18002 41370
rect 18014 41318 18066 41370
rect 18078 41318 18130 41370
rect 18142 41318 18194 41370
rect 18206 41318 18258 41370
rect 3976 41259 4028 41268
rect 3976 41225 3985 41259
rect 3985 41225 4019 41259
rect 4019 41225 4028 41259
rect 3976 41216 4028 41225
rect 4528 41216 4580 41268
rect 7564 41216 7616 41268
rect 7104 41148 7156 41200
rect 8484 41216 8536 41268
rect 9680 41216 9732 41268
rect 12256 41216 12308 41268
rect 12624 41216 12676 41268
rect 10968 41148 11020 41200
rect 13268 41216 13320 41268
rect 14372 41148 14424 41200
rect 17316 41259 17368 41268
rect 17316 41225 17325 41259
rect 17325 41225 17359 41259
rect 17359 41225 17368 41259
rect 17316 41216 17368 41225
rect 14556 41148 14608 41200
rect 16212 41148 16264 41200
rect 19340 41216 19392 41268
rect 22008 41216 22060 41268
rect 22560 41216 22612 41268
rect 22744 41259 22796 41268
rect 22744 41225 22753 41259
rect 22753 41225 22787 41259
rect 22787 41225 22796 41259
rect 22744 41216 22796 41225
rect 23848 41216 23900 41268
rect 24216 41148 24268 41200
rect 4252 41080 4304 41132
rect 6368 41012 6420 41064
rect 7840 41012 7892 41064
rect 9404 41055 9456 41064
rect 9404 41021 9413 41055
rect 9413 41021 9447 41055
rect 9447 41021 9456 41055
rect 9404 41012 9456 41021
rect 10876 41012 10928 41064
rect 15476 41080 15528 41132
rect 17224 41123 17276 41132
rect 17224 41089 17233 41123
rect 17233 41089 17267 41123
rect 17267 41089 17276 41123
rect 17224 41080 17276 41089
rect 18420 41123 18472 41132
rect 18420 41089 18429 41123
rect 18429 41089 18463 41123
rect 18463 41089 18472 41123
rect 18420 41080 18472 41089
rect 11888 41055 11940 41064
rect 11888 41021 11897 41055
rect 11897 41021 11931 41055
rect 11931 41021 11940 41055
rect 11888 41012 11940 41021
rect 14832 41012 14884 41064
rect 17408 41055 17460 41064
rect 17408 41021 17417 41055
rect 17417 41021 17451 41055
rect 17451 41021 17460 41055
rect 17408 41012 17460 41021
rect 23388 41080 23440 41132
rect 20536 41055 20588 41064
rect 20536 41021 20545 41055
rect 20545 41021 20579 41055
rect 20579 41021 20588 41055
rect 20536 41012 20588 41021
rect 21364 41012 21416 41064
rect 21732 41012 21784 41064
rect 22192 41055 22244 41064
rect 22192 41021 22201 41055
rect 22201 41021 22235 41055
rect 22235 41021 22244 41055
rect 22192 41012 22244 41021
rect 22560 41012 22612 41064
rect 24124 41012 24176 41064
rect 24952 41055 25004 41064
rect 24952 41021 24961 41055
rect 24961 41021 24995 41055
rect 24995 41021 25004 41055
rect 24952 41012 25004 41021
rect 11336 40944 11388 40996
rect 4252 40876 4304 40928
rect 8576 40919 8628 40928
rect 8576 40885 8585 40919
rect 8585 40885 8619 40919
rect 8619 40885 8628 40919
rect 8576 40876 8628 40885
rect 11152 40919 11204 40928
rect 11152 40885 11161 40919
rect 11161 40885 11195 40919
rect 11195 40885 11204 40919
rect 11152 40876 11204 40885
rect 11888 40876 11940 40928
rect 13636 40876 13688 40928
rect 13820 40876 13872 40928
rect 14464 40876 14516 40928
rect 16856 40919 16908 40928
rect 16856 40885 16865 40919
rect 16865 40885 16899 40919
rect 16899 40885 16908 40919
rect 16856 40876 16908 40885
rect 17224 40876 17276 40928
rect 21548 40944 21600 40996
rect 19984 40876 20036 40928
rect 20536 40876 20588 40928
rect 26056 40944 26108 40996
rect 25320 40876 25372 40928
rect 2950 40774 3002 40826
rect 3014 40774 3066 40826
rect 3078 40774 3130 40826
rect 3142 40774 3194 40826
rect 3206 40774 3258 40826
rect 12950 40774 13002 40826
rect 13014 40774 13066 40826
rect 13078 40774 13130 40826
rect 13142 40774 13194 40826
rect 13206 40774 13258 40826
rect 22950 40774 23002 40826
rect 23014 40774 23066 40826
rect 23078 40774 23130 40826
rect 23142 40774 23194 40826
rect 23206 40774 23258 40826
rect 8576 40672 8628 40724
rect 9864 40672 9916 40724
rect 14372 40672 14424 40724
rect 15660 40672 15712 40724
rect 17500 40672 17552 40724
rect 3332 40604 3384 40656
rect 7840 40536 7892 40588
rect 11244 40536 11296 40588
rect 12164 40536 12216 40588
rect 5908 40468 5960 40520
rect 6368 40511 6420 40520
rect 6368 40477 6377 40511
rect 6377 40477 6411 40511
rect 6411 40477 6420 40511
rect 6368 40468 6420 40477
rect 13452 40536 13504 40588
rect 13360 40468 13412 40520
rect 13636 40468 13688 40520
rect 6736 40400 6788 40452
rect 4160 40332 4212 40384
rect 6552 40332 6604 40384
rect 7104 40400 7156 40452
rect 17868 40604 17920 40656
rect 20996 40604 21048 40656
rect 21640 40604 21692 40656
rect 24216 40604 24268 40656
rect 24768 40604 24820 40656
rect 16028 40579 16080 40588
rect 16028 40545 16037 40579
rect 16037 40545 16071 40579
rect 16071 40545 16080 40579
rect 16028 40536 16080 40545
rect 16672 40536 16724 40588
rect 15660 40468 15712 40520
rect 19156 40536 19208 40588
rect 20076 40536 20128 40588
rect 20720 40536 20772 40588
rect 21456 40536 21508 40588
rect 22284 40536 22336 40588
rect 24952 40536 25004 40588
rect 23388 40511 23440 40520
rect 23388 40477 23397 40511
rect 23397 40477 23431 40511
rect 23431 40477 23440 40511
rect 23388 40468 23440 40477
rect 8576 40332 8628 40384
rect 10232 40332 10284 40384
rect 16396 40400 16448 40452
rect 18696 40400 18748 40452
rect 21364 40400 21416 40452
rect 13360 40332 13412 40384
rect 14004 40332 14056 40384
rect 15476 40332 15528 40384
rect 16672 40332 16724 40384
rect 18328 40332 18380 40384
rect 18604 40332 18656 40384
rect 20168 40375 20220 40384
rect 20168 40341 20177 40375
rect 20177 40341 20211 40375
rect 20211 40341 20220 40375
rect 20168 40332 20220 40341
rect 21640 40332 21692 40384
rect 22836 40332 22888 40384
rect 24216 40375 24268 40384
rect 24216 40341 24225 40375
rect 24225 40341 24259 40375
rect 24259 40341 24268 40375
rect 24216 40332 24268 40341
rect 24768 40332 24820 40384
rect 7950 40230 8002 40282
rect 8014 40230 8066 40282
rect 8078 40230 8130 40282
rect 8142 40230 8194 40282
rect 8206 40230 8258 40282
rect 17950 40230 18002 40282
rect 18014 40230 18066 40282
rect 18078 40230 18130 40282
rect 18142 40230 18194 40282
rect 18206 40230 18258 40282
rect 7564 40128 7616 40180
rect 10048 40128 10100 40180
rect 6368 40060 6420 40112
rect 9404 40060 9456 40112
rect 14280 40128 14332 40180
rect 4068 39992 4120 40044
rect 7104 39924 7156 39976
rect 9680 39992 9732 40044
rect 13728 40060 13780 40112
rect 14372 40060 14424 40112
rect 20352 40128 20404 40180
rect 20536 40128 20588 40180
rect 20996 40171 21048 40180
rect 20996 40137 21005 40171
rect 21005 40137 21039 40171
rect 21039 40137 21048 40171
rect 20996 40128 21048 40137
rect 16396 40060 16448 40112
rect 16948 40060 17000 40112
rect 21732 40128 21784 40180
rect 22652 40128 22704 40180
rect 10232 39992 10284 40044
rect 12164 40035 12216 40044
rect 12164 40001 12173 40035
rect 12173 40001 12207 40035
rect 12207 40001 12216 40035
rect 12164 39992 12216 40001
rect 23664 40060 23716 40112
rect 12440 39967 12492 39976
rect 12440 39933 12449 39967
rect 12449 39933 12483 39967
rect 12483 39933 12492 39967
rect 12440 39924 12492 39933
rect 13820 39924 13872 39976
rect 14372 39967 14424 39976
rect 14372 39933 14381 39967
rect 14381 39933 14415 39967
rect 14415 39933 14424 39967
rect 14372 39924 14424 39933
rect 16948 39924 17000 39976
rect 7380 39788 7432 39840
rect 8208 39788 8260 39840
rect 10232 39831 10284 39840
rect 10232 39797 10241 39831
rect 10241 39797 10275 39831
rect 10275 39797 10284 39831
rect 10232 39788 10284 39797
rect 11336 39788 11388 39840
rect 11796 39788 11848 39840
rect 13912 39831 13964 39840
rect 13912 39797 13921 39831
rect 13921 39797 13955 39831
rect 13955 39797 13964 39831
rect 13912 39788 13964 39797
rect 15200 39831 15252 39840
rect 15200 39797 15209 39831
rect 15209 39797 15243 39831
rect 15243 39797 15252 39831
rect 15200 39788 15252 39797
rect 19708 39788 19760 39840
rect 21824 39992 21876 40044
rect 20720 39924 20772 39976
rect 22008 39924 22060 39976
rect 24584 39992 24636 40044
rect 19892 39856 19944 39908
rect 20076 39856 20128 39908
rect 20444 39788 20496 39840
rect 22652 39924 22704 39976
rect 23572 39924 23624 39976
rect 23664 39924 23716 39976
rect 24216 39924 24268 39976
rect 24952 39924 25004 39976
rect 25044 39967 25096 39976
rect 25044 39933 25053 39967
rect 25053 39933 25087 39967
rect 25087 39933 25096 39967
rect 25044 39924 25096 39933
rect 25320 39967 25372 39976
rect 25320 39933 25329 39967
rect 25329 39933 25363 39967
rect 25363 39933 25372 39967
rect 25320 39924 25372 39933
rect 2950 39686 3002 39738
rect 3014 39686 3066 39738
rect 3078 39686 3130 39738
rect 3142 39686 3194 39738
rect 3206 39686 3258 39738
rect 12950 39686 13002 39738
rect 13014 39686 13066 39738
rect 13078 39686 13130 39738
rect 13142 39686 13194 39738
rect 13206 39686 13258 39738
rect 22950 39686 23002 39738
rect 23014 39686 23066 39738
rect 23078 39686 23130 39738
rect 23142 39686 23194 39738
rect 23206 39686 23258 39738
rect 8392 39627 8444 39636
rect 8392 39593 8401 39627
rect 8401 39593 8435 39627
rect 8435 39593 8444 39627
rect 8392 39584 8444 39593
rect 6736 39516 6788 39568
rect 9864 39516 9916 39568
rect 14464 39584 14516 39636
rect 19524 39627 19576 39636
rect 19524 39593 19533 39627
rect 19533 39593 19567 39627
rect 19567 39593 19576 39627
rect 19524 39584 19576 39593
rect 20812 39584 20864 39636
rect 20996 39584 21048 39636
rect 22744 39584 22796 39636
rect 23204 39584 23256 39636
rect 23388 39584 23440 39636
rect 6920 39448 6972 39500
rect 7380 39380 7432 39432
rect 10692 39448 10744 39500
rect 8208 39380 8260 39432
rect 11888 39491 11940 39500
rect 11888 39457 11897 39491
rect 11897 39457 11931 39491
rect 11931 39457 11940 39491
rect 11888 39448 11940 39457
rect 12164 39491 12216 39500
rect 12164 39457 12173 39491
rect 12173 39457 12207 39491
rect 12207 39457 12216 39491
rect 12164 39448 12216 39457
rect 13636 39516 13688 39568
rect 13912 39448 13964 39500
rect 9312 39312 9364 39364
rect 9956 39312 10008 39364
rect 10508 39312 10560 39364
rect 8484 39244 8536 39296
rect 9864 39287 9916 39296
rect 9864 39253 9873 39287
rect 9873 39253 9907 39287
rect 9907 39253 9916 39287
rect 9864 39244 9916 39253
rect 12256 39380 12308 39432
rect 15200 39380 15252 39432
rect 18420 39516 18472 39568
rect 25044 39516 25096 39568
rect 17592 39491 17644 39500
rect 17592 39457 17601 39491
rect 17601 39457 17635 39491
rect 17635 39457 17644 39491
rect 17592 39448 17644 39457
rect 17684 39491 17736 39500
rect 17684 39457 17693 39491
rect 17693 39457 17727 39491
rect 17727 39457 17736 39491
rect 17684 39448 17736 39457
rect 20812 39448 20864 39500
rect 18788 39380 18840 39432
rect 21640 39448 21692 39500
rect 22836 39380 22888 39432
rect 19248 39312 19300 39364
rect 20628 39312 20680 39364
rect 11244 39244 11296 39296
rect 12624 39287 12676 39296
rect 12624 39253 12633 39287
rect 12633 39253 12667 39287
rect 12667 39253 12676 39287
rect 12624 39244 12676 39253
rect 14648 39287 14700 39296
rect 14648 39253 14657 39287
rect 14657 39253 14691 39287
rect 14691 39253 14700 39287
rect 14648 39244 14700 39253
rect 15936 39244 15988 39296
rect 16580 39244 16632 39296
rect 19800 39244 19852 39296
rect 19892 39287 19944 39296
rect 19892 39253 19901 39287
rect 19901 39253 19935 39287
rect 19935 39253 19944 39287
rect 19892 39244 19944 39253
rect 20076 39244 20128 39296
rect 22468 39312 22520 39364
rect 21916 39287 21968 39296
rect 21916 39253 21925 39287
rect 21925 39253 21959 39287
rect 21959 39253 21968 39287
rect 21916 39244 21968 39253
rect 22100 39244 22152 39296
rect 23388 39380 23440 39432
rect 24676 39448 24728 39500
rect 25412 39380 25464 39432
rect 23204 39312 23256 39364
rect 25136 39312 25188 39364
rect 24032 39244 24084 39296
rect 24676 39244 24728 39296
rect 7950 39142 8002 39194
rect 8014 39142 8066 39194
rect 8078 39142 8130 39194
rect 8142 39142 8194 39194
rect 8206 39142 8258 39194
rect 17950 39142 18002 39194
rect 18014 39142 18066 39194
rect 18078 39142 18130 39194
rect 18142 39142 18194 39194
rect 18206 39142 18258 39194
rect 4988 38972 5040 39024
rect 6736 39040 6788 39092
rect 9772 39083 9824 39092
rect 9772 39049 9781 39083
rect 9781 39049 9815 39083
rect 9815 39049 9824 39083
rect 9772 39040 9824 39049
rect 12348 39040 12400 39092
rect 12900 39083 12952 39092
rect 12900 39049 12909 39083
rect 12909 39049 12943 39083
rect 12943 39049 12952 39083
rect 12900 39040 12952 39049
rect 13728 39040 13780 39092
rect 14372 39040 14424 39092
rect 15476 39040 15528 39092
rect 16856 39040 16908 39092
rect 17592 39040 17644 39092
rect 17868 39040 17920 39092
rect 20168 39083 20220 39092
rect 20168 39049 20177 39083
rect 20177 39049 20211 39083
rect 20211 39049 20220 39083
rect 20168 39040 20220 39049
rect 20628 39040 20680 39092
rect 6552 38972 6604 39024
rect 10324 38972 10376 39024
rect 10508 38972 10560 39024
rect 14740 38972 14792 39024
rect 18604 38972 18656 39024
rect 19064 38972 19116 39024
rect 1216 38904 1268 38956
rect 12164 38947 12216 38956
rect 12164 38913 12173 38947
rect 12173 38913 12207 38947
rect 12207 38913 12216 38947
rect 12164 38904 12216 38913
rect 3976 38700 4028 38752
rect 4988 38836 5040 38888
rect 8576 38879 8628 38888
rect 8576 38845 8585 38879
rect 8585 38845 8619 38879
rect 8619 38845 8628 38879
rect 8576 38836 8628 38845
rect 10416 38879 10468 38888
rect 10416 38845 10425 38879
rect 10425 38845 10459 38879
rect 10459 38845 10468 38879
rect 10416 38836 10468 38845
rect 11060 38836 11112 38888
rect 11796 38836 11848 38888
rect 11980 38836 12032 38888
rect 12256 38836 12308 38888
rect 14096 38904 14148 38956
rect 15200 38904 15252 38956
rect 12440 38768 12492 38820
rect 5908 38700 5960 38752
rect 11336 38700 11388 38752
rect 12256 38700 12308 38752
rect 12348 38700 12400 38752
rect 12900 38700 12952 38752
rect 15568 38879 15620 38888
rect 15568 38845 15577 38879
rect 15577 38845 15611 38879
rect 15611 38845 15620 38879
rect 15568 38836 15620 38845
rect 18604 38836 18656 38888
rect 17316 38768 17368 38820
rect 19524 38836 19576 38888
rect 19616 38836 19668 38888
rect 21364 38904 21416 38956
rect 22008 38972 22060 39024
rect 22652 38972 22704 39024
rect 24308 38972 24360 39024
rect 25044 38972 25096 39024
rect 22100 38904 22152 38956
rect 20168 38836 20220 38888
rect 21824 38836 21876 38888
rect 22008 38836 22060 38888
rect 22468 38836 22520 38888
rect 14924 38700 14976 38752
rect 15292 38700 15344 38752
rect 17408 38700 17460 38752
rect 18972 38700 19024 38752
rect 23388 38768 23440 38820
rect 20536 38700 20588 38752
rect 22008 38743 22060 38752
rect 22008 38709 22017 38743
rect 22017 38709 22051 38743
rect 22051 38709 22060 38743
rect 22008 38700 22060 38709
rect 22100 38700 22152 38752
rect 22376 38700 22428 38752
rect 2950 38598 3002 38650
rect 3014 38598 3066 38650
rect 3078 38598 3130 38650
rect 3142 38598 3194 38650
rect 3206 38598 3258 38650
rect 12950 38598 13002 38650
rect 13014 38598 13066 38650
rect 13078 38598 13130 38650
rect 13142 38598 13194 38650
rect 13206 38598 13258 38650
rect 22950 38598 23002 38650
rect 23014 38598 23066 38650
rect 23078 38598 23130 38650
rect 23142 38598 23194 38650
rect 23206 38598 23258 38650
rect 6920 38496 6972 38548
rect 8300 38496 8352 38548
rect 9312 38496 9364 38548
rect 8116 38428 8168 38480
rect 11336 38496 11388 38548
rect 12072 38496 12124 38548
rect 12716 38496 12768 38548
rect 12992 38496 13044 38548
rect 16580 38496 16632 38548
rect 16764 38496 16816 38548
rect 22744 38496 22796 38548
rect 5908 38360 5960 38412
rect 7840 38360 7892 38412
rect 7196 38292 7248 38344
rect 8116 38335 8168 38344
rect 8116 38301 8125 38335
rect 8125 38301 8159 38335
rect 8159 38301 8168 38335
rect 8116 38292 8168 38301
rect 8576 38292 8628 38344
rect 9588 38360 9640 38412
rect 9864 38360 9916 38412
rect 10140 38403 10192 38412
rect 10140 38369 10149 38403
rect 10149 38369 10183 38403
rect 10183 38369 10192 38403
rect 10140 38360 10192 38369
rect 11520 38360 11572 38412
rect 6092 38224 6144 38276
rect 10140 38224 10192 38276
rect 11060 38335 11112 38344
rect 11060 38301 11069 38335
rect 11069 38301 11103 38335
rect 11103 38301 11112 38335
rect 11060 38292 11112 38301
rect 15568 38360 15620 38412
rect 15844 38403 15896 38412
rect 15844 38369 15853 38403
rect 15853 38369 15887 38403
rect 15887 38369 15896 38403
rect 15844 38360 15896 38369
rect 22928 38428 22980 38480
rect 25964 38496 26016 38548
rect 19984 38360 20036 38412
rect 22100 38360 22152 38412
rect 22652 38360 22704 38412
rect 25136 38428 25188 38480
rect 23296 38403 23348 38412
rect 23296 38369 23305 38403
rect 23305 38369 23339 38403
rect 23339 38369 23348 38403
rect 23296 38360 23348 38369
rect 19432 38292 19484 38344
rect 22284 38335 22336 38344
rect 22284 38301 22293 38335
rect 22293 38301 22327 38335
rect 22327 38301 22336 38335
rect 22284 38292 22336 38301
rect 23388 38292 23440 38344
rect 25412 38292 25464 38344
rect 11244 38224 11296 38276
rect 12072 38224 12124 38276
rect 15292 38224 15344 38276
rect 17500 38224 17552 38276
rect 6552 38156 6604 38208
rect 8300 38156 8352 38208
rect 9864 38199 9916 38208
rect 9864 38165 9873 38199
rect 9873 38165 9907 38199
rect 9907 38165 9916 38199
rect 9864 38156 9916 38165
rect 10968 38199 11020 38208
rect 10968 38165 10977 38199
rect 10977 38165 11011 38199
rect 11011 38165 11020 38199
rect 10968 38156 11020 38165
rect 12256 38156 12308 38208
rect 12624 38156 12676 38208
rect 14464 38199 14516 38208
rect 14464 38165 14473 38199
rect 14473 38165 14507 38199
rect 14507 38165 14516 38199
rect 14464 38156 14516 38165
rect 16120 38156 16172 38208
rect 16488 38156 16540 38208
rect 18604 38156 18656 38208
rect 19340 38156 19392 38208
rect 20720 38156 20772 38208
rect 21088 38199 21140 38208
rect 21088 38165 21097 38199
rect 21097 38165 21131 38199
rect 21131 38165 21140 38199
rect 22468 38224 22520 38276
rect 21088 38156 21140 38165
rect 21548 38156 21600 38208
rect 22836 38156 22888 38208
rect 23756 38199 23808 38208
rect 23756 38165 23765 38199
rect 23765 38165 23799 38199
rect 23799 38165 23808 38199
rect 23756 38156 23808 38165
rect 24492 38199 24544 38208
rect 24492 38165 24501 38199
rect 24501 38165 24535 38199
rect 24535 38165 24544 38199
rect 24492 38156 24544 38165
rect 24768 38156 24820 38208
rect 7950 38054 8002 38106
rect 8014 38054 8066 38106
rect 8078 38054 8130 38106
rect 8142 38054 8194 38106
rect 8206 38054 8258 38106
rect 17950 38054 18002 38106
rect 18014 38054 18066 38106
rect 18078 38054 18130 38106
rect 18142 38054 18194 38106
rect 18206 38054 18258 38106
rect 10876 37995 10928 38004
rect 10876 37961 10885 37995
rect 10885 37961 10919 37995
rect 10919 37961 10928 37995
rect 10876 37952 10928 37961
rect 12164 37952 12216 38004
rect 12900 37952 12952 38004
rect 15200 37952 15252 38004
rect 15384 37995 15436 38004
rect 15384 37961 15393 37995
rect 15393 37961 15427 37995
rect 15427 37961 15436 37995
rect 15384 37952 15436 37961
rect 16120 37995 16172 38004
rect 16120 37961 16129 37995
rect 16129 37961 16163 37995
rect 16163 37961 16172 37995
rect 16120 37952 16172 37961
rect 9312 37884 9364 37936
rect 10416 37884 10468 37936
rect 10692 37884 10744 37936
rect 15568 37884 15620 37936
rect 8300 37816 8352 37868
rect 9680 37859 9732 37868
rect 9680 37825 9689 37859
rect 9689 37825 9723 37859
rect 9723 37825 9732 37859
rect 9680 37816 9732 37825
rect 10508 37859 10560 37868
rect 10508 37825 10517 37859
rect 10517 37825 10551 37859
rect 10551 37825 10560 37859
rect 10508 37816 10560 37825
rect 7380 37748 7432 37800
rect 9404 37748 9456 37800
rect 10416 37791 10468 37800
rect 10416 37757 10425 37791
rect 10425 37757 10459 37791
rect 10459 37757 10468 37791
rect 10416 37748 10468 37757
rect 12992 37791 13044 37800
rect 12992 37757 13001 37791
rect 13001 37757 13035 37791
rect 13035 37757 13044 37791
rect 12992 37748 13044 37757
rect 15200 37816 15252 37868
rect 19524 37952 19576 38004
rect 22192 37952 22244 38004
rect 22376 37995 22428 38004
rect 22376 37961 22385 37995
rect 22385 37961 22419 37995
rect 22419 37961 22428 37995
rect 22376 37952 22428 37961
rect 18604 37884 18656 37936
rect 22100 37884 22152 37936
rect 10876 37680 10928 37732
rect 7472 37612 7524 37664
rect 10968 37612 11020 37664
rect 12808 37680 12860 37732
rect 13360 37748 13412 37800
rect 13728 37748 13780 37800
rect 15660 37680 15712 37732
rect 11520 37655 11572 37664
rect 11520 37621 11529 37655
rect 11529 37621 11563 37655
rect 11563 37621 11572 37655
rect 11520 37612 11572 37621
rect 12348 37612 12400 37664
rect 14924 37655 14976 37664
rect 14924 37621 14933 37655
rect 14933 37621 14967 37655
rect 14967 37621 14976 37655
rect 14924 37612 14976 37621
rect 17316 37791 17368 37800
rect 17316 37757 17325 37791
rect 17325 37757 17359 37791
rect 17359 37757 17368 37791
rect 17316 37748 17368 37757
rect 18052 37748 18104 37800
rect 19156 37816 19208 37868
rect 19892 37816 19944 37868
rect 21548 37816 21600 37868
rect 23388 37884 23440 37936
rect 18788 37791 18840 37800
rect 18788 37757 18797 37791
rect 18797 37757 18831 37791
rect 18831 37757 18840 37791
rect 18788 37748 18840 37757
rect 19432 37791 19484 37800
rect 19432 37757 19441 37791
rect 19441 37757 19475 37791
rect 19475 37757 19484 37791
rect 19432 37748 19484 37757
rect 19708 37680 19760 37732
rect 20812 37748 20864 37800
rect 23848 37748 23900 37800
rect 24124 37748 24176 37800
rect 20628 37680 20680 37732
rect 22468 37680 22520 37732
rect 24492 37680 24544 37732
rect 18420 37612 18472 37664
rect 19892 37655 19944 37664
rect 19892 37621 19901 37655
rect 19901 37621 19935 37655
rect 19935 37621 19944 37655
rect 19892 37612 19944 37621
rect 22652 37612 22704 37664
rect 22928 37612 22980 37664
rect 23480 37655 23532 37664
rect 23480 37621 23510 37655
rect 23510 37621 23532 37655
rect 23480 37612 23532 37621
rect 25136 37612 25188 37664
rect 25320 37655 25372 37664
rect 25320 37621 25329 37655
rect 25329 37621 25363 37655
rect 25363 37621 25372 37655
rect 25320 37612 25372 37621
rect 2950 37510 3002 37562
rect 3014 37510 3066 37562
rect 3078 37510 3130 37562
rect 3142 37510 3194 37562
rect 3206 37510 3258 37562
rect 12950 37510 13002 37562
rect 13014 37510 13066 37562
rect 13078 37510 13130 37562
rect 13142 37510 13194 37562
rect 13206 37510 13258 37562
rect 22950 37510 23002 37562
rect 23014 37510 23066 37562
rect 23078 37510 23130 37562
rect 23142 37510 23194 37562
rect 23206 37510 23258 37562
rect 5908 37408 5960 37460
rect 7472 37408 7524 37460
rect 8300 37408 8352 37460
rect 9128 37408 9180 37460
rect 10416 37408 10468 37460
rect 10784 37408 10836 37460
rect 12624 37408 12676 37460
rect 12808 37451 12860 37460
rect 12808 37417 12817 37451
rect 12817 37417 12851 37451
rect 12851 37417 12860 37451
rect 12808 37408 12860 37417
rect 6920 37272 6972 37324
rect 7196 37272 7248 37324
rect 10784 37272 10836 37324
rect 10876 37315 10928 37324
rect 10876 37281 10885 37315
rect 10885 37281 10919 37315
rect 10919 37281 10928 37315
rect 10876 37272 10928 37281
rect 11428 37272 11480 37324
rect 12072 37272 12124 37324
rect 12624 37272 12676 37324
rect 15844 37272 15896 37324
rect 18052 37340 18104 37392
rect 17776 37315 17828 37324
rect 17776 37281 17785 37315
rect 17785 37281 17819 37315
rect 17819 37281 17828 37315
rect 17776 37272 17828 37281
rect 20904 37408 20956 37460
rect 20996 37408 21048 37460
rect 23848 37408 23900 37460
rect 25504 37408 25556 37460
rect 25688 37340 25740 37392
rect 18420 37315 18472 37324
rect 18420 37281 18429 37315
rect 18429 37281 18463 37315
rect 18463 37281 18472 37315
rect 18420 37272 18472 37281
rect 22284 37272 22336 37324
rect 5264 37247 5316 37256
rect 5264 37213 5273 37247
rect 5273 37213 5307 37247
rect 5307 37213 5316 37247
rect 5264 37204 5316 37213
rect 9956 37204 10008 37256
rect 10048 37204 10100 37256
rect 15292 37204 15344 37256
rect 19432 37204 19484 37256
rect 19524 37247 19576 37256
rect 19524 37213 19533 37247
rect 19533 37213 19567 37247
rect 19567 37213 19576 37247
rect 19524 37204 19576 37213
rect 24400 37272 24452 37324
rect 6552 37136 6604 37188
rect 7104 37136 7156 37188
rect 7748 37111 7800 37120
rect 7748 37077 7757 37111
rect 7757 37077 7791 37111
rect 7791 37077 7800 37111
rect 7748 37068 7800 37077
rect 11244 37136 11296 37188
rect 10876 37068 10928 37120
rect 17500 37136 17552 37188
rect 17960 37136 18012 37188
rect 15476 37111 15528 37120
rect 15476 37077 15485 37111
rect 15485 37077 15519 37111
rect 15519 37077 15528 37111
rect 16028 37111 16080 37120
rect 15476 37068 15528 37077
rect 16028 37077 16037 37111
rect 16037 37077 16071 37111
rect 16071 37077 16080 37111
rect 16028 37068 16080 37077
rect 16304 37068 16356 37120
rect 19064 37136 19116 37188
rect 20720 37136 20772 37188
rect 21640 37136 21692 37188
rect 25320 37247 25372 37256
rect 25320 37213 25329 37247
rect 25329 37213 25363 37247
rect 25363 37213 25372 37247
rect 25320 37204 25372 37213
rect 24952 37136 25004 37188
rect 20444 37068 20496 37120
rect 23020 37068 23072 37120
rect 23848 37111 23900 37120
rect 23848 37077 23857 37111
rect 23857 37077 23891 37111
rect 23891 37077 23900 37111
rect 23848 37068 23900 37077
rect 24124 37068 24176 37120
rect 7950 36966 8002 37018
rect 8014 36966 8066 37018
rect 8078 36966 8130 37018
rect 8142 36966 8194 37018
rect 8206 36966 8258 37018
rect 17950 36966 18002 37018
rect 18014 36966 18066 37018
rect 18078 36966 18130 37018
rect 18142 36966 18194 37018
rect 18206 36966 18258 37018
rect 5172 36907 5224 36916
rect 5172 36873 5181 36907
rect 5181 36873 5215 36907
rect 5215 36873 5224 36907
rect 5172 36864 5224 36873
rect 9128 36864 9180 36916
rect 9312 36907 9364 36916
rect 9312 36873 9321 36907
rect 9321 36873 9355 36907
rect 9355 36873 9364 36907
rect 9312 36864 9364 36873
rect 9496 36864 9548 36916
rect 10508 36864 10560 36916
rect 12072 36907 12124 36916
rect 12072 36873 12081 36907
rect 12081 36873 12115 36907
rect 12115 36873 12124 36907
rect 12072 36864 12124 36873
rect 12164 36907 12216 36916
rect 12164 36873 12173 36907
rect 12173 36873 12207 36907
rect 12207 36873 12216 36907
rect 12164 36864 12216 36873
rect 12440 36864 12492 36916
rect 14464 36864 14516 36916
rect 15292 36907 15344 36916
rect 15292 36873 15301 36907
rect 15301 36873 15335 36907
rect 15335 36873 15344 36907
rect 15292 36864 15344 36873
rect 16488 36864 16540 36916
rect 18236 36864 18288 36916
rect 18328 36864 18380 36916
rect 19248 36864 19300 36916
rect 22008 36864 22060 36916
rect 8300 36796 8352 36848
rect 13544 36796 13596 36848
rect 15384 36796 15436 36848
rect 16304 36839 16356 36848
rect 16304 36805 16313 36839
rect 16313 36805 16347 36839
rect 16347 36805 16356 36839
rect 16304 36796 16356 36805
rect 17316 36796 17368 36848
rect 1308 36728 1360 36780
rect 5356 36728 5408 36780
rect 10140 36771 10192 36780
rect 10140 36737 10149 36771
rect 10149 36737 10183 36771
rect 10183 36737 10192 36771
rect 10140 36728 10192 36737
rect 10968 36728 11020 36780
rect 16764 36728 16816 36780
rect 4988 36592 5040 36644
rect 7564 36703 7616 36712
rect 7564 36669 7573 36703
rect 7573 36669 7607 36703
rect 7607 36669 7616 36703
rect 7564 36660 7616 36669
rect 9404 36660 9456 36712
rect 9496 36660 9548 36712
rect 11612 36660 11664 36712
rect 11244 36592 11296 36644
rect 1952 36524 2004 36576
rect 9588 36524 9640 36576
rect 11888 36592 11940 36644
rect 15844 36703 15896 36712
rect 15844 36669 15853 36703
rect 15853 36669 15887 36703
rect 15887 36669 15896 36703
rect 15844 36660 15896 36669
rect 16304 36660 16356 36712
rect 19064 36728 19116 36780
rect 18512 36660 18564 36712
rect 19156 36660 19208 36712
rect 19432 36796 19484 36848
rect 23848 36864 23900 36916
rect 23020 36839 23072 36848
rect 23020 36805 23029 36839
rect 23029 36805 23063 36839
rect 23063 36805 23072 36839
rect 23020 36796 23072 36805
rect 24400 36796 24452 36848
rect 22192 36728 22244 36780
rect 22284 36728 22336 36780
rect 24768 36728 24820 36780
rect 21732 36660 21784 36712
rect 23020 36660 23072 36712
rect 15200 36592 15252 36644
rect 20720 36592 20772 36644
rect 16856 36524 16908 36576
rect 18512 36524 18564 36576
rect 19156 36567 19208 36576
rect 19156 36533 19165 36567
rect 19165 36533 19199 36567
rect 19199 36533 19208 36567
rect 19156 36524 19208 36533
rect 23204 36524 23256 36576
rect 24492 36567 24544 36576
rect 24492 36533 24501 36567
rect 24501 36533 24535 36567
rect 24535 36533 24544 36567
rect 24492 36524 24544 36533
rect 2950 36422 3002 36474
rect 3014 36422 3066 36474
rect 3078 36422 3130 36474
rect 3142 36422 3194 36474
rect 3206 36422 3258 36474
rect 12950 36422 13002 36474
rect 13014 36422 13066 36474
rect 13078 36422 13130 36474
rect 13142 36422 13194 36474
rect 13206 36422 13258 36474
rect 22950 36422 23002 36474
rect 23014 36422 23066 36474
rect 23078 36422 23130 36474
rect 23142 36422 23194 36474
rect 23206 36422 23258 36474
rect 6092 36363 6144 36372
rect 6092 36329 6101 36363
rect 6101 36329 6135 36363
rect 6135 36329 6144 36363
rect 6092 36320 6144 36329
rect 8300 36320 8352 36372
rect 9312 36320 9364 36372
rect 15660 36320 15712 36372
rect 19340 36320 19392 36372
rect 19616 36363 19668 36372
rect 19616 36329 19625 36363
rect 19625 36329 19659 36363
rect 19659 36329 19668 36363
rect 19616 36320 19668 36329
rect 20444 36320 20496 36372
rect 9036 36252 9088 36304
rect 7012 36184 7064 36236
rect 7564 36184 7616 36236
rect 10508 36227 10560 36236
rect 10508 36193 10517 36227
rect 10517 36193 10551 36227
rect 10551 36193 10560 36227
rect 10508 36184 10560 36193
rect 15016 36184 15068 36236
rect 16028 36227 16080 36236
rect 16028 36193 16037 36227
rect 16037 36193 16071 36227
rect 16071 36193 16080 36227
rect 16028 36184 16080 36193
rect 10232 36116 10284 36168
rect 15200 36116 15252 36168
rect 17132 36295 17184 36304
rect 17132 36261 17141 36295
rect 17141 36261 17175 36295
rect 17175 36261 17184 36295
rect 17132 36252 17184 36261
rect 17224 36252 17276 36304
rect 21824 36320 21876 36372
rect 22836 36320 22888 36372
rect 22560 36252 22612 36304
rect 16304 36159 16356 36168
rect 16304 36125 16313 36159
rect 16313 36125 16347 36159
rect 16347 36125 16356 36159
rect 16304 36116 16356 36125
rect 6552 36048 6604 36100
rect 7380 35980 7432 36032
rect 9680 36048 9732 36100
rect 10876 36048 10928 36100
rect 11152 36048 11204 36100
rect 17592 36159 17644 36168
rect 17592 36125 17601 36159
rect 17601 36125 17635 36159
rect 17635 36125 17644 36159
rect 17592 36116 17644 36125
rect 18696 36116 18748 36168
rect 19432 36116 19484 36168
rect 20812 36184 20864 36236
rect 21088 36184 21140 36236
rect 23480 36320 23532 36372
rect 24492 36320 24544 36372
rect 23848 36252 23900 36304
rect 25044 36252 25096 36304
rect 23756 36184 23808 36236
rect 20444 36116 20496 36168
rect 21456 36116 21508 36168
rect 25320 36159 25372 36168
rect 25320 36125 25329 36159
rect 25329 36125 25363 36159
rect 25363 36125 25372 36159
rect 25320 36116 25372 36125
rect 20904 36048 20956 36100
rect 13360 35980 13412 36032
rect 14556 35980 14608 36032
rect 14740 36023 14792 36032
rect 14740 35989 14749 36023
rect 14749 35989 14783 36023
rect 14783 35989 14792 36023
rect 14740 35980 14792 35989
rect 16580 35980 16632 36032
rect 18420 35980 18472 36032
rect 20996 36023 21048 36032
rect 20996 35989 21005 36023
rect 21005 35989 21039 36023
rect 21039 35989 21048 36023
rect 20996 35980 21048 35989
rect 21456 35980 21508 36032
rect 21824 36023 21876 36032
rect 21824 35989 21833 36023
rect 21833 35989 21867 36023
rect 21867 35989 21876 36023
rect 21824 35980 21876 35989
rect 22100 35980 22152 36032
rect 23112 35980 23164 36032
rect 23296 35980 23348 36032
rect 23664 36023 23716 36032
rect 23664 35989 23673 36023
rect 23673 35989 23707 36023
rect 23707 35989 23716 36023
rect 23664 35980 23716 35989
rect 24584 35980 24636 36032
rect 7950 35878 8002 35930
rect 8014 35878 8066 35930
rect 8078 35878 8130 35930
rect 8142 35878 8194 35930
rect 8206 35878 8258 35930
rect 17950 35878 18002 35930
rect 18014 35878 18066 35930
rect 18078 35878 18130 35930
rect 18142 35878 18194 35930
rect 18206 35878 18258 35930
rect 7196 35776 7248 35828
rect 9404 35819 9456 35828
rect 9404 35785 9413 35819
rect 9413 35785 9447 35819
rect 9447 35785 9456 35819
rect 9404 35776 9456 35785
rect 11888 35776 11940 35828
rect 14188 35819 14240 35828
rect 14188 35785 14197 35819
rect 14197 35785 14231 35819
rect 14231 35785 14240 35819
rect 14188 35776 14240 35785
rect 16856 35819 16908 35828
rect 16856 35785 16865 35819
rect 16865 35785 16899 35819
rect 16899 35785 16908 35819
rect 16856 35776 16908 35785
rect 19708 35776 19760 35828
rect 20260 35776 20312 35828
rect 20812 35776 20864 35828
rect 23480 35776 23532 35828
rect 6552 35708 6604 35760
rect 9312 35708 9364 35760
rect 12164 35751 12216 35760
rect 12164 35717 12173 35751
rect 12173 35717 12207 35751
rect 12207 35717 12216 35751
rect 12164 35708 12216 35717
rect 15016 35708 15068 35760
rect 15384 35708 15436 35760
rect 18880 35708 18932 35760
rect 18972 35751 19024 35760
rect 18972 35717 18981 35751
rect 18981 35717 19015 35751
rect 19015 35717 19024 35751
rect 18972 35708 19024 35717
rect 19616 35708 19668 35760
rect 24400 35708 24452 35760
rect 4528 35615 4580 35624
rect 4528 35581 4537 35615
rect 4537 35581 4571 35615
rect 4571 35581 4580 35615
rect 4528 35572 4580 35581
rect 10232 35572 10284 35624
rect 11152 35615 11204 35624
rect 11152 35581 11161 35615
rect 11161 35581 11195 35615
rect 11195 35581 11204 35615
rect 11152 35572 11204 35581
rect 13820 35640 13872 35692
rect 13452 35572 13504 35624
rect 14372 35640 14424 35692
rect 5264 35436 5316 35488
rect 10232 35436 10284 35488
rect 10692 35436 10744 35488
rect 11244 35436 11296 35488
rect 11520 35479 11572 35488
rect 11520 35445 11529 35479
rect 11529 35445 11563 35479
rect 11563 35445 11572 35479
rect 11520 35436 11572 35445
rect 11704 35436 11756 35488
rect 14740 35615 14792 35624
rect 14740 35581 14749 35615
rect 14749 35581 14783 35615
rect 14783 35581 14792 35615
rect 14740 35572 14792 35581
rect 15660 35572 15712 35624
rect 14832 35504 14884 35556
rect 18696 35683 18748 35692
rect 18696 35649 18705 35683
rect 18705 35649 18739 35683
rect 18739 35649 18748 35683
rect 18696 35640 18748 35649
rect 19984 35572 20036 35624
rect 13820 35436 13872 35488
rect 18696 35436 18748 35488
rect 19524 35436 19576 35488
rect 19616 35436 19668 35488
rect 23848 35572 23900 35624
rect 25044 35615 25096 35624
rect 25044 35581 25053 35615
rect 25053 35581 25087 35615
rect 25087 35581 25096 35615
rect 25044 35572 25096 35581
rect 20352 35436 20404 35488
rect 22744 35436 22796 35488
rect 23940 35436 23992 35488
rect 25228 35436 25280 35488
rect 2950 35334 3002 35386
rect 3014 35334 3066 35386
rect 3078 35334 3130 35386
rect 3142 35334 3194 35386
rect 3206 35334 3258 35386
rect 12950 35334 13002 35386
rect 13014 35334 13066 35386
rect 13078 35334 13130 35386
rect 13142 35334 13194 35386
rect 13206 35334 13258 35386
rect 22950 35334 23002 35386
rect 23014 35334 23066 35386
rect 23078 35334 23130 35386
rect 23142 35334 23194 35386
rect 23206 35334 23258 35386
rect 4528 35232 4580 35284
rect 7656 35275 7708 35284
rect 7656 35241 7665 35275
rect 7665 35241 7699 35275
rect 7699 35241 7708 35275
rect 7656 35232 7708 35241
rect 10324 35275 10376 35284
rect 10324 35241 10333 35275
rect 10333 35241 10367 35275
rect 10367 35241 10376 35275
rect 10324 35232 10376 35241
rect 13728 35232 13780 35284
rect 14004 35232 14056 35284
rect 10784 35164 10836 35216
rect 6092 35096 6144 35148
rect 9404 35096 9456 35148
rect 7012 35071 7064 35080
rect 7012 35037 7021 35071
rect 7021 35037 7055 35071
rect 7055 35037 7064 35071
rect 7012 35028 7064 35037
rect 11704 35096 11756 35148
rect 12164 35096 12216 35148
rect 14096 35096 14148 35148
rect 10508 35028 10560 35080
rect 13728 35071 13780 35080
rect 13728 35037 13737 35071
rect 13737 35037 13771 35071
rect 13771 35037 13780 35071
rect 13728 35028 13780 35037
rect 7104 34960 7156 35012
rect 13176 34960 13228 35012
rect 13820 34960 13872 35012
rect 15936 35232 15988 35284
rect 16028 35232 16080 35284
rect 22744 35232 22796 35284
rect 23664 35232 23716 35284
rect 14648 35164 14700 35216
rect 18788 35164 18840 35216
rect 19616 35164 19668 35216
rect 20168 35164 20220 35216
rect 24124 35164 24176 35216
rect 17316 35096 17368 35148
rect 14740 35028 14792 35080
rect 16948 35028 17000 35080
rect 18880 35096 18932 35148
rect 18604 35028 18656 35080
rect 21732 35139 21784 35148
rect 21732 35105 21741 35139
rect 21741 35105 21775 35139
rect 21775 35105 21784 35139
rect 21732 35096 21784 35105
rect 21916 35096 21968 35148
rect 25044 35096 25096 35148
rect 20444 35028 20496 35080
rect 22284 35028 22336 35080
rect 6552 34892 6604 34944
rect 7288 34935 7340 34944
rect 7288 34901 7297 34935
rect 7297 34901 7331 34935
rect 7331 34901 7340 34935
rect 7288 34892 7340 34901
rect 7840 34892 7892 34944
rect 9036 34892 9088 34944
rect 9864 34935 9916 34944
rect 9864 34901 9873 34935
rect 9873 34901 9907 34935
rect 9907 34901 9916 34935
rect 9864 34892 9916 34901
rect 12164 34892 12216 34944
rect 14004 34892 14056 34944
rect 20168 34960 20220 35012
rect 25412 35028 25464 35080
rect 18696 34892 18748 34944
rect 20260 34892 20312 34944
rect 20720 34892 20772 34944
rect 22744 34892 22796 34944
rect 23204 34892 23256 34944
rect 24400 34892 24452 34944
rect 24768 34892 24820 34944
rect 7950 34790 8002 34842
rect 8014 34790 8066 34842
rect 8078 34790 8130 34842
rect 8142 34790 8194 34842
rect 8206 34790 8258 34842
rect 17950 34790 18002 34842
rect 18014 34790 18066 34842
rect 18078 34790 18130 34842
rect 18142 34790 18194 34842
rect 18206 34790 18258 34842
rect 2688 34688 2740 34740
rect 4988 34688 5040 34740
rect 5816 34688 5868 34740
rect 6552 34688 6604 34740
rect 7196 34688 7248 34740
rect 8484 34688 8536 34740
rect 7288 34620 7340 34672
rect 11152 34688 11204 34740
rect 1584 34595 1636 34604
rect 1584 34561 1593 34595
rect 1593 34561 1627 34595
rect 1627 34561 1636 34595
rect 1584 34552 1636 34561
rect 5264 34527 5316 34536
rect 5264 34493 5273 34527
rect 5273 34493 5307 34527
rect 5307 34493 5316 34527
rect 6736 34527 6788 34536
rect 5264 34484 5316 34493
rect 6736 34493 6745 34527
rect 6745 34493 6779 34527
rect 6779 34493 6788 34527
rect 6736 34484 6788 34493
rect 7012 34484 7064 34536
rect 7656 34484 7708 34536
rect 9772 34620 9824 34672
rect 13176 34620 13228 34672
rect 13728 34688 13780 34740
rect 14004 34688 14056 34740
rect 16028 34688 16080 34740
rect 16856 34688 16908 34740
rect 14280 34620 14332 34672
rect 18236 34620 18288 34672
rect 18972 34688 19024 34740
rect 19340 34620 19392 34672
rect 19524 34620 19576 34672
rect 10048 34484 10100 34536
rect 19064 34552 19116 34604
rect 19248 34552 19300 34604
rect 12808 34484 12860 34536
rect 13452 34416 13504 34468
rect 4988 34391 5040 34400
rect 4988 34357 5009 34391
rect 5009 34357 5040 34391
rect 4988 34348 5040 34357
rect 11704 34391 11756 34400
rect 11704 34357 11713 34391
rect 11713 34357 11747 34391
rect 11747 34357 11756 34391
rect 11704 34348 11756 34357
rect 14556 34348 14608 34400
rect 16764 34484 16816 34536
rect 19432 34484 19484 34536
rect 19708 34552 19760 34604
rect 22376 34731 22428 34740
rect 22376 34697 22385 34731
rect 22385 34697 22419 34731
rect 22419 34697 22428 34731
rect 22376 34688 22428 34697
rect 22468 34731 22520 34740
rect 22468 34697 22477 34731
rect 22477 34697 22511 34731
rect 22511 34697 22520 34731
rect 22468 34688 22520 34697
rect 23204 34731 23256 34740
rect 23204 34697 23213 34731
rect 23213 34697 23247 34731
rect 23247 34697 23256 34731
rect 23204 34688 23256 34697
rect 20260 34527 20312 34536
rect 20260 34493 20269 34527
rect 20269 34493 20303 34527
rect 20303 34493 20312 34527
rect 20260 34484 20312 34493
rect 25228 34552 25280 34604
rect 25320 34595 25372 34604
rect 25320 34561 25329 34595
rect 25329 34561 25363 34595
rect 25363 34561 25372 34595
rect 25320 34552 25372 34561
rect 22284 34484 22336 34536
rect 20168 34416 20220 34468
rect 23664 34484 23716 34536
rect 19064 34391 19116 34400
rect 19064 34357 19073 34391
rect 19073 34357 19107 34391
rect 19107 34357 19116 34391
rect 19064 34348 19116 34357
rect 22008 34391 22060 34400
rect 22008 34357 22017 34391
rect 22017 34357 22051 34391
rect 22051 34357 22060 34391
rect 22008 34348 22060 34357
rect 22468 34348 22520 34400
rect 2950 34246 3002 34298
rect 3014 34246 3066 34298
rect 3078 34246 3130 34298
rect 3142 34246 3194 34298
rect 3206 34246 3258 34298
rect 12950 34246 13002 34298
rect 13014 34246 13066 34298
rect 13078 34246 13130 34298
rect 13142 34246 13194 34298
rect 13206 34246 13258 34298
rect 22950 34246 23002 34298
rect 23014 34246 23066 34298
rect 23078 34246 23130 34298
rect 23142 34246 23194 34298
rect 23206 34246 23258 34298
rect 7288 34144 7340 34196
rect 8484 34144 8536 34196
rect 9128 34187 9180 34196
rect 9128 34153 9137 34187
rect 9137 34153 9171 34187
rect 9171 34153 9180 34187
rect 9128 34144 9180 34153
rect 10968 34144 11020 34196
rect 20720 34144 20772 34196
rect 21640 34144 21692 34196
rect 4712 34008 4764 34060
rect 4988 34008 5040 34060
rect 9588 34051 9640 34060
rect 9588 34017 9597 34051
rect 9597 34017 9631 34051
rect 9631 34017 9640 34051
rect 9588 34008 9640 34017
rect 6736 33940 6788 33992
rect 7748 33940 7800 33992
rect 9220 33940 9272 33992
rect 22284 34008 22336 34060
rect 23480 34008 23532 34060
rect 13360 33940 13412 33992
rect 20260 33940 20312 33992
rect 23572 33983 23624 33992
rect 23572 33949 23581 33983
rect 23581 33949 23615 33983
rect 23615 33949 23624 33983
rect 23572 33940 23624 33949
rect 24676 33940 24728 33992
rect 5816 33872 5868 33924
rect 7288 33872 7340 33924
rect 15660 33872 15712 33924
rect 19524 33872 19576 33924
rect 20628 33872 20680 33924
rect 22652 33872 22704 33924
rect 24860 33872 24912 33924
rect 12348 33804 12400 33856
rect 13728 33804 13780 33856
rect 18236 33804 18288 33856
rect 18788 33847 18840 33856
rect 18788 33813 18797 33847
rect 18797 33813 18831 33847
rect 18831 33813 18840 33847
rect 18788 33804 18840 33813
rect 18972 33847 19024 33856
rect 18972 33813 18981 33847
rect 18981 33813 19015 33847
rect 19015 33813 19024 33847
rect 18972 33804 19024 33813
rect 22468 33804 22520 33856
rect 24400 33804 24452 33856
rect 24676 33804 24728 33856
rect 25320 33847 25372 33856
rect 25320 33813 25329 33847
rect 25329 33813 25363 33847
rect 25363 33813 25372 33847
rect 25320 33804 25372 33813
rect 7950 33702 8002 33754
rect 8014 33702 8066 33754
rect 8078 33702 8130 33754
rect 8142 33702 8194 33754
rect 8206 33702 8258 33754
rect 17950 33702 18002 33754
rect 18014 33702 18066 33754
rect 18078 33702 18130 33754
rect 18142 33702 18194 33754
rect 18206 33702 18258 33754
rect 7564 33600 7616 33652
rect 8484 33532 8536 33584
rect 9496 33643 9548 33652
rect 9496 33609 9505 33643
rect 9505 33609 9539 33643
rect 9539 33609 9548 33643
rect 9496 33600 9548 33609
rect 9956 33643 10008 33652
rect 9956 33609 9965 33643
rect 9965 33609 9999 33643
rect 9999 33609 10008 33643
rect 9956 33600 10008 33609
rect 11980 33600 12032 33652
rect 12256 33600 12308 33652
rect 13820 33600 13872 33652
rect 13912 33643 13964 33652
rect 13912 33609 13921 33643
rect 13921 33609 13955 33643
rect 13955 33609 13964 33643
rect 13912 33600 13964 33609
rect 14924 33643 14976 33652
rect 14924 33609 14933 33643
rect 14933 33609 14967 33643
rect 14967 33609 14976 33643
rect 14924 33600 14976 33609
rect 19616 33600 19668 33652
rect 21916 33600 21968 33652
rect 22652 33600 22704 33652
rect 25504 33600 25556 33652
rect 10692 33532 10744 33584
rect 11704 33532 11756 33584
rect 9772 33464 9824 33516
rect 9956 33464 10008 33516
rect 7748 33439 7800 33448
rect 7748 33405 7757 33439
rect 7757 33405 7791 33439
rect 7791 33405 7800 33439
rect 7748 33396 7800 33405
rect 9220 33396 9272 33448
rect 10416 33439 10468 33448
rect 10416 33405 10425 33439
rect 10425 33405 10459 33439
rect 10459 33405 10468 33439
rect 10416 33396 10468 33405
rect 10784 33396 10836 33448
rect 9036 33328 9088 33380
rect 9496 33328 9548 33380
rect 6460 33260 6512 33312
rect 11888 33464 11940 33516
rect 13912 33464 13964 33516
rect 11520 33396 11572 33448
rect 12072 33396 12124 33448
rect 12532 33439 12584 33448
rect 12532 33405 12541 33439
rect 12541 33405 12575 33439
rect 12575 33405 12584 33439
rect 12532 33396 12584 33405
rect 15568 33532 15620 33584
rect 15016 33507 15068 33516
rect 15016 33473 15025 33507
rect 15025 33473 15059 33507
rect 15059 33473 15068 33507
rect 15016 33464 15068 33473
rect 14096 33396 14148 33448
rect 23480 33507 23532 33516
rect 23480 33473 23489 33507
rect 23489 33473 23523 33507
rect 23523 33473 23532 33507
rect 23480 33464 23532 33473
rect 24860 33464 24912 33516
rect 13544 33328 13596 33380
rect 23756 33439 23808 33448
rect 23756 33405 23765 33439
rect 23765 33405 23799 33439
rect 23799 33405 23808 33439
rect 23756 33396 23808 33405
rect 23296 33328 23348 33380
rect 13452 33303 13504 33312
rect 13452 33269 13461 33303
rect 13461 33269 13495 33303
rect 13495 33269 13504 33303
rect 13452 33260 13504 33269
rect 16028 33260 16080 33312
rect 2950 33158 3002 33210
rect 3014 33158 3066 33210
rect 3078 33158 3130 33210
rect 3142 33158 3194 33210
rect 3206 33158 3258 33210
rect 12950 33158 13002 33210
rect 13014 33158 13066 33210
rect 13078 33158 13130 33210
rect 13142 33158 13194 33210
rect 13206 33158 13258 33210
rect 22950 33158 23002 33210
rect 23014 33158 23066 33210
rect 23078 33158 23130 33210
rect 23142 33158 23194 33210
rect 23206 33158 23258 33210
rect 7288 33099 7340 33108
rect 7288 33065 7297 33099
rect 7297 33065 7331 33099
rect 7331 33065 7340 33099
rect 7288 33056 7340 33065
rect 9312 33056 9364 33108
rect 9496 33056 9548 33108
rect 10140 33056 10192 33108
rect 15016 33056 15068 33108
rect 16948 33056 17000 33108
rect 17684 33056 17736 33108
rect 19524 33056 19576 33108
rect 21732 33056 21784 33108
rect 22560 33056 22612 33108
rect 23112 33056 23164 33108
rect 16672 32988 16724 33040
rect 7748 32920 7800 32972
rect 9220 32963 9272 32972
rect 9220 32929 9229 32963
rect 9229 32929 9263 32963
rect 9263 32929 9272 32963
rect 9220 32920 9272 32929
rect 9312 32920 9364 32972
rect 11612 32920 11664 32972
rect 12164 32963 12216 32972
rect 12164 32929 12173 32963
rect 12173 32929 12207 32963
rect 12207 32929 12216 32963
rect 12164 32920 12216 32929
rect 8300 32852 8352 32904
rect 13636 32920 13688 32972
rect 16856 32963 16908 32972
rect 16856 32929 16865 32963
rect 16865 32929 16899 32963
rect 16899 32929 16908 32963
rect 16856 32920 16908 32929
rect 18328 32988 18380 33040
rect 20168 32988 20220 33040
rect 12716 32852 12768 32904
rect 14556 32852 14608 32904
rect 15108 32852 15160 32904
rect 20720 32920 20772 32972
rect 6092 32784 6144 32836
rect 7104 32784 7156 32836
rect 8484 32784 8536 32836
rect 9772 32784 9824 32836
rect 15752 32784 15804 32836
rect 16120 32784 16172 32836
rect 9496 32759 9548 32768
rect 9496 32725 9505 32759
rect 9505 32725 9539 32759
rect 9539 32725 9548 32759
rect 9496 32716 9548 32725
rect 9588 32716 9640 32768
rect 13360 32716 13412 32768
rect 14004 32716 14056 32768
rect 16212 32716 16264 32768
rect 18144 32716 18196 32768
rect 18788 32716 18840 32768
rect 21916 32920 21968 32972
rect 22284 32920 22336 32972
rect 22560 32920 22612 32972
rect 22836 32920 22888 32972
rect 23296 32852 23348 32904
rect 25320 32895 25372 32904
rect 25320 32861 25329 32895
rect 25329 32861 25363 32895
rect 25363 32861 25372 32895
rect 25320 32852 25372 32861
rect 22468 32784 22520 32836
rect 23204 32784 23256 32836
rect 22652 32759 22704 32768
rect 22652 32725 22661 32759
rect 22661 32725 22695 32759
rect 22695 32725 22704 32759
rect 22652 32716 22704 32725
rect 23112 32759 23164 32768
rect 23112 32725 23121 32759
rect 23121 32725 23155 32759
rect 23155 32725 23164 32759
rect 23112 32716 23164 32725
rect 23664 32716 23716 32768
rect 7950 32614 8002 32666
rect 8014 32614 8066 32666
rect 8078 32614 8130 32666
rect 8142 32614 8194 32666
rect 8206 32614 8258 32666
rect 17950 32614 18002 32666
rect 18014 32614 18066 32666
rect 18078 32614 18130 32666
rect 18142 32614 18194 32666
rect 18206 32614 18258 32666
rect 7104 32555 7156 32564
rect 7104 32521 7113 32555
rect 7113 32521 7147 32555
rect 7147 32521 7156 32555
rect 7104 32512 7156 32521
rect 9496 32512 9548 32564
rect 9588 32512 9640 32564
rect 11244 32555 11296 32564
rect 11244 32521 11253 32555
rect 11253 32521 11287 32555
rect 11287 32521 11296 32555
rect 11244 32512 11296 32521
rect 12716 32555 12768 32564
rect 12716 32521 12725 32555
rect 12725 32521 12759 32555
rect 12759 32521 12768 32555
rect 12716 32512 12768 32521
rect 13360 32555 13412 32564
rect 13360 32521 13369 32555
rect 13369 32521 13403 32555
rect 13403 32521 13412 32555
rect 13360 32512 13412 32521
rect 14924 32512 14976 32564
rect 19064 32512 19116 32564
rect 19708 32512 19760 32564
rect 20904 32512 20956 32564
rect 21272 32512 21324 32564
rect 22100 32512 22152 32564
rect 8484 32444 8536 32496
rect 13728 32444 13780 32496
rect 17040 32444 17092 32496
rect 18512 32487 18564 32496
rect 18512 32453 18521 32487
rect 18521 32453 18555 32487
rect 18555 32453 18564 32487
rect 18512 32444 18564 32453
rect 19800 32444 19852 32496
rect 1308 32376 1360 32428
rect 16856 32376 16908 32428
rect 4988 32351 5040 32360
rect 4988 32317 4997 32351
rect 4997 32317 5031 32351
rect 5031 32317 5040 32351
rect 4988 32308 5040 32317
rect 7472 32351 7524 32360
rect 7472 32317 7481 32351
rect 7481 32317 7515 32351
rect 7515 32317 7524 32351
rect 7472 32308 7524 32317
rect 7748 32308 7800 32360
rect 9128 32351 9180 32360
rect 9128 32317 9137 32351
rect 9137 32317 9171 32351
rect 9171 32317 9180 32351
rect 9128 32308 9180 32317
rect 9404 32351 9456 32360
rect 9404 32317 9413 32351
rect 9413 32317 9447 32351
rect 9447 32317 9456 32351
rect 9404 32308 9456 32317
rect 11796 32308 11848 32360
rect 12532 32308 12584 32360
rect 13728 32308 13780 32360
rect 14464 32308 14516 32360
rect 14556 32308 14608 32360
rect 15936 32351 15988 32360
rect 15936 32317 15945 32351
rect 15945 32317 15979 32351
rect 15979 32317 15988 32351
rect 15936 32308 15988 32317
rect 18880 32376 18932 32428
rect 19984 32376 20036 32428
rect 6920 32240 6972 32292
rect 2596 32172 2648 32224
rect 9588 32172 9640 32224
rect 16948 32240 17000 32292
rect 11796 32172 11848 32224
rect 12716 32172 12768 32224
rect 14556 32172 14608 32224
rect 17316 32240 17368 32292
rect 17592 32215 17644 32224
rect 17592 32181 17601 32215
rect 17601 32181 17635 32215
rect 17635 32181 17644 32215
rect 17592 32172 17644 32181
rect 17868 32240 17920 32292
rect 21180 32351 21232 32360
rect 21180 32317 21189 32351
rect 21189 32317 21223 32351
rect 21223 32317 21232 32351
rect 21180 32308 21232 32317
rect 22376 32308 22428 32360
rect 25136 32512 25188 32564
rect 22928 32444 22980 32496
rect 23296 32376 23348 32428
rect 25320 32419 25372 32428
rect 25320 32385 25329 32419
rect 25329 32385 25363 32419
rect 25363 32385 25372 32419
rect 25320 32376 25372 32385
rect 23204 32351 23256 32360
rect 23204 32317 23213 32351
rect 23213 32317 23247 32351
rect 23247 32317 23256 32351
rect 23204 32308 23256 32317
rect 19984 32240 20036 32292
rect 20628 32215 20680 32224
rect 20628 32181 20637 32215
rect 20637 32181 20671 32215
rect 20671 32181 20680 32215
rect 20628 32172 20680 32181
rect 23940 32172 23992 32224
rect 24492 32172 24544 32224
rect 2950 32070 3002 32122
rect 3014 32070 3066 32122
rect 3078 32070 3130 32122
rect 3142 32070 3194 32122
rect 3206 32070 3258 32122
rect 12950 32070 13002 32122
rect 13014 32070 13066 32122
rect 13078 32070 13130 32122
rect 13142 32070 13194 32122
rect 13206 32070 13258 32122
rect 22950 32070 23002 32122
rect 23014 32070 23066 32122
rect 23078 32070 23130 32122
rect 23142 32070 23194 32122
rect 23206 32070 23258 32122
rect 6092 31968 6144 32020
rect 7288 31968 7340 32020
rect 10784 31968 10836 32020
rect 11244 32011 11296 32020
rect 11244 31977 11253 32011
rect 11253 31977 11287 32011
rect 11287 31977 11296 32011
rect 11244 31968 11296 31977
rect 12348 32011 12400 32020
rect 12348 31977 12357 32011
rect 12357 31977 12391 32011
rect 12391 31977 12400 32011
rect 12348 31968 12400 31977
rect 15936 31968 15988 32020
rect 7840 31900 7892 31952
rect 17684 32011 17736 32020
rect 17684 31977 17693 32011
rect 17693 31977 17727 32011
rect 17727 31977 17736 32011
rect 17684 31968 17736 31977
rect 8300 31832 8352 31884
rect 9220 31832 9272 31884
rect 11612 31832 11664 31884
rect 6920 31807 6972 31816
rect 6920 31773 6929 31807
rect 6929 31773 6963 31807
rect 6963 31773 6972 31807
rect 6920 31764 6972 31773
rect 7564 31764 7616 31816
rect 9036 31764 9088 31816
rect 9496 31764 9548 31816
rect 10968 31764 11020 31816
rect 16948 31875 17000 31884
rect 16948 31841 16957 31875
rect 16957 31841 16991 31875
rect 16991 31841 17000 31875
rect 16948 31832 17000 31841
rect 17040 31832 17092 31884
rect 19248 31900 19300 31952
rect 19800 31968 19852 32020
rect 19984 31968 20036 32020
rect 20444 31968 20496 32020
rect 20720 31968 20772 32020
rect 21088 31900 21140 31952
rect 22284 31900 22336 31952
rect 22376 31900 22428 31952
rect 22744 31900 22796 31952
rect 23388 31900 23440 31952
rect 7104 31696 7156 31748
rect 10600 31739 10652 31748
rect 10600 31705 10609 31739
rect 10609 31705 10643 31739
rect 10643 31705 10652 31739
rect 10600 31696 10652 31705
rect 12716 31739 12768 31748
rect 12716 31705 12725 31739
rect 12725 31705 12759 31739
rect 12759 31705 12768 31739
rect 12716 31696 12768 31705
rect 13728 31696 13780 31748
rect 16212 31696 16264 31748
rect 16672 31739 16724 31748
rect 16672 31705 16681 31739
rect 16681 31705 16715 31739
rect 16715 31705 16724 31739
rect 16672 31696 16724 31705
rect 18328 31696 18380 31748
rect 20352 31832 20404 31884
rect 22468 31832 22520 31884
rect 23296 31832 23348 31884
rect 22192 31807 22244 31816
rect 22192 31773 22201 31807
rect 22201 31773 22235 31807
rect 22235 31773 22244 31807
rect 22192 31764 22244 31773
rect 22744 31764 22796 31816
rect 20444 31696 20496 31748
rect 25596 31900 25648 31952
rect 25412 31764 25464 31816
rect 7840 31671 7892 31680
rect 7840 31637 7849 31671
rect 7849 31637 7883 31671
rect 7883 31637 7892 31671
rect 7840 31628 7892 31637
rect 9956 31628 10008 31680
rect 14464 31628 14516 31680
rect 19616 31628 19668 31680
rect 19892 31671 19944 31680
rect 19892 31637 19901 31671
rect 19901 31637 19935 31671
rect 19935 31637 19944 31671
rect 19892 31628 19944 31637
rect 20904 31628 20956 31680
rect 21180 31628 21232 31680
rect 21364 31628 21416 31680
rect 7950 31526 8002 31578
rect 8014 31526 8066 31578
rect 8078 31526 8130 31578
rect 8142 31526 8194 31578
rect 8206 31526 8258 31578
rect 17950 31526 18002 31578
rect 18014 31526 18066 31578
rect 18078 31526 18130 31578
rect 18142 31526 18194 31578
rect 18206 31526 18258 31578
rect 4988 31424 5040 31476
rect 5356 31424 5408 31476
rect 7656 31424 7708 31476
rect 7840 31424 7892 31476
rect 9864 31424 9916 31476
rect 10232 31424 10284 31476
rect 10508 31424 10560 31476
rect 10600 31424 10652 31476
rect 15384 31424 15436 31476
rect 16856 31424 16908 31476
rect 17592 31424 17644 31476
rect 19616 31424 19668 31476
rect 19892 31424 19944 31476
rect 20444 31467 20496 31476
rect 20444 31433 20453 31467
rect 20453 31433 20487 31467
rect 20487 31433 20496 31467
rect 20444 31424 20496 31433
rect 20996 31424 21048 31476
rect 23296 31424 23348 31476
rect 24860 31424 24912 31476
rect 17408 31356 17460 31408
rect 6828 31288 6880 31340
rect 7104 31288 7156 31340
rect 10048 31288 10100 31340
rect 11244 31288 11296 31340
rect 12256 31288 12308 31340
rect 18696 31288 18748 31340
rect 20536 31288 20588 31340
rect 23388 31331 23440 31340
rect 23388 31297 23397 31331
rect 23397 31297 23431 31331
rect 23431 31297 23440 31331
rect 23388 31288 23440 31297
rect 25320 31331 25372 31340
rect 25320 31297 25329 31331
rect 25329 31297 25363 31331
rect 25363 31297 25372 31331
rect 25320 31288 25372 31297
rect 4712 31263 4764 31272
rect 4712 31229 4721 31263
rect 4721 31229 4755 31263
rect 4755 31229 4764 31263
rect 4712 31220 4764 31229
rect 4804 31263 4856 31272
rect 4804 31229 4813 31263
rect 4813 31229 4847 31263
rect 4847 31229 4856 31263
rect 4804 31220 4856 31229
rect 4160 31152 4212 31204
rect 9864 31263 9916 31272
rect 9864 31229 9873 31263
rect 9873 31229 9907 31263
rect 9907 31229 9916 31263
rect 10600 31263 10652 31272
rect 9864 31220 9916 31229
rect 10600 31229 10609 31263
rect 10609 31229 10643 31263
rect 10643 31229 10652 31263
rect 10600 31220 10652 31229
rect 10876 31220 10928 31272
rect 17776 31263 17828 31272
rect 17776 31229 17785 31263
rect 17785 31229 17819 31263
rect 17819 31229 17828 31263
rect 17776 31220 17828 31229
rect 18052 31220 18104 31272
rect 7380 31152 7432 31204
rect 21272 31152 21324 31204
rect 21364 31152 21416 31204
rect 24308 31152 24360 31204
rect 6368 31084 6420 31136
rect 10048 31084 10100 31136
rect 12532 31084 12584 31136
rect 13360 31084 13412 31136
rect 17224 31127 17276 31136
rect 17224 31093 17233 31127
rect 17233 31093 17267 31127
rect 17267 31093 17276 31127
rect 17224 31084 17276 31093
rect 20904 31084 20956 31136
rect 21640 31084 21692 31136
rect 25044 31084 25096 31136
rect 2950 30982 3002 31034
rect 3014 30982 3066 31034
rect 3078 30982 3130 31034
rect 3142 30982 3194 31034
rect 3206 30982 3258 31034
rect 12950 30982 13002 31034
rect 13014 30982 13066 31034
rect 13078 30982 13130 31034
rect 13142 30982 13194 31034
rect 13206 30982 13258 31034
rect 22950 30982 23002 31034
rect 23014 30982 23066 31034
rect 23078 30982 23130 31034
rect 23142 30982 23194 31034
rect 23206 30982 23258 31034
rect 7748 30880 7800 30932
rect 10784 30880 10836 30932
rect 7288 30787 7340 30796
rect 7288 30753 7297 30787
rect 7297 30753 7331 30787
rect 7331 30753 7340 30787
rect 7288 30744 7340 30753
rect 10968 30744 11020 30796
rect 12808 30880 12860 30932
rect 17408 30880 17460 30932
rect 21180 30880 21232 30932
rect 24860 30880 24912 30932
rect 25320 30880 25372 30932
rect 16488 30812 16540 30864
rect 17684 30812 17736 30864
rect 7472 30719 7524 30728
rect 7472 30685 7481 30719
rect 7481 30685 7515 30719
rect 7515 30685 7524 30719
rect 7472 30676 7524 30685
rect 13820 30744 13872 30796
rect 14280 30719 14332 30728
rect 14280 30685 14289 30719
rect 14289 30685 14323 30719
rect 14323 30685 14332 30719
rect 14280 30676 14332 30685
rect 16948 30744 17000 30796
rect 17316 30744 17368 30796
rect 18144 30787 18196 30796
rect 18144 30753 18153 30787
rect 18153 30753 18187 30787
rect 18187 30753 18196 30787
rect 18144 30744 18196 30753
rect 18328 30787 18380 30796
rect 18328 30753 18337 30787
rect 18337 30753 18371 30787
rect 18371 30753 18380 30787
rect 18328 30744 18380 30753
rect 20720 30744 20772 30796
rect 22560 30744 22612 30796
rect 18052 30719 18104 30728
rect 18052 30685 18061 30719
rect 18061 30685 18095 30719
rect 18095 30685 18104 30719
rect 18052 30676 18104 30685
rect 19984 30676 20036 30728
rect 20812 30676 20864 30728
rect 21548 30676 21600 30728
rect 24584 30719 24636 30728
rect 24584 30685 24593 30719
rect 24593 30685 24627 30719
rect 24627 30685 24636 30719
rect 24584 30676 24636 30685
rect 10692 30608 10744 30660
rect 12256 30608 12308 30660
rect 13360 30651 13412 30660
rect 13360 30617 13369 30651
rect 13369 30617 13403 30651
rect 13403 30617 13412 30651
rect 13360 30608 13412 30617
rect 14464 30608 14516 30660
rect 14556 30651 14608 30660
rect 14556 30617 14565 30651
rect 14565 30617 14599 30651
rect 14599 30617 14608 30651
rect 14556 30608 14608 30617
rect 16120 30608 16172 30660
rect 6644 30540 6696 30592
rect 7012 30540 7064 30592
rect 12808 30540 12860 30592
rect 13544 30540 13596 30592
rect 16028 30583 16080 30592
rect 16028 30549 16037 30583
rect 16037 30549 16071 30583
rect 16071 30549 16080 30583
rect 16028 30540 16080 30549
rect 16304 30540 16356 30592
rect 17316 30540 17368 30592
rect 17684 30583 17736 30592
rect 17684 30549 17693 30583
rect 17693 30549 17727 30583
rect 17727 30549 17736 30583
rect 17684 30540 17736 30549
rect 22468 30608 22520 30660
rect 24860 30608 24912 30660
rect 18972 30540 19024 30592
rect 19432 30583 19484 30592
rect 19432 30549 19441 30583
rect 19441 30549 19475 30583
rect 19475 30549 19484 30583
rect 19432 30540 19484 30549
rect 19616 30540 19668 30592
rect 20812 30583 20864 30592
rect 20812 30549 20821 30583
rect 20821 30549 20855 30583
rect 20855 30549 20864 30583
rect 20812 30540 20864 30549
rect 23480 30540 23532 30592
rect 23572 30540 23624 30592
rect 24584 30540 24636 30592
rect 24768 30583 24820 30592
rect 24768 30549 24777 30583
rect 24777 30549 24811 30583
rect 24811 30549 24820 30583
rect 24768 30540 24820 30549
rect 7950 30438 8002 30490
rect 8014 30438 8066 30490
rect 8078 30438 8130 30490
rect 8142 30438 8194 30490
rect 8206 30438 8258 30490
rect 17950 30438 18002 30490
rect 18014 30438 18066 30490
rect 18078 30438 18130 30490
rect 18142 30438 18194 30490
rect 18206 30438 18258 30490
rect 7564 30336 7616 30388
rect 9128 30268 9180 30320
rect 15844 30336 15896 30388
rect 16120 30379 16172 30388
rect 16120 30345 16129 30379
rect 16129 30345 16163 30379
rect 16163 30345 16172 30379
rect 16120 30336 16172 30345
rect 16304 30336 16356 30388
rect 16488 30336 16540 30388
rect 10232 30268 10284 30320
rect 12992 30311 13044 30320
rect 12992 30277 13001 30311
rect 13001 30277 13035 30311
rect 13035 30277 13044 30311
rect 12992 30268 13044 30277
rect 15660 30268 15712 30320
rect 19432 30336 19484 30388
rect 18512 30268 18564 30320
rect 22284 30311 22336 30320
rect 22284 30277 22293 30311
rect 22293 30277 22327 30311
rect 22327 30277 22336 30311
rect 22284 30268 22336 30277
rect 22376 30311 22428 30320
rect 22376 30277 22385 30311
rect 22385 30277 22419 30311
rect 22419 30277 22428 30311
rect 22376 30268 22428 30277
rect 23664 30268 23716 30320
rect 24860 30336 24912 30388
rect 9496 30200 9548 30252
rect 11244 30200 11296 30252
rect 15016 30200 15068 30252
rect 9588 30132 9640 30184
rect 10968 30132 11020 30184
rect 14372 30132 14424 30184
rect 15384 30175 15436 30184
rect 15384 30141 15393 30175
rect 15393 30141 15427 30175
rect 15427 30141 15436 30175
rect 15384 30132 15436 30141
rect 16580 30200 16632 30252
rect 15752 30132 15804 30184
rect 10416 30064 10468 30116
rect 16856 30132 16908 30184
rect 18880 30243 18932 30252
rect 18880 30209 18889 30243
rect 18889 30209 18923 30243
rect 18923 30209 18932 30243
rect 18880 30200 18932 30209
rect 19064 30175 19116 30184
rect 19064 30141 19073 30175
rect 19073 30141 19107 30175
rect 19107 30141 19116 30175
rect 19064 30132 19116 30141
rect 19984 30175 20036 30184
rect 19984 30141 19993 30175
rect 19993 30141 20027 30175
rect 20027 30141 20036 30175
rect 19984 30132 20036 30141
rect 23572 30200 23624 30252
rect 20812 30132 20864 30184
rect 22192 30175 22244 30184
rect 22192 30141 22201 30175
rect 22201 30141 22235 30175
rect 22235 30141 22244 30175
rect 22192 30132 22244 30141
rect 22836 30132 22888 30184
rect 23756 30132 23808 30184
rect 24584 30132 24636 30184
rect 22560 30064 22612 30116
rect 14832 30039 14884 30048
rect 14832 30005 14841 30039
rect 14841 30005 14875 30039
rect 14875 30005 14884 30039
rect 14832 29996 14884 30005
rect 15844 29996 15896 30048
rect 16120 29996 16172 30048
rect 16212 29996 16264 30048
rect 20444 30039 20496 30048
rect 20444 30005 20453 30039
rect 20453 30005 20487 30039
rect 20487 30005 20496 30039
rect 20444 29996 20496 30005
rect 23388 29996 23440 30048
rect 2950 29894 3002 29946
rect 3014 29894 3066 29946
rect 3078 29894 3130 29946
rect 3142 29894 3194 29946
rect 3206 29894 3258 29946
rect 12950 29894 13002 29946
rect 13014 29894 13066 29946
rect 13078 29894 13130 29946
rect 13142 29894 13194 29946
rect 13206 29894 13258 29946
rect 22950 29894 23002 29946
rect 23014 29894 23066 29946
rect 23078 29894 23130 29946
rect 23142 29894 23194 29946
rect 23206 29894 23258 29946
rect 4344 29792 4396 29844
rect 1308 29656 1360 29708
rect 3976 29699 4028 29708
rect 3976 29665 3985 29699
rect 3985 29665 4019 29699
rect 4019 29665 4028 29699
rect 3976 29656 4028 29665
rect 1768 29631 1820 29640
rect 1768 29597 1777 29631
rect 1777 29597 1811 29631
rect 1811 29597 1820 29631
rect 1768 29588 1820 29597
rect 9036 29792 9088 29844
rect 12808 29792 12860 29844
rect 9588 29656 9640 29708
rect 10692 29699 10744 29708
rect 10692 29665 10701 29699
rect 10701 29665 10735 29699
rect 10735 29665 10744 29699
rect 10692 29656 10744 29665
rect 10876 29656 10928 29708
rect 9404 29588 9456 29640
rect 10968 29631 11020 29640
rect 10968 29597 10977 29631
rect 10977 29597 11011 29631
rect 11011 29597 11020 29631
rect 10968 29588 11020 29597
rect 15108 29792 15160 29844
rect 19064 29792 19116 29844
rect 25136 29835 25188 29844
rect 25136 29801 25145 29835
rect 25145 29801 25179 29835
rect 25179 29801 25188 29835
rect 25136 29792 25188 29801
rect 15016 29724 15068 29776
rect 16488 29724 16540 29776
rect 19248 29724 19300 29776
rect 21180 29724 21232 29776
rect 13452 29656 13504 29708
rect 17592 29656 17644 29708
rect 18236 29699 18288 29708
rect 18236 29665 18245 29699
rect 18245 29665 18279 29699
rect 18279 29665 18288 29699
rect 18236 29656 18288 29665
rect 19892 29699 19944 29708
rect 19892 29665 19901 29699
rect 19901 29665 19935 29699
rect 19935 29665 19944 29699
rect 19892 29656 19944 29665
rect 19984 29699 20036 29708
rect 19984 29665 19993 29699
rect 19993 29665 20027 29699
rect 20027 29665 20036 29699
rect 19984 29656 20036 29665
rect 20168 29656 20220 29708
rect 22284 29699 22336 29708
rect 22284 29665 22293 29699
rect 22293 29665 22327 29699
rect 22327 29665 22336 29699
rect 22284 29656 22336 29665
rect 22468 29656 22520 29708
rect 22744 29656 22796 29708
rect 23756 29724 23808 29776
rect 23388 29656 23440 29708
rect 19800 29631 19852 29640
rect 19800 29597 19809 29631
rect 19809 29597 19843 29631
rect 19843 29597 19852 29631
rect 19800 29588 19852 29597
rect 22008 29588 22060 29640
rect 23664 29588 23716 29640
rect 25320 29631 25372 29640
rect 25320 29597 25329 29631
rect 25329 29597 25363 29631
rect 25363 29597 25372 29631
rect 25320 29588 25372 29597
rect 3516 29520 3568 29572
rect 5816 29563 5868 29572
rect 5816 29529 5825 29563
rect 5825 29529 5859 29563
rect 5859 29529 5868 29563
rect 5816 29520 5868 29529
rect 8760 29563 8812 29572
rect 8760 29529 8769 29563
rect 8769 29529 8803 29563
rect 8803 29529 8812 29563
rect 8760 29520 8812 29529
rect 12348 29520 12400 29572
rect 12624 29520 12676 29572
rect 22100 29520 22152 29572
rect 10140 29452 10192 29504
rect 10324 29452 10376 29504
rect 10968 29452 11020 29504
rect 12164 29495 12216 29504
rect 12164 29461 12173 29495
rect 12173 29461 12207 29495
rect 12207 29461 12216 29495
rect 12164 29452 12216 29461
rect 12256 29495 12308 29504
rect 12256 29461 12265 29495
rect 12265 29461 12299 29495
rect 12299 29461 12308 29495
rect 12256 29452 12308 29461
rect 13084 29452 13136 29504
rect 13728 29495 13780 29504
rect 13728 29461 13737 29495
rect 13737 29461 13771 29495
rect 13771 29461 13780 29495
rect 13728 29452 13780 29461
rect 19432 29495 19484 29504
rect 19432 29461 19441 29495
rect 19441 29461 19475 29495
rect 19475 29461 19484 29495
rect 19432 29452 19484 29461
rect 20996 29452 21048 29504
rect 22744 29495 22796 29504
rect 22744 29461 22753 29495
rect 22753 29461 22787 29495
rect 22787 29461 22796 29495
rect 22744 29452 22796 29461
rect 23572 29495 23624 29504
rect 23572 29461 23581 29495
rect 23581 29461 23615 29495
rect 23615 29461 23624 29495
rect 23572 29452 23624 29461
rect 23940 29495 23992 29504
rect 23940 29461 23949 29495
rect 23949 29461 23983 29495
rect 23983 29461 23992 29495
rect 23940 29452 23992 29461
rect 7950 29350 8002 29402
rect 8014 29350 8066 29402
rect 8078 29350 8130 29402
rect 8142 29350 8194 29402
rect 8206 29350 8258 29402
rect 17950 29350 18002 29402
rect 18014 29350 18066 29402
rect 18078 29350 18130 29402
rect 18142 29350 18194 29402
rect 18206 29350 18258 29402
rect 8208 29291 8260 29300
rect 8208 29257 8217 29291
rect 8217 29257 8251 29291
rect 8251 29257 8260 29291
rect 8208 29248 8260 29257
rect 10876 29248 10928 29300
rect 12164 29248 12216 29300
rect 12900 29248 12952 29300
rect 13084 29291 13136 29300
rect 13084 29257 13093 29291
rect 13093 29257 13127 29291
rect 13127 29257 13136 29291
rect 13084 29248 13136 29257
rect 14648 29248 14700 29300
rect 18420 29248 18472 29300
rect 19800 29291 19852 29300
rect 9220 29180 9272 29232
rect 9588 29180 9640 29232
rect 10048 29180 10100 29232
rect 10324 29180 10376 29232
rect 13360 29223 13412 29232
rect 13360 29189 13369 29223
rect 13369 29189 13403 29223
rect 13403 29189 13412 29223
rect 13360 29180 13412 29189
rect 16212 29180 16264 29232
rect 19800 29257 19809 29291
rect 19809 29257 19843 29291
rect 19843 29257 19852 29291
rect 19800 29248 19852 29257
rect 25320 29248 25372 29300
rect 19340 29180 19392 29232
rect 9956 29087 10008 29096
rect 9956 29053 9965 29087
rect 9965 29053 9999 29087
rect 9999 29053 10008 29087
rect 9956 29044 10008 29053
rect 10048 29044 10100 29096
rect 16764 29112 16816 29164
rect 24676 29180 24728 29232
rect 24124 29155 24176 29164
rect 24124 29121 24133 29155
rect 24133 29121 24167 29155
rect 24167 29121 24176 29155
rect 24124 29112 24176 29121
rect 17500 29044 17552 29096
rect 18788 29044 18840 29096
rect 10416 28976 10468 29028
rect 12900 29019 12952 29028
rect 12900 28985 12909 29019
rect 12909 28985 12943 29019
rect 12943 28985 12952 29019
rect 12900 28976 12952 28985
rect 9864 28908 9916 28960
rect 12164 28908 12216 28960
rect 13360 28908 13412 28960
rect 15200 28976 15252 29028
rect 16764 29019 16816 29028
rect 16764 28985 16773 29019
rect 16773 28985 16807 29019
rect 16807 28985 16816 29019
rect 16764 28976 16816 28985
rect 17408 28976 17460 29028
rect 17776 28951 17828 28960
rect 17776 28917 17785 28951
rect 17785 28917 17819 28951
rect 17819 28917 17828 28951
rect 17776 28908 17828 28917
rect 18604 28908 18656 28960
rect 22192 29087 22244 29096
rect 22192 29053 22201 29087
rect 22201 29053 22235 29087
rect 22235 29053 22244 29087
rect 22192 29044 22244 29053
rect 24584 29019 24636 29028
rect 24584 28985 24593 29019
rect 24593 28985 24627 29019
rect 24627 28985 24636 29019
rect 24584 28976 24636 28985
rect 2950 28806 3002 28858
rect 3014 28806 3066 28858
rect 3078 28806 3130 28858
rect 3142 28806 3194 28858
rect 3206 28806 3258 28858
rect 12950 28806 13002 28858
rect 13014 28806 13066 28858
rect 13078 28806 13130 28858
rect 13142 28806 13194 28858
rect 13206 28806 13258 28858
rect 22950 28806 23002 28858
rect 23014 28806 23066 28858
rect 23078 28806 23130 28858
rect 23142 28806 23194 28858
rect 23206 28806 23258 28858
rect 4252 28704 4304 28756
rect 7380 28704 7432 28756
rect 1952 28568 2004 28620
rect 8024 28611 8076 28620
rect 8024 28577 8033 28611
rect 8033 28577 8067 28611
rect 8067 28577 8076 28611
rect 8024 28568 8076 28577
rect 4068 28364 4120 28416
rect 5724 28432 5776 28484
rect 7472 28432 7524 28484
rect 6920 28364 6972 28416
rect 7564 28364 7616 28416
rect 8208 28432 8260 28484
rect 9772 28704 9824 28756
rect 12624 28704 12676 28756
rect 14188 28704 14240 28756
rect 8576 28636 8628 28688
rect 9220 28636 9272 28688
rect 10784 28636 10836 28688
rect 16672 28704 16724 28756
rect 17592 28704 17644 28756
rect 21088 28704 21140 28756
rect 23572 28704 23624 28756
rect 25228 28704 25280 28756
rect 9956 28568 10008 28620
rect 10968 28568 11020 28620
rect 12808 28568 12860 28620
rect 13636 28568 13688 28620
rect 14280 28568 14332 28620
rect 17776 28568 17828 28620
rect 19524 28611 19576 28620
rect 19524 28577 19533 28611
rect 19533 28577 19567 28611
rect 19567 28577 19576 28611
rect 19524 28568 19576 28577
rect 19708 28636 19760 28688
rect 8944 28500 8996 28552
rect 9496 28500 9548 28552
rect 16580 28500 16632 28552
rect 17132 28500 17184 28552
rect 19248 28500 19300 28552
rect 20628 28500 20680 28552
rect 21180 28568 21232 28620
rect 22100 28568 22152 28620
rect 24676 28568 24728 28620
rect 12532 28432 12584 28484
rect 13820 28364 13872 28416
rect 20536 28432 20588 28484
rect 22192 28543 22244 28552
rect 22192 28509 22201 28543
rect 22201 28509 22235 28543
rect 22235 28509 22244 28543
rect 22192 28500 22244 28509
rect 17040 28407 17092 28416
rect 17040 28373 17049 28407
rect 17049 28373 17083 28407
rect 17083 28373 17092 28407
rect 17040 28364 17092 28373
rect 17500 28407 17552 28416
rect 17500 28373 17509 28407
rect 17509 28373 17543 28407
rect 17543 28373 17552 28407
rect 17500 28364 17552 28373
rect 18696 28407 18748 28416
rect 18696 28373 18705 28407
rect 18705 28373 18739 28407
rect 18739 28373 18748 28407
rect 18696 28364 18748 28373
rect 19984 28364 20036 28416
rect 20904 28407 20956 28416
rect 20904 28373 20913 28407
rect 20913 28373 20947 28407
rect 20947 28373 20956 28407
rect 20904 28364 20956 28373
rect 21364 28407 21416 28416
rect 21364 28373 21373 28407
rect 21373 28373 21407 28407
rect 21407 28373 21416 28407
rect 21364 28364 21416 28373
rect 25412 28500 25464 28552
rect 24860 28364 24912 28416
rect 7950 28262 8002 28314
rect 8014 28262 8066 28314
rect 8078 28262 8130 28314
rect 8142 28262 8194 28314
rect 8206 28262 8258 28314
rect 17950 28262 18002 28314
rect 18014 28262 18066 28314
rect 18078 28262 18130 28314
rect 18142 28262 18194 28314
rect 18206 28262 18258 28314
rect 6276 28024 6328 28076
rect 7840 28160 7892 28212
rect 8576 28203 8628 28212
rect 8576 28169 8585 28203
rect 8585 28169 8619 28203
rect 8619 28169 8628 28203
rect 8576 28160 8628 28169
rect 9864 28160 9916 28212
rect 10968 28067 11020 28076
rect 10968 28033 10977 28067
rect 10977 28033 11011 28067
rect 11011 28033 11020 28067
rect 10968 28024 11020 28033
rect 12532 28160 12584 28212
rect 16580 28160 16632 28212
rect 12624 28024 12676 28076
rect 16764 28092 16816 28144
rect 17316 28203 17368 28212
rect 17316 28169 17325 28203
rect 17325 28169 17359 28203
rect 17359 28169 17368 28203
rect 17316 28160 17368 28169
rect 17500 28160 17552 28212
rect 18604 28160 18656 28212
rect 20444 28160 20496 28212
rect 22652 28160 22704 28212
rect 17868 28092 17920 28144
rect 6920 27956 6972 28008
rect 7288 27956 7340 28008
rect 7840 27956 7892 28008
rect 10048 27956 10100 28008
rect 10600 27956 10652 28008
rect 12072 27956 12124 28008
rect 12348 27999 12400 28008
rect 12348 27965 12357 27999
rect 12357 27965 12391 27999
rect 12391 27965 12400 27999
rect 12348 27956 12400 27965
rect 12440 27999 12492 28008
rect 12440 27965 12449 27999
rect 12449 27965 12483 27999
rect 12483 27965 12492 27999
rect 12440 27956 12492 27965
rect 13360 27956 13412 28008
rect 14740 27999 14792 28008
rect 14740 27965 14749 27999
rect 14749 27965 14783 27999
rect 14783 27965 14792 27999
rect 14740 27956 14792 27965
rect 13452 27888 13504 27940
rect 10692 27820 10744 27872
rect 11980 27820 12032 27872
rect 14004 27820 14056 27872
rect 15936 28024 15988 28076
rect 18052 28024 18104 28076
rect 18604 28024 18656 28076
rect 20904 28092 20956 28144
rect 24400 28092 24452 28144
rect 25412 28203 25464 28212
rect 25412 28169 25421 28203
rect 25421 28169 25455 28203
rect 25455 28169 25464 28203
rect 25412 28160 25464 28169
rect 25504 28092 25556 28144
rect 20444 28067 20496 28076
rect 20444 28033 20453 28067
rect 20453 28033 20487 28067
rect 20487 28033 20496 28067
rect 20444 28024 20496 28033
rect 18788 27956 18840 28008
rect 15936 27888 15988 27940
rect 16488 27888 16540 27940
rect 21640 27888 21692 27940
rect 23940 28067 23992 28076
rect 23940 28033 23949 28067
rect 23949 28033 23983 28067
rect 23983 28033 23992 28067
rect 23940 28024 23992 28033
rect 24676 27956 24728 28008
rect 23940 27888 23992 27940
rect 24216 27888 24268 27940
rect 20076 27820 20128 27872
rect 20536 27820 20588 27872
rect 24124 27863 24176 27872
rect 24124 27829 24133 27863
rect 24133 27829 24167 27863
rect 24167 27829 24176 27863
rect 24124 27820 24176 27829
rect 2950 27718 3002 27770
rect 3014 27718 3066 27770
rect 3078 27718 3130 27770
rect 3142 27718 3194 27770
rect 3206 27718 3258 27770
rect 12950 27718 13002 27770
rect 13014 27718 13066 27770
rect 13078 27718 13130 27770
rect 13142 27718 13194 27770
rect 13206 27718 13258 27770
rect 22950 27718 23002 27770
rect 23014 27718 23066 27770
rect 23078 27718 23130 27770
rect 23142 27718 23194 27770
rect 23206 27718 23258 27770
rect 7656 27616 7708 27668
rect 1308 27480 1360 27532
rect 2688 27480 2740 27532
rect 5540 27480 5592 27532
rect 8024 27523 8076 27532
rect 8024 27489 8033 27523
rect 8033 27489 8067 27523
rect 8067 27489 8076 27523
rect 8024 27480 8076 27489
rect 8576 27548 8628 27600
rect 10048 27548 10100 27600
rect 10324 27548 10376 27600
rect 10968 27616 11020 27668
rect 11980 27616 12032 27668
rect 12348 27616 12400 27668
rect 19340 27616 19392 27668
rect 19524 27616 19576 27668
rect 14556 27480 14608 27532
rect 16028 27480 16080 27532
rect 16672 27548 16724 27600
rect 18972 27548 19024 27600
rect 20720 27616 20772 27668
rect 21088 27616 21140 27668
rect 23940 27548 23992 27600
rect 1952 27412 2004 27464
rect 13360 27412 13412 27464
rect 14924 27412 14976 27464
rect 3976 27344 4028 27396
rect 7472 27344 7524 27396
rect 6920 27276 6972 27328
rect 7840 27344 7892 27396
rect 8576 27276 8628 27328
rect 10600 27276 10652 27328
rect 11520 27276 11572 27328
rect 12440 27276 12492 27328
rect 17040 27412 17092 27464
rect 19248 27480 19300 27532
rect 23572 27480 23624 27532
rect 18052 27412 18104 27464
rect 18328 27412 18380 27464
rect 19800 27412 19852 27464
rect 21456 27412 21508 27464
rect 22284 27455 22336 27464
rect 22284 27421 22293 27455
rect 22293 27421 22327 27455
rect 22327 27421 22336 27455
rect 22284 27412 22336 27421
rect 24308 27412 24360 27464
rect 14280 27319 14332 27328
rect 14280 27285 14289 27319
rect 14289 27285 14323 27319
rect 14323 27285 14332 27319
rect 14280 27276 14332 27285
rect 14464 27276 14516 27328
rect 14832 27276 14884 27328
rect 15476 27276 15528 27328
rect 15568 27319 15620 27328
rect 15568 27285 15577 27319
rect 15577 27285 15611 27319
rect 15611 27285 15620 27319
rect 15568 27276 15620 27285
rect 15936 27319 15988 27328
rect 15936 27285 15945 27319
rect 15945 27285 15979 27319
rect 15979 27285 15988 27319
rect 15936 27276 15988 27285
rect 16488 27276 16540 27328
rect 16764 27319 16816 27328
rect 16764 27285 16773 27319
rect 16773 27285 16807 27319
rect 16807 27285 16816 27319
rect 16764 27276 16816 27285
rect 17224 27319 17276 27328
rect 17224 27285 17233 27319
rect 17233 27285 17267 27319
rect 17267 27285 17276 27319
rect 17224 27276 17276 27285
rect 18420 27276 18472 27328
rect 18696 27319 18748 27328
rect 18696 27285 18705 27319
rect 18705 27285 18739 27319
rect 18739 27285 18748 27319
rect 18696 27276 18748 27285
rect 20076 27276 20128 27328
rect 22836 27344 22888 27396
rect 23296 27276 23348 27328
rect 23572 27276 23624 27328
rect 23940 27344 23992 27396
rect 24400 27276 24452 27328
rect 7950 27174 8002 27226
rect 8014 27174 8066 27226
rect 8078 27174 8130 27226
rect 8142 27174 8194 27226
rect 8206 27174 8258 27226
rect 17950 27174 18002 27226
rect 18014 27174 18066 27226
rect 18078 27174 18130 27226
rect 18142 27174 18194 27226
rect 18206 27174 18258 27226
rect 1768 27072 1820 27124
rect 3516 27072 3568 27124
rect 10876 27072 10928 27124
rect 6000 27004 6052 27056
rect 11520 27004 11572 27056
rect 2228 26979 2280 26988
rect 2228 26945 2237 26979
rect 2237 26945 2271 26979
rect 2271 26945 2280 26979
rect 2228 26936 2280 26945
rect 3332 26979 3384 26988
rect 3332 26945 3376 26979
rect 3376 26945 3384 26979
rect 3332 26936 3384 26945
rect 7196 26936 7248 26988
rect 8668 26936 8720 26988
rect 8852 26936 8904 26988
rect 7748 26911 7800 26920
rect 7748 26877 7757 26911
rect 7757 26877 7791 26911
rect 7791 26877 7800 26911
rect 7748 26868 7800 26877
rect 8300 26868 8352 26920
rect 7288 26800 7340 26852
rect 10508 26868 10560 26920
rect 15384 27072 15436 27124
rect 15752 27115 15804 27124
rect 15752 27081 15761 27115
rect 15761 27081 15795 27115
rect 15795 27081 15804 27115
rect 15752 27072 15804 27081
rect 16304 27072 16356 27124
rect 12532 27004 12584 27056
rect 13820 27047 13872 27056
rect 13820 27013 13829 27047
rect 13829 27013 13863 27047
rect 13863 27013 13872 27047
rect 13820 27004 13872 27013
rect 14924 27004 14976 27056
rect 18420 27115 18472 27124
rect 18420 27081 18429 27115
rect 18429 27081 18463 27115
rect 18463 27081 18472 27115
rect 18420 27072 18472 27081
rect 18604 27072 18656 27124
rect 19248 27072 19300 27124
rect 22284 27072 22336 27124
rect 20352 27004 20404 27056
rect 23572 27004 23624 27056
rect 13452 26979 13504 26988
rect 13452 26945 13461 26979
rect 13461 26945 13495 26979
rect 13495 26945 13504 26979
rect 13452 26936 13504 26945
rect 11980 26868 12032 26920
rect 12532 26868 12584 26920
rect 12808 26868 12860 26920
rect 13636 26800 13688 26852
rect 7196 26775 7248 26784
rect 7196 26741 7205 26775
rect 7205 26741 7239 26775
rect 7239 26741 7248 26775
rect 7196 26732 7248 26741
rect 10324 26732 10376 26784
rect 11520 26732 11572 26784
rect 14648 26775 14700 26784
rect 14648 26741 14657 26775
rect 14657 26741 14691 26775
rect 14691 26741 14700 26775
rect 14648 26732 14700 26741
rect 15936 26936 15988 26988
rect 16396 26979 16448 26988
rect 16396 26945 16405 26979
rect 16405 26945 16439 26979
rect 16439 26945 16448 26979
rect 16396 26936 16448 26945
rect 17316 26936 17368 26988
rect 18604 26936 18656 26988
rect 25412 27115 25464 27124
rect 25412 27081 25421 27115
rect 25421 27081 25455 27115
rect 25455 27081 25464 27115
rect 25412 27072 25464 27081
rect 24768 27047 24820 27056
rect 24768 27013 24777 27047
rect 24777 27013 24811 27047
rect 24811 27013 24820 27047
rect 24768 27004 24820 27013
rect 15476 26800 15528 26852
rect 17408 26800 17460 26852
rect 18788 26868 18840 26920
rect 24860 26868 24912 26920
rect 19892 26800 19944 26852
rect 24308 26800 24360 26852
rect 16304 26732 16356 26784
rect 16488 26732 16540 26784
rect 18328 26732 18380 26784
rect 24400 26732 24452 26784
rect 2950 26630 3002 26682
rect 3014 26630 3066 26682
rect 3078 26630 3130 26682
rect 3142 26630 3194 26682
rect 3206 26630 3258 26682
rect 12950 26630 13002 26682
rect 13014 26630 13066 26682
rect 13078 26630 13130 26682
rect 13142 26630 13194 26682
rect 13206 26630 13258 26682
rect 22950 26630 23002 26682
rect 23014 26630 23066 26682
rect 23078 26630 23130 26682
rect 23142 26630 23194 26682
rect 23206 26630 23258 26682
rect 7656 26528 7708 26580
rect 2596 26392 2648 26444
rect 6000 26392 6052 26444
rect 6276 26435 6328 26444
rect 6276 26401 6285 26435
rect 6285 26401 6319 26435
rect 6319 26401 6328 26435
rect 6276 26392 6328 26401
rect 6920 26392 6972 26444
rect 7840 26392 7892 26444
rect 8576 26528 8628 26580
rect 11980 26528 12032 26580
rect 13912 26528 13964 26580
rect 15016 26528 15068 26580
rect 15936 26528 15988 26580
rect 16028 26528 16080 26580
rect 16212 26528 16264 26580
rect 16488 26528 16540 26580
rect 10508 26392 10560 26444
rect 12624 26392 12676 26444
rect 8392 26324 8444 26376
rect 9036 26324 9088 26376
rect 3884 26256 3936 26308
rect 8576 26256 8628 26308
rect 9680 26367 9732 26376
rect 9680 26333 9689 26367
rect 9689 26333 9723 26367
rect 9723 26333 9732 26367
rect 9680 26324 9732 26333
rect 10600 26367 10652 26376
rect 10600 26333 10609 26367
rect 10609 26333 10643 26367
rect 10643 26333 10652 26367
rect 10600 26324 10652 26333
rect 13728 26460 13780 26512
rect 19524 26460 19576 26512
rect 22836 26528 22888 26580
rect 23296 26528 23348 26580
rect 20812 26460 20864 26512
rect 13544 26324 13596 26376
rect 14556 26367 14608 26376
rect 14556 26333 14565 26367
rect 14565 26333 14599 26367
rect 14599 26333 14608 26367
rect 14556 26324 14608 26333
rect 15936 26324 15988 26376
rect 16672 26324 16724 26376
rect 17592 26435 17644 26444
rect 17592 26401 17601 26435
rect 17601 26401 17635 26435
rect 17635 26401 17644 26435
rect 17592 26392 17644 26401
rect 18604 26392 18656 26444
rect 20076 26392 20128 26444
rect 24400 26460 24452 26512
rect 24676 26460 24728 26512
rect 21456 26367 21508 26376
rect 21456 26333 21465 26367
rect 21465 26333 21499 26367
rect 21499 26333 21508 26367
rect 21456 26324 21508 26333
rect 25412 26392 25464 26444
rect 24492 26324 24544 26376
rect 10048 26256 10100 26308
rect 14464 26256 14516 26308
rect 17040 26256 17092 26308
rect 17132 26299 17184 26308
rect 17132 26265 17141 26299
rect 17141 26265 17175 26299
rect 17175 26265 17184 26299
rect 17132 26256 17184 26265
rect 16304 26188 16356 26240
rect 19708 26256 19760 26308
rect 21732 26299 21784 26308
rect 21732 26265 21741 26299
rect 21741 26265 21775 26299
rect 21775 26265 21784 26299
rect 21732 26256 21784 26265
rect 23112 26256 23164 26308
rect 23572 26256 23624 26308
rect 25228 26256 25280 26308
rect 7950 26086 8002 26138
rect 8014 26086 8066 26138
rect 8078 26086 8130 26138
rect 8142 26086 8194 26138
rect 8206 26086 8258 26138
rect 17950 26086 18002 26138
rect 18014 26086 18066 26138
rect 18078 26086 18130 26138
rect 18142 26086 18194 26138
rect 18206 26086 18258 26138
rect 2228 25984 2280 26036
rect 4068 25984 4120 26036
rect 8300 25984 8352 26036
rect 8668 26027 8720 26036
rect 8668 25993 8677 26027
rect 8677 25993 8711 26027
rect 8711 25993 8720 26027
rect 8668 25984 8720 25993
rect 10324 26027 10376 26036
rect 10324 25993 10333 26027
rect 10333 25993 10367 26027
rect 10367 25993 10376 26027
rect 10324 25984 10376 25993
rect 13912 26027 13964 26036
rect 13912 25993 13921 26027
rect 13921 25993 13955 26027
rect 13955 25993 13964 26027
rect 13912 25984 13964 25993
rect 18696 25984 18748 26036
rect 23388 25984 23440 26036
rect 10416 25916 10468 25968
rect 11980 25916 12032 25968
rect 13268 25916 13320 25968
rect 16672 25916 16724 25968
rect 19616 25959 19668 25968
rect 19616 25925 19625 25959
rect 19625 25925 19659 25959
rect 19659 25925 19668 25959
rect 19616 25916 19668 25925
rect 22468 25959 22520 25968
rect 22468 25925 22477 25959
rect 22477 25925 22511 25959
rect 22511 25925 22520 25959
rect 22468 25916 22520 25925
rect 22652 25916 22704 25968
rect 23112 25959 23164 25968
rect 23112 25925 23121 25959
rect 23121 25925 23155 25959
rect 23155 25925 23164 25959
rect 23112 25916 23164 25925
rect 23572 25959 23624 25968
rect 23572 25925 23581 25959
rect 23581 25925 23615 25959
rect 23615 25925 23624 25959
rect 23572 25916 23624 25925
rect 24032 25916 24084 25968
rect 25044 25959 25096 25968
rect 25044 25925 25053 25959
rect 25053 25925 25087 25959
rect 25087 25925 25096 25959
rect 25044 25916 25096 25925
rect 2872 25848 2924 25900
rect 13544 25891 13596 25900
rect 13544 25857 13553 25891
rect 13553 25857 13587 25891
rect 13587 25857 13596 25891
rect 13544 25848 13596 25857
rect 13912 25848 13964 25900
rect 14188 25848 14240 25900
rect 22284 25848 22336 25900
rect 4252 25780 4304 25832
rect 7564 25823 7616 25832
rect 7564 25789 7573 25823
rect 7573 25789 7607 25823
rect 7607 25789 7616 25823
rect 7564 25780 7616 25789
rect 3332 25712 3384 25764
rect 7840 25780 7892 25832
rect 12624 25780 12676 25832
rect 13636 25780 13688 25832
rect 16948 25823 17000 25832
rect 16948 25789 16957 25823
rect 16957 25789 16991 25823
rect 16991 25789 17000 25823
rect 16948 25780 17000 25789
rect 17224 25823 17276 25832
rect 17224 25789 17233 25823
rect 17233 25789 17267 25823
rect 17267 25789 17276 25823
rect 17224 25780 17276 25789
rect 18604 25780 18656 25832
rect 20168 25780 20220 25832
rect 20444 25823 20496 25832
rect 20444 25789 20453 25823
rect 20453 25789 20487 25823
rect 20487 25789 20496 25823
rect 20444 25780 20496 25789
rect 22560 25823 22612 25832
rect 22560 25789 22569 25823
rect 22569 25789 22603 25823
rect 22603 25789 22612 25823
rect 22560 25780 22612 25789
rect 4712 25644 4764 25696
rect 7012 25644 7064 25696
rect 8852 25712 8904 25764
rect 18512 25712 18564 25764
rect 22284 25712 22336 25764
rect 23296 25712 23348 25764
rect 24768 25712 24820 25764
rect 11704 25644 11756 25696
rect 12808 25644 12860 25696
rect 13452 25644 13504 25696
rect 16120 25687 16172 25696
rect 16120 25653 16129 25687
rect 16129 25653 16163 25687
rect 16163 25653 16172 25687
rect 16120 25644 16172 25653
rect 16304 25644 16356 25696
rect 18788 25644 18840 25696
rect 21548 25644 21600 25696
rect 2950 25542 3002 25594
rect 3014 25542 3066 25594
rect 3078 25542 3130 25594
rect 3142 25542 3194 25594
rect 3206 25542 3258 25594
rect 12950 25542 13002 25594
rect 13014 25542 13066 25594
rect 13078 25542 13130 25594
rect 13142 25542 13194 25594
rect 13206 25542 13258 25594
rect 22950 25542 23002 25594
rect 23014 25542 23066 25594
rect 23078 25542 23130 25594
rect 23142 25542 23194 25594
rect 23206 25542 23258 25594
rect 3608 25483 3660 25492
rect 3608 25449 3617 25483
rect 3617 25449 3651 25483
rect 3651 25449 3660 25483
rect 3608 25440 3660 25449
rect 4160 25483 4212 25492
rect 4160 25449 4169 25483
rect 4169 25449 4203 25483
rect 4203 25449 4212 25483
rect 4160 25440 4212 25449
rect 16120 25440 16172 25492
rect 16672 25440 16724 25492
rect 8392 25415 8444 25424
rect 8392 25381 8401 25415
rect 8401 25381 8435 25415
rect 8435 25381 8444 25415
rect 8392 25372 8444 25381
rect 13820 25372 13872 25424
rect 20904 25440 20956 25492
rect 1308 25304 1360 25356
rect 3332 25304 3384 25356
rect 5724 25304 5776 25356
rect 6000 25304 6052 25356
rect 6276 25304 6328 25356
rect 7656 25304 7708 25356
rect 1768 25279 1820 25288
rect 1768 25245 1777 25279
rect 1777 25245 1811 25279
rect 1811 25245 1820 25279
rect 1768 25236 1820 25245
rect 3608 25236 3660 25288
rect 4344 25236 4396 25288
rect 15568 25347 15620 25356
rect 15568 25313 15577 25347
rect 15577 25313 15611 25347
rect 15611 25313 15620 25347
rect 15568 25304 15620 25313
rect 15660 25347 15712 25356
rect 15660 25313 15669 25347
rect 15669 25313 15703 25347
rect 15703 25313 15712 25347
rect 15660 25304 15712 25313
rect 16580 25304 16632 25356
rect 17040 25304 17092 25356
rect 17500 25304 17552 25356
rect 17684 25236 17736 25288
rect 21456 25304 21508 25356
rect 22008 25304 22060 25356
rect 23480 25440 23532 25492
rect 23848 25440 23900 25492
rect 25044 25372 25096 25424
rect 22836 25304 22888 25356
rect 23388 25236 23440 25288
rect 16120 25168 16172 25220
rect 19340 25168 19392 25220
rect 22652 25168 22704 25220
rect 24124 25236 24176 25288
rect 7932 25100 7984 25152
rect 9128 25143 9180 25152
rect 9128 25109 9137 25143
rect 9137 25109 9171 25143
rect 9171 25109 9180 25143
rect 9128 25100 9180 25109
rect 12532 25100 12584 25152
rect 15108 25143 15160 25152
rect 15108 25109 15117 25143
rect 15117 25109 15151 25143
rect 15151 25109 15160 25143
rect 15108 25100 15160 25109
rect 16304 25143 16356 25152
rect 16304 25109 16313 25143
rect 16313 25109 16347 25143
rect 16347 25109 16356 25143
rect 16304 25100 16356 25109
rect 21088 25100 21140 25152
rect 21732 25100 21784 25152
rect 24124 25100 24176 25152
rect 7950 24998 8002 25050
rect 8014 24998 8066 25050
rect 8078 24998 8130 25050
rect 8142 24998 8194 25050
rect 8206 24998 8258 25050
rect 17950 24998 18002 25050
rect 18014 24998 18066 25050
rect 18078 24998 18130 25050
rect 18142 24998 18194 25050
rect 18206 24998 18258 25050
rect 8392 24896 8444 24948
rect 4068 24828 4120 24880
rect 2228 24803 2280 24812
rect 2228 24769 2237 24803
rect 2237 24769 2271 24803
rect 2271 24769 2280 24803
rect 2228 24760 2280 24769
rect 6276 24760 6328 24812
rect 12532 24939 12584 24948
rect 12532 24905 12541 24939
rect 12541 24905 12575 24939
rect 12575 24905 12584 24939
rect 12532 24896 12584 24905
rect 15016 24896 15068 24948
rect 19432 24896 19484 24948
rect 20444 24896 20496 24948
rect 22744 24896 22796 24948
rect 9588 24760 9640 24812
rect 10692 24803 10744 24812
rect 10692 24769 10701 24803
rect 10701 24769 10735 24803
rect 10735 24769 10744 24803
rect 10692 24760 10744 24769
rect 10784 24803 10836 24812
rect 10784 24769 10793 24803
rect 10793 24769 10827 24803
rect 10827 24769 10836 24803
rect 10784 24760 10836 24769
rect 11428 24760 11480 24812
rect 11888 24803 11940 24812
rect 11888 24769 11897 24803
rect 11897 24769 11931 24803
rect 11931 24769 11940 24803
rect 14556 24828 14608 24880
rect 11888 24760 11940 24769
rect 4160 24692 4212 24744
rect 5724 24692 5776 24744
rect 7472 24735 7524 24744
rect 7472 24701 7481 24735
rect 7481 24701 7515 24735
rect 7515 24701 7524 24735
rect 7472 24692 7524 24701
rect 7840 24692 7892 24744
rect 12624 24760 12676 24812
rect 1952 24624 2004 24676
rect 9772 24624 9824 24676
rect 10968 24624 11020 24676
rect 14188 24692 14240 24744
rect 16120 24760 16172 24812
rect 16672 24803 16724 24812
rect 16672 24769 16681 24803
rect 16681 24769 16715 24803
rect 16715 24769 16724 24803
rect 16672 24760 16724 24769
rect 18420 24803 18472 24812
rect 18420 24769 18429 24803
rect 18429 24769 18463 24803
rect 18463 24769 18472 24803
rect 18420 24760 18472 24769
rect 19524 24803 19576 24812
rect 19524 24769 19533 24803
rect 19533 24769 19567 24803
rect 19567 24769 19576 24803
rect 19524 24760 19576 24769
rect 21364 24760 21416 24812
rect 24584 24760 24636 24812
rect 13820 24624 13872 24676
rect 5632 24556 5684 24608
rect 13636 24556 13688 24608
rect 16212 24692 16264 24744
rect 16580 24692 16632 24744
rect 17224 24692 17276 24744
rect 18604 24735 18656 24744
rect 18604 24701 18613 24735
rect 18613 24701 18647 24735
rect 18647 24701 18656 24735
rect 18604 24692 18656 24701
rect 19340 24735 19392 24744
rect 19340 24701 19349 24735
rect 19349 24701 19383 24735
rect 19383 24701 19392 24735
rect 19340 24692 19392 24701
rect 22100 24735 22152 24744
rect 22100 24701 22109 24735
rect 22109 24701 22143 24735
rect 22143 24701 22152 24735
rect 22100 24692 22152 24701
rect 16948 24624 17000 24676
rect 22192 24624 22244 24676
rect 22836 24624 22888 24676
rect 23480 24735 23532 24744
rect 23480 24701 23489 24735
rect 23489 24701 23523 24735
rect 23523 24701 23532 24735
rect 23480 24692 23532 24701
rect 24860 24692 24912 24744
rect 25412 24692 25464 24744
rect 16672 24556 16724 24608
rect 17592 24556 17644 24608
rect 18328 24556 18380 24608
rect 19892 24556 19944 24608
rect 22744 24599 22796 24608
rect 22744 24565 22753 24599
rect 22753 24565 22787 24599
rect 22787 24565 22796 24599
rect 22744 24556 22796 24565
rect 2950 24454 3002 24506
rect 3014 24454 3066 24506
rect 3078 24454 3130 24506
rect 3142 24454 3194 24506
rect 3206 24454 3258 24506
rect 12950 24454 13002 24506
rect 13014 24454 13066 24506
rect 13078 24454 13130 24506
rect 13142 24454 13194 24506
rect 13206 24454 13258 24506
rect 22950 24454 23002 24506
rect 23014 24454 23066 24506
rect 23078 24454 23130 24506
rect 23142 24454 23194 24506
rect 23206 24454 23258 24506
rect 2872 24395 2924 24404
rect 2872 24361 2881 24395
rect 2881 24361 2915 24395
rect 2915 24361 2924 24395
rect 2872 24352 2924 24361
rect 3148 24395 3200 24404
rect 3148 24361 3157 24395
rect 3157 24361 3191 24395
rect 3191 24361 3200 24395
rect 3148 24352 3200 24361
rect 4068 24352 4120 24404
rect 5632 24352 5684 24404
rect 7380 24352 7432 24404
rect 7564 24352 7616 24404
rect 7656 24216 7708 24268
rect 10784 24352 10836 24404
rect 10968 24352 11020 24404
rect 11336 24352 11388 24404
rect 12440 24352 12492 24404
rect 10968 24216 11020 24268
rect 17500 24352 17552 24404
rect 24400 24352 24452 24404
rect 24584 24352 24636 24404
rect 17224 24284 17276 24336
rect 13452 24216 13504 24268
rect 14648 24216 14700 24268
rect 3608 24148 3660 24200
rect 4068 24191 4120 24200
rect 4068 24157 4086 24191
rect 4086 24157 4120 24191
rect 4068 24148 4120 24157
rect 7472 24148 7524 24200
rect 10876 24191 10928 24200
rect 10876 24157 10885 24191
rect 10885 24157 10919 24191
rect 10919 24157 10928 24191
rect 10876 24148 10928 24157
rect 13636 24148 13688 24200
rect 16304 24216 16356 24268
rect 18972 24284 19024 24336
rect 18512 24216 18564 24268
rect 19984 24259 20036 24268
rect 19984 24225 19993 24259
rect 19993 24225 20027 24259
rect 20027 24225 20036 24259
rect 19984 24216 20036 24225
rect 21088 24216 21140 24268
rect 21180 24216 21232 24268
rect 21456 24216 21508 24268
rect 24860 24216 24912 24268
rect 16212 24148 16264 24200
rect 19892 24191 19944 24200
rect 19892 24157 19901 24191
rect 19901 24157 19935 24191
rect 19935 24157 19944 24191
rect 19892 24148 19944 24157
rect 4528 24080 4580 24132
rect 9036 24080 9088 24132
rect 9588 24080 9640 24132
rect 11336 24080 11388 24132
rect 12440 24080 12492 24132
rect 3976 24012 4028 24064
rect 9864 24012 9916 24064
rect 11612 24012 11664 24064
rect 13544 24012 13596 24064
rect 18880 24080 18932 24132
rect 13820 24012 13872 24064
rect 15936 24012 15988 24064
rect 17132 24012 17184 24064
rect 18512 24055 18564 24064
rect 18512 24021 18521 24055
rect 18521 24021 18555 24055
rect 18555 24021 18564 24055
rect 18512 24012 18564 24021
rect 18788 24012 18840 24064
rect 20720 24055 20772 24064
rect 20720 24021 20729 24055
rect 20729 24021 20763 24055
rect 20763 24021 20772 24055
rect 20720 24012 20772 24021
rect 21088 24055 21140 24064
rect 21088 24021 21097 24055
rect 21097 24021 21131 24055
rect 21131 24021 21140 24055
rect 21088 24012 21140 24021
rect 21272 24080 21324 24132
rect 24492 24148 24544 24200
rect 24492 24012 24544 24064
rect 24676 24055 24728 24064
rect 24676 24021 24685 24055
rect 24685 24021 24719 24055
rect 24719 24021 24728 24055
rect 24676 24012 24728 24021
rect 7950 23910 8002 23962
rect 8014 23910 8066 23962
rect 8078 23910 8130 23962
rect 8142 23910 8194 23962
rect 8206 23910 8258 23962
rect 17950 23910 18002 23962
rect 18014 23910 18066 23962
rect 18078 23910 18130 23962
rect 18142 23910 18194 23962
rect 18206 23910 18258 23962
rect 4160 23740 4212 23792
rect 5632 23808 5684 23860
rect 6736 23808 6788 23860
rect 9128 23808 9180 23860
rect 9404 23808 9456 23860
rect 13544 23851 13596 23860
rect 13544 23817 13553 23851
rect 13553 23817 13587 23851
rect 13587 23817 13596 23851
rect 13544 23808 13596 23817
rect 15936 23851 15988 23860
rect 15936 23817 15945 23851
rect 15945 23817 15979 23851
rect 15979 23817 15988 23851
rect 15936 23808 15988 23817
rect 16856 23808 16908 23860
rect 17868 23808 17920 23860
rect 21088 23808 21140 23860
rect 5448 23740 5500 23792
rect 9036 23740 9088 23792
rect 11980 23740 12032 23792
rect 14004 23740 14056 23792
rect 25136 23783 25188 23792
rect 25136 23749 25145 23783
rect 25145 23749 25179 23783
rect 25179 23749 25188 23783
rect 25136 23740 25188 23749
rect 6276 23672 6328 23724
rect 7288 23672 7340 23724
rect 5356 23604 5408 23656
rect 5632 23604 5684 23656
rect 6644 23604 6696 23656
rect 6736 23536 6788 23588
rect 7012 23536 7064 23588
rect 9772 23647 9824 23656
rect 9772 23613 9781 23647
rect 9781 23613 9815 23647
rect 9815 23613 9824 23647
rect 9772 23604 9824 23613
rect 13728 23672 13780 23724
rect 23940 23672 23992 23724
rect 24124 23715 24176 23724
rect 24124 23681 24133 23715
rect 24133 23681 24167 23715
rect 24167 23681 24176 23715
rect 24124 23672 24176 23681
rect 11336 23604 11388 23656
rect 9864 23536 9916 23588
rect 13636 23604 13688 23656
rect 16028 23604 16080 23656
rect 16580 23604 16632 23656
rect 23388 23604 23440 23656
rect 3148 23468 3200 23520
rect 4160 23468 4212 23520
rect 5724 23468 5776 23520
rect 6552 23468 6604 23520
rect 9588 23468 9640 23520
rect 10692 23468 10744 23520
rect 14832 23468 14884 23520
rect 15752 23468 15804 23520
rect 20444 23468 20496 23520
rect 2950 23366 3002 23418
rect 3014 23366 3066 23418
rect 3078 23366 3130 23418
rect 3142 23366 3194 23418
rect 3206 23366 3258 23418
rect 12950 23366 13002 23418
rect 13014 23366 13066 23418
rect 13078 23366 13130 23418
rect 13142 23366 13194 23418
rect 13206 23366 13258 23418
rect 22950 23366 23002 23418
rect 23014 23366 23066 23418
rect 23078 23366 23130 23418
rect 23142 23366 23194 23418
rect 23206 23366 23258 23418
rect 4252 23264 4304 23316
rect 9036 23307 9088 23316
rect 9036 23273 9045 23307
rect 9045 23273 9079 23307
rect 9079 23273 9088 23307
rect 9036 23264 9088 23273
rect 8300 23196 8352 23248
rect 9404 23264 9456 23316
rect 13176 23264 13228 23316
rect 13728 23307 13780 23316
rect 13728 23273 13737 23307
rect 13737 23273 13771 23307
rect 13771 23273 13780 23307
rect 13728 23264 13780 23273
rect 18604 23264 18656 23316
rect 18880 23307 18932 23316
rect 18880 23273 18889 23307
rect 18889 23273 18923 23307
rect 18923 23273 18932 23307
rect 18880 23264 18932 23273
rect 20168 23307 20220 23316
rect 20168 23273 20177 23307
rect 20177 23273 20211 23307
rect 20211 23273 20220 23307
rect 20168 23264 20220 23273
rect 9312 23196 9364 23248
rect 12072 23196 12124 23248
rect 17132 23196 17184 23248
rect 2780 23103 2832 23112
rect 2780 23069 2789 23103
rect 2789 23069 2823 23103
rect 2823 23069 2832 23103
rect 2780 23060 2832 23069
rect 6368 23128 6420 23180
rect 7012 23171 7064 23180
rect 7012 23137 7021 23171
rect 7021 23137 7055 23171
rect 7055 23137 7064 23171
rect 7012 23128 7064 23137
rect 7288 23171 7340 23180
rect 7288 23137 7297 23171
rect 7297 23137 7331 23171
rect 7331 23137 7340 23171
rect 7288 23128 7340 23137
rect 940 22992 992 23044
rect 6736 22992 6788 23044
rect 7104 22992 7156 23044
rect 9128 23128 9180 23180
rect 9588 23128 9640 23180
rect 9772 23128 9824 23180
rect 10232 23171 10284 23180
rect 10232 23137 10241 23171
rect 10241 23137 10275 23171
rect 10275 23137 10284 23171
rect 10232 23128 10284 23137
rect 8668 23060 8720 23112
rect 12624 23128 12676 23180
rect 13636 23128 13688 23180
rect 15292 23128 15344 23180
rect 17040 23128 17092 23180
rect 17408 23171 17460 23180
rect 17408 23137 17417 23171
rect 17417 23137 17451 23171
rect 17451 23137 17460 23171
rect 17408 23128 17460 23137
rect 18972 23128 19024 23180
rect 21272 23128 21324 23180
rect 12992 23060 13044 23112
rect 16948 23060 17000 23112
rect 21916 23103 21968 23112
rect 21916 23069 21925 23103
rect 21925 23069 21959 23103
rect 21959 23069 21968 23103
rect 21916 23060 21968 23069
rect 12532 22992 12584 23044
rect 22376 23264 22428 23316
rect 24400 23264 24452 23316
rect 24860 23128 24912 23180
rect 25412 23128 25464 23180
rect 24308 23060 24360 23112
rect 25044 23060 25096 23112
rect 5632 22924 5684 22976
rect 6828 22924 6880 22976
rect 8392 22967 8444 22976
rect 8392 22933 8401 22967
rect 8401 22933 8435 22967
rect 8435 22933 8444 22967
rect 8392 22924 8444 22933
rect 9588 22967 9640 22976
rect 9588 22933 9597 22967
rect 9597 22933 9631 22967
rect 9631 22933 9640 22967
rect 9588 22924 9640 22933
rect 11060 22924 11112 22976
rect 12440 22924 12492 22976
rect 13176 22924 13228 22976
rect 13728 22924 13780 22976
rect 15384 22924 15436 22976
rect 24584 22967 24636 22976
rect 24584 22933 24593 22967
rect 24593 22933 24627 22967
rect 24627 22933 24636 22967
rect 24584 22924 24636 22933
rect 25504 22924 25556 22976
rect 7950 22822 8002 22874
rect 8014 22822 8066 22874
rect 8078 22822 8130 22874
rect 8142 22822 8194 22874
rect 8206 22822 8258 22874
rect 17950 22822 18002 22874
rect 18014 22822 18066 22874
rect 18078 22822 18130 22874
rect 18142 22822 18194 22874
rect 18206 22822 18258 22874
rect 1768 22720 1820 22772
rect 2228 22720 2280 22772
rect 3884 22720 3936 22772
rect 7288 22652 7340 22704
rect 8392 22720 8444 22772
rect 10508 22720 10560 22772
rect 11060 22720 11112 22772
rect 12256 22720 12308 22772
rect 12992 22720 13044 22772
rect 13452 22720 13504 22772
rect 9128 22652 9180 22704
rect 9864 22652 9916 22704
rect 10692 22652 10744 22704
rect 12532 22695 12584 22704
rect 12532 22661 12541 22695
rect 12541 22661 12575 22695
rect 12575 22661 12584 22695
rect 12532 22652 12584 22661
rect 13544 22652 13596 22704
rect 14556 22720 14608 22772
rect 15660 22720 15712 22772
rect 21088 22720 21140 22772
rect 21456 22720 21508 22772
rect 22192 22720 22244 22772
rect 13728 22652 13780 22704
rect 16120 22695 16172 22704
rect 16120 22661 16129 22695
rect 16129 22661 16163 22695
rect 16163 22661 16172 22695
rect 16120 22652 16172 22661
rect 17868 22652 17920 22704
rect 2136 22627 2188 22636
rect 2136 22593 2145 22627
rect 2145 22593 2179 22627
rect 2179 22593 2188 22627
rect 2136 22584 2188 22593
rect 2872 22584 2924 22636
rect 3332 22584 3384 22636
rect 3884 22627 3936 22636
rect 3884 22593 3928 22627
rect 3928 22593 3936 22627
rect 3884 22584 3936 22593
rect 5540 22627 5592 22636
rect 5540 22593 5549 22627
rect 5549 22593 5583 22627
rect 5583 22593 5592 22627
rect 5540 22584 5592 22593
rect 7748 22584 7800 22636
rect 10876 22584 10928 22636
rect 11244 22584 11296 22636
rect 13360 22627 13412 22636
rect 13360 22593 13369 22627
rect 13369 22593 13403 22627
rect 13403 22593 13412 22627
rect 13360 22584 13412 22593
rect 21640 22652 21692 22704
rect 24492 22720 24544 22772
rect 4896 22516 4948 22568
rect 5724 22559 5776 22568
rect 5724 22525 5733 22559
rect 5733 22525 5767 22559
rect 5767 22525 5776 22559
rect 5724 22516 5776 22525
rect 8668 22559 8720 22568
rect 8668 22525 8677 22559
rect 8677 22525 8711 22559
rect 8711 22525 8720 22559
rect 8668 22516 8720 22525
rect 12624 22516 12676 22568
rect 13176 22516 13228 22568
rect 22376 22584 22428 22636
rect 22836 22584 22888 22636
rect 24492 22584 24544 22636
rect 25320 22627 25372 22636
rect 25320 22593 25329 22627
rect 25329 22593 25363 22627
rect 25363 22593 25372 22627
rect 25320 22584 25372 22593
rect 11520 22448 11572 22500
rect 4160 22380 4212 22432
rect 17500 22516 17552 22568
rect 20812 22559 20864 22568
rect 20812 22525 20821 22559
rect 20821 22525 20855 22559
rect 20855 22525 20864 22559
rect 20812 22516 20864 22525
rect 18972 22448 19024 22500
rect 18420 22380 18472 22432
rect 18696 22380 18748 22432
rect 21916 22516 21968 22568
rect 21272 22448 21324 22500
rect 21640 22448 21692 22500
rect 23940 22380 23992 22432
rect 24308 22380 24360 22432
rect 2950 22278 3002 22330
rect 3014 22278 3066 22330
rect 3078 22278 3130 22330
rect 3142 22278 3194 22330
rect 3206 22278 3258 22330
rect 12950 22278 13002 22330
rect 13014 22278 13066 22330
rect 13078 22278 13130 22330
rect 13142 22278 13194 22330
rect 13206 22278 13258 22330
rect 22950 22278 23002 22330
rect 23014 22278 23066 22330
rect 23078 22278 23130 22330
rect 23142 22278 23194 22330
rect 23206 22278 23258 22330
rect 5540 22176 5592 22228
rect 12164 22176 12216 22228
rect 12532 22176 12584 22228
rect 13544 22176 13596 22228
rect 15936 22176 15988 22228
rect 17408 22219 17460 22228
rect 17408 22185 17417 22219
rect 17417 22185 17451 22219
rect 17451 22185 17460 22219
rect 17408 22176 17460 22185
rect 3424 22108 3476 22160
rect 5264 22108 5316 22160
rect 6828 22083 6880 22092
rect 6828 22049 6837 22083
rect 6837 22049 6871 22083
rect 6871 22049 6880 22083
rect 6828 22040 6880 22049
rect 8392 22040 8444 22092
rect 11336 22083 11388 22092
rect 11336 22049 11345 22083
rect 11345 22049 11379 22083
rect 11379 22049 11388 22083
rect 11336 22040 11388 22049
rect 11888 22040 11940 22092
rect 12992 22040 13044 22092
rect 13544 22040 13596 22092
rect 17316 22108 17368 22160
rect 19708 22176 19760 22228
rect 22376 22176 22428 22228
rect 25320 22176 25372 22228
rect 16948 22040 17000 22092
rect 18696 22083 18748 22092
rect 18696 22049 18705 22083
rect 18705 22049 18739 22083
rect 18739 22049 18748 22083
rect 18696 22040 18748 22049
rect 22100 22108 22152 22160
rect 24308 22108 24360 22160
rect 24492 22108 24544 22160
rect 22836 22040 22888 22092
rect 24860 22040 24912 22092
rect 25044 22040 25096 22092
rect 2872 22015 2924 22024
rect 2872 21981 2881 22015
rect 2881 21981 2915 22015
rect 2915 21981 2924 22015
rect 2872 21972 2924 21981
rect 6552 22015 6604 22024
rect 6552 21981 6561 22015
rect 6561 21981 6595 22015
rect 6595 21981 6604 22015
rect 6552 21972 6604 21981
rect 9588 21972 9640 22024
rect 14280 21972 14332 22024
rect 10508 21947 10560 21956
rect 10508 21913 10517 21947
rect 10517 21913 10551 21947
rect 10551 21913 10560 21947
rect 10508 21904 10560 21913
rect 11520 21904 11572 21956
rect 12164 21904 12216 21956
rect 1768 21836 1820 21888
rect 2780 21836 2832 21888
rect 7288 21836 7340 21888
rect 7380 21879 7432 21888
rect 7380 21845 7389 21879
rect 7389 21845 7423 21879
rect 7423 21845 7432 21879
rect 7380 21836 7432 21845
rect 7840 21879 7892 21888
rect 7840 21845 7849 21879
rect 7849 21845 7883 21879
rect 7883 21845 7892 21879
rect 7840 21836 7892 21845
rect 9036 21836 9088 21888
rect 12992 21836 13044 21888
rect 13728 21836 13780 21888
rect 13820 21879 13872 21888
rect 13820 21845 13829 21879
rect 13829 21845 13863 21879
rect 13863 21845 13872 21879
rect 13820 21836 13872 21845
rect 14280 21879 14332 21888
rect 14280 21845 14289 21879
rect 14289 21845 14323 21879
rect 14323 21845 14332 21879
rect 14280 21836 14332 21845
rect 14372 21836 14424 21888
rect 14648 21836 14700 21888
rect 14740 21879 14792 21888
rect 14740 21845 14749 21879
rect 14749 21845 14783 21879
rect 14783 21845 14792 21879
rect 14740 21836 14792 21845
rect 20720 21972 20772 22024
rect 24216 21972 24268 22024
rect 16028 21904 16080 21956
rect 16212 21904 16264 21956
rect 17776 21904 17828 21956
rect 17316 21836 17368 21888
rect 19800 21879 19852 21888
rect 19800 21845 19809 21879
rect 19809 21845 19843 21879
rect 19843 21845 19852 21879
rect 19800 21836 19852 21845
rect 22376 21904 22428 21956
rect 7950 21734 8002 21786
rect 8014 21734 8066 21786
rect 8078 21734 8130 21786
rect 8142 21734 8194 21786
rect 8206 21734 8258 21786
rect 17950 21734 18002 21786
rect 18014 21734 18066 21786
rect 18078 21734 18130 21786
rect 18142 21734 18194 21786
rect 18206 21734 18258 21786
rect 2136 21632 2188 21684
rect 6460 21632 6512 21684
rect 7380 21632 7432 21684
rect 7748 21675 7800 21684
rect 7748 21641 7757 21675
rect 7757 21641 7791 21675
rect 7791 21641 7800 21675
rect 7748 21632 7800 21641
rect 9404 21632 9456 21684
rect 11060 21675 11112 21684
rect 11060 21641 11069 21675
rect 11069 21641 11103 21675
rect 11103 21641 11112 21675
rect 11060 21632 11112 21641
rect 11520 21632 11572 21684
rect 15200 21632 15252 21684
rect 17776 21675 17828 21684
rect 17776 21641 17785 21675
rect 17785 21641 17819 21675
rect 17819 21641 17828 21675
rect 17776 21632 17828 21641
rect 18420 21632 18472 21684
rect 19800 21632 19852 21684
rect 25044 21675 25096 21684
rect 25044 21641 25053 21675
rect 25053 21641 25087 21675
rect 25087 21641 25096 21675
rect 25044 21632 25096 21641
rect 6828 21564 6880 21616
rect 4160 21496 4212 21548
rect 4344 21496 4396 21548
rect 2780 21428 2832 21480
rect 3976 21428 4028 21480
rect 4068 21360 4120 21412
rect 6920 21360 6972 21412
rect 3424 21292 3476 21344
rect 5724 21292 5776 21344
rect 8116 21539 8168 21548
rect 8116 21505 8125 21539
rect 8125 21505 8159 21539
rect 8159 21505 8168 21539
rect 8116 21496 8168 21505
rect 9956 21564 10008 21616
rect 12164 21564 12216 21616
rect 12624 21564 12676 21616
rect 13544 21496 13596 21548
rect 19340 21564 19392 21616
rect 19432 21564 19484 21616
rect 21640 21564 21692 21616
rect 24860 21564 24912 21616
rect 15476 21539 15528 21548
rect 15476 21505 15485 21539
rect 15485 21505 15519 21539
rect 15519 21505 15528 21539
rect 15476 21496 15528 21505
rect 18512 21496 18564 21548
rect 22100 21496 22152 21548
rect 22836 21496 22888 21548
rect 10232 21428 10284 21480
rect 8484 21360 8536 21412
rect 12716 21428 12768 21480
rect 12900 21471 12952 21480
rect 12900 21437 12909 21471
rect 12909 21437 12943 21471
rect 12943 21437 12952 21471
rect 12900 21428 12952 21437
rect 14372 21471 14424 21480
rect 14372 21437 14381 21471
rect 14381 21437 14415 21471
rect 14415 21437 14424 21471
rect 14372 21428 14424 21437
rect 11428 21360 11480 21412
rect 9128 21292 9180 21344
rect 12164 21292 12216 21344
rect 14004 21360 14056 21412
rect 14648 21428 14700 21480
rect 20076 21428 20128 21480
rect 24400 21471 24452 21480
rect 24400 21437 24409 21471
rect 24409 21437 24443 21471
rect 24443 21437 24452 21471
rect 24400 21428 24452 21437
rect 17868 21360 17920 21412
rect 14740 21292 14792 21344
rect 16212 21292 16264 21344
rect 19432 21360 19484 21412
rect 18512 21292 18564 21344
rect 19616 21335 19668 21344
rect 19616 21301 19625 21335
rect 19625 21301 19659 21335
rect 19659 21301 19668 21335
rect 19616 21292 19668 21301
rect 20720 21292 20772 21344
rect 22836 21292 22888 21344
rect 25044 21428 25096 21480
rect 2950 21190 3002 21242
rect 3014 21190 3066 21242
rect 3078 21190 3130 21242
rect 3142 21190 3194 21242
rect 3206 21190 3258 21242
rect 12950 21190 13002 21242
rect 13014 21190 13066 21242
rect 13078 21190 13130 21242
rect 13142 21190 13194 21242
rect 13206 21190 13258 21242
rect 22950 21190 23002 21242
rect 23014 21190 23066 21242
rect 23078 21190 23130 21242
rect 23142 21190 23194 21242
rect 23206 21190 23258 21242
rect 2872 21131 2924 21140
rect 2872 21097 2881 21131
rect 2881 21097 2915 21131
rect 2915 21097 2924 21131
rect 2872 21088 2924 21097
rect 7288 21088 7340 21140
rect 8116 21088 8168 21140
rect 12348 21088 12400 21140
rect 12624 21131 12676 21140
rect 12624 21097 12633 21131
rect 12633 21097 12667 21131
rect 12667 21097 12676 21131
rect 12624 21088 12676 21097
rect 12716 21088 12768 21140
rect 14004 21088 14056 21140
rect 16212 21088 16264 21140
rect 24308 21088 24360 21140
rect 7012 21020 7064 21072
rect 3424 20995 3476 21004
rect 3424 20961 3433 20995
rect 3433 20961 3467 20995
rect 3467 20961 3476 20995
rect 3424 20952 3476 20961
rect 5264 20995 5316 21004
rect 5264 20961 5273 20995
rect 5273 20961 5307 20995
rect 5307 20961 5316 20995
rect 5264 20952 5316 20961
rect 5816 20952 5868 21004
rect 6276 20952 6328 21004
rect 11704 21020 11756 21072
rect 3884 20884 3936 20936
rect 4068 20884 4120 20936
rect 4988 20927 5040 20936
rect 4988 20893 4997 20927
rect 4997 20893 5031 20927
rect 5031 20893 5040 20927
rect 4988 20884 5040 20893
rect 6368 20884 6420 20936
rect 7104 20884 7156 20936
rect 10324 20952 10376 21004
rect 10784 20995 10836 21004
rect 10784 20961 10793 20995
rect 10793 20961 10827 20995
rect 10827 20961 10836 20995
rect 10784 20952 10836 20961
rect 22192 21020 22244 21072
rect 13360 20952 13412 21004
rect 14556 20995 14608 21004
rect 14556 20961 14565 20995
rect 14565 20961 14599 20995
rect 14599 20961 14608 20995
rect 14556 20952 14608 20961
rect 18604 20995 18656 21004
rect 18604 20961 18613 20995
rect 18613 20961 18647 20995
rect 18647 20961 18656 20995
rect 18604 20952 18656 20961
rect 19616 20952 19668 21004
rect 22100 20952 22152 21004
rect 7748 20816 7800 20868
rect 13544 20927 13596 20936
rect 13544 20893 13553 20927
rect 13553 20893 13587 20927
rect 13587 20893 13596 20927
rect 13544 20884 13596 20893
rect 18512 20927 18564 20936
rect 18512 20893 18521 20927
rect 18521 20893 18555 20927
rect 18555 20893 18564 20927
rect 18512 20884 18564 20893
rect 4344 20791 4396 20800
rect 4344 20757 4353 20791
rect 4353 20757 4387 20791
rect 4387 20757 4396 20791
rect 4344 20748 4396 20757
rect 6920 20748 6972 20800
rect 7288 20791 7340 20800
rect 7288 20757 7297 20791
rect 7297 20757 7331 20791
rect 7331 20757 7340 20791
rect 7288 20748 7340 20757
rect 8300 20748 8352 20800
rect 8944 20748 8996 20800
rect 9956 20748 10008 20800
rect 11612 20816 11664 20868
rect 12072 20816 12124 20868
rect 16212 20816 16264 20868
rect 17224 20816 17276 20868
rect 21824 20884 21876 20936
rect 24860 21020 24912 21072
rect 20720 20816 20772 20868
rect 21272 20816 21324 20868
rect 12348 20748 12400 20800
rect 16028 20791 16080 20800
rect 16028 20757 16037 20791
rect 16037 20757 16071 20791
rect 16071 20757 16080 20791
rect 16028 20748 16080 20757
rect 16856 20791 16908 20800
rect 16856 20757 16865 20791
rect 16865 20757 16899 20791
rect 16899 20757 16908 20791
rect 16856 20748 16908 20757
rect 17132 20748 17184 20800
rect 20904 20748 20956 20800
rect 23756 20816 23808 20868
rect 7950 20646 8002 20698
rect 8014 20646 8066 20698
rect 8078 20646 8130 20698
rect 8142 20646 8194 20698
rect 8206 20646 8258 20698
rect 17950 20646 18002 20698
rect 18014 20646 18066 20698
rect 18078 20646 18130 20698
rect 18142 20646 18194 20698
rect 18206 20646 18258 20698
rect 1768 20451 1820 20460
rect 1768 20417 1777 20451
rect 1777 20417 1811 20451
rect 1811 20417 1820 20451
rect 1768 20408 1820 20417
rect 4988 20544 5040 20596
rect 5448 20544 5500 20596
rect 4252 20476 4304 20528
rect 1308 20340 1360 20392
rect 5724 20204 5776 20256
rect 7012 20408 7064 20460
rect 7196 20408 7248 20460
rect 10324 20587 10376 20596
rect 10324 20553 10333 20587
rect 10333 20553 10367 20587
rect 10367 20553 10376 20587
rect 10324 20544 10376 20553
rect 12440 20544 12492 20596
rect 14740 20587 14792 20596
rect 14740 20553 14749 20587
rect 14749 20553 14783 20587
rect 14783 20553 14792 20587
rect 14740 20544 14792 20553
rect 15108 20544 15160 20596
rect 16396 20587 16448 20596
rect 16396 20553 16405 20587
rect 16405 20553 16439 20587
rect 16439 20553 16448 20587
rect 16396 20544 16448 20553
rect 16856 20544 16908 20596
rect 9864 20476 9916 20528
rect 11980 20476 12032 20528
rect 13452 20476 13504 20528
rect 13636 20408 13688 20460
rect 16764 20408 16816 20460
rect 8300 20340 8352 20392
rect 9864 20340 9916 20392
rect 10968 20340 11020 20392
rect 11704 20340 11756 20392
rect 6368 20204 6420 20256
rect 7012 20247 7064 20256
rect 7012 20213 7021 20247
rect 7021 20213 7055 20247
rect 7055 20213 7064 20247
rect 7012 20204 7064 20213
rect 7104 20204 7156 20256
rect 7840 20272 7892 20324
rect 10140 20272 10192 20324
rect 10692 20272 10744 20324
rect 16028 20340 16080 20392
rect 18880 20476 18932 20528
rect 21272 20544 21324 20596
rect 21824 20544 21876 20596
rect 22376 20587 22428 20596
rect 22376 20553 22385 20587
rect 22385 20553 22419 20587
rect 22419 20553 22428 20587
rect 22376 20544 22428 20553
rect 22744 20544 22796 20596
rect 19432 20476 19484 20528
rect 18696 20451 18748 20460
rect 18696 20417 18705 20451
rect 18705 20417 18739 20451
rect 18739 20417 18748 20451
rect 18696 20408 18748 20417
rect 20720 20340 20772 20392
rect 24400 20544 24452 20596
rect 24860 20544 24912 20596
rect 25044 20451 25096 20460
rect 25044 20417 25053 20451
rect 25053 20417 25087 20451
rect 25087 20417 25096 20451
rect 25044 20408 25096 20417
rect 24216 20340 24268 20392
rect 20628 20272 20680 20324
rect 10416 20204 10468 20256
rect 14372 20247 14424 20256
rect 14372 20213 14381 20247
rect 14381 20213 14415 20247
rect 14415 20213 14424 20247
rect 14372 20204 14424 20213
rect 15660 20204 15712 20256
rect 18236 20204 18288 20256
rect 2950 20102 3002 20154
rect 3014 20102 3066 20154
rect 3078 20102 3130 20154
rect 3142 20102 3194 20154
rect 3206 20102 3258 20154
rect 12950 20102 13002 20154
rect 13014 20102 13066 20154
rect 13078 20102 13130 20154
rect 13142 20102 13194 20154
rect 13206 20102 13258 20154
rect 22950 20102 23002 20154
rect 23014 20102 23066 20154
rect 23078 20102 23130 20154
rect 23142 20102 23194 20154
rect 23206 20102 23258 20154
rect 5356 20000 5408 20052
rect 7104 20000 7156 20052
rect 8392 20000 8444 20052
rect 6828 19864 6880 19916
rect 7380 19864 7432 19916
rect 9128 20043 9180 20052
rect 9128 20009 9137 20043
rect 9137 20009 9171 20043
rect 9171 20009 9180 20043
rect 9128 20000 9180 20009
rect 9956 20000 10008 20052
rect 12532 20000 12584 20052
rect 24216 20000 24268 20052
rect 24860 20000 24912 20052
rect 19800 19932 19852 19984
rect 11980 19907 12032 19916
rect 11980 19873 11989 19907
rect 11989 19873 12023 19907
rect 12023 19873 12032 19907
rect 11980 19864 12032 19873
rect 18328 19907 18380 19916
rect 18328 19873 18337 19907
rect 18337 19873 18371 19907
rect 18371 19873 18380 19907
rect 18328 19864 18380 19873
rect 20720 19864 20772 19916
rect 25136 19864 25188 19916
rect 3332 19796 3384 19848
rect 8484 19796 8536 19848
rect 10416 19796 10468 19848
rect 11704 19839 11756 19848
rect 11704 19805 11713 19839
rect 11713 19805 11747 19839
rect 11747 19805 11756 19839
rect 11704 19796 11756 19805
rect 14188 19796 14240 19848
rect 17224 19839 17276 19848
rect 17224 19805 17233 19839
rect 17233 19805 17267 19839
rect 17267 19805 17276 19839
rect 17224 19796 17276 19805
rect 18236 19839 18288 19848
rect 18236 19805 18245 19839
rect 18245 19805 18279 19839
rect 18279 19805 18288 19839
rect 18236 19796 18288 19805
rect 20996 19796 21048 19848
rect 21088 19796 21140 19848
rect 24768 19796 24820 19848
rect 6368 19728 6420 19780
rect 7656 19728 7708 19780
rect 10784 19728 10836 19780
rect 13084 19728 13136 19780
rect 20444 19728 20496 19780
rect 22652 19728 22704 19780
rect 1860 19660 1912 19712
rect 6184 19660 6236 19712
rect 6736 19660 6788 19712
rect 7472 19703 7524 19712
rect 7472 19669 7481 19703
rect 7481 19669 7515 19703
rect 7515 19669 7524 19703
rect 7472 19660 7524 19669
rect 7840 19703 7892 19712
rect 7840 19669 7849 19703
rect 7849 19669 7883 19703
rect 7883 19669 7892 19703
rect 7840 19660 7892 19669
rect 9588 19703 9640 19712
rect 9588 19669 9597 19703
rect 9597 19669 9631 19703
rect 9631 19669 9640 19703
rect 9588 19660 9640 19669
rect 10600 19660 10652 19712
rect 17040 19660 17092 19712
rect 17500 19660 17552 19712
rect 19892 19660 19944 19712
rect 21732 19660 21784 19712
rect 7950 19558 8002 19610
rect 8014 19558 8066 19610
rect 8078 19558 8130 19610
rect 8142 19558 8194 19610
rect 8206 19558 8258 19610
rect 17950 19558 18002 19610
rect 18014 19558 18066 19610
rect 18078 19558 18130 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 4896 19499 4948 19508
rect 4896 19465 4905 19499
rect 4905 19465 4939 19499
rect 4939 19465 4948 19499
rect 4896 19456 4948 19465
rect 5724 19456 5776 19508
rect 6368 19388 6420 19440
rect 6460 19320 6512 19372
rect 6828 19320 6880 19372
rect 9404 19456 9456 19508
rect 11888 19456 11940 19508
rect 13084 19499 13136 19508
rect 13084 19465 13093 19499
rect 13093 19465 13127 19499
rect 13127 19465 13136 19499
rect 13084 19456 13136 19465
rect 19248 19456 19300 19508
rect 11612 19388 11664 19440
rect 12716 19388 12768 19440
rect 13912 19388 13964 19440
rect 19156 19388 19208 19440
rect 22100 19388 22152 19440
rect 24860 19388 24912 19440
rect 9680 19320 9732 19372
rect 12440 19320 12492 19372
rect 6920 19252 6972 19304
rect 9956 19252 10008 19304
rect 10324 19252 10376 19304
rect 13544 19295 13596 19304
rect 8760 19184 8812 19236
rect 13544 19261 13553 19295
rect 13553 19261 13587 19295
rect 13587 19261 13596 19295
rect 13544 19252 13596 19261
rect 13360 19184 13412 19236
rect 14832 19320 14884 19372
rect 18788 19363 18840 19372
rect 18788 19329 18797 19363
rect 18797 19329 18831 19363
rect 18831 19329 18840 19363
rect 18788 19320 18840 19329
rect 22284 19320 22336 19372
rect 23388 19363 23440 19372
rect 23388 19329 23397 19363
rect 23397 19329 23431 19363
rect 23431 19329 23440 19363
rect 23388 19320 23440 19329
rect 24492 19320 24544 19372
rect 25228 19363 25280 19372
rect 25228 19329 25237 19363
rect 25237 19329 25271 19363
rect 25271 19329 25280 19363
rect 25228 19320 25280 19329
rect 18512 19184 18564 19236
rect 9864 19116 9916 19168
rect 17408 19159 17460 19168
rect 17408 19125 17417 19159
rect 17417 19125 17451 19159
rect 17451 19125 17460 19159
rect 17408 19116 17460 19125
rect 18788 19116 18840 19168
rect 2950 19014 3002 19066
rect 3014 19014 3066 19066
rect 3078 19014 3130 19066
rect 3142 19014 3194 19066
rect 3206 19014 3258 19066
rect 12950 19014 13002 19066
rect 13014 19014 13066 19066
rect 13078 19014 13130 19066
rect 13142 19014 13194 19066
rect 13206 19014 13258 19066
rect 22950 19014 23002 19066
rect 23014 19014 23066 19066
rect 23078 19014 23130 19066
rect 23142 19014 23194 19066
rect 23206 19014 23258 19066
rect 3976 18955 4028 18964
rect 3976 18921 3985 18955
rect 3985 18921 4019 18955
rect 4019 18921 4028 18955
rect 3976 18912 4028 18921
rect 8300 18912 8352 18964
rect 11428 18912 11480 18964
rect 12624 18912 12676 18964
rect 9772 18887 9824 18896
rect 9772 18853 9781 18887
rect 9781 18853 9815 18887
rect 9815 18853 9824 18887
rect 9772 18844 9824 18853
rect 9956 18844 10008 18896
rect 12072 18844 12124 18896
rect 6920 18776 6972 18828
rect 7932 18776 7984 18828
rect 8668 18776 8720 18828
rect 12808 18776 12860 18828
rect 14004 18844 14056 18896
rect 2780 18708 2832 18760
rect 4160 18751 4212 18760
rect 4160 18717 4169 18751
rect 4169 18717 4203 18751
rect 4203 18717 4212 18751
rect 4160 18708 4212 18717
rect 8576 18751 8628 18760
rect 8576 18717 8585 18751
rect 8585 18717 8619 18751
rect 8619 18717 8628 18751
rect 8576 18708 8628 18717
rect 12532 18708 12584 18760
rect 15660 18776 15712 18828
rect 19064 18912 19116 18964
rect 22560 18912 22612 18964
rect 23204 18912 23256 18964
rect 24216 18955 24268 18964
rect 24216 18921 24225 18955
rect 24225 18921 24259 18955
rect 24259 18921 24268 18955
rect 24216 18912 24268 18921
rect 19984 18844 20036 18896
rect 20536 18844 20588 18896
rect 17592 18776 17644 18828
rect 19616 18819 19668 18828
rect 19616 18785 19625 18819
rect 19625 18785 19659 18819
rect 19659 18785 19668 18819
rect 19616 18776 19668 18785
rect 20444 18776 20496 18828
rect 13544 18708 13596 18760
rect 21548 18708 21600 18760
rect 9772 18640 9824 18692
rect 13728 18640 13780 18692
rect 1768 18572 1820 18624
rect 7656 18572 7708 18624
rect 7932 18572 7984 18624
rect 9220 18615 9272 18624
rect 9220 18581 9229 18615
rect 9229 18581 9263 18615
rect 9263 18581 9272 18615
rect 9220 18572 9272 18581
rect 10140 18572 10192 18624
rect 11796 18572 11848 18624
rect 13544 18572 13596 18624
rect 14188 18572 14240 18624
rect 20352 18572 20404 18624
rect 21456 18615 21508 18624
rect 21456 18581 21465 18615
rect 21465 18581 21499 18615
rect 21499 18581 21508 18615
rect 21456 18572 21508 18581
rect 22836 18776 22888 18828
rect 24308 18708 24360 18760
rect 22560 18572 22612 18624
rect 22744 18572 22796 18624
rect 23664 18640 23716 18692
rect 24216 18572 24268 18624
rect 7950 18470 8002 18522
rect 8014 18470 8066 18522
rect 8078 18470 8130 18522
rect 8142 18470 8194 18522
rect 8206 18470 8258 18522
rect 17950 18470 18002 18522
rect 18014 18470 18066 18522
rect 18078 18470 18130 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 11244 18368 11296 18420
rect 12440 18411 12492 18420
rect 12440 18377 12449 18411
rect 12449 18377 12483 18411
rect 12483 18377 12492 18411
rect 12440 18368 12492 18377
rect 13636 18411 13688 18420
rect 13636 18377 13645 18411
rect 13645 18377 13679 18411
rect 13679 18377 13688 18411
rect 13636 18368 13688 18377
rect 17776 18368 17828 18420
rect 1860 18232 1912 18284
rect 8300 18232 8352 18284
rect 9772 18232 9824 18284
rect 17132 18343 17184 18352
rect 17132 18309 17141 18343
rect 17141 18309 17175 18343
rect 17175 18309 17184 18343
rect 17132 18300 17184 18309
rect 21824 18368 21876 18420
rect 22744 18368 22796 18420
rect 22928 18368 22980 18420
rect 23204 18368 23256 18420
rect 12440 18232 12492 18284
rect 13912 18232 13964 18284
rect 18788 18232 18840 18284
rect 22008 18232 22060 18284
rect 22836 18300 22888 18352
rect 24216 18300 24268 18352
rect 1308 18164 1360 18216
rect 6276 18164 6328 18216
rect 6828 18164 6880 18216
rect 8576 18164 8628 18216
rect 11152 18207 11204 18216
rect 11152 18173 11161 18207
rect 11161 18173 11195 18207
rect 11195 18173 11204 18207
rect 11152 18164 11204 18173
rect 12716 18164 12768 18216
rect 13360 18164 13412 18216
rect 13820 18164 13872 18216
rect 12440 18096 12492 18148
rect 17776 18164 17828 18216
rect 18512 18164 18564 18216
rect 20076 18164 20128 18216
rect 23296 18164 23348 18216
rect 2136 18028 2188 18080
rect 7288 18028 7340 18080
rect 10692 18028 10744 18080
rect 13912 18028 13964 18080
rect 18512 18028 18564 18080
rect 21824 18028 21876 18080
rect 2950 17926 3002 17978
rect 3014 17926 3066 17978
rect 3078 17926 3130 17978
rect 3142 17926 3194 17978
rect 3206 17926 3258 17978
rect 12950 17926 13002 17978
rect 13014 17926 13066 17978
rect 13078 17926 13130 17978
rect 13142 17926 13194 17978
rect 13206 17926 13258 17978
rect 22950 17926 23002 17978
rect 23014 17926 23066 17978
rect 23078 17926 23130 17978
rect 23142 17926 23194 17978
rect 23206 17926 23258 17978
rect 4344 17824 4396 17876
rect 6920 17799 6972 17808
rect 6920 17765 6929 17799
rect 6929 17765 6963 17799
rect 6963 17765 6972 17799
rect 6920 17756 6972 17765
rect 8300 17824 8352 17876
rect 6276 17688 6328 17740
rect 7656 17731 7708 17740
rect 7656 17697 7665 17731
rect 7665 17697 7699 17731
rect 7699 17697 7708 17731
rect 7656 17688 7708 17697
rect 8208 17620 8260 17672
rect 5724 17552 5776 17604
rect 6552 17552 6604 17604
rect 4804 17527 4856 17536
rect 4804 17493 4813 17527
rect 4813 17493 4847 17527
rect 4847 17493 4856 17527
rect 4804 17484 4856 17493
rect 4896 17484 4948 17536
rect 11888 17824 11940 17876
rect 12808 17824 12860 17876
rect 13728 17824 13780 17876
rect 15292 17824 15344 17876
rect 18328 17824 18380 17876
rect 18972 17867 19024 17876
rect 18972 17833 18981 17867
rect 18981 17833 19015 17867
rect 19015 17833 19024 17867
rect 18972 17824 19024 17833
rect 11520 17731 11572 17740
rect 8392 17620 8444 17672
rect 9312 17620 9364 17672
rect 11520 17697 11529 17731
rect 11529 17697 11563 17731
rect 11563 17697 11572 17731
rect 11520 17688 11572 17697
rect 11980 17688 12032 17740
rect 13636 17688 13688 17740
rect 13912 17688 13964 17740
rect 15476 17688 15528 17740
rect 16856 17688 16908 17740
rect 17776 17731 17828 17740
rect 17776 17697 17785 17731
rect 17785 17697 17819 17731
rect 17819 17697 17828 17731
rect 17776 17688 17828 17697
rect 17868 17688 17920 17740
rect 14280 17620 14332 17672
rect 10600 17552 10652 17604
rect 11152 17552 11204 17604
rect 8300 17527 8352 17536
rect 8300 17493 8309 17527
rect 8309 17493 8343 17527
rect 8343 17493 8352 17527
rect 8300 17484 8352 17493
rect 9128 17527 9180 17536
rect 9128 17493 9137 17527
rect 9137 17493 9171 17527
rect 9171 17493 9180 17527
rect 9128 17484 9180 17493
rect 12532 17527 12584 17536
rect 12532 17493 12541 17527
rect 12541 17493 12575 17527
rect 12575 17493 12584 17527
rect 12532 17484 12584 17493
rect 16488 17552 16540 17604
rect 18604 17620 18656 17672
rect 22008 17688 22060 17740
rect 23388 17731 23440 17740
rect 23388 17697 23397 17731
rect 23397 17697 23431 17731
rect 23431 17697 23440 17731
rect 23388 17688 23440 17697
rect 18328 17595 18380 17604
rect 18328 17561 18337 17595
rect 18337 17561 18371 17595
rect 18371 17561 18380 17595
rect 18328 17552 18380 17561
rect 18880 17552 18932 17604
rect 17868 17484 17920 17536
rect 18696 17484 18748 17536
rect 24676 17620 24728 17672
rect 19064 17552 19116 17604
rect 20720 17552 20772 17604
rect 22100 17552 22152 17604
rect 21180 17527 21232 17536
rect 21180 17493 21189 17527
rect 21189 17493 21223 17527
rect 21223 17493 21232 17527
rect 21180 17484 21232 17493
rect 21824 17484 21876 17536
rect 7950 17382 8002 17434
rect 8014 17382 8066 17434
rect 8078 17382 8130 17434
rect 8142 17382 8194 17434
rect 8206 17382 8258 17434
rect 17950 17382 18002 17434
rect 18014 17382 18066 17434
rect 18078 17382 18130 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 4160 17280 4212 17332
rect 7840 17280 7892 17332
rect 9588 17280 9640 17332
rect 5724 17212 5776 17264
rect 4804 17144 4856 17196
rect 12072 17323 12124 17332
rect 12072 17289 12081 17323
rect 12081 17289 12115 17323
rect 12115 17289 12124 17323
rect 12072 17280 12124 17289
rect 12164 17323 12216 17332
rect 12164 17289 12173 17323
rect 12173 17289 12207 17323
rect 12207 17289 12216 17323
rect 12164 17280 12216 17289
rect 12716 17280 12768 17332
rect 6920 17144 6972 17196
rect 8760 17144 8812 17196
rect 6092 17076 6144 17128
rect 6552 17076 6604 17128
rect 4068 16940 4120 16992
rect 9128 16940 9180 16992
rect 12716 17144 12768 17196
rect 10692 17119 10744 17128
rect 10692 17085 10701 17119
rect 10701 17085 10735 17119
rect 10735 17085 10744 17119
rect 10692 17076 10744 17085
rect 11060 17076 11112 17128
rect 13728 17280 13780 17332
rect 16672 17323 16724 17332
rect 16672 17289 16681 17323
rect 16681 17289 16715 17323
rect 16715 17289 16724 17323
rect 16672 17280 16724 17289
rect 19064 17323 19116 17332
rect 19064 17289 19073 17323
rect 19073 17289 19107 17323
rect 19107 17289 19116 17323
rect 19064 17280 19116 17289
rect 19616 17280 19668 17332
rect 14372 17212 14424 17264
rect 20720 17212 20772 17264
rect 21916 17212 21968 17264
rect 23296 17280 23348 17332
rect 24216 17280 24268 17332
rect 13912 17144 13964 17196
rect 18696 17144 18748 17196
rect 13728 17119 13780 17128
rect 13728 17085 13737 17119
rect 13737 17085 13771 17119
rect 13771 17085 13780 17119
rect 13728 17076 13780 17085
rect 16856 17076 16908 17128
rect 17592 17119 17644 17128
rect 17592 17085 17601 17119
rect 17601 17085 17635 17119
rect 17635 17085 17644 17119
rect 17592 17076 17644 17085
rect 20720 17076 20772 17128
rect 21180 17119 21232 17128
rect 21180 17085 21189 17119
rect 21189 17085 21223 17119
rect 21223 17085 21232 17119
rect 21180 17076 21232 17085
rect 21548 17076 21600 17128
rect 22008 17119 22060 17128
rect 22008 17085 22017 17119
rect 22017 17085 22051 17119
rect 22051 17085 22060 17119
rect 22008 17076 22060 17085
rect 11796 16940 11848 16992
rect 12440 16940 12492 16992
rect 16120 17008 16172 17060
rect 14740 16940 14792 16992
rect 18328 16940 18380 16992
rect 2950 16838 3002 16890
rect 3014 16838 3066 16890
rect 3078 16838 3130 16890
rect 3142 16838 3194 16890
rect 3206 16838 3258 16890
rect 12950 16838 13002 16890
rect 13014 16838 13066 16890
rect 13078 16838 13130 16890
rect 13142 16838 13194 16890
rect 13206 16838 13258 16890
rect 22950 16838 23002 16890
rect 23014 16838 23066 16890
rect 23078 16838 23130 16890
rect 23142 16838 23194 16890
rect 23206 16838 23258 16890
rect 6092 16736 6144 16788
rect 6920 16736 6972 16788
rect 2780 16600 2832 16652
rect 6276 16600 6328 16652
rect 4068 16532 4120 16584
rect 7840 16736 7892 16788
rect 11428 16779 11480 16788
rect 11428 16745 11437 16779
rect 11437 16745 11471 16779
rect 11471 16745 11480 16779
rect 11428 16736 11480 16745
rect 14924 16736 14976 16788
rect 15384 16736 15436 16788
rect 16212 16779 16264 16788
rect 16212 16745 16221 16779
rect 16221 16745 16255 16779
rect 16255 16745 16264 16779
rect 16212 16736 16264 16745
rect 18512 16736 18564 16788
rect 18788 16736 18840 16788
rect 21548 16736 21600 16788
rect 9864 16668 9916 16720
rect 9588 16643 9640 16652
rect 9588 16609 9597 16643
rect 9597 16609 9631 16643
rect 9631 16609 9640 16643
rect 9588 16600 9640 16609
rect 8852 16532 8904 16584
rect 10784 16643 10836 16652
rect 10784 16609 10793 16643
rect 10793 16609 10827 16643
rect 10827 16609 10836 16643
rect 10784 16600 10836 16609
rect 11704 16668 11756 16720
rect 10600 16532 10652 16584
rect 15476 16668 15528 16720
rect 19984 16600 20036 16652
rect 21180 16600 21232 16652
rect 22560 16600 22612 16652
rect 24216 16736 24268 16788
rect 7748 16396 7800 16448
rect 9128 16439 9180 16448
rect 9128 16405 9137 16439
rect 9137 16405 9171 16439
rect 9171 16405 9180 16439
rect 9128 16396 9180 16405
rect 10508 16464 10560 16516
rect 11428 16464 11480 16516
rect 11244 16396 11296 16448
rect 15752 16575 15804 16584
rect 15752 16541 15761 16575
rect 15761 16541 15795 16575
rect 15795 16541 15804 16575
rect 15752 16532 15804 16541
rect 22008 16532 22060 16584
rect 13636 16439 13688 16448
rect 13636 16405 13645 16439
rect 13645 16405 13679 16439
rect 13679 16405 13688 16439
rect 13636 16396 13688 16405
rect 15200 16396 15252 16448
rect 20260 16439 20312 16448
rect 20260 16405 20269 16439
rect 20269 16405 20303 16439
rect 20303 16405 20312 16439
rect 20260 16396 20312 16405
rect 21364 16396 21416 16448
rect 21640 16439 21692 16448
rect 21640 16405 21649 16439
rect 21649 16405 21683 16439
rect 21683 16405 21692 16439
rect 21640 16396 21692 16405
rect 21824 16396 21876 16448
rect 7950 16294 8002 16346
rect 8014 16294 8066 16346
rect 8078 16294 8130 16346
rect 8142 16294 8194 16346
rect 8206 16294 8258 16346
rect 17950 16294 18002 16346
rect 18014 16294 18066 16346
rect 18078 16294 18130 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 6460 16192 6512 16244
rect 9128 16192 9180 16244
rect 12532 16192 12584 16244
rect 16948 16192 17000 16244
rect 17776 16192 17828 16244
rect 1768 16099 1820 16108
rect 1768 16065 1777 16099
rect 1777 16065 1811 16099
rect 1811 16065 1820 16099
rect 1768 16056 1820 16065
rect 7840 16056 7892 16108
rect 9220 16124 9272 16176
rect 16212 16167 16264 16176
rect 16212 16133 16221 16167
rect 16221 16133 16255 16167
rect 16255 16133 16264 16167
rect 16212 16124 16264 16133
rect 19248 16124 19300 16176
rect 1308 15988 1360 16040
rect 8484 15988 8536 16040
rect 9404 16056 9456 16108
rect 11704 16056 11756 16108
rect 12808 16056 12860 16108
rect 9312 16031 9364 16040
rect 9312 15997 9321 16031
rect 9321 15997 9355 16031
rect 9355 15997 9364 16031
rect 9312 15988 9364 15997
rect 10876 16031 10928 16040
rect 10876 15997 10885 16031
rect 10885 15997 10919 16031
rect 10919 15997 10928 16031
rect 10876 15988 10928 15997
rect 8760 15895 8812 15904
rect 8760 15861 8769 15895
rect 8769 15861 8803 15895
rect 8803 15861 8812 15895
rect 8760 15852 8812 15861
rect 8852 15852 8904 15904
rect 14832 15895 14884 15904
rect 14832 15861 14841 15895
rect 14841 15861 14875 15895
rect 14875 15861 14884 15895
rect 14832 15852 14884 15861
rect 19800 16056 19852 16108
rect 23664 16056 23716 16108
rect 23940 16099 23992 16108
rect 23940 16065 23949 16099
rect 23949 16065 23983 16099
rect 23983 16065 23992 16099
rect 23940 16056 23992 16065
rect 15292 16031 15344 16040
rect 15292 15997 15301 16031
rect 15301 15997 15335 16031
rect 15335 15997 15344 16031
rect 15292 15988 15344 15997
rect 15476 16031 15528 16040
rect 15476 15997 15485 16031
rect 15485 15997 15519 16031
rect 15519 15997 15528 16031
rect 15476 15988 15528 15997
rect 19524 16031 19576 16040
rect 19524 15997 19533 16031
rect 19533 15997 19567 16031
rect 19567 15997 19576 16031
rect 19524 15988 19576 15997
rect 16028 15963 16080 15972
rect 16028 15929 16037 15963
rect 16037 15929 16071 15963
rect 16071 15929 16080 15963
rect 16028 15920 16080 15929
rect 16580 15920 16632 15972
rect 24860 16056 24912 16108
rect 24768 16031 24820 16040
rect 24768 15997 24777 16031
rect 24777 15997 24811 16031
rect 24811 15997 24820 16031
rect 24768 15988 24820 15997
rect 16672 15852 16724 15904
rect 19432 15852 19484 15904
rect 19800 15852 19852 15904
rect 23940 15920 23992 15972
rect 23664 15852 23716 15904
rect 2950 15750 3002 15802
rect 3014 15750 3066 15802
rect 3078 15750 3130 15802
rect 3142 15750 3194 15802
rect 3206 15750 3258 15802
rect 12950 15750 13002 15802
rect 13014 15750 13066 15802
rect 13078 15750 13130 15802
rect 13142 15750 13194 15802
rect 13206 15750 13258 15802
rect 22950 15750 23002 15802
rect 23014 15750 23066 15802
rect 23078 15750 23130 15802
rect 23142 15750 23194 15802
rect 23206 15750 23258 15802
rect 6552 15648 6604 15700
rect 7288 15648 7340 15700
rect 9312 15648 9364 15700
rect 10508 15648 10560 15700
rect 11060 15648 11112 15700
rect 11888 15648 11940 15700
rect 12808 15691 12860 15700
rect 12808 15657 12817 15691
rect 12817 15657 12851 15691
rect 12851 15657 12860 15691
rect 12808 15648 12860 15657
rect 17592 15648 17644 15700
rect 7932 15580 7984 15632
rect 10600 15512 10652 15564
rect 11244 15512 11296 15564
rect 16856 15512 16908 15564
rect 18328 15512 18380 15564
rect 6920 15376 6972 15428
rect 7380 15376 7432 15428
rect 6276 15308 6328 15360
rect 6828 15308 6880 15360
rect 14464 15487 14516 15496
rect 14464 15453 14473 15487
rect 14473 15453 14507 15487
rect 14507 15453 14516 15487
rect 14464 15444 14516 15453
rect 17776 15444 17828 15496
rect 19984 15512 20036 15564
rect 20260 15512 20312 15564
rect 23296 15512 23348 15564
rect 24860 15512 24912 15564
rect 9680 15376 9732 15428
rect 11244 15376 11296 15428
rect 16120 15376 16172 15428
rect 16672 15376 16724 15428
rect 17868 15376 17920 15428
rect 19800 15419 19852 15428
rect 19800 15385 19809 15419
rect 19809 15385 19843 15419
rect 19843 15385 19852 15419
rect 19800 15376 19852 15385
rect 14648 15308 14700 15360
rect 18512 15351 18564 15360
rect 18512 15317 18521 15351
rect 18521 15317 18555 15351
rect 18555 15317 18564 15351
rect 18512 15308 18564 15317
rect 20536 15444 20588 15496
rect 21824 15487 21876 15496
rect 21824 15453 21833 15487
rect 21833 15453 21867 15487
rect 21867 15453 21876 15487
rect 21824 15444 21876 15453
rect 22652 15487 22704 15496
rect 22652 15453 22661 15487
rect 22661 15453 22695 15487
rect 22695 15453 22704 15487
rect 22652 15444 22704 15453
rect 22008 15376 22060 15428
rect 20996 15308 21048 15360
rect 23296 15308 23348 15360
rect 7950 15206 8002 15258
rect 8014 15206 8066 15258
rect 8078 15206 8130 15258
rect 8142 15206 8194 15258
rect 8206 15206 8258 15258
rect 17950 15206 18002 15258
rect 18014 15206 18066 15258
rect 18078 15206 18130 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 10876 15104 10928 15156
rect 14832 15104 14884 15156
rect 15292 15104 15344 15156
rect 16212 15104 16264 15156
rect 11244 15036 11296 15088
rect 12256 15036 12308 15088
rect 12808 15036 12860 15088
rect 15936 15036 15988 15088
rect 18512 15147 18564 15156
rect 18512 15113 18521 15147
rect 18521 15113 18555 15147
rect 18555 15113 18564 15147
rect 18512 15104 18564 15113
rect 19524 15147 19576 15156
rect 19524 15113 19533 15147
rect 19533 15113 19567 15147
rect 19567 15113 19576 15147
rect 19524 15104 19576 15113
rect 20352 15104 20404 15156
rect 12440 14968 12492 15020
rect 14924 14968 14976 15020
rect 15108 14968 15160 15020
rect 20628 14968 20680 15020
rect 24584 15104 24636 15156
rect 24860 15036 24912 15088
rect 22100 15011 22152 15020
rect 22100 14977 22109 15011
rect 22109 14977 22143 15011
rect 22143 14977 22152 15011
rect 22100 14968 22152 14977
rect 23756 14968 23808 15020
rect 9864 14900 9916 14952
rect 10600 14943 10652 14952
rect 10600 14909 10609 14943
rect 10609 14909 10643 14943
rect 10643 14909 10652 14943
rect 10600 14900 10652 14909
rect 12256 14900 12308 14952
rect 13636 14943 13688 14952
rect 13636 14909 13645 14943
rect 13645 14909 13679 14943
rect 13679 14909 13688 14943
rect 13636 14900 13688 14909
rect 17132 14943 17184 14952
rect 17132 14909 17141 14943
rect 17141 14909 17175 14943
rect 17175 14909 17184 14943
rect 17132 14900 17184 14909
rect 8852 14807 8904 14816
rect 8852 14773 8861 14807
rect 8861 14773 8895 14807
rect 8895 14773 8904 14807
rect 8852 14764 8904 14773
rect 11060 14832 11112 14884
rect 16396 14832 16448 14884
rect 16488 14832 16540 14884
rect 18420 14832 18472 14884
rect 22836 14900 22888 14952
rect 24676 14943 24728 14952
rect 24676 14909 24685 14943
rect 24685 14909 24719 14943
rect 24719 14909 24728 14943
rect 24676 14900 24728 14909
rect 15936 14764 15988 14816
rect 20352 14807 20404 14816
rect 20352 14773 20361 14807
rect 20361 14773 20395 14807
rect 20395 14773 20404 14807
rect 20352 14764 20404 14773
rect 21272 14807 21324 14816
rect 21272 14773 21281 14807
rect 21281 14773 21315 14807
rect 21315 14773 21324 14807
rect 21272 14764 21324 14773
rect 2950 14662 3002 14714
rect 3014 14662 3066 14714
rect 3078 14662 3130 14714
rect 3142 14662 3194 14714
rect 3206 14662 3258 14714
rect 12950 14662 13002 14714
rect 13014 14662 13066 14714
rect 13078 14662 13130 14714
rect 13142 14662 13194 14714
rect 13206 14662 13258 14714
rect 22950 14662 23002 14714
rect 23014 14662 23066 14714
rect 23078 14662 23130 14714
rect 23142 14662 23194 14714
rect 23206 14662 23258 14714
rect 9588 14560 9640 14612
rect 10508 14603 10560 14612
rect 10508 14569 10517 14603
rect 10517 14569 10551 14603
rect 10551 14569 10560 14603
rect 10508 14560 10560 14569
rect 11336 14560 11388 14612
rect 11612 14560 11664 14612
rect 16120 14560 16172 14612
rect 18052 14560 18104 14612
rect 19156 14560 19208 14612
rect 8852 14424 8904 14476
rect 9036 14424 9088 14476
rect 9864 14467 9916 14476
rect 9864 14433 9873 14467
rect 9873 14433 9907 14467
rect 9907 14433 9916 14467
rect 9864 14424 9916 14433
rect 10968 14424 11020 14476
rect 6920 14356 6972 14408
rect 7196 14356 7248 14408
rect 8576 14399 8628 14408
rect 8576 14365 8585 14399
rect 8585 14365 8619 14399
rect 8619 14365 8628 14399
rect 8576 14356 8628 14365
rect 12256 14399 12308 14408
rect 12256 14365 12265 14399
rect 12265 14365 12299 14399
rect 12299 14365 12308 14399
rect 12256 14356 12308 14365
rect 11244 14288 11296 14340
rect 13176 14424 13228 14476
rect 15108 14492 15160 14544
rect 13360 14467 13412 14476
rect 13360 14433 13369 14467
rect 13369 14433 13403 14467
rect 13403 14433 13412 14467
rect 13360 14424 13412 14433
rect 14004 14288 14056 14340
rect 15108 14288 15160 14340
rect 6920 14220 6972 14272
rect 9036 14220 9088 14272
rect 13084 14220 13136 14272
rect 14740 14220 14792 14272
rect 19800 14424 19852 14476
rect 16856 14356 16908 14408
rect 17500 14399 17552 14408
rect 17500 14365 17509 14399
rect 17509 14365 17543 14399
rect 17543 14365 17552 14399
rect 17500 14356 17552 14365
rect 18052 14399 18104 14408
rect 18052 14365 18061 14399
rect 18061 14365 18095 14399
rect 18095 14365 18104 14399
rect 18052 14356 18104 14365
rect 21456 14356 21508 14408
rect 16488 14331 16540 14340
rect 16488 14297 16497 14331
rect 16497 14297 16531 14331
rect 16531 14297 16540 14331
rect 16488 14288 16540 14297
rect 18972 14288 19024 14340
rect 21732 14288 21784 14340
rect 22928 14288 22980 14340
rect 16580 14220 16632 14272
rect 17316 14263 17368 14272
rect 17316 14229 17325 14263
rect 17325 14229 17359 14263
rect 17359 14229 17368 14263
rect 17316 14220 17368 14229
rect 17592 14220 17644 14272
rect 22560 14220 22612 14272
rect 7950 14118 8002 14170
rect 8014 14118 8066 14170
rect 8078 14118 8130 14170
rect 8142 14118 8194 14170
rect 8206 14118 8258 14170
rect 17950 14118 18002 14170
rect 18014 14118 18066 14170
rect 18078 14118 18130 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 7196 14016 7248 14068
rect 8484 14059 8536 14068
rect 8484 14025 8493 14059
rect 8493 14025 8527 14059
rect 8527 14025 8536 14059
rect 8484 14016 8536 14025
rect 10784 14016 10836 14068
rect 10968 13948 11020 14000
rect 11244 13991 11296 14000
rect 11244 13957 11253 13991
rect 11253 13957 11287 13991
rect 11287 13957 11296 13991
rect 11244 13948 11296 13957
rect 12716 14059 12768 14068
rect 12716 14025 12725 14059
rect 12725 14025 12759 14059
rect 12759 14025 12768 14059
rect 12716 14016 12768 14025
rect 13084 14059 13136 14068
rect 13084 14025 13093 14059
rect 13093 14025 13127 14059
rect 13127 14025 13136 14059
rect 13084 14016 13136 14025
rect 13176 14059 13228 14068
rect 13176 14025 13185 14059
rect 13185 14025 13219 14059
rect 13219 14025 13228 14059
rect 13176 14016 13228 14025
rect 17040 14016 17092 14068
rect 18604 14059 18656 14068
rect 18604 14025 18613 14059
rect 18613 14025 18647 14059
rect 18647 14025 18656 14059
rect 18604 14016 18656 14025
rect 20996 14059 21048 14068
rect 20996 14025 21005 14059
rect 21005 14025 21039 14059
rect 21039 14025 21048 14059
rect 20996 14016 21048 14025
rect 21916 14016 21968 14068
rect 22744 14016 22796 14068
rect 16028 13991 16080 14000
rect 16028 13957 16037 13991
rect 16037 13957 16071 13991
rect 16071 13957 16080 13991
rect 16028 13948 16080 13957
rect 16304 13948 16356 14000
rect 16580 13948 16632 14000
rect 17592 13948 17644 14000
rect 19708 13948 19760 14000
rect 22836 13948 22888 14000
rect 25136 13991 25188 14000
rect 25136 13957 25145 13991
rect 25145 13957 25179 13991
rect 25179 13957 25188 13991
rect 25136 13948 25188 13957
rect 2780 13923 2832 13932
rect 2780 13889 2789 13923
rect 2789 13889 2823 13923
rect 2823 13889 2832 13923
rect 2780 13880 2832 13889
rect 1768 13855 1820 13864
rect 1768 13821 1777 13855
rect 1777 13821 1811 13855
rect 1811 13821 1820 13855
rect 1768 13812 1820 13821
rect 6828 13812 6880 13864
rect 8576 13812 8628 13864
rect 6920 13744 6972 13796
rect 7840 13744 7892 13796
rect 12164 13812 12216 13864
rect 13176 13812 13228 13864
rect 12532 13744 12584 13796
rect 15752 13812 15804 13864
rect 21824 13880 21876 13932
rect 22008 13923 22060 13932
rect 22008 13889 22017 13923
rect 22017 13889 22051 13923
rect 22051 13889 22060 13923
rect 22008 13880 22060 13889
rect 15936 13812 15988 13864
rect 16856 13855 16908 13864
rect 16856 13821 16865 13855
rect 16865 13821 16899 13855
rect 16899 13821 16908 13855
rect 16856 13812 16908 13821
rect 17132 13855 17184 13864
rect 17132 13821 17141 13855
rect 17141 13821 17175 13855
rect 17175 13821 17184 13855
rect 17132 13812 17184 13821
rect 19064 13855 19116 13864
rect 19064 13821 19073 13855
rect 19073 13821 19107 13855
rect 19107 13821 19116 13855
rect 19064 13812 19116 13821
rect 14464 13744 14516 13796
rect 21364 13812 21416 13864
rect 22928 13880 22980 13932
rect 20904 13744 20956 13796
rect 23388 13812 23440 13864
rect 16028 13676 16080 13728
rect 17868 13676 17920 13728
rect 21364 13676 21416 13728
rect 21732 13676 21784 13728
rect 2950 13574 3002 13626
rect 3014 13574 3066 13626
rect 3078 13574 3130 13626
rect 3142 13574 3194 13626
rect 3206 13574 3258 13626
rect 12950 13574 13002 13626
rect 13014 13574 13066 13626
rect 13078 13574 13130 13626
rect 13142 13574 13194 13626
rect 13206 13574 13258 13626
rect 22950 13574 23002 13626
rect 23014 13574 23066 13626
rect 23078 13574 23130 13626
rect 23142 13574 23194 13626
rect 23206 13574 23258 13626
rect 8484 13472 8536 13524
rect 12440 13472 12492 13524
rect 13544 13472 13596 13524
rect 14188 13515 14240 13524
rect 14188 13481 14197 13515
rect 14197 13481 14231 13515
rect 14231 13481 14240 13515
rect 14188 13472 14240 13481
rect 14740 13472 14792 13524
rect 14556 13404 14608 13456
rect 7104 13379 7156 13388
rect 7104 13345 7113 13379
rect 7113 13345 7147 13379
rect 7147 13345 7156 13379
rect 7104 13336 7156 13345
rect 7656 13336 7708 13388
rect 12440 13336 12492 13388
rect 6828 13311 6880 13320
rect 6828 13277 6837 13311
rect 6837 13277 6871 13311
rect 6871 13277 6880 13311
rect 6828 13268 6880 13277
rect 8484 13200 8536 13252
rect 9036 13200 9088 13252
rect 8576 13175 8628 13184
rect 8576 13141 8585 13175
rect 8585 13141 8619 13175
rect 8619 13141 8628 13175
rect 8576 13132 8628 13141
rect 14096 13336 14148 13388
rect 15568 13472 15620 13524
rect 21088 13472 21140 13524
rect 18604 13404 18656 13456
rect 19340 13447 19392 13456
rect 19340 13413 19349 13447
rect 19349 13413 19383 13447
rect 19383 13413 19392 13447
rect 19340 13404 19392 13413
rect 21180 13404 21232 13456
rect 18420 13379 18472 13388
rect 18420 13345 18429 13379
rect 18429 13345 18463 13379
rect 18463 13345 18472 13379
rect 18420 13336 18472 13345
rect 21548 13336 21600 13388
rect 22836 13336 22888 13388
rect 19064 13268 19116 13320
rect 19616 13268 19668 13320
rect 19340 13200 19392 13252
rect 15016 13175 15068 13184
rect 15016 13141 15025 13175
rect 15025 13141 15059 13175
rect 15059 13141 15068 13175
rect 15016 13132 15068 13141
rect 17224 13132 17276 13184
rect 18512 13132 18564 13184
rect 20904 13132 20956 13184
rect 23296 13268 23348 13320
rect 21364 13132 21416 13184
rect 21640 13132 21692 13184
rect 23848 13175 23900 13184
rect 23848 13141 23857 13175
rect 23857 13141 23891 13175
rect 23891 13141 23900 13175
rect 23848 13132 23900 13141
rect 7950 13030 8002 13082
rect 8014 13030 8066 13082
rect 8078 13030 8130 13082
rect 8142 13030 8194 13082
rect 8206 13030 8258 13082
rect 17950 13030 18002 13082
rect 18014 13030 18066 13082
rect 18078 13030 18130 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 8300 12928 8352 12980
rect 11796 12971 11848 12980
rect 11796 12937 11805 12971
rect 11805 12937 11839 12971
rect 11839 12937 11848 12971
rect 11796 12928 11848 12937
rect 12808 12928 12860 12980
rect 13452 12928 13504 12980
rect 7564 12860 7616 12912
rect 8484 12860 8536 12912
rect 9588 12860 9640 12912
rect 14004 12860 14056 12912
rect 7288 12792 7340 12844
rect 13452 12792 13504 12844
rect 13544 12835 13596 12844
rect 13544 12801 13553 12835
rect 13553 12801 13587 12835
rect 13587 12801 13596 12835
rect 13544 12792 13596 12801
rect 16856 12928 16908 12980
rect 17040 12928 17092 12980
rect 17224 12971 17276 12980
rect 17224 12937 17233 12971
rect 17233 12937 17267 12971
rect 17267 12937 17276 12971
rect 17224 12928 17276 12937
rect 14464 12903 14516 12912
rect 14464 12869 14473 12903
rect 14473 12869 14507 12903
rect 14507 12869 14516 12903
rect 14464 12860 14516 12869
rect 16304 12903 16356 12912
rect 16304 12869 16313 12903
rect 16313 12869 16347 12903
rect 16347 12869 16356 12903
rect 16304 12860 16356 12869
rect 21364 12928 21416 12980
rect 20904 12860 20956 12912
rect 24860 12860 24912 12912
rect 8576 12724 8628 12776
rect 8852 12724 8904 12776
rect 11336 12724 11388 12776
rect 14096 12724 14148 12776
rect 15660 12724 15712 12776
rect 18420 12835 18472 12844
rect 18420 12801 18429 12835
rect 18429 12801 18463 12835
rect 18463 12801 18472 12835
rect 18420 12792 18472 12801
rect 22100 12835 22152 12844
rect 22100 12801 22109 12835
rect 22109 12801 22143 12835
rect 22143 12801 22152 12835
rect 22100 12792 22152 12801
rect 23940 12835 23992 12844
rect 23940 12801 23949 12835
rect 23949 12801 23983 12835
rect 23983 12801 23992 12835
rect 23940 12792 23992 12801
rect 16488 12724 16540 12776
rect 19432 12724 19484 12776
rect 21456 12767 21508 12776
rect 21456 12733 21465 12767
rect 21465 12733 21499 12767
rect 21499 12733 21508 12767
rect 21456 12724 21508 12733
rect 24768 12767 24820 12776
rect 24768 12733 24777 12767
rect 24777 12733 24811 12767
rect 24811 12733 24820 12767
rect 24768 12724 24820 12733
rect 10968 12588 11020 12640
rect 14280 12588 14332 12640
rect 19524 12588 19576 12640
rect 19708 12588 19760 12640
rect 2950 12486 3002 12538
rect 3014 12486 3066 12538
rect 3078 12486 3130 12538
rect 3142 12486 3194 12538
rect 3206 12486 3258 12538
rect 12950 12486 13002 12538
rect 13014 12486 13066 12538
rect 13078 12486 13130 12538
rect 13142 12486 13194 12538
rect 13206 12486 13258 12538
rect 22950 12486 23002 12538
rect 23014 12486 23066 12538
rect 23078 12486 23130 12538
rect 23142 12486 23194 12538
rect 23206 12486 23258 12538
rect 12440 12384 12492 12436
rect 13452 12384 13504 12436
rect 14464 12384 14516 12436
rect 15568 12384 15620 12436
rect 3332 12316 3384 12368
rect 6736 12316 6788 12368
rect 10968 12316 11020 12368
rect 11244 12248 11296 12300
rect 15108 12248 15160 12300
rect 12808 12223 12860 12232
rect 12808 12189 12817 12223
rect 12817 12189 12851 12223
rect 12851 12189 12860 12223
rect 12808 12180 12860 12189
rect 15200 12180 15252 12232
rect 15384 12180 15436 12232
rect 17132 12427 17184 12436
rect 17132 12393 17141 12427
rect 17141 12393 17175 12427
rect 17175 12393 17184 12427
rect 17132 12384 17184 12393
rect 19984 12359 20036 12368
rect 19984 12325 19993 12359
rect 19993 12325 20027 12359
rect 20027 12325 20036 12359
rect 19984 12316 20036 12325
rect 16856 12248 16908 12300
rect 8852 12112 8904 12164
rect 9680 12112 9732 12164
rect 12624 12112 12676 12164
rect 13452 12112 13504 12164
rect 14188 12112 14240 12164
rect 11980 12044 12032 12096
rect 12716 12044 12768 12096
rect 14740 12087 14792 12096
rect 14740 12053 14749 12087
rect 14749 12053 14783 12087
rect 14783 12053 14792 12087
rect 14740 12044 14792 12053
rect 15660 12087 15712 12096
rect 15660 12053 15669 12087
rect 15669 12053 15703 12087
rect 15703 12053 15712 12087
rect 15660 12044 15712 12053
rect 22100 12384 22152 12436
rect 22652 12223 22704 12232
rect 22652 12189 22661 12223
rect 22661 12189 22695 12223
rect 22695 12189 22704 12223
rect 22652 12180 22704 12189
rect 22744 12180 22796 12232
rect 19248 12112 19300 12164
rect 24952 12112 25004 12164
rect 19064 12044 19116 12096
rect 19432 12044 19484 12096
rect 21364 12044 21416 12096
rect 24584 12087 24636 12096
rect 24584 12053 24593 12087
rect 24593 12053 24627 12087
rect 24627 12053 24636 12087
rect 24584 12044 24636 12053
rect 7950 11942 8002 11994
rect 8014 11942 8066 11994
rect 8078 11942 8130 11994
rect 8142 11942 8194 11994
rect 8206 11942 8258 11994
rect 17950 11942 18002 11994
rect 18014 11942 18066 11994
rect 18078 11942 18130 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 11980 11772 12032 11824
rect 13820 11840 13872 11892
rect 14372 11883 14424 11892
rect 14372 11849 14381 11883
rect 14381 11849 14415 11883
rect 14415 11849 14424 11883
rect 14372 11840 14424 11849
rect 14924 11883 14976 11892
rect 14924 11849 14933 11883
rect 14933 11849 14967 11883
rect 14967 11849 14976 11883
rect 14924 11840 14976 11849
rect 15384 11840 15436 11892
rect 18420 11840 18472 11892
rect 14464 11772 14516 11824
rect 17316 11772 17368 11824
rect 19340 11772 19392 11824
rect 22652 11883 22704 11892
rect 22652 11849 22661 11883
rect 22661 11849 22695 11883
rect 22695 11849 22704 11883
rect 22652 11840 22704 11849
rect 19616 11747 19668 11756
rect 19616 11713 19625 11747
rect 19625 11713 19659 11747
rect 19659 11713 19668 11747
rect 19616 11704 19668 11713
rect 22468 11747 22520 11756
rect 22468 11713 22477 11747
rect 22477 11713 22511 11747
rect 22511 11713 22520 11747
rect 22468 11704 22520 11713
rect 23664 11704 23716 11756
rect 11244 11636 11296 11688
rect 12256 11636 12308 11688
rect 13360 11636 13412 11688
rect 15384 11679 15436 11688
rect 15384 11645 15393 11679
rect 15393 11645 15427 11679
rect 15427 11645 15436 11679
rect 15384 11636 15436 11645
rect 15476 11679 15528 11688
rect 15476 11645 15485 11679
rect 15485 11645 15519 11679
rect 15519 11645 15528 11679
rect 15476 11636 15528 11645
rect 15568 11636 15620 11688
rect 24676 11679 24728 11688
rect 24676 11645 24685 11679
rect 24685 11645 24719 11679
rect 24719 11645 24728 11679
rect 24676 11636 24728 11645
rect 15844 11568 15896 11620
rect 19984 11568 20036 11620
rect 20352 11568 20404 11620
rect 23480 11568 23532 11620
rect 19064 11543 19116 11552
rect 19064 11509 19073 11543
rect 19073 11509 19107 11543
rect 19107 11509 19116 11543
rect 19064 11500 19116 11509
rect 23940 11500 23992 11552
rect 2950 11398 3002 11450
rect 3014 11398 3066 11450
rect 3078 11398 3130 11450
rect 3142 11398 3194 11450
rect 3206 11398 3258 11450
rect 12950 11398 13002 11450
rect 13014 11398 13066 11450
rect 13078 11398 13130 11450
rect 13142 11398 13194 11450
rect 13206 11398 13258 11450
rect 22950 11398 23002 11450
rect 23014 11398 23066 11450
rect 23078 11398 23130 11450
rect 23142 11398 23194 11450
rect 23206 11398 23258 11450
rect 11980 11296 12032 11348
rect 14004 11296 14056 11348
rect 22468 11296 22520 11348
rect 13452 11228 13504 11280
rect 11244 11203 11296 11212
rect 11244 11169 11253 11203
rect 11253 11169 11287 11203
rect 11287 11169 11296 11203
rect 11244 11160 11296 11169
rect 12532 11160 12584 11212
rect 13360 11160 13412 11212
rect 14556 11203 14608 11212
rect 14556 11169 14565 11203
rect 14565 11169 14599 11203
rect 14599 11169 14608 11203
rect 14556 11160 14608 11169
rect 15108 11160 15160 11212
rect 15568 11092 15620 11144
rect 15844 11135 15896 11144
rect 15844 11101 15853 11135
rect 15853 11101 15887 11135
rect 15887 11101 15896 11135
rect 15844 11092 15896 11101
rect 22008 11228 22060 11280
rect 22836 11228 22888 11280
rect 19248 11160 19300 11212
rect 19708 11203 19760 11212
rect 19708 11169 19717 11203
rect 19717 11169 19751 11203
rect 19751 11169 19760 11203
rect 19708 11160 19760 11169
rect 22560 11160 22612 11212
rect 21916 11092 21968 11144
rect 23388 11092 23440 11144
rect 11980 11024 12032 11076
rect 24216 11024 24268 11076
rect 16028 10956 16080 11008
rect 24032 10999 24084 11008
rect 24032 10965 24041 10999
rect 24041 10965 24075 10999
rect 24075 10965 24084 10999
rect 24032 10956 24084 10965
rect 7950 10854 8002 10906
rect 8014 10854 8066 10906
rect 8078 10854 8130 10906
rect 8142 10854 8194 10906
rect 8206 10854 8258 10906
rect 17950 10854 18002 10906
rect 18014 10854 18066 10906
rect 18078 10854 18130 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 13820 10752 13872 10804
rect 15844 10752 15896 10804
rect 16212 10752 16264 10804
rect 19248 10752 19300 10804
rect 19524 10727 19576 10736
rect 19524 10693 19533 10727
rect 19533 10693 19567 10727
rect 19567 10693 19576 10727
rect 19524 10684 19576 10693
rect 21088 10659 21140 10668
rect 21088 10625 21097 10659
rect 21097 10625 21131 10659
rect 21131 10625 21140 10659
rect 21088 10616 21140 10625
rect 23940 10659 23992 10668
rect 23940 10625 23949 10659
rect 23949 10625 23983 10659
rect 23983 10625 23992 10659
rect 23940 10616 23992 10625
rect 19064 10548 19116 10600
rect 21456 10548 21508 10600
rect 24768 10591 24820 10600
rect 24768 10557 24777 10591
rect 24777 10557 24811 10591
rect 24811 10557 24820 10591
rect 24768 10548 24820 10557
rect 21364 10480 21416 10532
rect 16028 10412 16080 10464
rect 24308 10412 24360 10464
rect 2950 10310 3002 10362
rect 3014 10310 3066 10362
rect 3078 10310 3130 10362
rect 3142 10310 3194 10362
rect 3206 10310 3258 10362
rect 12950 10310 13002 10362
rect 13014 10310 13066 10362
rect 13078 10310 13130 10362
rect 13142 10310 13194 10362
rect 13206 10310 13258 10362
rect 22950 10310 23002 10362
rect 23014 10310 23066 10362
rect 23078 10310 23130 10362
rect 23142 10310 23194 10362
rect 23206 10310 23258 10362
rect 24860 10072 24912 10124
rect 9404 10004 9456 10056
rect 19892 10004 19944 10056
rect 24584 10004 24636 10056
rect 12348 9936 12400 9988
rect 16488 9936 16540 9988
rect 23848 9936 23900 9988
rect 24124 9868 24176 9920
rect 7950 9766 8002 9818
rect 8014 9766 8066 9818
rect 8078 9766 8130 9818
rect 8142 9766 8194 9818
rect 8206 9766 8258 9818
rect 17950 9766 18002 9818
rect 18014 9766 18066 9818
rect 18078 9766 18130 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 2872 9596 2924 9648
rect 5632 9596 5684 9648
rect 5724 9596 5776 9648
rect 13544 9596 13596 9648
rect 22008 9571 22060 9580
rect 22008 9537 22017 9571
rect 22017 9537 22051 9571
rect 22051 9537 22060 9571
rect 22008 9528 22060 9537
rect 23940 9571 23992 9580
rect 23940 9537 23949 9571
rect 23949 9537 23983 9571
rect 23983 9537 23992 9571
rect 23940 9528 23992 9537
rect 24768 9503 24820 9512
rect 24768 9469 24777 9503
rect 24777 9469 24811 9503
rect 24811 9469 24820 9503
rect 24768 9460 24820 9469
rect 7104 9392 7156 9444
rect 7288 9435 7340 9444
rect 7288 9401 7297 9435
rect 7297 9401 7331 9435
rect 7331 9401 7340 9435
rect 7288 9392 7340 9401
rect 15200 9392 15252 9444
rect 24492 9324 24544 9376
rect 2950 9222 3002 9274
rect 3014 9222 3066 9274
rect 3078 9222 3130 9274
rect 3142 9222 3194 9274
rect 3206 9222 3258 9274
rect 12950 9222 13002 9274
rect 13014 9222 13066 9274
rect 13078 9222 13130 9274
rect 13142 9222 13194 9274
rect 13206 9222 13258 9274
rect 22950 9222 23002 9274
rect 23014 9222 23066 9274
rect 23078 9222 23130 9274
rect 23142 9222 23194 9274
rect 23206 9222 23258 9274
rect 15936 8916 15988 8968
rect 18604 8916 18656 8968
rect 22836 8916 22888 8968
rect 24860 8959 24912 8968
rect 24860 8925 24869 8959
rect 24869 8925 24903 8959
rect 24903 8925 24912 8959
rect 24860 8916 24912 8925
rect 25044 8916 25096 8968
rect 17776 8848 17828 8900
rect 20720 8848 20772 8900
rect 22744 8848 22796 8900
rect 25504 8848 25556 8900
rect 23296 8823 23348 8832
rect 23296 8789 23305 8823
rect 23305 8789 23339 8823
rect 23339 8789 23348 8823
rect 23296 8780 23348 8789
rect 24676 8823 24728 8832
rect 24676 8789 24685 8823
rect 24685 8789 24719 8823
rect 24719 8789 24728 8823
rect 24676 8780 24728 8789
rect 25228 8823 25280 8832
rect 25228 8789 25237 8823
rect 25237 8789 25271 8823
rect 25271 8789 25280 8823
rect 25228 8780 25280 8789
rect 7950 8678 8002 8730
rect 8014 8678 8066 8730
rect 8078 8678 8130 8730
rect 8142 8678 8194 8730
rect 8206 8678 8258 8730
rect 17950 8678 18002 8730
rect 18014 8678 18066 8730
rect 18078 8678 18130 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 6828 8576 6880 8628
rect 12624 8508 12676 8560
rect 7564 8440 7616 8492
rect 24676 8508 24728 8560
rect 25136 8551 25188 8560
rect 25136 8517 25145 8551
rect 25145 8517 25179 8551
rect 25179 8517 25188 8551
rect 25136 8508 25188 8517
rect 24032 8483 24084 8492
rect 24032 8449 24041 8483
rect 24041 8449 24075 8483
rect 24075 8449 24084 8483
rect 24032 8440 24084 8449
rect 2780 8372 2832 8424
rect 24584 8372 24636 8424
rect 2950 8134 3002 8186
rect 3014 8134 3066 8186
rect 3078 8134 3130 8186
rect 3142 8134 3194 8186
rect 3206 8134 3258 8186
rect 12950 8134 13002 8186
rect 13014 8134 13066 8186
rect 13078 8134 13130 8186
rect 13142 8134 13194 8186
rect 13206 8134 13258 8186
rect 22950 8134 23002 8186
rect 23014 8134 23066 8186
rect 23078 8134 23130 8186
rect 23142 8134 23194 8186
rect 23206 8134 23258 8186
rect 24952 7896 25004 7948
rect 18788 7828 18840 7880
rect 21272 7828 21324 7880
rect 24216 7828 24268 7880
rect 24308 7828 24360 7880
rect 20260 7760 20312 7812
rect 21088 7760 21140 7812
rect 24676 7735 24728 7744
rect 24676 7701 24685 7735
rect 24685 7701 24719 7735
rect 24719 7701 24728 7735
rect 24676 7692 24728 7701
rect 7950 7590 8002 7642
rect 8014 7590 8066 7642
rect 8078 7590 8130 7642
rect 8142 7590 8194 7642
rect 8206 7590 8258 7642
rect 17950 7590 18002 7642
rect 18014 7590 18066 7642
rect 18078 7590 18130 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 22744 7420 22796 7472
rect 21548 7352 21600 7404
rect 24124 7395 24176 7404
rect 24124 7361 24133 7395
rect 24133 7361 24167 7395
rect 24167 7361 24176 7395
rect 24124 7352 24176 7361
rect 20996 7327 21048 7336
rect 20996 7293 21005 7327
rect 21005 7293 21039 7327
rect 21039 7293 21048 7327
rect 20996 7284 21048 7293
rect 22468 7284 22520 7336
rect 24768 7327 24820 7336
rect 24768 7293 24777 7327
rect 24777 7293 24811 7327
rect 24811 7293 24820 7327
rect 24768 7284 24820 7293
rect 2950 7046 3002 7098
rect 3014 7046 3066 7098
rect 3078 7046 3130 7098
rect 3142 7046 3194 7098
rect 3206 7046 3258 7098
rect 12950 7046 13002 7098
rect 13014 7046 13066 7098
rect 13078 7046 13130 7098
rect 13142 7046 13194 7098
rect 13206 7046 13258 7098
rect 22950 7046 23002 7098
rect 23014 7046 23066 7098
rect 23078 7046 23130 7098
rect 23142 7046 23194 7098
rect 23206 7046 23258 7098
rect 24860 6808 24912 6860
rect 15292 6740 15344 6792
rect 19800 6740 19852 6792
rect 3424 6672 3476 6724
rect 7012 6672 7064 6724
rect 19708 6672 19760 6724
rect 3148 6604 3200 6656
rect 6276 6604 6328 6656
rect 22008 6715 22060 6724
rect 22008 6681 22017 6715
rect 22017 6681 22051 6715
rect 22051 6681 22060 6715
rect 22008 6672 22060 6681
rect 24492 6740 24544 6792
rect 7950 6502 8002 6554
rect 8014 6502 8066 6554
rect 8078 6502 8130 6554
rect 8142 6502 8194 6554
rect 8206 6502 8258 6554
rect 17950 6502 18002 6554
rect 18014 6502 18066 6554
rect 18078 6502 18130 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 21548 6400 21600 6452
rect 11980 6332 12032 6384
rect 17316 6264 17368 6316
rect 23388 6332 23440 6384
rect 20168 6264 20220 6316
rect 23296 6264 23348 6316
rect 24768 6239 24820 6248
rect 24768 6205 24777 6239
rect 24777 6205 24811 6239
rect 24811 6205 24820 6239
rect 24768 6196 24820 6205
rect 22100 6128 22152 6180
rect 16212 6060 16264 6112
rect 23940 6060 23992 6112
rect 2950 5958 3002 6010
rect 3014 5958 3066 6010
rect 3078 5958 3130 6010
rect 3142 5958 3194 6010
rect 3206 5958 3258 6010
rect 12950 5958 13002 6010
rect 13014 5958 13066 6010
rect 13078 5958 13130 6010
rect 13142 5958 13194 6010
rect 13206 5958 13258 6010
rect 22950 5958 23002 6010
rect 23014 5958 23066 6010
rect 23078 5958 23130 6010
rect 23142 5958 23194 6010
rect 23206 5958 23258 6010
rect 20168 5899 20220 5908
rect 20168 5865 20177 5899
rect 20177 5865 20211 5899
rect 20211 5865 20220 5899
rect 20168 5856 20220 5865
rect 20260 5788 20312 5840
rect 10876 5720 10928 5772
rect 15844 5720 15896 5772
rect 18880 5720 18932 5772
rect 19340 5720 19392 5772
rect 20628 5720 20680 5772
rect 19984 5695 20036 5704
rect 19984 5661 19993 5695
rect 19993 5661 20027 5695
rect 20027 5661 20036 5695
rect 19984 5652 20036 5661
rect 20720 5695 20772 5704
rect 20720 5661 20729 5695
rect 20729 5661 20763 5695
rect 20763 5661 20772 5695
rect 20720 5652 20772 5661
rect 21916 5584 21968 5636
rect 7564 5516 7616 5568
rect 13912 5516 13964 5568
rect 7950 5414 8002 5466
rect 8014 5414 8066 5466
rect 8078 5414 8130 5466
rect 8142 5414 8194 5466
rect 8206 5414 8258 5466
rect 17950 5414 18002 5466
rect 18014 5414 18066 5466
rect 18078 5414 18130 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 15752 5312 15804 5364
rect 16856 5312 16908 5364
rect 16212 5287 16264 5296
rect 16212 5253 16221 5287
rect 16221 5253 16255 5287
rect 16255 5253 16264 5287
rect 16212 5244 16264 5253
rect 16028 5219 16080 5228
rect 16028 5185 16037 5219
rect 16037 5185 16071 5219
rect 16071 5185 16080 5219
rect 16028 5176 16080 5185
rect 19800 5244 19852 5296
rect 19432 5176 19484 5228
rect 19708 5176 19760 5228
rect 24676 5176 24728 5228
rect 19524 5108 19576 5160
rect 22284 5108 22336 5160
rect 24768 5151 24820 5160
rect 24768 5117 24777 5151
rect 24777 5117 24811 5151
rect 24811 5117 24820 5151
rect 24768 5108 24820 5117
rect 20536 5040 20588 5092
rect 16948 4972 17000 5024
rect 18696 4972 18748 5024
rect 2950 4870 3002 4922
rect 3014 4870 3066 4922
rect 3078 4870 3130 4922
rect 3142 4870 3194 4922
rect 3206 4870 3258 4922
rect 12950 4870 13002 4922
rect 13014 4870 13066 4922
rect 13078 4870 13130 4922
rect 13142 4870 13194 4922
rect 13206 4870 13258 4922
rect 22950 4870 23002 4922
rect 23014 4870 23066 4922
rect 23078 4870 23130 4922
rect 23142 4870 23194 4922
rect 23206 4870 23258 4922
rect 3240 4768 3292 4820
rect 6368 4768 6420 4820
rect 25320 4811 25372 4820
rect 25320 4777 25329 4811
rect 25329 4777 25363 4811
rect 25363 4777 25372 4811
rect 25320 4768 25372 4777
rect 5172 4700 5224 4752
rect 10324 4700 10376 4752
rect 19892 4675 19944 4684
rect 19892 4641 19901 4675
rect 19901 4641 19935 4675
rect 19935 4641 19944 4675
rect 19892 4632 19944 4641
rect 21732 4675 21784 4684
rect 21732 4641 21741 4675
rect 21741 4641 21775 4675
rect 21775 4641 21784 4675
rect 21732 4632 21784 4641
rect 16396 4564 16448 4616
rect 19340 4564 19392 4616
rect 21180 4564 21232 4616
rect 18328 4539 18380 4548
rect 18328 4505 18337 4539
rect 18337 4505 18371 4539
rect 18371 4505 18380 4539
rect 18328 4496 18380 4505
rect 1400 4471 1452 4480
rect 1400 4437 1409 4471
rect 1409 4437 1443 4471
rect 1443 4437 1452 4471
rect 1400 4428 1452 4437
rect 7950 4326 8002 4378
rect 8014 4326 8066 4378
rect 8078 4326 8130 4378
rect 8142 4326 8194 4378
rect 8206 4326 8258 4378
rect 17950 4326 18002 4378
rect 18014 4326 18066 4378
rect 18078 4326 18130 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 8392 4224 8444 4276
rect 10048 4224 10100 4276
rect 5080 4156 5132 4208
rect 8944 4156 8996 4208
rect 13728 4156 13780 4208
rect 14648 4156 14700 4208
rect 21824 4156 21876 4208
rect 1124 4088 1176 4140
rect 1400 4088 1452 4140
rect 5724 3952 5776 4004
rect 7840 3952 7892 4004
rect 2688 3884 2740 3936
rect 2872 3927 2924 3936
rect 2872 3893 2881 3927
rect 2881 3893 2915 3927
rect 2915 3893 2924 3927
rect 2872 3884 2924 3893
rect 3332 3884 3384 3936
rect 5540 3927 5592 3936
rect 5540 3893 5549 3927
rect 5549 3893 5583 3927
rect 5583 3893 5592 3927
rect 5540 3884 5592 3893
rect 9220 4088 9272 4140
rect 12716 4088 12768 4140
rect 15200 4088 15252 4140
rect 18604 4088 18656 4140
rect 23480 4088 23532 4140
rect 12808 4020 12860 4072
rect 16212 4020 16264 4072
rect 18420 4020 18472 4072
rect 20260 4020 20312 4072
rect 12072 3952 12124 4004
rect 21364 3952 21416 4004
rect 8760 3884 8812 3936
rect 10968 3884 11020 3936
rect 11796 3884 11848 3936
rect 20996 3884 21048 3936
rect 25320 3884 25372 3936
rect 2950 3782 3002 3834
rect 3014 3782 3066 3834
rect 3078 3782 3130 3834
rect 3142 3782 3194 3834
rect 3206 3782 3258 3834
rect 12950 3782 13002 3834
rect 13014 3782 13066 3834
rect 13078 3782 13130 3834
rect 13142 3782 13194 3834
rect 13206 3782 13258 3834
rect 22950 3782 23002 3834
rect 23014 3782 23066 3834
rect 23078 3782 23130 3834
rect 23142 3782 23194 3834
rect 23206 3782 23258 3834
rect 2780 3680 2832 3732
rect 3424 3680 3476 3732
rect 5080 3723 5132 3732
rect 5080 3689 5089 3723
rect 5089 3689 5123 3723
rect 5123 3689 5132 3723
rect 5080 3680 5132 3689
rect 6644 3680 6696 3732
rect 7748 3680 7800 3732
rect 8392 3723 8444 3732
rect 8392 3689 8401 3723
rect 8401 3689 8435 3723
rect 8435 3689 8444 3723
rect 8392 3680 8444 3689
rect 13636 3680 13688 3732
rect 25228 3723 25280 3732
rect 25228 3689 25237 3723
rect 25237 3689 25271 3723
rect 25271 3689 25280 3723
rect 25228 3680 25280 3689
rect 4896 3612 4948 3664
rect 16028 3612 16080 3664
rect 19800 3612 19852 3664
rect 2780 3476 2832 3528
rect 2872 3476 2924 3528
rect 1492 3408 1544 3460
rect 5540 3476 5592 3528
rect 6276 3476 6328 3528
rect 7840 3476 7892 3528
rect 9588 3519 9640 3528
rect 9588 3485 9597 3519
rect 9597 3485 9631 3519
rect 9631 3485 9640 3519
rect 9588 3476 9640 3485
rect 9956 3476 10008 3528
rect 10692 3476 10744 3528
rect 13728 3519 13780 3528
rect 13728 3485 13737 3519
rect 13737 3485 13771 3519
rect 13771 3485 13780 3519
rect 13728 3476 13780 3485
rect 12532 3451 12584 3460
rect 12532 3417 12541 3451
rect 12541 3417 12575 3451
rect 12575 3417 12584 3451
rect 12532 3408 12584 3417
rect 14004 3544 14056 3596
rect 15476 3544 15528 3596
rect 17684 3544 17736 3596
rect 14280 3519 14332 3528
rect 14280 3485 14289 3519
rect 14289 3485 14323 3519
rect 14323 3485 14332 3519
rect 14280 3476 14332 3485
rect 15016 3476 15068 3528
rect 17776 3476 17828 3528
rect 21088 3476 21140 3528
rect 14740 3408 14792 3460
rect 19156 3408 19208 3460
rect 3700 3340 3752 3392
rect 3976 3340 4028 3392
rect 4436 3383 4488 3392
rect 4436 3349 4445 3383
rect 4445 3349 4479 3383
rect 4479 3349 4488 3383
rect 4436 3340 4488 3349
rect 4804 3340 4856 3392
rect 7380 3340 7432 3392
rect 11888 3340 11940 3392
rect 21456 3340 21508 3392
rect 23848 3476 23900 3528
rect 25044 3519 25096 3528
rect 25044 3485 25053 3519
rect 25053 3485 25087 3519
rect 25087 3485 25096 3519
rect 25044 3476 25096 3485
rect 7950 3238 8002 3290
rect 8014 3238 8066 3290
rect 8078 3238 8130 3290
rect 8142 3238 8194 3290
rect 8206 3238 8258 3290
rect 17950 3238 18002 3290
rect 18014 3238 18066 3290
rect 18078 3238 18130 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 2136 3179 2188 3188
rect 2136 3145 2145 3179
rect 2145 3145 2179 3179
rect 2179 3145 2188 3179
rect 2136 3136 2188 3145
rect 5172 3136 5224 3188
rect 5908 3179 5960 3188
rect 5908 3145 5917 3179
rect 5917 3145 5951 3179
rect 5951 3145 5960 3179
rect 5908 3136 5960 3145
rect 23848 3179 23900 3188
rect 23848 3145 23857 3179
rect 23857 3145 23891 3179
rect 23891 3145 23900 3179
rect 23848 3136 23900 3145
rect 10416 3068 10468 3120
rect 1860 3000 1912 3052
rect 3332 3000 3384 3052
rect 3700 3000 3752 3052
rect 4436 3000 4488 3052
rect 5172 3000 5224 3052
rect 5908 3000 5960 3052
rect 7564 3000 7616 3052
rect 8852 3043 8904 3052
rect 8852 3009 8861 3043
rect 8861 3009 8895 3043
rect 8895 3009 8904 3043
rect 8852 3000 8904 3009
rect 10324 3000 10376 3052
rect 10968 3000 11020 3052
rect 12256 3043 12308 3052
rect 12256 3009 12265 3043
rect 12265 3009 12299 3043
rect 12299 3009 12308 3043
rect 12256 3000 12308 3009
rect 14188 3043 14240 3052
rect 14188 3009 14197 3043
rect 14197 3009 14231 3043
rect 14231 3009 14240 3043
rect 14188 3000 14240 3009
rect 16488 3000 16540 3052
rect 16856 3043 16908 3052
rect 16856 3009 16865 3043
rect 16865 3009 16899 3043
rect 16899 3009 16908 3043
rect 16856 3000 16908 3009
rect 18696 3043 18748 3052
rect 18696 3009 18705 3043
rect 18705 3009 18739 3043
rect 18739 3009 18748 3043
rect 18696 3000 18748 3009
rect 22008 3000 22060 3052
rect 22836 3000 22888 3052
rect 4712 2932 4764 2984
rect 4620 2864 4672 2916
rect 8484 2932 8536 2984
rect 10876 2975 10928 2984
rect 10876 2941 10885 2975
rect 10885 2941 10919 2975
rect 10919 2941 10928 2975
rect 10876 2932 10928 2941
rect 11796 2932 11848 2984
rect 13636 2975 13688 2984
rect 13636 2941 13645 2975
rect 13645 2941 13679 2975
rect 13679 2941 13688 2975
rect 13636 2932 13688 2941
rect 14740 2932 14792 2984
rect 15844 2932 15896 2984
rect 16580 2864 16632 2916
rect 20536 2932 20588 2984
rect 23940 2932 23992 2984
rect 19984 2864 20036 2916
rect 21732 2864 21784 2916
rect 23572 2864 23624 2916
rect 25412 2864 25464 2916
rect 1492 2839 1544 2848
rect 1492 2805 1501 2839
rect 1501 2805 1535 2839
rect 1535 2805 1544 2839
rect 1492 2796 1544 2805
rect 1860 2796 1912 2848
rect 7012 2796 7064 2848
rect 7840 2796 7892 2848
rect 9588 2796 9640 2848
rect 9956 2839 10008 2848
rect 9956 2805 9965 2839
rect 9965 2805 9999 2839
rect 9999 2805 10008 2839
rect 9956 2796 10008 2805
rect 17316 2796 17368 2848
rect 18328 2796 18380 2848
rect 18788 2796 18840 2848
rect 19892 2796 19944 2848
rect 20996 2796 21048 2848
rect 22284 2796 22336 2848
rect 2950 2694 3002 2746
rect 3014 2694 3066 2746
rect 3078 2694 3130 2746
rect 3142 2694 3194 2746
rect 3206 2694 3258 2746
rect 12950 2694 13002 2746
rect 13014 2694 13066 2746
rect 13078 2694 13130 2746
rect 13142 2694 13194 2746
rect 13206 2694 13258 2746
rect 22950 2694 23002 2746
rect 23014 2694 23066 2746
rect 23078 2694 23130 2746
rect 23142 2694 23194 2746
rect 23206 2694 23258 2746
rect 2596 2456 2648 2508
rect 3976 2456 4028 2508
rect 2228 2388 2280 2440
rect 3148 2431 3200 2440
rect 3148 2397 3157 2431
rect 3157 2397 3191 2431
rect 3191 2397 3200 2431
rect 3148 2388 3200 2397
rect 10784 2592 10836 2644
rect 15384 2592 15436 2644
rect 24952 2592 25004 2644
rect 25412 2635 25464 2644
rect 25412 2601 25421 2635
rect 25421 2601 25455 2635
rect 25455 2601 25464 2635
rect 25412 2592 25464 2601
rect 6920 2456 6972 2508
rect 9496 2524 9548 2576
rect 11612 2524 11664 2576
rect 18972 2524 19024 2576
rect 12164 2456 12216 2508
rect 4068 2252 4120 2304
rect 5172 2252 5224 2304
rect 8300 2431 8352 2440
rect 8300 2397 8309 2431
rect 8309 2397 8343 2431
rect 8343 2397 8352 2431
rect 8300 2388 8352 2397
rect 7748 2320 7800 2372
rect 6644 2252 6696 2304
rect 6920 2252 6972 2304
rect 7656 2252 7708 2304
rect 8484 2252 8536 2304
rect 11060 2431 11112 2440
rect 11060 2397 11069 2431
rect 11069 2397 11103 2431
rect 11103 2397 11112 2431
rect 11060 2388 11112 2397
rect 11428 2388 11480 2440
rect 15108 2456 15160 2508
rect 12348 2431 12400 2440
rect 12348 2397 12357 2431
rect 12357 2397 12391 2431
rect 12391 2397 12400 2431
rect 12348 2388 12400 2397
rect 15660 2431 15712 2440
rect 15660 2397 15669 2431
rect 15669 2397 15703 2431
rect 15703 2397 15712 2431
rect 15660 2388 15712 2397
rect 15752 2388 15804 2440
rect 16948 2388 17000 2440
rect 13268 2363 13320 2372
rect 13268 2329 13277 2363
rect 13277 2329 13311 2363
rect 13311 2329 13320 2363
rect 13268 2320 13320 2329
rect 14372 2320 14424 2372
rect 17408 2320 17460 2372
rect 18512 2320 18564 2372
rect 24308 2388 24360 2440
rect 10968 2252 11020 2304
rect 7950 2150 8002 2202
rect 8014 2150 8066 2202
rect 8078 2150 8130 2202
rect 8142 2150 8194 2202
rect 8206 2150 8258 2202
rect 17950 2150 18002 2202
rect 18014 2150 18066 2202
rect 18078 2150 18130 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
rect 3148 2048 3200 2100
rect 9036 2048 9088 2100
rect 8300 1980 8352 2032
rect 15936 1980 15988 2032
<< metal2 >>
rect 938 56200 994 57000
rect 1306 56200 1362 57000
rect 1674 56200 1730 57000
rect 2042 56200 2098 57000
rect 2410 56200 2466 57000
rect 2778 56200 2834 57000
rect 3146 56200 3202 57000
rect 3514 56200 3570 57000
rect 3882 56200 3938 57000
rect 4250 56200 4306 57000
rect 4618 56200 4674 57000
rect 4986 56200 5042 57000
rect 5354 56200 5410 57000
rect 5722 56200 5778 57000
rect 6090 56200 6146 57000
rect 6458 56200 6514 57000
rect 6826 56200 6882 57000
rect 7194 56200 7250 57000
rect 7562 56200 7618 57000
rect 7930 56200 7986 57000
rect 8298 56200 8354 57000
rect 8666 56200 8722 57000
rect 9034 56200 9090 57000
rect 9402 56200 9458 57000
rect 9770 56200 9826 57000
rect 10138 56200 10194 57000
rect 10506 56200 10562 57000
rect 10874 56200 10930 57000
rect 11242 56200 11298 57000
rect 11610 56200 11666 57000
rect 11978 56200 12034 57000
rect 12346 56200 12402 57000
rect 12714 56200 12770 57000
rect 12820 56222 13032 56250
rect 952 52698 980 56200
rect 1214 52728 1270 52737
rect 940 52692 992 52698
rect 1214 52663 1270 52672
rect 940 52634 992 52640
rect 1228 52630 1256 52663
rect 1216 52624 1268 52630
rect 1216 52566 1268 52572
rect 1124 50856 1176 50862
rect 1124 50798 1176 50804
rect 1136 50454 1164 50798
rect 1124 50448 1176 50454
rect 1122 50416 1124 50425
rect 1176 50416 1178 50425
rect 1122 50351 1178 50360
rect 1320 49298 1348 56200
rect 1688 49910 1716 56200
rect 2056 50386 2084 56200
rect 2424 51474 2452 56200
rect 2792 55214 2820 56200
rect 3160 55214 3188 56200
rect 2792 55186 2912 55214
rect 3160 55186 3372 55214
rect 2778 55040 2834 55049
rect 2778 54975 2834 54984
rect 2792 53242 2820 54975
rect 2780 53236 2832 53242
rect 2780 53178 2832 53184
rect 2412 51468 2464 51474
rect 2412 51410 2464 51416
rect 2884 50998 2912 55186
rect 2950 53884 3258 53893
rect 2950 53882 2956 53884
rect 3012 53882 3036 53884
rect 3092 53882 3116 53884
rect 3172 53882 3196 53884
rect 3252 53882 3258 53884
rect 3012 53830 3014 53882
rect 3194 53830 3196 53882
rect 2950 53828 2956 53830
rect 3012 53828 3036 53830
rect 3092 53828 3116 53830
rect 3172 53828 3196 53830
rect 3252 53828 3258 53830
rect 2950 53819 3258 53828
rect 2950 52796 3258 52805
rect 2950 52794 2956 52796
rect 3012 52794 3036 52796
rect 3092 52794 3116 52796
rect 3172 52794 3196 52796
rect 3252 52794 3258 52796
rect 3012 52742 3014 52794
rect 3194 52742 3196 52794
rect 2950 52740 2956 52742
rect 3012 52740 3036 52742
rect 3092 52740 3116 52742
rect 3172 52740 3196 52742
rect 3252 52740 3258 52742
rect 2950 52731 3258 52740
rect 3344 52562 3372 55186
rect 3332 52556 3384 52562
rect 3332 52498 3384 52504
rect 3528 51950 3556 56200
rect 3792 53440 3844 53446
rect 3792 53382 3844 53388
rect 3804 52630 3832 53382
rect 3896 53258 3924 56200
rect 3896 53230 4200 53258
rect 4068 52896 4120 52902
rect 4068 52838 4120 52844
rect 3792 52624 3844 52630
rect 3792 52566 3844 52572
rect 3516 51944 3568 51950
rect 3516 51886 3568 51892
rect 2950 51708 3258 51717
rect 2950 51706 2956 51708
rect 3012 51706 3036 51708
rect 3092 51706 3116 51708
rect 3172 51706 3196 51708
rect 3252 51706 3258 51708
rect 3012 51654 3014 51706
rect 3194 51654 3196 51706
rect 2950 51652 2956 51654
rect 3012 51652 3036 51654
rect 3092 51652 3116 51654
rect 3172 51652 3196 51654
rect 3252 51652 3258 51654
rect 2950 51643 3258 51652
rect 2872 50992 2924 50998
rect 2872 50934 2924 50940
rect 2950 50620 3258 50629
rect 2950 50618 2956 50620
rect 3012 50618 3036 50620
rect 3092 50618 3116 50620
rect 3172 50618 3196 50620
rect 3252 50618 3258 50620
rect 3012 50566 3014 50618
rect 3194 50566 3196 50618
rect 2950 50564 2956 50566
rect 3012 50564 3036 50566
rect 3092 50564 3116 50566
rect 3172 50564 3196 50566
rect 3252 50564 3258 50566
rect 2950 50555 3258 50564
rect 2044 50380 2096 50386
rect 2044 50322 2096 50328
rect 3976 50312 4028 50318
rect 3976 50254 4028 50260
rect 1676 49904 1728 49910
rect 1676 49846 1728 49852
rect 3700 49836 3752 49842
rect 3700 49778 3752 49784
rect 2950 49532 3258 49541
rect 2950 49530 2956 49532
rect 3012 49530 3036 49532
rect 3092 49530 3116 49532
rect 3172 49530 3196 49532
rect 3252 49530 3258 49532
rect 3012 49478 3014 49530
rect 3194 49478 3196 49530
rect 2950 49476 2956 49478
rect 3012 49476 3036 49478
rect 3092 49476 3116 49478
rect 3172 49476 3196 49478
rect 3252 49476 3258 49478
rect 2950 49467 3258 49476
rect 1308 49292 1360 49298
rect 1308 49234 1360 49240
rect 3332 49224 3384 49230
rect 3332 49166 3384 49172
rect 2950 48444 3258 48453
rect 2950 48442 2956 48444
rect 3012 48442 3036 48444
rect 3092 48442 3116 48444
rect 3172 48442 3196 48444
rect 3252 48442 3258 48444
rect 3012 48390 3014 48442
rect 3194 48390 3196 48442
rect 2950 48388 2956 48390
rect 3012 48388 3036 48390
rect 3092 48388 3116 48390
rect 3172 48388 3196 48390
rect 3252 48388 3258 48390
rect 2950 48379 3258 48388
rect 1306 48104 1362 48113
rect 1306 48039 1308 48048
rect 1360 48039 1362 48048
rect 1308 48010 1360 48016
rect 2950 47356 3258 47365
rect 2950 47354 2956 47356
rect 3012 47354 3036 47356
rect 3092 47354 3116 47356
rect 3172 47354 3196 47356
rect 3252 47354 3258 47356
rect 3012 47302 3014 47354
rect 3194 47302 3196 47354
rect 2950 47300 2956 47302
rect 3012 47300 3036 47302
rect 3092 47300 3116 47302
rect 3172 47300 3196 47302
rect 3252 47300 3258 47302
rect 2950 47291 3258 47300
rect 2950 46268 3258 46277
rect 2950 46266 2956 46268
rect 3012 46266 3036 46268
rect 3092 46266 3116 46268
rect 3172 46266 3196 46268
rect 3252 46266 3258 46268
rect 3012 46214 3014 46266
rect 3194 46214 3196 46266
rect 2950 46212 2956 46214
rect 3012 46212 3036 46214
rect 3092 46212 3116 46214
rect 3172 46212 3196 46214
rect 3252 46212 3258 46214
rect 2950 46203 3258 46212
rect 1216 45960 1268 45966
rect 1216 45902 1268 45908
rect 1228 45801 1256 45902
rect 1214 45792 1270 45801
rect 1214 45727 1270 45736
rect 1228 45626 1256 45727
rect 1216 45620 1268 45626
rect 1216 45562 1268 45568
rect 2950 45180 3258 45189
rect 2950 45178 2956 45180
rect 3012 45178 3036 45180
rect 3092 45178 3116 45180
rect 3172 45178 3196 45180
rect 3252 45178 3258 45180
rect 3012 45126 3014 45178
rect 3194 45126 3196 45178
rect 2950 45124 2956 45126
rect 3012 45124 3036 45126
rect 3092 45124 3116 45126
rect 3172 45124 3196 45126
rect 3252 45124 3258 45126
rect 2950 45115 3258 45124
rect 2950 44092 3258 44101
rect 2950 44090 2956 44092
rect 3012 44090 3036 44092
rect 3092 44090 3116 44092
rect 3172 44090 3196 44092
rect 3252 44090 3258 44092
rect 3012 44038 3014 44090
rect 3194 44038 3196 44090
rect 2950 44036 2956 44038
rect 3012 44036 3036 44038
rect 3092 44036 3116 44038
rect 3172 44036 3196 44038
rect 3252 44036 3258 44038
rect 2950 44027 3258 44036
rect 1308 43784 1360 43790
rect 1308 43726 1360 43732
rect 1320 43489 1348 43726
rect 1768 43648 1820 43654
rect 1768 43590 1820 43596
rect 1306 43480 1362 43489
rect 1780 43450 1808 43590
rect 1306 43415 1362 43424
rect 1768 43444 1820 43450
rect 1768 43386 1820 43392
rect 2950 43004 3258 43013
rect 2950 43002 2956 43004
rect 3012 43002 3036 43004
rect 3092 43002 3116 43004
rect 3172 43002 3196 43004
rect 3252 43002 3258 43004
rect 3012 42950 3014 43002
rect 3194 42950 3196 43002
rect 2950 42948 2956 42950
rect 3012 42948 3036 42950
rect 3092 42948 3116 42950
rect 3172 42948 3196 42950
rect 3252 42948 3258 42950
rect 2950 42939 3258 42948
rect 2950 41916 3258 41925
rect 2950 41914 2956 41916
rect 3012 41914 3036 41916
rect 3092 41914 3116 41916
rect 3172 41914 3196 41916
rect 3252 41914 3258 41916
rect 3012 41862 3014 41914
rect 3194 41862 3196 41914
rect 2950 41860 2956 41862
rect 3012 41860 3036 41862
rect 3092 41860 3116 41862
rect 3172 41860 3196 41862
rect 3252 41860 3258 41862
rect 2950 41851 3258 41860
rect 1676 41540 1728 41546
rect 1676 41482 1728 41488
rect 1688 41177 1716 41482
rect 1674 41168 1730 41177
rect 1674 41103 1730 41112
rect 2950 40828 3258 40837
rect 2950 40826 2956 40828
rect 3012 40826 3036 40828
rect 3092 40826 3116 40828
rect 3172 40826 3196 40828
rect 3252 40826 3258 40828
rect 3012 40774 3014 40826
rect 3194 40774 3196 40826
rect 2950 40772 2956 40774
rect 3012 40772 3036 40774
rect 3092 40772 3116 40774
rect 3172 40772 3196 40774
rect 3252 40772 3258 40774
rect 2950 40763 3258 40772
rect 3344 40662 3372 49166
rect 3712 42294 3740 49778
rect 3700 42288 3752 42294
rect 3700 42230 3752 42236
rect 3608 41472 3660 41478
rect 3608 41414 3660 41420
rect 3332 40656 3384 40662
rect 3332 40598 3384 40604
rect 2950 39740 3258 39749
rect 2950 39738 2956 39740
rect 3012 39738 3036 39740
rect 3092 39738 3116 39740
rect 3172 39738 3196 39740
rect 3252 39738 3258 39740
rect 3012 39686 3014 39738
rect 3194 39686 3196 39738
rect 2950 39684 2956 39686
rect 3012 39684 3036 39686
rect 3092 39684 3116 39686
rect 3172 39684 3196 39686
rect 3252 39684 3258 39686
rect 2950 39675 3258 39684
rect 1216 38956 1268 38962
rect 1216 38898 1268 38904
rect 1228 38865 1256 38898
rect 1214 38856 1270 38865
rect 1214 38791 1270 38800
rect 2950 38652 3258 38661
rect 2950 38650 2956 38652
rect 3012 38650 3036 38652
rect 3092 38650 3116 38652
rect 3172 38650 3196 38652
rect 3252 38650 3258 38652
rect 3012 38598 3014 38650
rect 3194 38598 3196 38650
rect 2950 38596 2956 38598
rect 3012 38596 3036 38598
rect 3092 38596 3116 38598
rect 3172 38596 3196 38598
rect 3252 38596 3258 38598
rect 2950 38587 3258 38596
rect 2950 37564 3258 37573
rect 2950 37562 2956 37564
rect 3012 37562 3036 37564
rect 3092 37562 3116 37564
rect 3172 37562 3196 37564
rect 3252 37562 3258 37564
rect 3012 37510 3014 37562
rect 3194 37510 3196 37562
rect 2950 37508 2956 37510
rect 3012 37508 3036 37510
rect 3092 37508 3116 37510
rect 3172 37508 3196 37510
rect 3252 37508 3258 37510
rect 2950 37499 3258 37508
rect 1308 36780 1360 36786
rect 1308 36722 1360 36728
rect 1320 36553 1348 36722
rect 1952 36576 2004 36582
rect 1306 36544 1362 36553
rect 1952 36518 2004 36524
rect 1306 36479 1362 36488
rect 1584 34604 1636 34610
rect 1584 34546 1636 34552
rect 1596 34241 1624 34546
rect 1582 34232 1638 34241
rect 1582 34167 1638 34176
rect 1308 32428 1360 32434
rect 1308 32370 1360 32376
rect 1320 31929 1348 32370
rect 1306 31920 1362 31929
rect 1306 31855 1362 31864
rect 1308 29708 1360 29714
rect 1308 29650 1360 29656
rect 1320 29617 1348 29650
rect 1768 29640 1820 29646
rect 1306 29608 1362 29617
rect 1768 29582 1820 29588
rect 1306 29543 1362 29552
rect 1308 27532 1360 27538
rect 1308 27474 1360 27480
rect 1320 27305 1348 27474
rect 1306 27296 1362 27305
rect 1306 27231 1362 27240
rect 1780 27130 1808 29582
rect 1964 28626 1992 36518
rect 2950 36476 3258 36485
rect 2950 36474 2956 36476
rect 3012 36474 3036 36476
rect 3092 36474 3116 36476
rect 3172 36474 3196 36476
rect 3252 36474 3258 36476
rect 3012 36422 3014 36474
rect 3194 36422 3196 36474
rect 2950 36420 2956 36422
rect 3012 36420 3036 36422
rect 3092 36420 3116 36422
rect 3172 36420 3196 36422
rect 3252 36420 3258 36422
rect 2950 36411 3258 36420
rect 2950 35388 3258 35397
rect 2950 35386 2956 35388
rect 3012 35386 3036 35388
rect 3092 35386 3116 35388
rect 3172 35386 3196 35388
rect 3252 35386 3258 35388
rect 3012 35334 3014 35386
rect 3194 35334 3196 35386
rect 2950 35332 2956 35334
rect 3012 35332 3036 35334
rect 3092 35332 3116 35334
rect 3172 35332 3196 35334
rect 3252 35332 3258 35334
rect 2950 35323 3258 35332
rect 2688 34740 2740 34746
rect 2688 34682 2740 34688
rect 2596 32224 2648 32230
rect 2596 32166 2648 32172
rect 1952 28620 2004 28626
rect 1952 28562 2004 28568
rect 1952 27464 2004 27470
rect 1952 27406 2004 27412
rect 1768 27124 1820 27130
rect 1768 27066 1820 27072
rect 1308 25356 1360 25362
rect 1308 25298 1360 25304
rect 1320 24993 1348 25298
rect 1768 25288 1820 25294
rect 1768 25230 1820 25236
rect 1306 24984 1362 24993
rect 1306 24919 1362 24928
rect 940 23044 992 23050
rect 940 22986 992 22992
rect 952 22681 980 22986
rect 1780 22778 1808 25230
rect 1964 24682 1992 27406
rect 2228 26988 2280 26994
rect 2228 26930 2280 26936
rect 2240 26042 2268 26930
rect 2608 26450 2636 32166
rect 2700 27538 2728 34682
rect 2950 34300 3258 34309
rect 2950 34298 2956 34300
rect 3012 34298 3036 34300
rect 3092 34298 3116 34300
rect 3172 34298 3196 34300
rect 3252 34298 3258 34300
rect 3012 34246 3014 34298
rect 3194 34246 3196 34298
rect 2950 34244 2956 34246
rect 3012 34244 3036 34246
rect 3092 34244 3116 34246
rect 3172 34244 3196 34246
rect 3252 34244 3258 34246
rect 2950 34235 3258 34244
rect 2950 33212 3258 33221
rect 2950 33210 2956 33212
rect 3012 33210 3036 33212
rect 3092 33210 3116 33212
rect 3172 33210 3196 33212
rect 3252 33210 3258 33212
rect 3012 33158 3014 33210
rect 3194 33158 3196 33210
rect 2950 33156 2956 33158
rect 3012 33156 3036 33158
rect 3092 33156 3116 33158
rect 3172 33156 3196 33158
rect 3252 33156 3258 33158
rect 2950 33147 3258 33156
rect 2950 32124 3258 32133
rect 2950 32122 2956 32124
rect 3012 32122 3036 32124
rect 3092 32122 3116 32124
rect 3172 32122 3196 32124
rect 3252 32122 3258 32124
rect 3012 32070 3014 32122
rect 3194 32070 3196 32122
rect 2950 32068 2956 32070
rect 3012 32068 3036 32070
rect 3092 32068 3116 32070
rect 3172 32068 3196 32070
rect 3252 32068 3258 32070
rect 2950 32059 3258 32068
rect 2950 31036 3258 31045
rect 2950 31034 2956 31036
rect 3012 31034 3036 31036
rect 3092 31034 3116 31036
rect 3172 31034 3196 31036
rect 3252 31034 3258 31036
rect 3012 30982 3014 31034
rect 3194 30982 3196 31034
rect 2950 30980 2956 30982
rect 3012 30980 3036 30982
rect 3092 30980 3116 30982
rect 3172 30980 3196 30982
rect 3252 30980 3258 30982
rect 2950 30971 3258 30980
rect 2950 29948 3258 29957
rect 2950 29946 2956 29948
rect 3012 29946 3036 29948
rect 3092 29946 3116 29948
rect 3172 29946 3196 29948
rect 3252 29946 3258 29948
rect 3012 29894 3014 29946
rect 3194 29894 3196 29946
rect 2950 29892 2956 29894
rect 3012 29892 3036 29894
rect 3092 29892 3116 29894
rect 3172 29892 3196 29894
rect 3252 29892 3258 29894
rect 2950 29883 3258 29892
rect 3516 29572 3568 29578
rect 3516 29514 3568 29520
rect 2950 28860 3258 28869
rect 2950 28858 2956 28860
rect 3012 28858 3036 28860
rect 3092 28858 3116 28860
rect 3172 28858 3196 28860
rect 3252 28858 3258 28860
rect 3012 28806 3014 28858
rect 3194 28806 3196 28858
rect 2950 28804 2956 28806
rect 3012 28804 3036 28806
rect 3092 28804 3116 28806
rect 3172 28804 3196 28806
rect 3252 28804 3258 28806
rect 2950 28795 3258 28804
rect 2950 27772 3258 27781
rect 2950 27770 2956 27772
rect 3012 27770 3036 27772
rect 3092 27770 3116 27772
rect 3172 27770 3196 27772
rect 3252 27770 3258 27772
rect 3012 27718 3014 27770
rect 3194 27718 3196 27770
rect 2950 27716 2956 27718
rect 3012 27716 3036 27718
rect 3092 27716 3116 27718
rect 3172 27716 3196 27718
rect 3252 27716 3258 27718
rect 2950 27707 3258 27716
rect 2688 27532 2740 27538
rect 2688 27474 2740 27480
rect 3528 27130 3556 29514
rect 3516 27124 3568 27130
rect 3516 27066 3568 27072
rect 3332 26988 3384 26994
rect 3332 26930 3384 26936
rect 2950 26684 3258 26693
rect 2950 26682 2956 26684
rect 3012 26682 3036 26684
rect 3092 26682 3116 26684
rect 3172 26682 3196 26684
rect 3252 26682 3258 26684
rect 3012 26630 3014 26682
rect 3194 26630 3196 26682
rect 2950 26628 2956 26630
rect 3012 26628 3036 26630
rect 3092 26628 3116 26630
rect 3172 26628 3196 26630
rect 3252 26628 3258 26630
rect 2950 26619 3258 26628
rect 2596 26444 2648 26450
rect 2596 26386 2648 26392
rect 2228 26036 2280 26042
rect 2228 25978 2280 25984
rect 2872 25900 2924 25906
rect 2872 25842 2924 25848
rect 2228 24812 2280 24818
rect 2228 24754 2280 24760
rect 1952 24676 2004 24682
rect 1952 24618 2004 24624
rect 2240 22778 2268 24754
rect 2884 24410 2912 25842
rect 3344 25770 3372 26930
rect 3332 25764 3384 25770
rect 3332 25706 3384 25712
rect 2950 25596 3258 25605
rect 2950 25594 2956 25596
rect 3012 25594 3036 25596
rect 3092 25594 3116 25596
rect 3172 25594 3196 25596
rect 3252 25594 3258 25596
rect 3012 25542 3014 25594
rect 3194 25542 3196 25594
rect 2950 25540 2956 25542
rect 3012 25540 3036 25542
rect 3092 25540 3116 25542
rect 3172 25540 3196 25542
rect 3252 25540 3258 25542
rect 2950 25531 3258 25540
rect 3344 25362 3372 25706
rect 3620 25498 3648 41414
rect 3988 41274 4016 50254
rect 4080 49162 4108 52838
rect 4172 51474 4200 53230
rect 4264 53038 4292 56200
rect 4632 53650 4660 56200
rect 4620 53644 4672 53650
rect 4620 53586 4672 53592
rect 4252 53032 4304 53038
rect 4252 52974 4304 52980
rect 4344 52692 4396 52698
rect 4344 52634 4396 52640
rect 4160 51468 4212 51474
rect 4160 51410 4212 51416
rect 4160 50924 4212 50930
rect 4160 50866 4212 50872
rect 4068 49156 4120 49162
rect 4068 49098 4120 49104
rect 4068 48000 4120 48006
rect 4068 47942 4120 47948
rect 3976 41268 4028 41274
rect 3976 41210 4028 41216
rect 4080 40050 4108 47942
rect 4172 42770 4200 50866
rect 4356 50386 4384 52634
rect 4436 52556 4488 52562
rect 4436 52498 4488 52504
rect 4344 50380 4396 50386
rect 4344 50322 4396 50328
rect 4160 42764 4212 42770
rect 4160 42706 4212 42712
rect 4344 42220 4396 42226
rect 4344 42162 4396 42168
rect 4356 42022 4384 42162
rect 4344 42016 4396 42022
rect 4344 41958 4396 41964
rect 4252 41132 4304 41138
rect 4252 41074 4304 41080
rect 4264 40934 4292 41074
rect 4252 40928 4304 40934
rect 4252 40870 4304 40876
rect 4160 40384 4212 40390
rect 4160 40326 4212 40332
rect 4068 40044 4120 40050
rect 4068 39986 4120 39992
rect 3976 38752 4028 38758
rect 3976 38694 4028 38700
rect 3988 29714 4016 38694
rect 4172 31210 4200 40326
rect 4160 31204 4212 31210
rect 4160 31146 4212 31152
rect 3976 29708 4028 29714
rect 3976 29650 4028 29656
rect 4264 28762 4292 40870
rect 4356 29850 4384 41958
rect 4448 41818 4476 52498
rect 4528 52488 4580 52494
rect 4528 52430 4580 52436
rect 4436 41812 4488 41818
rect 4436 41754 4488 41760
rect 4540 41274 4568 52430
rect 5000 52086 5028 56200
rect 5368 54126 5396 56200
rect 5356 54120 5408 54126
rect 5356 54062 5408 54068
rect 5736 53038 5764 56200
rect 5908 54188 5960 54194
rect 5908 54130 5960 54136
rect 5816 53100 5868 53106
rect 5816 53042 5868 53048
rect 5724 53032 5776 53038
rect 5724 52974 5776 52980
rect 4988 52080 5040 52086
rect 4988 52022 5040 52028
rect 5356 52012 5408 52018
rect 5356 51954 5408 51960
rect 4988 43308 5040 43314
rect 4988 43250 5040 43256
rect 5172 43308 5224 43314
rect 5172 43250 5224 43256
rect 4528 41268 4580 41274
rect 4528 41210 4580 41216
rect 5000 39030 5028 43250
rect 4988 39024 5040 39030
rect 4988 38966 5040 38972
rect 4988 38888 5040 38894
rect 4988 38830 5040 38836
rect 5000 36650 5028 38830
rect 5184 36922 5212 43250
rect 5368 41818 5396 51954
rect 5828 45014 5856 53042
rect 5920 51610 5948 54130
rect 6000 52896 6052 52902
rect 6000 52838 6052 52844
rect 5908 51604 5960 51610
rect 5908 51546 5960 51552
rect 6012 51406 6040 52838
rect 6104 52562 6132 56200
rect 6184 53576 6236 53582
rect 6184 53518 6236 53524
rect 6092 52556 6144 52562
rect 6092 52498 6144 52504
rect 6000 51400 6052 51406
rect 6000 51342 6052 51348
rect 5816 45008 5868 45014
rect 5816 44950 5868 44956
rect 6196 43926 6224 53518
rect 6368 53168 6420 53174
rect 6368 53110 6420 53116
rect 6184 43920 6236 43926
rect 6184 43862 6236 43868
rect 6380 42770 6408 53110
rect 6472 52562 6500 56200
rect 6644 53576 6696 53582
rect 6644 53518 6696 53524
rect 6460 52556 6512 52562
rect 6460 52498 6512 52504
rect 6552 52488 6604 52494
rect 6552 52430 6604 52436
rect 6564 49994 6592 52430
rect 6656 50130 6684 53518
rect 6736 53100 6788 53106
rect 6736 53042 6788 53048
rect 6748 51456 6776 53042
rect 6840 52714 6868 56200
rect 7208 54126 7236 56200
rect 7196 54120 7248 54126
rect 7196 54062 7248 54068
rect 7576 53650 7604 56200
rect 7944 55214 7972 56200
rect 7852 55186 7972 55214
rect 7564 53644 7616 53650
rect 7564 53586 7616 53592
rect 7380 53576 7432 53582
rect 7380 53518 7432 53524
rect 6840 52686 7052 52714
rect 7024 52578 7052 52686
rect 6920 52556 6972 52562
rect 7024 52550 7144 52578
rect 6920 52498 6972 52504
rect 6932 51474 6960 52498
rect 7012 52012 7064 52018
rect 7012 51954 7064 51960
rect 6920 51468 6972 51474
rect 6748 51428 6868 51456
rect 6736 51332 6788 51338
rect 6736 51274 6788 51280
rect 6748 50998 6776 51274
rect 6736 50992 6788 50998
rect 6736 50934 6788 50940
rect 6656 50102 6776 50130
rect 6564 49966 6684 49994
rect 6552 49836 6604 49842
rect 6552 49778 6604 49784
rect 6564 43450 6592 49778
rect 6656 45558 6684 49966
rect 6644 45552 6696 45558
rect 6644 45494 6696 45500
rect 6748 44334 6776 50102
rect 6840 47258 6868 51428
rect 6920 51410 6972 51416
rect 6920 50788 6972 50794
rect 6920 50730 6972 50736
rect 6828 47252 6880 47258
rect 6828 47194 6880 47200
rect 6736 44328 6788 44334
rect 6736 44270 6788 44276
rect 6552 43444 6604 43450
rect 6552 43386 6604 43392
rect 6368 42764 6420 42770
rect 6368 42706 6420 42712
rect 6460 42628 6512 42634
rect 6460 42570 6512 42576
rect 5356 41812 5408 41818
rect 5356 41754 5408 41760
rect 6276 41472 6328 41478
rect 6276 41414 6328 41420
rect 5908 40520 5960 40526
rect 5908 40462 5960 40468
rect 5920 38758 5948 40462
rect 5908 38752 5960 38758
rect 5908 38694 5960 38700
rect 5920 38418 5948 38694
rect 5908 38412 5960 38418
rect 5908 38354 5960 38360
rect 6092 38276 6144 38282
rect 6092 38218 6144 38224
rect 5908 37460 5960 37466
rect 5908 37402 5960 37408
rect 5264 37256 5316 37262
rect 5264 37198 5316 37204
rect 5172 36916 5224 36922
rect 5172 36858 5224 36864
rect 4988 36644 5040 36650
rect 4988 36586 5040 36592
rect 4528 35624 4580 35630
rect 4528 35566 4580 35572
rect 4540 35290 4568 35566
rect 4528 35284 4580 35290
rect 4528 35226 4580 35232
rect 5000 34746 5028 36586
rect 5276 35494 5304 37198
rect 5356 36780 5408 36786
rect 5356 36722 5408 36728
rect 5264 35488 5316 35494
rect 5264 35430 5316 35436
rect 4988 34740 5040 34746
rect 4988 34682 5040 34688
rect 5276 34542 5304 35430
rect 5264 34536 5316 34542
rect 5264 34478 5316 34484
rect 4988 34400 5040 34406
rect 4988 34342 5040 34348
rect 5000 34066 5028 34342
rect 4712 34060 4764 34066
rect 4712 34002 4764 34008
rect 4988 34060 5040 34066
rect 4988 34002 5040 34008
rect 4724 31278 4752 34002
rect 4988 32360 5040 32366
rect 4988 32302 5040 32308
rect 5000 31482 5028 32302
rect 5368 31482 5396 36722
rect 5816 34740 5868 34746
rect 5816 34682 5868 34688
rect 5828 33930 5856 34682
rect 5816 33924 5868 33930
rect 5816 33866 5868 33872
rect 4988 31476 5040 31482
rect 4988 31418 5040 31424
rect 5356 31476 5408 31482
rect 5356 31418 5408 31424
rect 4712 31272 4764 31278
rect 4712 31214 4764 31220
rect 4804 31272 4856 31278
rect 4804 31214 4856 31220
rect 4344 29844 4396 29850
rect 4344 29786 4396 29792
rect 4252 28756 4304 28762
rect 4252 28698 4304 28704
rect 4068 28416 4120 28422
rect 4068 28358 4120 28364
rect 3976 27396 4028 27402
rect 3976 27338 4028 27344
rect 3884 26308 3936 26314
rect 3884 26250 3936 26256
rect 3608 25492 3660 25498
rect 3608 25434 3660 25440
rect 3332 25356 3384 25362
rect 3332 25298 3384 25304
rect 3344 24698 3372 25298
rect 3620 25294 3648 25434
rect 3608 25288 3660 25294
rect 3608 25230 3660 25236
rect 3344 24670 3464 24698
rect 2950 24508 3258 24517
rect 2950 24506 2956 24508
rect 3012 24506 3036 24508
rect 3092 24506 3116 24508
rect 3172 24506 3196 24508
rect 3252 24506 3258 24508
rect 3012 24454 3014 24506
rect 3194 24454 3196 24506
rect 2950 24452 2956 24454
rect 3012 24452 3036 24454
rect 3092 24452 3116 24454
rect 3172 24452 3196 24454
rect 3252 24452 3258 24454
rect 2950 24443 3258 24452
rect 2872 24404 2924 24410
rect 2872 24346 2924 24352
rect 3148 24404 3200 24410
rect 3148 24346 3200 24352
rect 2780 23112 2832 23118
rect 2780 23054 2832 23060
rect 1768 22772 1820 22778
rect 1768 22714 1820 22720
rect 2228 22772 2280 22778
rect 2228 22714 2280 22720
rect 938 22672 994 22681
rect 938 22607 994 22616
rect 2136 22636 2188 22642
rect 2136 22578 2188 22584
rect 1768 21888 1820 21894
rect 1768 21830 1820 21836
rect 1780 20466 1808 21830
rect 2148 21690 2176 22578
rect 2792 21894 2820 23054
rect 2884 22642 2912 24346
rect 3160 23526 3188 24346
rect 3148 23520 3200 23526
rect 3148 23462 3200 23468
rect 2950 23420 3258 23429
rect 2950 23418 2956 23420
rect 3012 23418 3036 23420
rect 3092 23418 3116 23420
rect 3172 23418 3196 23420
rect 3252 23418 3258 23420
rect 3012 23366 3014 23418
rect 3194 23366 3196 23418
rect 2950 23364 2956 23366
rect 3012 23364 3036 23366
rect 3092 23364 3116 23366
rect 3172 23364 3196 23366
rect 3252 23364 3258 23366
rect 2950 23355 3258 23364
rect 2872 22636 2924 22642
rect 2872 22578 2924 22584
rect 3332 22636 3384 22642
rect 3332 22578 3384 22584
rect 2950 22332 3258 22341
rect 2950 22330 2956 22332
rect 3012 22330 3036 22332
rect 3092 22330 3116 22332
rect 3172 22330 3196 22332
rect 3252 22330 3258 22332
rect 3012 22278 3014 22330
rect 3194 22278 3196 22330
rect 2950 22276 2956 22278
rect 3012 22276 3036 22278
rect 3092 22276 3116 22278
rect 3172 22276 3196 22278
rect 3252 22276 3258 22278
rect 2950 22267 3258 22276
rect 2872 22024 2924 22030
rect 2872 21966 2924 21972
rect 2780 21888 2832 21894
rect 2780 21830 2832 21836
rect 2136 21684 2188 21690
rect 2136 21626 2188 21632
rect 2780 21480 2832 21486
rect 2780 21422 2832 21428
rect 1768 20460 1820 20466
rect 1768 20402 1820 20408
rect 1308 20392 1360 20398
rect 1306 20360 1308 20369
rect 1360 20360 1362 20369
rect 1306 20295 1362 20304
rect 1860 19712 1912 19718
rect 1860 19654 1912 19660
rect 1768 18624 1820 18630
rect 1768 18566 1820 18572
rect 1308 18216 1360 18222
rect 1308 18158 1360 18164
rect 1320 18057 1348 18158
rect 1306 18048 1362 18057
rect 1306 17983 1362 17992
rect 1780 16114 1808 18566
rect 1872 18290 1900 19654
rect 2792 18766 2820 21422
rect 2884 21146 2912 21966
rect 2950 21244 3258 21253
rect 2950 21242 2956 21244
rect 3012 21242 3036 21244
rect 3092 21242 3116 21244
rect 3172 21242 3196 21244
rect 3252 21242 3258 21244
rect 3012 21190 3014 21242
rect 3194 21190 3196 21242
rect 2950 21188 2956 21190
rect 3012 21188 3036 21190
rect 3092 21188 3116 21190
rect 3172 21188 3196 21190
rect 3252 21188 3258 21190
rect 2950 21179 3258 21188
rect 2872 21140 2924 21146
rect 2872 21082 2924 21088
rect 2950 20156 3258 20165
rect 2950 20154 2956 20156
rect 3012 20154 3036 20156
rect 3092 20154 3116 20156
rect 3172 20154 3196 20156
rect 3252 20154 3258 20156
rect 3012 20102 3014 20154
rect 3194 20102 3196 20154
rect 2950 20100 2956 20102
rect 3012 20100 3036 20102
rect 3092 20100 3116 20102
rect 3172 20100 3196 20102
rect 3252 20100 3258 20102
rect 2950 20091 3258 20100
rect 3344 19854 3372 22578
rect 3436 22166 3464 24670
rect 3620 24206 3648 25230
rect 3608 24200 3660 24206
rect 3608 24142 3660 24148
rect 3896 22778 3924 26250
rect 3988 24070 4016 27338
rect 4080 26042 4108 28358
rect 4068 26036 4120 26042
rect 4068 25978 4120 25984
rect 4252 25832 4304 25838
rect 4252 25774 4304 25780
rect 4160 25492 4212 25498
rect 4160 25434 4212 25440
rect 4068 24880 4120 24886
rect 4068 24822 4120 24828
rect 4080 24410 4108 24822
rect 4172 24750 4200 25434
rect 4160 24744 4212 24750
rect 4160 24686 4212 24692
rect 4068 24404 4120 24410
rect 4068 24346 4120 24352
rect 4068 24200 4120 24206
rect 4068 24142 4120 24148
rect 3976 24064 4028 24070
rect 3976 24006 4028 24012
rect 3884 22772 3936 22778
rect 3884 22714 3936 22720
rect 3884 22636 3936 22642
rect 3884 22578 3936 22584
rect 3424 22160 3476 22166
rect 3424 22102 3476 22108
rect 3424 21344 3476 21350
rect 3424 21286 3476 21292
rect 3436 21010 3464 21286
rect 3424 21004 3476 21010
rect 3424 20946 3476 20952
rect 3896 20942 3924 22578
rect 3976 21480 4028 21486
rect 3976 21422 4028 21428
rect 3884 20936 3936 20942
rect 3884 20878 3936 20884
rect 3332 19848 3384 19854
rect 3332 19790 3384 19796
rect 2950 19068 3258 19077
rect 2950 19066 2956 19068
rect 3012 19066 3036 19068
rect 3092 19066 3116 19068
rect 3172 19066 3196 19068
rect 3252 19066 3258 19068
rect 3012 19014 3014 19066
rect 3194 19014 3196 19066
rect 2950 19012 2956 19014
rect 3012 19012 3036 19014
rect 3092 19012 3116 19014
rect 3172 19012 3196 19014
rect 3252 19012 3258 19014
rect 2950 19003 3258 19012
rect 3988 18970 4016 21422
rect 4080 21418 4108 24142
rect 4172 23798 4200 24686
rect 4160 23792 4212 23798
rect 4160 23734 4212 23740
rect 4160 23520 4212 23526
rect 4160 23462 4212 23468
rect 4172 23202 4200 23462
rect 4264 23322 4292 25774
rect 4712 25696 4764 25702
rect 4712 25638 4764 25644
rect 4344 25288 4396 25294
rect 4344 25230 4396 25236
rect 4252 23316 4304 23322
rect 4252 23258 4304 23264
rect 4172 23174 4292 23202
rect 4160 22432 4212 22438
rect 4160 22374 4212 22380
rect 4172 21554 4200 22374
rect 4160 21548 4212 21554
rect 4160 21490 4212 21496
rect 4068 21412 4120 21418
rect 4068 21354 4120 21360
rect 4068 20936 4120 20942
rect 4068 20878 4120 20884
rect 3976 18964 4028 18970
rect 3976 18906 4028 18912
rect 2780 18760 2832 18766
rect 2780 18702 2832 18708
rect 1860 18284 1912 18290
rect 1860 18226 1912 18232
rect 2136 18080 2188 18086
rect 2136 18022 2188 18028
rect 1768 16108 1820 16114
rect 1768 16050 1820 16056
rect 1308 16040 1360 16046
rect 1308 15982 1360 15988
rect 1320 15745 1348 15982
rect 1306 15736 1362 15745
rect 1306 15671 1362 15680
rect 1768 13864 1820 13870
rect 1768 13806 1820 13812
rect 1780 13433 1808 13806
rect 1766 13424 1822 13433
rect 1766 13359 1822 13368
rect 1400 4480 1452 4486
rect 1400 4422 1452 4428
rect 1412 4146 1440 4422
rect 1124 4140 1176 4146
rect 1124 4082 1176 4088
rect 1400 4140 1452 4146
rect 1400 4082 1452 4088
rect 1136 800 1164 4082
rect 1492 3460 1544 3466
rect 1492 3402 1544 3408
rect 1504 2854 1532 3402
rect 2148 3194 2176 18022
rect 2950 17980 3258 17989
rect 2950 17978 2956 17980
rect 3012 17978 3036 17980
rect 3092 17978 3116 17980
rect 3172 17978 3196 17980
rect 3252 17978 3258 17980
rect 3012 17926 3014 17978
rect 3194 17926 3196 17978
rect 2950 17924 2956 17926
rect 3012 17924 3036 17926
rect 3092 17924 3116 17926
rect 3172 17924 3196 17926
rect 3252 17924 3258 17926
rect 2950 17915 3258 17924
rect 4080 16998 4108 20878
rect 4264 20534 4292 23174
rect 4356 21554 4384 25230
rect 4528 24132 4580 24138
rect 4528 24074 4580 24080
rect 4540 22094 4568 24074
rect 4540 22066 4660 22094
rect 4344 21548 4396 21554
rect 4344 21490 4396 21496
rect 4356 20806 4384 21490
rect 4344 20800 4396 20806
rect 4344 20742 4396 20748
rect 4252 20528 4304 20534
rect 4252 20470 4304 20476
rect 4160 18760 4212 18766
rect 4160 18702 4212 18708
rect 4172 17338 4200 18702
rect 4356 17882 4384 20742
rect 4344 17876 4396 17882
rect 4344 17818 4396 17824
rect 4160 17332 4212 17338
rect 4160 17274 4212 17280
rect 4068 16992 4120 16998
rect 4068 16934 4120 16940
rect 2950 16892 3258 16901
rect 2950 16890 2956 16892
rect 3012 16890 3036 16892
rect 3092 16890 3116 16892
rect 3172 16890 3196 16892
rect 3252 16890 3258 16892
rect 3012 16838 3014 16890
rect 3194 16838 3196 16890
rect 2950 16836 2956 16838
rect 3012 16836 3036 16838
rect 3092 16836 3116 16838
rect 3172 16836 3196 16838
rect 3252 16836 3258 16838
rect 2950 16827 3258 16836
rect 2780 16652 2832 16658
rect 2780 16594 2832 16600
rect 2792 13938 2820 16594
rect 4080 16590 4108 16934
rect 4068 16584 4120 16590
rect 4068 16526 4120 16532
rect 2950 15804 3258 15813
rect 2950 15802 2956 15804
rect 3012 15802 3036 15804
rect 3092 15802 3116 15804
rect 3172 15802 3196 15804
rect 3252 15802 3258 15804
rect 3012 15750 3014 15802
rect 3194 15750 3196 15802
rect 2950 15748 2956 15750
rect 3012 15748 3036 15750
rect 3092 15748 3116 15750
rect 3172 15748 3196 15750
rect 3252 15748 3258 15750
rect 2950 15739 3258 15748
rect 2950 14716 3258 14725
rect 2950 14714 2956 14716
rect 3012 14714 3036 14716
rect 3092 14714 3116 14716
rect 3172 14714 3196 14716
rect 3252 14714 3258 14716
rect 3012 14662 3014 14714
rect 3194 14662 3196 14714
rect 2950 14660 2956 14662
rect 3012 14660 3036 14662
rect 3092 14660 3116 14662
rect 3172 14660 3196 14662
rect 3252 14660 3258 14662
rect 2950 14651 3258 14660
rect 2780 13932 2832 13938
rect 2780 13874 2832 13880
rect 2950 13628 3258 13637
rect 2950 13626 2956 13628
rect 3012 13626 3036 13628
rect 3092 13626 3116 13628
rect 3172 13626 3196 13628
rect 3252 13626 3258 13628
rect 3012 13574 3014 13626
rect 3194 13574 3196 13626
rect 2950 13572 2956 13574
rect 3012 13572 3036 13574
rect 3092 13572 3116 13574
rect 3172 13572 3196 13574
rect 3252 13572 3258 13574
rect 2950 13563 3258 13572
rect 2950 12540 3258 12549
rect 2950 12538 2956 12540
rect 3012 12538 3036 12540
rect 3092 12538 3116 12540
rect 3172 12538 3196 12540
rect 3252 12538 3258 12540
rect 3012 12486 3014 12538
rect 3194 12486 3196 12538
rect 2950 12484 2956 12486
rect 3012 12484 3036 12486
rect 3092 12484 3116 12486
rect 3172 12484 3196 12486
rect 3252 12484 3258 12486
rect 2950 12475 3258 12484
rect 3332 12368 3384 12374
rect 3332 12310 3384 12316
rect 2950 11452 3258 11461
rect 2950 11450 2956 11452
rect 3012 11450 3036 11452
rect 3092 11450 3116 11452
rect 3172 11450 3196 11452
rect 3252 11450 3258 11452
rect 3012 11398 3014 11450
rect 3194 11398 3196 11450
rect 2950 11396 2956 11398
rect 3012 11396 3036 11398
rect 3092 11396 3116 11398
rect 3172 11396 3196 11398
rect 3252 11396 3258 11398
rect 2950 11387 3258 11396
rect 3344 11121 3372 12310
rect 3330 11112 3386 11121
rect 3330 11047 3386 11056
rect 2950 10364 3258 10373
rect 2950 10362 2956 10364
rect 3012 10362 3036 10364
rect 3092 10362 3116 10364
rect 3172 10362 3196 10364
rect 3252 10362 3258 10364
rect 3012 10310 3014 10362
rect 3194 10310 3196 10362
rect 2950 10308 2956 10310
rect 3012 10308 3036 10310
rect 3092 10308 3116 10310
rect 3172 10308 3196 10310
rect 3252 10308 3258 10310
rect 2950 10299 3258 10308
rect 2872 9648 2924 9654
rect 2872 9590 2924 9596
rect 2884 8809 2912 9590
rect 2950 9276 3258 9285
rect 2950 9274 2956 9276
rect 3012 9274 3036 9276
rect 3092 9274 3116 9276
rect 3172 9274 3196 9276
rect 3252 9274 3258 9276
rect 3012 9222 3014 9274
rect 3194 9222 3196 9274
rect 2950 9220 2956 9222
rect 3012 9220 3036 9222
rect 3092 9220 3116 9222
rect 3172 9220 3196 9222
rect 3252 9220 3258 9222
rect 2950 9211 3258 9220
rect 2870 8800 2926 8809
rect 2870 8735 2926 8744
rect 2780 8424 2832 8430
rect 2780 8366 2832 8372
rect 2688 3936 2740 3942
rect 2688 3878 2740 3884
rect 2700 3618 2728 3878
rect 2792 3738 2820 8366
rect 2950 8188 3258 8197
rect 2950 8186 2956 8188
rect 3012 8186 3036 8188
rect 3092 8186 3116 8188
rect 3172 8186 3196 8188
rect 3252 8186 3258 8188
rect 3012 8134 3014 8186
rect 3194 8134 3196 8186
rect 2950 8132 2956 8134
rect 3012 8132 3036 8134
rect 3092 8132 3116 8134
rect 3172 8132 3196 8134
rect 3252 8132 3258 8134
rect 2950 8123 3258 8132
rect 2950 7100 3258 7109
rect 2950 7098 2956 7100
rect 3012 7098 3036 7100
rect 3092 7098 3116 7100
rect 3172 7098 3196 7100
rect 3252 7098 3258 7100
rect 3012 7046 3014 7098
rect 3194 7046 3196 7098
rect 2950 7044 2956 7046
rect 3012 7044 3036 7046
rect 3092 7044 3116 7046
rect 3172 7044 3196 7046
rect 3252 7044 3258 7046
rect 2950 7035 3258 7044
rect 3424 6724 3476 6730
rect 3424 6666 3476 6672
rect 3148 6656 3200 6662
rect 3148 6598 3200 6604
rect 3160 6497 3188 6598
rect 3146 6488 3202 6497
rect 3146 6423 3202 6432
rect 2950 6012 3258 6021
rect 2950 6010 2956 6012
rect 3012 6010 3036 6012
rect 3092 6010 3116 6012
rect 3172 6010 3196 6012
rect 3252 6010 3258 6012
rect 3012 5958 3014 6010
rect 3194 5958 3196 6010
rect 2950 5956 2956 5958
rect 3012 5956 3036 5958
rect 3092 5956 3116 5958
rect 3172 5956 3196 5958
rect 3252 5956 3258 5958
rect 2950 5947 3258 5956
rect 2950 4924 3258 4933
rect 2950 4922 2956 4924
rect 3012 4922 3036 4924
rect 3092 4922 3116 4924
rect 3172 4922 3196 4924
rect 3252 4922 3258 4924
rect 3012 4870 3014 4922
rect 3194 4870 3196 4922
rect 2950 4868 2956 4870
rect 3012 4868 3036 4870
rect 3092 4868 3116 4870
rect 3172 4868 3196 4870
rect 3252 4868 3258 4870
rect 2950 4859 3258 4868
rect 3240 4820 3292 4826
rect 3240 4762 3292 4768
rect 3252 4185 3280 4762
rect 3238 4176 3294 4185
rect 3238 4111 3294 4120
rect 2872 3936 2924 3942
rect 2872 3878 2924 3884
rect 3332 3936 3384 3942
rect 3332 3878 3384 3884
rect 2780 3732 2832 3738
rect 2780 3674 2832 3680
rect 2700 3590 2820 3618
rect 2792 3534 2820 3590
rect 2884 3534 2912 3878
rect 2950 3836 3258 3845
rect 2950 3834 2956 3836
rect 3012 3834 3036 3836
rect 3092 3834 3116 3836
rect 3172 3834 3196 3836
rect 3252 3834 3258 3836
rect 3012 3782 3014 3834
rect 3194 3782 3196 3834
rect 2950 3780 2956 3782
rect 3012 3780 3036 3782
rect 3092 3780 3116 3782
rect 3172 3780 3196 3782
rect 3252 3780 3258 3782
rect 2950 3771 3258 3780
rect 2780 3528 2832 3534
rect 2780 3470 2832 3476
rect 2872 3528 2924 3534
rect 2872 3470 2924 3476
rect 2136 3188 2188 3194
rect 2136 3130 2188 3136
rect 1860 3052 1912 3058
rect 1860 2994 1912 3000
rect 1872 2854 1900 2994
rect 1492 2848 1544 2854
rect 1492 2790 1544 2796
rect 1860 2848 1912 2854
rect 1860 2790 1912 2796
rect 1504 800 1532 2790
rect 1872 800 1900 2790
rect 2596 2508 2648 2514
rect 2596 2450 2648 2456
rect 2228 2440 2280 2446
rect 2228 2382 2280 2388
rect 2240 800 2268 2382
rect 2608 800 2636 2450
rect 2792 1873 2820 3470
rect 2884 2530 2912 3470
rect 3344 3058 3372 3878
rect 3436 3738 3464 6666
rect 3424 3732 3476 3738
rect 3424 3674 3476 3680
rect 3700 3392 3752 3398
rect 3700 3334 3752 3340
rect 3976 3392 4028 3398
rect 3976 3334 4028 3340
rect 4436 3392 4488 3398
rect 4436 3334 4488 3340
rect 3712 3058 3740 3334
rect 3332 3052 3384 3058
rect 3332 2994 3384 3000
rect 3700 3052 3752 3058
rect 3700 2994 3752 3000
rect 2950 2748 3258 2757
rect 2950 2746 2956 2748
rect 3012 2746 3036 2748
rect 3092 2746 3116 2748
rect 3172 2746 3196 2748
rect 3252 2746 3258 2748
rect 3012 2694 3014 2746
rect 3194 2694 3196 2746
rect 2950 2692 2956 2694
rect 3012 2692 3036 2694
rect 3092 2692 3116 2694
rect 3172 2692 3196 2694
rect 3252 2692 3258 2694
rect 2950 2683 3258 2692
rect 2884 2502 3004 2530
rect 2778 1864 2834 1873
rect 2778 1799 2834 1808
rect 2976 800 3004 2502
rect 3148 2440 3200 2446
rect 3148 2382 3200 2388
rect 3160 2106 3188 2382
rect 3148 2100 3200 2106
rect 3148 2042 3200 2048
rect 3344 800 3372 2994
rect 3712 800 3740 2994
rect 3988 2514 4016 3334
rect 4448 3058 4476 3334
rect 4436 3052 4488 3058
rect 4436 2994 4488 3000
rect 3976 2508 4028 2514
rect 3976 2450 4028 2456
rect 4068 2304 4120 2310
rect 4068 2246 4120 2252
rect 4080 800 4108 2246
rect 4448 800 4476 2994
rect 4632 2922 4660 22066
rect 4724 2990 4752 25638
rect 4816 17626 4844 31214
rect 5816 29572 5868 29578
rect 5816 29514 5868 29520
rect 5724 28484 5776 28490
rect 5724 28426 5776 28432
rect 5540 27532 5592 27538
rect 5540 27474 5592 27480
rect 5448 23792 5500 23798
rect 5448 23734 5500 23740
rect 5356 23656 5408 23662
rect 5460 23610 5488 23734
rect 5408 23604 5488 23610
rect 5356 23598 5488 23604
rect 5368 23582 5488 23598
rect 4896 22568 4948 22574
rect 4896 22510 4948 22516
rect 4908 19514 4936 22510
rect 5264 22160 5316 22166
rect 5264 22102 5316 22108
rect 5276 21010 5304 22102
rect 5264 21004 5316 21010
rect 5316 20964 5396 20992
rect 5264 20946 5316 20952
rect 4988 20936 5040 20942
rect 4988 20878 5040 20884
rect 5000 20602 5028 20878
rect 4988 20596 5040 20602
rect 4988 20538 5040 20544
rect 5368 20058 5396 20964
rect 5460 20602 5488 23582
rect 5552 22794 5580 27474
rect 5736 25362 5764 28426
rect 5724 25356 5776 25362
rect 5724 25298 5776 25304
rect 5724 24744 5776 24750
rect 5724 24686 5776 24692
rect 5632 24608 5684 24614
rect 5632 24550 5684 24556
rect 5644 24410 5672 24550
rect 5632 24404 5684 24410
rect 5632 24346 5684 24352
rect 5644 23866 5672 24346
rect 5632 23860 5684 23866
rect 5632 23802 5684 23808
rect 5632 23656 5684 23662
rect 5632 23598 5684 23604
rect 5644 22982 5672 23598
rect 5736 23526 5764 24686
rect 5724 23520 5776 23526
rect 5724 23462 5776 23468
rect 5632 22976 5684 22982
rect 5632 22918 5684 22924
rect 5552 22766 5672 22794
rect 5540 22636 5592 22642
rect 5540 22578 5592 22584
rect 5552 22234 5580 22578
rect 5540 22228 5592 22234
rect 5540 22170 5592 22176
rect 5448 20596 5500 20602
rect 5448 20538 5500 20544
rect 5356 20052 5408 20058
rect 5356 19994 5408 20000
rect 4896 19508 4948 19514
rect 4896 19450 4948 19456
rect 4816 17598 4936 17626
rect 4908 17542 4936 17598
rect 4804 17536 4856 17542
rect 4804 17478 4856 17484
rect 4896 17536 4948 17542
rect 4896 17478 4948 17484
rect 4816 17202 4844 17478
rect 4804 17196 4856 17202
rect 4804 17138 4856 17144
rect 4908 3670 4936 17478
rect 5644 9654 5672 22766
rect 5736 22574 5764 23462
rect 5724 22568 5776 22574
rect 5724 22510 5776 22516
rect 5724 21344 5776 21350
rect 5724 21286 5776 21292
rect 5736 20262 5764 21286
rect 5828 21010 5856 29514
rect 5816 21004 5868 21010
rect 5816 20946 5868 20952
rect 5724 20256 5776 20262
rect 5724 20198 5776 20204
rect 5736 19514 5764 20198
rect 5724 19508 5776 19514
rect 5724 19450 5776 19456
rect 5724 17604 5776 17610
rect 5724 17546 5776 17552
rect 5736 17270 5764 17546
rect 5724 17264 5776 17270
rect 5724 17206 5776 17212
rect 5632 9648 5684 9654
rect 5632 9590 5684 9596
rect 5724 9648 5776 9654
rect 5724 9590 5776 9596
rect 5172 4752 5224 4758
rect 5172 4694 5224 4700
rect 5080 4208 5132 4214
rect 5080 4150 5132 4156
rect 5092 3738 5120 4150
rect 5080 3732 5132 3738
rect 5080 3674 5132 3680
rect 4896 3664 4948 3670
rect 4896 3606 4948 3612
rect 4804 3392 4856 3398
rect 4804 3334 4856 3340
rect 4712 2984 4764 2990
rect 4712 2926 4764 2932
rect 4620 2916 4672 2922
rect 4620 2858 4672 2864
rect 4816 800 4844 3334
rect 5184 3194 5212 4694
rect 5736 4010 5764 9590
rect 5724 4004 5776 4010
rect 5724 3946 5776 3952
rect 5540 3936 5592 3942
rect 5540 3878 5592 3884
rect 5552 3534 5580 3878
rect 5540 3528 5592 3534
rect 5540 3470 5592 3476
rect 5172 3188 5224 3194
rect 5172 3130 5224 3136
rect 5172 3052 5224 3058
rect 5172 2994 5224 3000
rect 5184 2310 5212 2994
rect 5172 2304 5224 2310
rect 5172 2246 5224 2252
rect 5184 800 5212 2246
rect 5552 800 5580 3470
rect 5920 3194 5948 37402
rect 6104 36378 6132 38218
rect 6288 36632 6316 41414
rect 6368 41064 6420 41070
rect 6368 41006 6420 41012
rect 6380 40526 6408 41006
rect 6368 40520 6420 40526
rect 6368 40462 6420 40468
rect 6380 40118 6408 40462
rect 6368 40112 6420 40118
rect 6368 40054 6420 40060
rect 6288 36604 6408 36632
rect 6092 36372 6144 36378
rect 6092 36314 6144 36320
rect 6092 35148 6144 35154
rect 6092 35090 6144 35096
rect 6104 32842 6132 35090
rect 6092 32836 6144 32842
rect 6092 32778 6144 32784
rect 6104 32026 6132 32778
rect 6092 32020 6144 32026
rect 6092 31962 6144 31968
rect 6380 31142 6408 36604
rect 6472 33318 6500 42570
rect 6828 42560 6880 42566
rect 6828 42502 6880 42508
rect 6644 41608 6696 41614
rect 6644 41550 6696 41556
rect 6552 40384 6604 40390
rect 6552 40326 6604 40332
rect 6564 39030 6592 40326
rect 6552 39024 6604 39030
rect 6552 38966 6604 38972
rect 6564 38214 6592 38966
rect 6552 38208 6604 38214
rect 6552 38150 6604 38156
rect 6564 37194 6592 38150
rect 6552 37188 6604 37194
rect 6552 37130 6604 37136
rect 6564 36106 6592 37130
rect 6552 36100 6604 36106
rect 6552 36042 6604 36048
rect 6564 35766 6592 36042
rect 6552 35760 6604 35766
rect 6552 35702 6604 35708
rect 6564 34950 6592 35702
rect 6552 34944 6604 34950
rect 6552 34886 6604 34892
rect 6564 34746 6592 34886
rect 6552 34740 6604 34746
rect 6552 34682 6604 34688
rect 6460 33312 6512 33318
rect 6460 33254 6512 33260
rect 6368 31136 6420 31142
rect 6368 31078 6420 31084
rect 6656 30598 6684 41550
rect 6736 40452 6788 40458
rect 6736 40394 6788 40400
rect 6748 39574 6776 40394
rect 6736 39568 6788 39574
rect 6736 39510 6788 39516
rect 6748 39098 6776 39510
rect 6736 39092 6788 39098
rect 6736 39034 6788 39040
rect 6736 34536 6788 34542
rect 6736 34478 6788 34484
rect 6748 33998 6776 34478
rect 6736 33992 6788 33998
rect 6736 33934 6788 33940
rect 6840 31346 6868 42502
rect 6932 42362 6960 50730
rect 7024 49978 7052 51954
rect 7116 51950 7144 52550
rect 7196 52080 7248 52086
rect 7196 52022 7248 52028
rect 7104 51944 7156 51950
rect 7104 51886 7156 51892
rect 7104 51400 7156 51406
rect 7104 51342 7156 51348
rect 7012 49972 7064 49978
rect 7012 49914 7064 49920
rect 7116 46714 7144 51342
rect 7104 46708 7156 46714
rect 7104 46650 7156 46656
rect 7104 45280 7156 45286
rect 7104 45222 7156 45228
rect 6920 42356 6972 42362
rect 6920 42298 6972 42304
rect 7116 41414 7144 45222
rect 7208 44538 7236 52022
rect 7392 49978 7420 53518
rect 7852 52562 7880 55186
rect 7950 54428 8258 54437
rect 7950 54426 7956 54428
rect 8012 54426 8036 54428
rect 8092 54426 8116 54428
rect 8172 54426 8196 54428
rect 8252 54426 8258 54428
rect 8012 54374 8014 54426
rect 8194 54374 8196 54426
rect 7950 54372 7956 54374
rect 8012 54372 8036 54374
rect 8092 54372 8116 54374
rect 8172 54372 8196 54374
rect 8252 54372 8258 54374
rect 7950 54363 8258 54372
rect 8312 53650 8340 56200
rect 8484 54256 8536 54262
rect 8484 54198 8536 54204
rect 8300 53644 8352 53650
rect 8300 53586 8352 53592
rect 7950 53340 8258 53349
rect 7950 53338 7956 53340
rect 8012 53338 8036 53340
rect 8092 53338 8116 53340
rect 8172 53338 8196 53340
rect 8252 53338 8258 53340
rect 8012 53286 8014 53338
rect 8194 53286 8196 53338
rect 7950 53284 7956 53286
rect 8012 53284 8036 53286
rect 8092 53284 8116 53286
rect 8172 53284 8196 53286
rect 8252 53284 8258 53286
rect 7950 53275 8258 53284
rect 7840 52556 7892 52562
rect 7840 52498 7892 52504
rect 7950 52252 8258 52261
rect 7950 52250 7956 52252
rect 8012 52250 8036 52252
rect 8092 52250 8116 52252
rect 8172 52250 8196 52252
rect 8252 52250 8258 52252
rect 8012 52198 8014 52250
rect 8194 52198 8196 52250
rect 7950 52196 7956 52198
rect 8012 52196 8036 52198
rect 8092 52196 8116 52198
rect 8172 52196 8196 52198
rect 8252 52196 8258 52198
rect 7950 52187 8258 52196
rect 7748 51400 7800 51406
rect 7748 51342 7800 51348
rect 7760 51074 7788 51342
rect 7950 51164 8258 51173
rect 7950 51162 7956 51164
rect 8012 51162 8036 51164
rect 8092 51162 8116 51164
rect 8172 51162 8196 51164
rect 8252 51162 8258 51164
rect 8012 51110 8014 51162
rect 8194 51110 8196 51162
rect 7950 51108 7956 51110
rect 8012 51108 8036 51110
rect 8092 51108 8116 51110
rect 8172 51108 8196 51110
rect 8252 51108 8258 51110
rect 7950 51099 8258 51108
rect 7760 51046 7880 51074
rect 7748 50244 7800 50250
rect 7748 50186 7800 50192
rect 7380 49972 7432 49978
rect 7380 49914 7432 49920
rect 7656 49904 7708 49910
rect 7656 49846 7708 49852
rect 7380 49836 7432 49842
rect 7380 49778 7432 49784
rect 7288 46572 7340 46578
rect 7288 46514 7340 46520
rect 7196 44532 7248 44538
rect 7196 44474 7248 44480
rect 7300 41818 7328 46514
rect 7392 42566 7420 49778
rect 7472 44872 7524 44878
rect 7472 44814 7524 44820
rect 7380 42560 7432 42566
rect 7380 42502 7432 42508
rect 7380 42356 7432 42362
rect 7380 42298 7432 42304
rect 7288 41812 7340 41818
rect 7288 41754 7340 41760
rect 7116 41386 7236 41414
rect 7104 41200 7156 41206
rect 7104 41142 7156 41148
rect 7116 40458 7144 41142
rect 7104 40452 7156 40458
rect 7104 40394 7156 40400
rect 7104 39976 7156 39982
rect 7104 39918 7156 39924
rect 6920 39500 6972 39506
rect 6920 39442 6972 39448
rect 6932 38554 6960 39442
rect 6920 38548 6972 38554
rect 6920 38490 6972 38496
rect 6932 37330 6960 38490
rect 6920 37324 6972 37330
rect 6920 37266 6972 37272
rect 7116 37194 7144 39918
rect 7208 38350 7236 41386
rect 7392 39846 7420 42298
rect 7380 39840 7432 39846
rect 7380 39782 7432 39788
rect 7380 39432 7432 39438
rect 7380 39374 7432 39380
rect 7196 38344 7248 38350
rect 7196 38286 7248 38292
rect 7392 37806 7420 39374
rect 7380 37800 7432 37806
rect 7380 37742 7432 37748
rect 7196 37324 7248 37330
rect 7196 37266 7248 37272
rect 7104 37188 7156 37194
rect 7104 37130 7156 37136
rect 7012 36236 7064 36242
rect 7012 36178 7064 36184
rect 7024 35086 7052 36178
rect 7012 35080 7064 35086
rect 7012 35022 7064 35028
rect 7024 34542 7052 35022
rect 7116 35018 7144 37130
rect 7208 35834 7236 37266
rect 7392 36038 7420 37742
rect 7484 37670 7512 44814
rect 7564 42696 7616 42702
rect 7564 42638 7616 42644
rect 7576 41414 7604 42638
rect 7668 42566 7696 49846
rect 7760 44538 7788 50186
rect 7748 44532 7800 44538
rect 7748 44474 7800 44480
rect 7748 44396 7800 44402
rect 7748 44338 7800 44344
rect 7656 42560 7708 42566
rect 7656 42502 7708 42508
rect 7576 41386 7696 41414
rect 7564 41268 7616 41274
rect 7564 41210 7616 41216
rect 7576 40186 7604 41210
rect 7564 40180 7616 40186
rect 7564 40122 7616 40128
rect 7472 37664 7524 37670
rect 7472 37606 7524 37612
rect 7484 37466 7512 37606
rect 7472 37460 7524 37466
rect 7472 37402 7524 37408
rect 7564 36712 7616 36718
rect 7564 36654 7616 36660
rect 7576 36242 7604 36654
rect 7564 36236 7616 36242
rect 7564 36178 7616 36184
rect 7380 36032 7432 36038
rect 7380 35974 7432 35980
rect 7196 35828 7248 35834
rect 7196 35770 7248 35776
rect 7104 35012 7156 35018
rect 7104 34954 7156 34960
rect 7116 34626 7144 34954
rect 7208 34746 7236 35770
rect 7288 34944 7340 34950
rect 7288 34886 7340 34892
rect 7196 34740 7248 34746
rect 7196 34682 7248 34688
rect 7300 34678 7328 34886
rect 7288 34672 7340 34678
rect 7116 34598 7236 34626
rect 7288 34614 7340 34620
rect 7012 34536 7064 34542
rect 7012 34478 7064 34484
rect 7104 32836 7156 32842
rect 7104 32778 7156 32784
rect 7116 32570 7144 32778
rect 7104 32564 7156 32570
rect 7104 32506 7156 32512
rect 6920 32292 6972 32298
rect 6920 32234 6972 32240
rect 6932 31822 6960 32234
rect 6920 31816 6972 31822
rect 6920 31758 6972 31764
rect 7116 31754 7144 32506
rect 7208 31793 7236 34598
rect 7300 34202 7328 34614
rect 7288 34196 7340 34202
rect 7288 34138 7340 34144
rect 7288 33924 7340 33930
rect 7288 33866 7340 33872
rect 7300 33114 7328 33866
rect 7288 33108 7340 33114
rect 7288 33050 7340 33056
rect 7392 32994 7420 35974
rect 7668 35290 7696 41386
rect 7760 37126 7788 44338
rect 7852 43926 7880 51046
rect 8300 50924 8352 50930
rect 8300 50866 8352 50872
rect 7950 50076 8258 50085
rect 7950 50074 7956 50076
rect 8012 50074 8036 50076
rect 8092 50074 8116 50076
rect 8172 50074 8196 50076
rect 8252 50074 8258 50076
rect 8012 50022 8014 50074
rect 8194 50022 8196 50074
rect 7950 50020 7956 50022
rect 8012 50020 8036 50022
rect 8092 50020 8116 50022
rect 8172 50020 8196 50022
rect 8252 50020 8258 50022
rect 7950 50011 8258 50020
rect 7950 48988 8258 48997
rect 7950 48986 7956 48988
rect 8012 48986 8036 48988
rect 8092 48986 8116 48988
rect 8172 48986 8196 48988
rect 8252 48986 8258 48988
rect 8012 48934 8014 48986
rect 8194 48934 8196 48986
rect 7950 48932 7956 48934
rect 8012 48932 8036 48934
rect 8092 48932 8116 48934
rect 8172 48932 8196 48934
rect 8252 48932 8258 48934
rect 7950 48923 8258 48932
rect 7950 47900 8258 47909
rect 7950 47898 7956 47900
rect 8012 47898 8036 47900
rect 8092 47898 8116 47900
rect 8172 47898 8196 47900
rect 8252 47898 8258 47900
rect 8012 47846 8014 47898
rect 8194 47846 8196 47898
rect 7950 47844 7956 47846
rect 8012 47844 8036 47846
rect 8092 47844 8116 47846
rect 8172 47844 8196 47846
rect 8252 47844 8258 47846
rect 7950 47835 8258 47844
rect 7950 46812 8258 46821
rect 7950 46810 7956 46812
rect 8012 46810 8036 46812
rect 8092 46810 8116 46812
rect 8172 46810 8196 46812
rect 8252 46810 8258 46812
rect 8012 46758 8014 46810
rect 8194 46758 8196 46810
rect 7950 46756 7956 46758
rect 8012 46756 8036 46758
rect 8092 46756 8116 46758
rect 8172 46756 8196 46758
rect 8252 46756 8258 46758
rect 7950 46747 8258 46756
rect 7950 45724 8258 45733
rect 7950 45722 7956 45724
rect 8012 45722 8036 45724
rect 8092 45722 8116 45724
rect 8172 45722 8196 45724
rect 8252 45722 8258 45724
rect 8012 45670 8014 45722
rect 8194 45670 8196 45722
rect 7950 45668 7956 45670
rect 8012 45668 8036 45670
rect 8092 45668 8116 45670
rect 8172 45668 8196 45670
rect 8252 45668 8258 45670
rect 7950 45659 8258 45668
rect 8312 45286 8340 50866
rect 8392 45484 8444 45490
rect 8392 45426 8444 45432
rect 8300 45280 8352 45286
rect 8300 45222 8352 45228
rect 7950 44636 8258 44645
rect 7950 44634 7956 44636
rect 8012 44634 8036 44636
rect 8092 44634 8116 44636
rect 8172 44634 8196 44636
rect 8252 44634 8258 44636
rect 8012 44582 8014 44634
rect 8194 44582 8196 44634
rect 7950 44580 7956 44582
rect 8012 44580 8036 44582
rect 8092 44580 8116 44582
rect 8172 44580 8196 44582
rect 8252 44580 8258 44582
rect 7950 44571 8258 44580
rect 8300 44328 8352 44334
rect 8300 44270 8352 44276
rect 7840 43920 7892 43926
rect 7840 43862 7892 43868
rect 7950 43548 8258 43557
rect 7950 43546 7956 43548
rect 8012 43546 8036 43548
rect 8092 43546 8116 43548
rect 8172 43546 8196 43548
rect 8252 43546 8258 43548
rect 8012 43494 8014 43546
rect 8194 43494 8196 43546
rect 7950 43492 7956 43494
rect 8012 43492 8036 43494
rect 8092 43492 8116 43494
rect 8172 43492 8196 43494
rect 8252 43492 8258 43494
rect 7950 43483 8258 43492
rect 8312 42770 8340 44270
rect 8300 42764 8352 42770
rect 8300 42706 8352 42712
rect 7950 42460 8258 42469
rect 7950 42458 7956 42460
rect 8012 42458 8036 42460
rect 8092 42458 8116 42460
rect 8172 42458 8196 42460
rect 8252 42458 8258 42460
rect 8012 42406 8014 42458
rect 8194 42406 8196 42458
rect 7950 42404 7956 42406
rect 8012 42404 8036 42406
rect 8092 42404 8116 42406
rect 8172 42404 8196 42406
rect 8252 42404 8258 42406
rect 7950 42395 8258 42404
rect 8300 41608 8352 41614
rect 8300 41550 8352 41556
rect 7950 41372 8258 41381
rect 7950 41370 7956 41372
rect 8012 41370 8036 41372
rect 8092 41370 8116 41372
rect 8172 41370 8196 41372
rect 8252 41370 8258 41372
rect 8012 41318 8014 41370
rect 8194 41318 8196 41370
rect 7950 41316 7956 41318
rect 8012 41316 8036 41318
rect 8092 41316 8116 41318
rect 8172 41316 8196 41318
rect 8252 41316 8258 41318
rect 7950 41307 8258 41316
rect 7840 41064 7892 41070
rect 7840 41006 7892 41012
rect 7852 40594 7880 41006
rect 7840 40588 7892 40594
rect 7840 40530 7892 40536
rect 7852 38418 7880 40530
rect 7950 40284 8258 40293
rect 7950 40282 7956 40284
rect 8012 40282 8036 40284
rect 8092 40282 8116 40284
rect 8172 40282 8196 40284
rect 8252 40282 8258 40284
rect 8012 40230 8014 40282
rect 8194 40230 8196 40282
rect 7950 40228 7956 40230
rect 8012 40228 8036 40230
rect 8092 40228 8116 40230
rect 8172 40228 8196 40230
rect 8252 40228 8258 40230
rect 7950 40219 8258 40228
rect 8208 39840 8260 39846
rect 8208 39782 8260 39788
rect 8220 39438 8248 39782
rect 8208 39432 8260 39438
rect 8208 39374 8260 39380
rect 7950 39196 8258 39205
rect 7950 39194 7956 39196
rect 8012 39194 8036 39196
rect 8092 39194 8116 39196
rect 8172 39194 8196 39196
rect 8252 39194 8258 39196
rect 8012 39142 8014 39194
rect 8194 39142 8196 39194
rect 7950 39140 7956 39142
rect 8012 39140 8036 39142
rect 8092 39140 8116 39142
rect 8172 39140 8196 39142
rect 8252 39140 8258 39142
rect 7950 39131 8258 39140
rect 8312 38554 8340 41550
rect 8404 39642 8432 45426
rect 8496 44470 8524 54198
rect 8680 53038 8708 56200
rect 9048 53582 9076 56200
rect 9416 54126 9444 56200
rect 9404 54120 9456 54126
rect 9404 54062 9456 54068
rect 9036 53576 9088 53582
rect 9036 53518 9088 53524
rect 9680 53576 9732 53582
rect 9680 53518 9732 53524
rect 9128 53100 9180 53106
rect 9128 53042 9180 53048
rect 9404 53100 9456 53106
rect 9404 53042 9456 53048
rect 8668 53032 8720 53038
rect 8668 52974 8720 52980
rect 8576 50924 8628 50930
rect 8576 50866 8628 50872
rect 8588 45354 8616 50866
rect 8668 50312 8720 50318
rect 8668 50254 8720 50260
rect 8576 45348 8628 45354
rect 8576 45290 8628 45296
rect 8484 44464 8536 44470
rect 8484 44406 8536 44412
rect 8680 43450 8708 50254
rect 9036 49156 9088 49162
rect 9036 49098 9088 49104
rect 8760 44736 8812 44742
rect 8760 44678 8812 44684
rect 8772 44402 8800 44678
rect 9048 44538 9076 49098
rect 9036 44532 9088 44538
rect 9036 44474 9088 44480
rect 8760 44396 8812 44402
rect 8760 44338 8812 44344
rect 8668 43444 8720 43450
rect 8668 43386 8720 43392
rect 8484 43104 8536 43110
rect 8484 43046 8536 43052
rect 8496 42702 8524 43046
rect 8484 42696 8536 42702
rect 8484 42638 8536 42644
rect 8576 42288 8628 42294
rect 8576 42230 8628 42236
rect 8484 42152 8536 42158
rect 8484 42094 8536 42100
rect 8496 41682 8524 42094
rect 8484 41676 8536 41682
rect 8484 41618 8536 41624
rect 8496 41274 8524 41618
rect 8484 41268 8536 41274
rect 8484 41210 8536 41216
rect 8588 40934 8616 42230
rect 8680 42022 8708 43386
rect 8668 42016 8720 42022
rect 8668 41958 8720 41964
rect 8576 40928 8628 40934
rect 8576 40870 8628 40876
rect 8588 40730 8616 40870
rect 8576 40724 8628 40730
rect 8576 40666 8628 40672
rect 8588 40390 8616 40666
rect 8576 40384 8628 40390
rect 8576 40326 8628 40332
rect 8392 39636 8444 39642
rect 8392 39578 8444 39584
rect 8484 39296 8536 39302
rect 8484 39238 8536 39244
rect 8300 38548 8352 38554
rect 8300 38490 8352 38496
rect 8116 38480 8168 38486
rect 8116 38422 8168 38428
rect 7840 38412 7892 38418
rect 7840 38354 7892 38360
rect 8128 38350 8156 38422
rect 8116 38344 8168 38350
rect 8116 38286 8168 38292
rect 8300 38208 8352 38214
rect 8300 38150 8352 38156
rect 7950 38108 8258 38117
rect 7950 38106 7956 38108
rect 8012 38106 8036 38108
rect 8092 38106 8116 38108
rect 8172 38106 8196 38108
rect 8252 38106 8258 38108
rect 8012 38054 8014 38106
rect 8194 38054 8196 38106
rect 7950 38052 7956 38054
rect 8012 38052 8036 38054
rect 8092 38052 8116 38054
rect 8172 38052 8196 38054
rect 8252 38052 8258 38054
rect 7950 38043 8258 38052
rect 8312 37874 8340 38150
rect 8300 37868 8352 37874
rect 8300 37810 8352 37816
rect 8312 37466 8340 37810
rect 8300 37460 8352 37466
rect 8300 37402 8352 37408
rect 7748 37120 7800 37126
rect 7748 37062 7800 37068
rect 7950 37020 8258 37029
rect 7950 37018 7956 37020
rect 8012 37018 8036 37020
rect 8092 37018 8116 37020
rect 8172 37018 8196 37020
rect 8252 37018 8258 37020
rect 8012 36966 8014 37018
rect 8194 36966 8196 37018
rect 7950 36964 7956 36966
rect 8012 36964 8036 36966
rect 8092 36964 8116 36966
rect 8172 36964 8196 36966
rect 8252 36964 8258 36966
rect 7950 36955 8258 36964
rect 8312 36854 8340 37402
rect 8300 36848 8352 36854
rect 8300 36790 8352 36796
rect 8312 36378 8340 36790
rect 8300 36372 8352 36378
rect 8300 36314 8352 36320
rect 7950 35932 8258 35941
rect 7950 35930 7956 35932
rect 8012 35930 8036 35932
rect 8092 35930 8116 35932
rect 8172 35930 8196 35932
rect 8252 35930 8258 35932
rect 8012 35878 8014 35930
rect 8194 35878 8196 35930
rect 7950 35876 7956 35878
rect 8012 35876 8036 35878
rect 8092 35876 8116 35878
rect 8172 35876 8196 35878
rect 8252 35876 8258 35878
rect 7950 35867 8258 35876
rect 7656 35284 7708 35290
rect 7656 35226 7708 35232
rect 7840 34944 7892 34950
rect 7840 34886 7892 34892
rect 7656 34536 7708 34542
rect 7656 34478 7708 34484
rect 7564 33652 7616 33658
rect 7564 33594 7616 33600
rect 7300 32966 7420 32994
rect 7300 32026 7328 32966
rect 7472 32360 7524 32366
rect 7472 32302 7524 32308
rect 7288 32020 7340 32026
rect 7288 31962 7340 31968
rect 7194 31784 7250 31793
rect 7104 31748 7156 31754
rect 7194 31719 7250 31728
rect 7104 31690 7156 31696
rect 6828 31340 6880 31346
rect 6828 31282 6880 31288
rect 7104 31340 7156 31346
rect 7104 31282 7156 31288
rect 6644 30592 6696 30598
rect 6644 30534 6696 30540
rect 7012 30592 7064 30598
rect 7012 30534 7064 30540
rect 6920 28416 6972 28422
rect 6920 28358 6972 28364
rect 6276 28076 6328 28082
rect 6276 28018 6328 28024
rect 6000 27056 6052 27062
rect 6000 26998 6052 27004
rect 6012 26450 6040 26998
rect 6288 26450 6316 28018
rect 6932 28014 6960 28358
rect 6920 28008 6972 28014
rect 6920 27950 6972 27956
rect 6920 27328 6972 27334
rect 6920 27270 6972 27276
rect 6932 26450 6960 27270
rect 6000 26444 6052 26450
rect 6276 26444 6328 26450
rect 6052 26404 6224 26432
rect 6000 26386 6052 26392
rect 6000 25356 6052 25362
rect 6000 25298 6052 25304
rect 6012 12434 6040 25298
rect 6196 19718 6224 26404
rect 6276 26386 6328 26392
rect 6920 26444 6972 26450
rect 6920 26386 6972 26392
rect 6288 25362 6316 26386
rect 7024 25702 7052 30534
rect 7116 27282 7144 31282
rect 7300 30802 7328 31962
rect 7378 31784 7434 31793
rect 7378 31719 7434 31728
rect 7392 31210 7420 31719
rect 7380 31204 7432 31210
rect 7380 31146 7432 31152
rect 7288 30796 7340 30802
rect 7288 30738 7340 30744
rect 7484 30734 7512 32302
rect 7576 31906 7604 33594
rect 7668 32212 7696 34478
rect 7748 33992 7800 33998
rect 7748 33934 7800 33940
rect 7760 33454 7788 33934
rect 7748 33448 7800 33454
rect 7748 33390 7800 33396
rect 7760 32978 7788 33390
rect 7748 32972 7800 32978
rect 7748 32914 7800 32920
rect 7760 32366 7788 32914
rect 7748 32360 7800 32366
rect 7748 32302 7800 32308
rect 7668 32184 7788 32212
rect 7576 31878 7696 31906
rect 7564 31816 7616 31822
rect 7564 31758 7616 31764
rect 7472 30728 7524 30734
rect 7472 30670 7524 30676
rect 7576 30394 7604 31758
rect 7668 31482 7696 31878
rect 7656 31476 7708 31482
rect 7656 31418 7708 31424
rect 7760 30938 7788 32184
rect 7852 31958 7880 34886
rect 7950 34844 8258 34853
rect 7950 34842 7956 34844
rect 8012 34842 8036 34844
rect 8092 34842 8116 34844
rect 8172 34842 8196 34844
rect 8252 34842 8258 34844
rect 8012 34790 8014 34842
rect 8194 34790 8196 34842
rect 7950 34788 7956 34790
rect 8012 34788 8036 34790
rect 8092 34788 8116 34790
rect 8172 34788 8196 34790
rect 8252 34788 8258 34790
rect 7950 34779 8258 34788
rect 8496 34746 8524 39238
rect 8576 38888 8628 38894
rect 8576 38830 8628 38836
rect 8588 38350 8616 38830
rect 8576 38344 8628 38350
rect 8576 38286 8628 38292
rect 8772 35873 8800 44338
rect 9140 43994 9168 53042
rect 9416 50454 9444 53042
rect 9496 52488 9548 52494
rect 9496 52430 9548 52436
rect 9588 52488 9640 52494
rect 9588 52430 9640 52436
rect 9404 50448 9456 50454
rect 9404 50390 9456 50396
rect 9404 49292 9456 49298
rect 9404 49234 9456 49240
rect 9220 44532 9272 44538
rect 9220 44474 9272 44480
rect 9128 43988 9180 43994
rect 9128 43930 9180 43936
rect 9128 43648 9180 43654
rect 9128 43590 9180 43596
rect 9036 42696 9088 42702
rect 9036 42638 9088 42644
rect 9048 36310 9076 42638
rect 9140 37466 9168 43590
rect 9232 42770 9260 44474
rect 9416 44402 9444 49234
rect 9404 44396 9456 44402
rect 9404 44338 9456 44344
rect 9220 42764 9272 42770
rect 9220 42706 9272 42712
rect 9232 41414 9260 42706
rect 9416 42362 9444 44338
rect 9508 43926 9536 52430
rect 9600 49910 9628 52430
rect 9692 51950 9720 53518
rect 9784 52562 9812 56200
rect 9864 54188 9916 54194
rect 9864 54130 9916 54136
rect 9772 52556 9824 52562
rect 9772 52498 9824 52504
rect 9680 51944 9732 51950
rect 9680 51886 9732 51892
rect 9876 51066 9904 54130
rect 10152 53038 10180 56200
rect 10520 53650 10548 56200
rect 10888 54262 10916 56200
rect 10876 54256 10928 54262
rect 10876 54198 10928 54204
rect 10508 53644 10560 53650
rect 10508 53586 10560 53592
rect 11060 53576 11112 53582
rect 11060 53518 11112 53524
rect 10692 53100 10744 53106
rect 10692 53042 10744 53048
rect 10140 53032 10192 53038
rect 10140 52974 10192 52980
rect 10140 52012 10192 52018
rect 10140 51954 10192 51960
rect 9864 51060 9916 51066
rect 9864 51002 9916 51008
rect 9956 50924 10008 50930
rect 9956 50866 10008 50872
rect 9588 49904 9640 49910
rect 9588 49846 9640 49852
rect 9864 45960 9916 45966
rect 9864 45902 9916 45908
rect 9772 45484 9824 45490
rect 9772 45426 9824 45432
rect 9680 44736 9732 44742
rect 9678 44704 9680 44713
rect 9732 44704 9734 44713
rect 9678 44639 9734 44648
rect 9496 43920 9548 43926
rect 9496 43862 9548 43868
rect 9680 42696 9732 42702
rect 9680 42638 9732 42644
rect 9496 42628 9548 42634
rect 9496 42570 9548 42576
rect 9404 42356 9456 42362
rect 9404 42298 9456 42304
rect 9232 41386 9352 41414
rect 9324 39522 9352 41386
rect 9416 41070 9444 42298
rect 9404 41064 9456 41070
rect 9404 41006 9456 41012
rect 9416 40118 9444 41006
rect 9404 40112 9456 40118
rect 9404 40054 9456 40060
rect 9324 39494 9444 39522
rect 9312 39364 9364 39370
rect 9312 39306 9364 39312
rect 9324 38554 9352 39306
rect 9312 38548 9364 38554
rect 9312 38490 9364 38496
rect 9312 37936 9364 37942
rect 9312 37878 9364 37884
rect 9128 37460 9180 37466
rect 9128 37402 9180 37408
rect 9324 36922 9352 37878
rect 9416 37806 9444 39494
rect 9404 37800 9456 37806
rect 9404 37742 9456 37748
rect 9508 36922 9536 42570
rect 9588 41472 9640 41478
rect 9588 41414 9640 41420
rect 9600 38418 9628 41414
rect 9692 41274 9720 42638
rect 9680 41268 9732 41274
rect 9680 41210 9732 41216
rect 9680 40044 9732 40050
rect 9680 39986 9732 39992
rect 9588 38412 9640 38418
rect 9588 38354 9640 38360
rect 9692 37874 9720 39986
rect 9784 39098 9812 45426
rect 9876 42566 9904 45902
rect 9968 45354 9996 50866
rect 10048 49224 10100 49230
rect 10048 49166 10100 49172
rect 9956 45348 10008 45354
rect 9956 45290 10008 45296
rect 10060 44538 10088 49166
rect 10152 45082 10180 51954
rect 10704 51066 10732 53042
rect 10692 51060 10744 51066
rect 10692 51002 10744 51008
rect 10968 47048 11020 47054
rect 10968 46990 11020 46996
rect 10140 45076 10192 45082
rect 10140 45018 10192 45024
rect 10692 44872 10744 44878
rect 10692 44814 10744 44820
rect 10048 44532 10100 44538
rect 10048 44474 10100 44480
rect 10060 43382 10088 44474
rect 10704 43790 10732 44814
rect 10508 43784 10560 43790
rect 10692 43784 10744 43790
rect 10560 43732 10640 43738
rect 10508 43726 10640 43732
rect 10692 43726 10744 43732
rect 10520 43710 10640 43726
rect 10048 43376 10100 43382
rect 10048 43318 10100 43324
rect 9864 42560 9916 42566
rect 9864 42502 9916 42508
rect 9876 41414 9904 42502
rect 10060 42362 10088 43318
rect 10048 42356 10100 42362
rect 10048 42298 10100 42304
rect 9876 41386 9996 41414
rect 9864 40724 9916 40730
rect 9864 40666 9916 40672
rect 9876 39574 9904 40666
rect 9864 39568 9916 39574
rect 9864 39510 9916 39516
rect 9968 39370 9996 41386
rect 10232 40384 10284 40390
rect 10232 40326 10284 40332
rect 10048 40180 10100 40186
rect 10048 40122 10100 40128
rect 9956 39364 10008 39370
rect 9956 39306 10008 39312
rect 9864 39296 9916 39302
rect 9864 39238 9916 39244
rect 9772 39092 9824 39098
rect 9772 39034 9824 39040
rect 9876 38418 9904 39238
rect 9864 38412 9916 38418
rect 9864 38354 9916 38360
rect 9864 38208 9916 38214
rect 9864 38150 9916 38156
rect 9680 37868 9732 37874
rect 9680 37810 9732 37816
rect 9876 36961 9904 38150
rect 10060 37262 10088 40122
rect 10244 40050 10272 40326
rect 10232 40044 10284 40050
rect 10232 39986 10284 39992
rect 10244 39846 10272 39986
rect 10232 39840 10284 39846
rect 10232 39782 10284 39788
rect 10140 38412 10192 38418
rect 10140 38354 10192 38360
rect 10152 38282 10180 38354
rect 10140 38276 10192 38282
rect 10140 38218 10192 38224
rect 9956 37256 10008 37262
rect 9956 37198 10008 37204
rect 10048 37256 10100 37262
rect 10048 37198 10100 37204
rect 9862 36952 9918 36961
rect 9128 36916 9180 36922
rect 9128 36858 9180 36864
rect 9312 36916 9364 36922
rect 9312 36858 9364 36864
rect 9496 36916 9548 36922
rect 9862 36887 9918 36896
rect 9496 36858 9548 36864
rect 9036 36304 9088 36310
rect 8956 36252 9036 36258
rect 8956 36246 9088 36252
rect 8956 36230 9076 36246
rect 8758 35864 8814 35873
rect 8758 35799 8814 35808
rect 8484 34740 8536 34746
rect 8484 34682 8536 34688
rect 8484 34196 8536 34202
rect 8484 34138 8536 34144
rect 7950 33756 8258 33765
rect 7950 33754 7956 33756
rect 8012 33754 8036 33756
rect 8092 33754 8116 33756
rect 8172 33754 8196 33756
rect 8252 33754 8258 33756
rect 8012 33702 8014 33754
rect 8194 33702 8196 33754
rect 7950 33700 7956 33702
rect 8012 33700 8036 33702
rect 8092 33700 8116 33702
rect 8172 33700 8196 33702
rect 8252 33700 8258 33702
rect 7950 33691 8258 33700
rect 8496 33590 8524 34138
rect 8484 33584 8536 33590
rect 8484 33526 8536 33532
rect 8300 32904 8352 32910
rect 8300 32846 8352 32852
rect 7950 32668 8258 32677
rect 7950 32666 7956 32668
rect 8012 32666 8036 32668
rect 8092 32666 8116 32668
rect 8172 32666 8196 32668
rect 8252 32666 8258 32668
rect 8012 32614 8014 32666
rect 8194 32614 8196 32666
rect 7950 32612 7956 32614
rect 8012 32612 8036 32614
rect 8092 32612 8116 32614
rect 8172 32612 8196 32614
rect 8252 32612 8258 32614
rect 7950 32603 8258 32612
rect 7840 31952 7892 31958
rect 7840 31894 7892 31900
rect 8312 31890 8340 32846
rect 8496 32842 8524 33526
rect 8484 32836 8536 32842
rect 8484 32778 8536 32784
rect 8496 32502 8524 32778
rect 8484 32496 8536 32502
rect 8484 32438 8536 32444
rect 8300 31884 8352 31890
rect 8300 31826 8352 31832
rect 7840 31680 7892 31686
rect 7840 31622 7892 31628
rect 7852 31482 7880 31622
rect 7950 31580 8258 31589
rect 7950 31578 7956 31580
rect 8012 31578 8036 31580
rect 8092 31578 8116 31580
rect 8172 31578 8196 31580
rect 8252 31578 8258 31580
rect 8012 31526 8014 31578
rect 8194 31526 8196 31578
rect 7950 31524 7956 31526
rect 8012 31524 8036 31526
rect 8092 31524 8116 31526
rect 8172 31524 8196 31526
rect 8252 31524 8258 31526
rect 7950 31515 8258 31524
rect 7840 31476 7892 31482
rect 7840 31418 7892 31424
rect 7748 30932 7800 30938
rect 7748 30874 7800 30880
rect 7950 30492 8258 30501
rect 7950 30490 7956 30492
rect 8012 30490 8036 30492
rect 8092 30490 8116 30492
rect 8172 30490 8196 30492
rect 8252 30490 8258 30492
rect 8012 30438 8014 30490
rect 8194 30438 8196 30490
rect 7950 30436 7956 30438
rect 8012 30436 8036 30438
rect 8092 30436 8116 30438
rect 8172 30436 8196 30438
rect 8252 30436 8258 30438
rect 7950 30427 8258 30436
rect 7564 30388 7616 30394
rect 7564 30330 7616 30336
rect 8772 29578 8800 35799
rect 8760 29572 8812 29578
rect 8760 29514 8812 29520
rect 7950 29404 8258 29413
rect 7950 29402 7956 29404
rect 8012 29402 8036 29404
rect 8092 29402 8116 29404
rect 8172 29402 8196 29404
rect 8252 29402 8258 29404
rect 8012 29350 8014 29402
rect 8194 29350 8196 29402
rect 7950 29348 7956 29350
rect 8012 29348 8036 29350
rect 8092 29348 8116 29350
rect 8172 29348 8196 29350
rect 8252 29348 8258 29350
rect 7950 29339 8258 29348
rect 8208 29300 8260 29306
rect 8208 29242 8260 29248
rect 7380 28756 7432 28762
rect 7380 28698 7432 28704
rect 7288 28008 7340 28014
rect 7288 27950 7340 27956
rect 7116 27254 7236 27282
rect 7208 26994 7236 27254
rect 7196 26988 7248 26994
rect 7196 26930 7248 26936
rect 7208 26790 7236 26930
rect 7300 26858 7328 27950
rect 7288 26852 7340 26858
rect 7288 26794 7340 26800
rect 7196 26784 7248 26790
rect 7196 26726 7248 26732
rect 7012 25696 7064 25702
rect 7012 25638 7064 25644
rect 6276 25356 6328 25362
rect 6276 25298 6328 25304
rect 6288 24818 6316 25298
rect 6276 24812 6328 24818
rect 6276 24754 6328 24760
rect 6288 23730 6316 24754
rect 6736 23860 6788 23866
rect 6736 23802 6788 23808
rect 6276 23724 6328 23730
rect 6276 23666 6328 23672
rect 6644 23656 6696 23662
rect 6644 23598 6696 23604
rect 6552 23520 6604 23526
rect 6552 23462 6604 23468
rect 6368 23180 6420 23186
rect 6368 23122 6420 23128
rect 6380 22094 6408 23122
rect 6380 22066 6500 22094
rect 6472 21690 6500 22066
rect 6564 22030 6592 23462
rect 6552 22024 6604 22030
rect 6552 21966 6604 21972
rect 6460 21684 6512 21690
rect 6460 21626 6512 21632
rect 6276 21004 6328 21010
rect 6276 20946 6328 20952
rect 6184 19712 6236 19718
rect 6184 19654 6236 19660
rect 6288 19258 6316 20946
rect 6368 20936 6420 20942
rect 6368 20878 6420 20884
rect 6380 20262 6408 20878
rect 6368 20256 6420 20262
rect 6368 20198 6420 20204
rect 6380 19786 6408 20198
rect 6368 19780 6420 19786
rect 6368 19722 6420 19728
rect 6380 19446 6408 19722
rect 6368 19440 6420 19446
rect 6368 19382 6420 19388
rect 6460 19372 6512 19378
rect 6460 19314 6512 19320
rect 6288 19230 6408 19258
rect 6276 18216 6328 18222
rect 6276 18158 6328 18164
rect 6288 17746 6316 18158
rect 6276 17740 6328 17746
rect 6276 17682 6328 17688
rect 6092 17128 6144 17134
rect 6092 17070 6144 17076
rect 6104 16794 6132 17070
rect 6092 16788 6144 16794
rect 6092 16730 6144 16736
rect 6288 16658 6316 17682
rect 6276 16652 6328 16658
rect 6276 16594 6328 16600
rect 6288 15366 6316 16594
rect 6276 15360 6328 15366
rect 6276 15302 6328 15308
rect 6380 12434 6408 19230
rect 6472 16250 6500 19314
rect 6552 17604 6604 17610
rect 6552 17546 6604 17552
rect 6564 17134 6592 17546
rect 6552 17128 6604 17134
rect 6552 17070 6604 17076
rect 6460 16244 6512 16250
rect 6460 16186 6512 16192
rect 6564 15706 6592 17070
rect 6552 15700 6604 15706
rect 6552 15642 6604 15648
rect 6012 12406 6224 12434
rect 6380 12406 6500 12434
rect 6196 6914 6224 12406
rect 6472 6914 6500 12406
rect 6196 6886 6316 6914
rect 6288 6662 6316 6886
rect 6380 6886 6500 6914
rect 6276 6656 6328 6662
rect 6276 6598 6328 6604
rect 6380 4826 6408 6886
rect 6368 4820 6420 4826
rect 6368 4762 6420 4768
rect 6656 3738 6684 23598
rect 6748 23594 6776 23802
rect 6736 23588 6788 23594
rect 6736 23530 6788 23536
rect 7012 23588 7064 23594
rect 7012 23530 7064 23536
rect 6748 23050 6776 23530
rect 7024 23186 7052 23530
rect 7012 23180 7064 23186
rect 7012 23122 7064 23128
rect 6736 23044 6788 23050
rect 6736 22986 6788 22992
rect 6828 22976 6880 22982
rect 6828 22918 6880 22924
rect 6840 22098 6868 22918
rect 6828 22092 6880 22098
rect 6828 22034 6880 22040
rect 6840 21622 6868 22034
rect 6828 21616 6880 21622
rect 6828 21558 6880 21564
rect 6920 21412 6972 21418
rect 6920 21354 6972 21360
rect 6932 20806 6960 21354
rect 7024 21078 7052 23122
rect 7104 23044 7156 23050
rect 7104 22986 7156 22992
rect 7012 21072 7064 21078
rect 7012 21014 7064 21020
rect 7116 20942 7144 22986
rect 7104 20936 7156 20942
rect 7104 20878 7156 20884
rect 6920 20800 6972 20806
rect 6920 20742 6972 20748
rect 6828 19916 6880 19922
rect 6828 19858 6880 19864
rect 6736 19712 6788 19718
rect 6736 19654 6788 19660
rect 6748 12374 6776 19654
rect 6840 19378 6868 19858
rect 6828 19372 6880 19378
rect 6828 19314 6880 19320
rect 6840 18222 6868 19314
rect 6932 19310 6960 20742
rect 7208 20466 7236 26726
rect 7392 24410 7420 28698
rect 8024 28620 8076 28626
rect 7852 28580 8024 28608
rect 7472 28484 7524 28490
rect 7472 28426 7524 28432
rect 7484 27402 7512 28426
rect 7564 28416 7616 28422
rect 7564 28358 7616 28364
rect 7472 27396 7524 27402
rect 7472 27338 7524 27344
rect 7576 25838 7604 28358
rect 7852 28218 7880 28580
rect 8024 28562 8076 28568
rect 8220 28490 8248 29242
rect 8576 28688 8628 28694
rect 8576 28630 8628 28636
rect 8208 28484 8260 28490
rect 8208 28426 8260 28432
rect 7950 28316 8258 28325
rect 7950 28314 7956 28316
rect 8012 28314 8036 28316
rect 8092 28314 8116 28316
rect 8172 28314 8196 28316
rect 8252 28314 8258 28316
rect 8012 28262 8014 28314
rect 8194 28262 8196 28314
rect 7950 28260 7956 28262
rect 8012 28260 8036 28262
rect 8092 28260 8116 28262
rect 8172 28260 8196 28262
rect 8252 28260 8258 28262
rect 7950 28251 8258 28260
rect 8588 28218 8616 28630
rect 8956 28558 8984 36230
rect 9036 34944 9088 34950
rect 9036 34886 9088 34892
rect 9048 33386 9076 34886
rect 9140 34202 9168 36858
rect 9404 36712 9456 36718
rect 9404 36654 9456 36660
rect 9496 36712 9548 36718
rect 9496 36654 9548 36660
rect 9312 36372 9364 36378
rect 9312 36314 9364 36320
rect 9324 35766 9352 36314
rect 9416 35834 9444 36654
rect 9404 35828 9456 35834
rect 9404 35770 9456 35776
rect 9312 35760 9364 35766
rect 9312 35702 9364 35708
rect 9416 35154 9444 35770
rect 9404 35148 9456 35154
rect 9404 35090 9456 35096
rect 9128 34196 9180 34202
rect 9128 34138 9180 34144
rect 9220 33992 9272 33998
rect 9220 33934 9272 33940
rect 9232 33454 9260 33934
rect 9508 33658 9536 36654
rect 9588 36576 9640 36582
rect 9588 36518 9640 36524
rect 9600 34066 9628 36518
rect 9680 36100 9732 36106
rect 9680 36042 9732 36048
rect 9588 34060 9640 34066
rect 9588 34002 9640 34008
rect 9496 33652 9548 33658
rect 9496 33594 9548 33600
rect 9508 33538 9536 33594
rect 9416 33510 9536 33538
rect 9220 33448 9272 33454
rect 9220 33390 9272 33396
rect 9036 33380 9088 33386
rect 9036 33322 9088 33328
rect 9232 32978 9260 33390
rect 9312 33108 9364 33114
rect 9312 33050 9364 33056
rect 9324 32978 9352 33050
rect 9220 32972 9272 32978
rect 9220 32914 9272 32920
rect 9312 32972 9364 32978
rect 9312 32914 9364 32920
rect 9128 32360 9180 32366
rect 9128 32302 9180 32308
rect 9036 31816 9088 31822
rect 9036 31758 9088 31764
rect 9048 29850 9076 31758
rect 9140 30326 9168 32302
rect 9232 31890 9260 32914
rect 9416 32366 9444 33510
rect 9496 33380 9548 33386
rect 9496 33322 9548 33328
rect 9508 33114 9536 33322
rect 9496 33108 9548 33114
rect 9496 33050 9548 33056
rect 9496 32768 9548 32774
rect 9496 32710 9548 32716
rect 9588 32768 9640 32774
rect 9588 32710 9640 32716
rect 9508 32570 9536 32710
rect 9600 32570 9628 32710
rect 9496 32564 9548 32570
rect 9496 32506 9548 32512
rect 9588 32564 9640 32570
rect 9588 32506 9640 32512
rect 9404 32360 9456 32366
rect 9600 32348 9628 32506
rect 9404 32302 9456 32308
rect 9508 32320 9628 32348
rect 9220 31884 9272 31890
rect 9220 31826 9272 31832
rect 9508 31822 9536 32320
rect 9588 32224 9640 32230
rect 9588 32166 9640 32172
rect 9496 31816 9548 31822
rect 9496 31758 9548 31764
rect 9128 30320 9180 30326
rect 9128 30262 9180 30268
rect 9496 30252 9548 30258
rect 9496 30194 9548 30200
rect 9036 29844 9088 29850
rect 9036 29786 9088 29792
rect 9404 29640 9456 29646
rect 9404 29582 9456 29588
rect 9220 29232 9272 29238
rect 9220 29174 9272 29180
rect 9232 28694 9260 29174
rect 9220 28688 9272 28694
rect 9220 28630 9272 28636
rect 8944 28552 8996 28558
rect 8944 28494 8996 28500
rect 7840 28212 7892 28218
rect 7840 28154 7892 28160
rect 8576 28212 8628 28218
rect 8576 28154 8628 28160
rect 7852 28098 7880 28154
rect 7852 28070 8064 28098
rect 7840 28008 7892 28014
rect 7840 27950 7892 27956
rect 7656 27668 7708 27674
rect 7656 27610 7708 27616
rect 7668 26586 7696 27610
rect 7852 27402 7880 27950
rect 8036 27538 8064 28070
rect 8588 27606 8616 28154
rect 8576 27600 8628 27606
rect 8576 27542 8628 27548
rect 8024 27532 8076 27538
rect 8024 27474 8076 27480
rect 7840 27396 7892 27402
rect 7840 27338 7892 27344
rect 7748 26920 7800 26926
rect 7852 26908 7880 27338
rect 8588 27334 8616 27542
rect 8576 27328 8628 27334
rect 8576 27270 8628 27276
rect 7950 27228 8258 27237
rect 7950 27226 7956 27228
rect 8012 27226 8036 27228
rect 8092 27226 8116 27228
rect 8172 27226 8196 27228
rect 8252 27226 8258 27228
rect 8012 27174 8014 27226
rect 8194 27174 8196 27226
rect 7950 27172 7956 27174
rect 8012 27172 8036 27174
rect 8092 27172 8116 27174
rect 8172 27172 8196 27174
rect 8252 27172 8258 27174
rect 7950 27163 8258 27172
rect 7800 26880 7880 26908
rect 8300 26920 8352 26926
rect 7748 26862 7800 26868
rect 8300 26862 8352 26868
rect 7656 26580 7708 26586
rect 7656 26522 7708 26528
rect 7564 25832 7616 25838
rect 7564 25774 7616 25780
rect 7668 25362 7696 26522
rect 7840 26444 7892 26450
rect 7840 26386 7892 26392
rect 7852 25838 7880 26386
rect 7950 26140 8258 26149
rect 7950 26138 7956 26140
rect 8012 26138 8036 26140
rect 8092 26138 8116 26140
rect 8172 26138 8196 26140
rect 8252 26138 8258 26140
rect 8012 26086 8014 26138
rect 8194 26086 8196 26138
rect 7950 26084 7956 26086
rect 8012 26084 8036 26086
rect 8092 26084 8116 26086
rect 8172 26084 8196 26086
rect 8252 26084 8258 26086
rect 7950 26075 8258 26084
rect 8312 26042 8340 26862
rect 8588 26586 8616 27270
rect 8668 26988 8720 26994
rect 8668 26930 8720 26936
rect 8852 26988 8904 26994
rect 8852 26930 8904 26936
rect 8576 26580 8628 26586
rect 8576 26522 8628 26528
rect 8392 26376 8444 26382
rect 8392 26318 8444 26324
rect 8300 26036 8352 26042
rect 8300 25978 8352 25984
rect 7840 25832 7892 25838
rect 7840 25774 7892 25780
rect 8404 25430 8432 26318
rect 8576 26308 8628 26314
rect 8576 26250 8628 26256
rect 8392 25424 8444 25430
rect 8392 25366 8444 25372
rect 7656 25356 7708 25362
rect 7656 25298 7708 25304
rect 7472 24744 7524 24750
rect 7472 24686 7524 24692
rect 7380 24404 7432 24410
rect 7380 24346 7432 24352
rect 7484 24206 7512 24686
rect 7564 24404 7616 24410
rect 7564 24346 7616 24352
rect 7472 24200 7524 24206
rect 7472 24142 7524 24148
rect 7288 23724 7340 23730
rect 7288 23666 7340 23672
rect 7300 23186 7328 23666
rect 7288 23180 7340 23186
rect 7288 23122 7340 23128
rect 7300 22710 7328 23122
rect 7288 22704 7340 22710
rect 7288 22646 7340 22652
rect 7576 22094 7604 24346
rect 7668 24274 7696 25298
rect 7932 25152 7984 25158
rect 7852 25112 7932 25140
rect 7852 24750 7880 25112
rect 7932 25094 7984 25100
rect 7950 25052 8258 25061
rect 7950 25050 7956 25052
rect 8012 25050 8036 25052
rect 8092 25050 8116 25052
rect 8172 25050 8196 25052
rect 8252 25050 8258 25052
rect 8012 24998 8014 25050
rect 8194 24998 8196 25050
rect 7950 24996 7956 24998
rect 8012 24996 8036 24998
rect 8092 24996 8116 24998
rect 8172 24996 8196 24998
rect 8252 24996 8258 24998
rect 7950 24987 8258 24996
rect 8404 24954 8432 25366
rect 8392 24948 8444 24954
rect 8392 24890 8444 24896
rect 7840 24744 7892 24750
rect 7840 24686 7892 24692
rect 7656 24268 7708 24274
rect 7656 24210 7708 24216
rect 7950 23964 8258 23973
rect 7950 23962 7956 23964
rect 8012 23962 8036 23964
rect 8092 23962 8116 23964
rect 8172 23962 8196 23964
rect 8252 23962 8258 23964
rect 8012 23910 8014 23962
rect 8194 23910 8196 23962
rect 7950 23908 7956 23910
rect 8012 23908 8036 23910
rect 8092 23908 8116 23910
rect 8172 23908 8196 23910
rect 8252 23908 8258 23910
rect 7950 23899 8258 23908
rect 8300 23248 8352 23254
rect 8300 23190 8352 23196
rect 7950 22876 8258 22885
rect 7950 22874 7956 22876
rect 8012 22874 8036 22876
rect 8092 22874 8116 22876
rect 8172 22874 8196 22876
rect 8252 22874 8258 22876
rect 8012 22822 8014 22874
rect 8194 22822 8196 22874
rect 7950 22820 7956 22822
rect 8012 22820 8036 22822
rect 8092 22820 8116 22822
rect 8172 22820 8196 22822
rect 8252 22820 8258 22822
rect 7950 22811 8258 22820
rect 7748 22636 7800 22642
rect 7748 22578 7800 22584
rect 7576 22066 7696 22094
rect 7288 21888 7340 21894
rect 7288 21830 7340 21836
rect 7380 21888 7432 21894
rect 7380 21830 7432 21836
rect 7300 21146 7328 21830
rect 7392 21690 7420 21830
rect 7380 21684 7432 21690
rect 7380 21626 7432 21632
rect 7288 21140 7340 21146
rect 7288 21082 7340 21088
rect 7288 20800 7340 20806
rect 7288 20742 7340 20748
rect 7012 20460 7064 20466
rect 7012 20402 7064 20408
rect 7196 20460 7248 20466
rect 7196 20402 7248 20408
rect 7024 20262 7052 20402
rect 7012 20256 7064 20262
rect 7012 20198 7064 20204
rect 7104 20256 7156 20262
rect 7104 20198 7156 20204
rect 6920 19304 6972 19310
rect 6920 19246 6972 19252
rect 6920 18828 6972 18834
rect 6920 18770 6972 18776
rect 6828 18216 6880 18222
rect 6828 18158 6880 18164
rect 6932 17814 6960 18770
rect 6920 17808 6972 17814
rect 6920 17750 6972 17756
rect 6932 17202 6960 17750
rect 6920 17196 6972 17202
rect 6920 17138 6972 17144
rect 6932 16794 6960 17138
rect 6920 16788 6972 16794
rect 6920 16730 6972 16736
rect 6932 15434 6960 16730
rect 6920 15428 6972 15434
rect 6920 15370 6972 15376
rect 6828 15360 6880 15366
rect 6828 15302 6880 15308
rect 6840 13870 6868 15302
rect 6932 14414 6960 15370
rect 6920 14408 6972 14414
rect 6920 14350 6972 14356
rect 6920 14272 6972 14278
rect 6920 14214 6972 14220
rect 6828 13864 6880 13870
rect 6828 13806 6880 13812
rect 6840 13326 6868 13806
rect 6932 13802 6960 14214
rect 6920 13796 6972 13802
rect 6920 13738 6972 13744
rect 6828 13320 6880 13326
rect 6828 13262 6880 13268
rect 6736 12368 6788 12374
rect 6736 12310 6788 12316
rect 6840 8634 6868 13262
rect 6828 8628 6880 8634
rect 6828 8570 6880 8576
rect 7024 6730 7052 20198
rect 7116 20058 7144 20198
rect 7104 20052 7156 20058
rect 7104 19994 7156 20000
rect 7300 18086 7328 20742
rect 7380 19916 7432 19922
rect 7380 19858 7432 19864
rect 7288 18080 7340 18086
rect 7288 18022 7340 18028
rect 7288 15700 7340 15706
rect 7392 15688 7420 19858
rect 7668 19786 7696 22066
rect 7760 21690 7788 22578
rect 7840 21888 7892 21894
rect 7840 21830 7892 21836
rect 7748 21684 7800 21690
rect 7748 21626 7800 21632
rect 7748 20868 7800 20874
rect 7748 20810 7800 20816
rect 7656 19780 7708 19786
rect 7656 19722 7708 19728
rect 7472 19712 7524 19718
rect 7472 19654 7524 19660
rect 7340 15660 7420 15688
rect 7288 15642 7340 15648
rect 7392 15434 7420 15660
rect 7380 15428 7432 15434
rect 7380 15370 7432 15376
rect 7196 14408 7248 14414
rect 7196 14350 7248 14356
rect 7208 14074 7236 14350
rect 7196 14068 7248 14074
rect 7196 14010 7248 14016
rect 7104 13388 7156 13394
rect 7104 13330 7156 13336
rect 7116 9450 7144 13330
rect 7484 13138 7512 19654
rect 7656 18624 7708 18630
rect 7656 18566 7708 18572
rect 7668 17746 7696 18566
rect 7656 17740 7708 17746
rect 7656 17682 7708 17688
rect 7668 13394 7696 17682
rect 7760 16454 7788 20810
rect 7852 20330 7880 21830
rect 7950 21788 8258 21797
rect 7950 21786 7956 21788
rect 8012 21786 8036 21788
rect 8092 21786 8116 21788
rect 8172 21786 8196 21788
rect 8252 21786 8258 21788
rect 8012 21734 8014 21786
rect 8194 21734 8196 21786
rect 7950 21732 7956 21734
rect 8012 21732 8036 21734
rect 8092 21732 8116 21734
rect 8172 21732 8196 21734
rect 8252 21732 8258 21734
rect 7950 21723 8258 21732
rect 8116 21548 8168 21554
rect 8116 21490 8168 21496
rect 8128 21146 8156 21490
rect 8116 21140 8168 21146
rect 8116 21082 8168 21088
rect 8312 20806 8340 23190
rect 8392 22976 8444 22982
rect 8392 22918 8444 22924
rect 8404 22778 8432 22918
rect 8392 22772 8444 22778
rect 8392 22714 8444 22720
rect 8392 22092 8444 22098
rect 8392 22034 8444 22040
rect 8300 20800 8352 20806
rect 8300 20742 8352 20748
rect 7950 20700 8258 20709
rect 7950 20698 7956 20700
rect 8012 20698 8036 20700
rect 8092 20698 8116 20700
rect 8172 20698 8196 20700
rect 8252 20698 8258 20700
rect 8012 20646 8014 20698
rect 8194 20646 8196 20698
rect 7950 20644 7956 20646
rect 8012 20644 8036 20646
rect 8092 20644 8116 20646
rect 8172 20644 8196 20646
rect 8252 20644 8258 20646
rect 7950 20635 8258 20644
rect 8300 20392 8352 20398
rect 8300 20334 8352 20340
rect 7840 20324 7892 20330
rect 7840 20266 7892 20272
rect 7840 19712 7892 19718
rect 7840 19654 7892 19660
rect 7852 17338 7880 19654
rect 7950 19612 8258 19621
rect 7950 19610 7956 19612
rect 8012 19610 8036 19612
rect 8092 19610 8116 19612
rect 8172 19610 8196 19612
rect 8252 19610 8258 19612
rect 8012 19558 8014 19610
rect 8194 19558 8196 19610
rect 7950 19556 7956 19558
rect 8012 19556 8036 19558
rect 8092 19556 8116 19558
rect 8172 19556 8196 19558
rect 8252 19556 8258 19558
rect 7950 19547 8258 19556
rect 8312 18970 8340 20334
rect 8404 20058 8432 22034
rect 8484 21412 8536 21418
rect 8484 21354 8536 21360
rect 8392 20052 8444 20058
rect 8392 19994 8444 20000
rect 8496 19854 8524 21354
rect 8484 19848 8536 19854
rect 8484 19790 8536 19796
rect 8588 19496 8616 26250
rect 8680 26042 8708 26930
rect 8668 26036 8720 26042
rect 8668 25978 8720 25984
rect 8864 25770 8892 26930
rect 9036 26376 9088 26382
rect 9036 26318 9088 26324
rect 8852 25764 8904 25770
rect 8852 25706 8904 25712
rect 9048 24138 9076 26318
rect 9128 25152 9180 25158
rect 9128 25094 9180 25100
rect 9036 24132 9088 24138
rect 9036 24074 9088 24080
rect 9140 23866 9168 25094
rect 9416 23866 9444 29582
rect 9508 29322 9536 30194
rect 9600 30190 9628 32166
rect 9588 30184 9640 30190
rect 9588 30126 9640 30132
rect 9600 29714 9628 30126
rect 9588 29708 9640 29714
rect 9588 29650 9640 29656
rect 9508 29294 9628 29322
rect 9600 29238 9628 29294
rect 9588 29232 9640 29238
rect 9588 29174 9640 29180
rect 9496 28552 9548 28558
rect 9496 28494 9548 28500
rect 9128 23860 9180 23866
rect 9128 23802 9180 23808
rect 9404 23860 9456 23866
rect 9404 23802 9456 23808
rect 9036 23792 9088 23798
rect 9036 23734 9088 23740
rect 9048 23322 9076 23734
rect 9416 23322 9444 23802
rect 9036 23316 9088 23322
rect 9036 23258 9088 23264
rect 9404 23316 9456 23322
rect 9404 23258 9456 23264
rect 9312 23248 9364 23254
rect 9312 23190 9364 23196
rect 9128 23180 9180 23186
rect 9128 23122 9180 23128
rect 8668 23112 8720 23118
rect 8668 23054 8720 23060
rect 8680 22574 8708 23054
rect 9140 22710 9168 23122
rect 9128 22704 9180 22710
rect 9128 22646 9180 22652
rect 8668 22568 8720 22574
rect 8668 22510 8720 22516
rect 8496 19468 8616 19496
rect 8300 18964 8352 18970
rect 8300 18906 8352 18912
rect 7932 18828 7984 18834
rect 7932 18770 7984 18776
rect 7944 18630 7972 18770
rect 7932 18624 7984 18630
rect 7932 18566 7984 18572
rect 7950 18524 8258 18533
rect 7950 18522 7956 18524
rect 8012 18522 8036 18524
rect 8092 18522 8116 18524
rect 8172 18522 8196 18524
rect 8252 18522 8258 18524
rect 8012 18470 8014 18522
rect 8194 18470 8196 18522
rect 7950 18468 7956 18470
rect 8012 18468 8036 18470
rect 8092 18468 8116 18470
rect 8172 18468 8196 18470
rect 8252 18468 8258 18470
rect 7950 18459 8258 18468
rect 8300 18284 8352 18290
rect 8300 18226 8352 18232
rect 8312 17882 8340 18226
rect 8300 17876 8352 17882
rect 8300 17818 8352 17824
rect 8208 17672 8260 17678
rect 8392 17672 8444 17678
rect 8260 17620 8392 17626
rect 8208 17614 8444 17620
rect 8220 17598 8432 17614
rect 8300 17536 8352 17542
rect 8300 17478 8352 17484
rect 7950 17436 8258 17445
rect 7950 17434 7956 17436
rect 8012 17434 8036 17436
rect 8092 17434 8116 17436
rect 8172 17434 8196 17436
rect 8252 17434 8258 17436
rect 8012 17382 8014 17434
rect 8194 17382 8196 17434
rect 7950 17380 7956 17382
rect 8012 17380 8036 17382
rect 8092 17380 8116 17382
rect 8172 17380 8196 17382
rect 8252 17380 8258 17382
rect 7950 17371 8258 17380
rect 7840 17332 7892 17338
rect 7840 17274 7892 17280
rect 7840 16788 7892 16794
rect 7840 16730 7892 16736
rect 7748 16448 7800 16454
rect 7748 16390 7800 16396
rect 7852 16232 7880 16730
rect 7950 16348 8258 16357
rect 7950 16346 7956 16348
rect 8012 16346 8036 16348
rect 8092 16346 8116 16348
rect 8172 16346 8196 16348
rect 8252 16346 8258 16348
rect 8012 16294 8014 16346
rect 8194 16294 8196 16346
rect 7950 16292 7956 16294
rect 8012 16292 8036 16294
rect 8092 16292 8116 16294
rect 8172 16292 8196 16294
rect 8252 16292 8258 16294
rect 7950 16283 8258 16292
rect 7852 16204 7972 16232
rect 7840 16108 7892 16114
rect 7840 16050 7892 16056
rect 7852 13802 7880 16050
rect 7944 15638 7972 16204
rect 7932 15632 7984 15638
rect 7932 15574 7984 15580
rect 7950 15260 8258 15269
rect 7950 15258 7956 15260
rect 8012 15258 8036 15260
rect 8092 15258 8116 15260
rect 8172 15258 8196 15260
rect 8252 15258 8258 15260
rect 8012 15206 8014 15258
rect 8194 15206 8196 15258
rect 7950 15204 7956 15206
rect 8012 15204 8036 15206
rect 8092 15204 8116 15206
rect 8172 15204 8196 15206
rect 8252 15204 8258 15206
rect 7950 15195 8258 15204
rect 7950 14172 8258 14181
rect 7950 14170 7956 14172
rect 8012 14170 8036 14172
rect 8092 14170 8116 14172
rect 8172 14170 8196 14172
rect 8252 14170 8258 14172
rect 8012 14118 8014 14170
rect 8194 14118 8196 14170
rect 7950 14116 7956 14118
rect 8012 14116 8036 14118
rect 8092 14116 8116 14118
rect 8172 14116 8196 14118
rect 8252 14116 8258 14118
rect 7950 14107 8258 14116
rect 7840 13796 7892 13802
rect 7840 13738 7892 13744
rect 7656 13388 7708 13394
rect 7656 13330 7708 13336
rect 7484 13110 7696 13138
rect 7564 12912 7616 12918
rect 7564 12854 7616 12860
rect 7288 12844 7340 12850
rect 7288 12786 7340 12792
rect 7300 9450 7328 12786
rect 7104 9444 7156 9450
rect 7104 9386 7156 9392
rect 7288 9444 7340 9450
rect 7288 9386 7340 9392
rect 7576 8498 7604 12854
rect 7564 8492 7616 8498
rect 7564 8434 7616 8440
rect 7012 6724 7064 6730
rect 7012 6666 7064 6672
rect 7564 5568 7616 5574
rect 7564 5510 7616 5516
rect 6644 3732 6696 3738
rect 6644 3674 6696 3680
rect 6276 3528 6328 3534
rect 6276 3470 6328 3476
rect 5908 3188 5960 3194
rect 5908 3130 5960 3136
rect 5908 3052 5960 3058
rect 5908 2994 5960 3000
rect 5920 800 5948 2994
rect 6288 800 6316 3470
rect 7380 3392 7432 3398
rect 7380 3334 7432 3340
rect 7012 2848 7064 2854
rect 7012 2790 7064 2796
rect 6920 2508 6972 2514
rect 6920 2450 6972 2456
rect 6932 2310 6960 2450
rect 6644 2304 6696 2310
rect 6644 2246 6696 2252
rect 6920 2304 6972 2310
rect 6920 2246 6972 2252
rect 6656 800 6684 2246
rect 7024 800 7052 2790
rect 7392 800 7420 3334
rect 7576 3058 7604 5510
rect 7564 3052 7616 3058
rect 7564 2994 7616 3000
rect 7668 2310 7696 13110
rect 7950 13084 8258 13093
rect 7950 13082 7956 13084
rect 8012 13082 8036 13084
rect 8092 13082 8116 13084
rect 8172 13082 8196 13084
rect 8252 13082 8258 13084
rect 8012 13030 8014 13082
rect 8194 13030 8196 13082
rect 7950 13028 7956 13030
rect 8012 13028 8036 13030
rect 8092 13028 8116 13030
rect 8172 13028 8196 13030
rect 8252 13028 8258 13030
rect 7950 13019 8258 13028
rect 8312 12986 8340 17478
rect 8496 16046 8524 19468
rect 8680 18834 8708 22510
rect 9036 21888 9088 21894
rect 9036 21830 9088 21836
rect 8944 20800 8996 20806
rect 8944 20742 8996 20748
rect 8760 19236 8812 19242
rect 8760 19178 8812 19184
rect 8668 18828 8720 18834
rect 8668 18770 8720 18776
rect 8576 18760 8628 18766
rect 8576 18702 8628 18708
rect 8588 18222 8616 18702
rect 8576 18216 8628 18222
rect 8576 18158 8628 18164
rect 8772 17320 8800 19178
rect 8680 17292 8800 17320
rect 8484 16040 8536 16046
rect 8484 15982 8536 15988
rect 8576 14408 8628 14414
rect 8576 14350 8628 14356
rect 8484 14068 8536 14074
rect 8484 14010 8536 14016
rect 8496 13530 8524 14010
rect 8588 13870 8616 14350
rect 8576 13864 8628 13870
rect 8576 13806 8628 13812
rect 8484 13524 8536 13530
rect 8484 13466 8536 13472
rect 8496 13258 8524 13466
rect 8484 13252 8536 13258
rect 8484 13194 8536 13200
rect 8300 12980 8352 12986
rect 8300 12922 8352 12928
rect 8496 12918 8524 13194
rect 8576 13184 8628 13190
rect 8576 13126 8628 13132
rect 8484 12912 8536 12918
rect 8484 12854 8536 12860
rect 8588 12782 8616 13126
rect 8576 12776 8628 12782
rect 8576 12718 8628 12724
rect 8680 12434 8708 17292
rect 8760 17196 8812 17202
rect 8760 17138 8812 17144
rect 8772 15910 8800 17138
rect 8852 16584 8904 16590
rect 8852 16526 8904 16532
rect 8864 15910 8892 16526
rect 8760 15904 8812 15910
rect 8760 15846 8812 15852
rect 8852 15904 8904 15910
rect 8852 15846 8904 15852
rect 8864 14822 8892 15846
rect 8852 14816 8904 14822
rect 8852 14758 8904 14764
rect 8864 14482 8892 14758
rect 8852 14476 8904 14482
rect 8852 14418 8904 14424
rect 8852 12776 8904 12782
rect 8852 12718 8904 12724
rect 8588 12406 8708 12434
rect 7950 11996 8258 12005
rect 7950 11994 7956 11996
rect 8012 11994 8036 11996
rect 8092 11994 8116 11996
rect 8172 11994 8196 11996
rect 8252 11994 8258 11996
rect 8012 11942 8014 11994
rect 8194 11942 8196 11994
rect 7950 11940 7956 11942
rect 8012 11940 8036 11942
rect 8092 11940 8116 11942
rect 8172 11940 8196 11942
rect 8252 11940 8258 11942
rect 7950 11931 8258 11940
rect 7950 10908 8258 10917
rect 7950 10906 7956 10908
rect 8012 10906 8036 10908
rect 8092 10906 8116 10908
rect 8172 10906 8196 10908
rect 8252 10906 8258 10908
rect 8012 10854 8014 10906
rect 8194 10854 8196 10906
rect 7950 10852 7956 10854
rect 8012 10852 8036 10854
rect 8092 10852 8116 10854
rect 8172 10852 8196 10854
rect 8252 10852 8258 10854
rect 7950 10843 8258 10852
rect 7950 9820 8258 9829
rect 7950 9818 7956 9820
rect 8012 9818 8036 9820
rect 8092 9818 8116 9820
rect 8172 9818 8196 9820
rect 8252 9818 8258 9820
rect 8012 9766 8014 9818
rect 8194 9766 8196 9818
rect 7950 9764 7956 9766
rect 8012 9764 8036 9766
rect 8092 9764 8116 9766
rect 8172 9764 8196 9766
rect 8252 9764 8258 9766
rect 7950 9755 8258 9764
rect 7950 8732 8258 8741
rect 7950 8730 7956 8732
rect 8012 8730 8036 8732
rect 8092 8730 8116 8732
rect 8172 8730 8196 8732
rect 8252 8730 8258 8732
rect 8012 8678 8014 8730
rect 8194 8678 8196 8730
rect 7950 8676 7956 8678
rect 8012 8676 8036 8678
rect 8092 8676 8116 8678
rect 8172 8676 8196 8678
rect 8252 8676 8258 8678
rect 7950 8667 8258 8676
rect 7950 7644 8258 7653
rect 7950 7642 7956 7644
rect 8012 7642 8036 7644
rect 8092 7642 8116 7644
rect 8172 7642 8196 7644
rect 8252 7642 8258 7644
rect 8012 7590 8014 7642
rect 8194 7590 8196 7642
rect 7950 7588 7956 7590
rect 8012 7588 8036 7590
rect 8092 7588 8116 7590
rect 8172 7588 8196 7590
rect 8252 7588 8258 7590
rect 7950 7579 8258 7588
rect 8588 6914 8616 12406
rect 8864 12170 8892 12718
rect 8852 12164 8904 12170
rect 8852 12106 8904 12112
rect 8588 6886 8892 6914
rect 7950 6556 8258 6565
rect 7950 6554 7956 6556
rect 8012 6554 8036 6556
rect 8092 6554 8116 6556
rect 8172 6554 8196 6556
rect 8252 6554 8258 6556
rect 8012 6502 8014 6554
rect 8194 6502 8196 6554
rect 7950 6500 7956 6502
rect 8012 6500 8036 6502
rect 8092 6500 8116 6502
rect 8172 6500 8196 6502
rect 8252 6500 8258 6502
rect 7950 6491 8258 6500
rect 7838 5808 7894 5817
rect 7838 5743 7894 5752
rect 7746 5672 7802 5681
rect 7746 5607 7802 5616
rect 7760 3738 7788 5607
rect 7852 4010 7880 5743
rect 7950 5468 8258 5477
rect 7950 5466 7956 5468
rect 8012 5466 8036 5468
rect 8092 5466 8116 5468
rect 8172 5466 8196 5468
rect 8252 5466 8258 5468
rect 8012 5414 8014 5466
rect 8194 5414 8196 5466
rect 7950 5412 7956 5414
rect 8012 5412 8036 5414
rect 8092 5412 8116 5414
rect 8172 5412 8196 5414
rect 8252 5412 8258 5414
rect 7950 5403 8258 5412
rect 7950 4380 8258 4389
rect 7950 4378 7956 4380
rect 8012 4378 8036 4380
rect 8092 4378 8116 4380
rect 8172 4378 8196 4380
rect 8252 4378 8258 4380
rect 8012 4326 8014 4378
rect 8194 4326 8196 4378
rect 7950 4324 7956 4326
rect 8012 4324 8036 4326
rect 8092 4324 8116 4326
rect 8172 4324 8196 4326
rect 8252 4324 8258 4326
rect 7950 4315 8258 4324
rect 8392 4276 8444 4282
rect 8392 4218 8444 4224
rect 7840 4004 7892 4010
rect 7840 3946 7892 3952
rect 8404 3738 8432 4218
rect 8760 3936 8812 3942
rect 8760 3878 8812 3884
rect 7748 3732 7800 3738
rect 7748 3674 7800 3680
rect 8392 3732 8444 3738
rect 8392 3674 8444 3680
rect 7840 3528 7892 3534
rect 7840 3470 7892 3476
rect 7852 2854 7880 3470
rect 7950 3292 8258 3301
rect 7950 3290 7956 3292
rect 8012 3290 8036 3292
rect 8092 3290 8116 3292
rect 8172 3290 8196 3292
rect 8252 3290 8258 3292
rect 8012 3238 8014 3290
rect 8194 3238 8196 3290
rect 7950 3236 7956 3238
rect 8012 3236 8036 3238
rect 8092 3236 8116 3238
rect 8172 3236 8196 3238
rect 8252 3236 8258 3238
rect 7950 3227 8258 3236
rect 8484 2984 8536 2990
rect 8484 2926 8536 2932
rect 7840 2848 7892 2854
rect 7840 2790 7892 2796
rect 7748 2372 7800 2378
rect 7748 2314 7800 2320
rect 7656 2304 7708 2310
rect 7656 2246 7708 2252
rect 7760 800 7788 2314
rect 1122 0 1178 800
rect 1490 0 1546 800
rect 1858 0 1914 800
rect 2226 0 2282 800
rect 2594 0 2650 800
rect 2962 0 3018 800
rect 3330 0 3386 800
rect 3698 0 3754 800
rect 4066 0 4122 800
rect 4434 0 4490 800
rect 4802 0 4858 800
rect 5170 0 5226 800
rect 5538 0 5594 800
rect 5906 0 5962 800
rect 6274 0 6330 800
rect 6642 0 6698 800
rect 7010 0 7066 800
rect 7378 0 7434 800
rect 7746 0 7802 800
rect 7852 762 7880 2790
rect 8300 2440 8352 2446
rect 8300 2382 8352 2388
rect 7950 2204 8258 2213
rect 7950 2202 7956 2204
rect 8012 2202 8036 2204
rect 8092 2202 8116 2204
rect 8172 2202 8196 2204
rect 8252 2202 8258 2204
rect 8012 2150 8014 2202
rect 8194 2150 8196 2202
rect 7950 2148 7956 2150
rect 8012 2148 8036 2150
rect 8092 2148 8116 2150
rect 8172 2148 8196 2150
rect 8252 2148 8258 2150
rect 7950 2139 8258 2148
rect 8312 2038 8340 2382
rect 8496 2310 8524 2926
rect 8772 2904 8800 3878
rect 8864 3058 8892 6886
rect 8956 4214 8984 20742
rect 9048 14482 9076 21830
rect 9128 21344 9180 21350
rect 9128 21286 9180 21292
rect 9140 20058 9168 21286
rect 9128 20052 9180 20058
rect 9128 19994 9180 20000
rect 9220 18624 9272 18630
rect 9220 18566 9272 18572
rect 9128 17536 9180 17542
rect 9128 17478 9180 17484
rect 9140 16998 9168 17478
rect 9128 16992 9180 16998
rect 9128 16934 9180 16940
rect 9128 16448 9180 16454
rect 9128 16390 9180 16396
rect 9140 16250 9168 16390
rect 9128 16244 9180 16250
rect 9128 16186 9180 16192
rect 9232 16182 9260 18566
rect 9324 17678 9352 23190
rect 9404 21684 9456 21690
rect 9404 21626 9456 21632
rect 9416 19514 9444 21626
rect 9404 19508 9456 19514
rect 9404 19450 9456 19456
rect 9312 17672 9364 17678
rect 9312 17614 9364 17620
rect 9220 16176 9272 16182
rect 9220 16118 9272 16124
rect 9404 16108 9456 16114
rect 9404 16050 9456 16056
rect 9312 16040 9364 16046
rect 9312 15982 9364 15988
rect 9324 15706 9352 15982
rect 9312 15700 9364 15706
rect 9312 15642 9364 15648
rect 9036 14476 9088 14482
rect 9036 14418 9088 14424
rect 9036 14272 9088 14278
rect 9036 14214 9088 14220
rect 9048 13258 9076 14214
rect 9036 13252 9088 13258
rect 9036 13194 9088 13200
rect 8944 4208 8996 4214
rect 8944 4150 8996 4156
rect 8852 3052 8904 3058
rect 8852 2994 8904 3000
rect 8772 2876 8892 2904
rect 8484 2304 8536 2310
rect 8484 2246 8536 2252
rect 8300 2032 8352 2038
rect 8300 1974 8352 1980
rect 8036 870 8156 898
rect 8036 762 8064 870
rect 8128 800 8156 870
rect 8496 800 8524 2246
rect 8864 800 8892 2876
rect 9048 2106 9076 13194
rect 9416 10062 9444 16050
rect 9404 10056 9456 10062
rect 9404 9998 9456 10004
rect 9220 4140 9272 4146
rect 9220 4082 9272 4088
rect 9036 2100 9088 2106
rect 9036 2042 9088 2048
rect 9232 800 9260 4082
rect 9508 2582 9536 28494
rect 9692 26382 9720 36042
rect 9864 34944 9916 34950
rect 9864 34886 9916 34892
rect 9772 34672 9824 34678
rect 9772 34614 9824 34620
rect 9784 33522 9812 34614
rect 9772 33516 9824 33522
rect 9772 33458 9824 33464
rect 9772 32836 9824 32842
rect 9772 32778 9824 32784
rect 9784 28762 9812 32778
rect 9876 31482 9904 34886
rect 9968 33658 9996 37198
rect 10152 36938 10180 38218
rect 10060 36910 10180 36938
rect 10060 34542 10088 36910
rect 10140 36780 10192 36786
rect 10140 36722 10192 36728
rect 10048 34536 10100 34542
rect 10048 34478 10100 34484
rect 9956 33652 10008 33658
rect 9956 33594 10008 33600
rect 9956 33516 10008 33522
rect 9956 33458 10008 33464
rect 9968 31686 9996 33458
rect 10152 33114 10180 36722
rect 10244 36174 10272 39782
rect 10508 39364 10560 39370
rect 10508 39306 10560 39312
rect 10520 39030 10548 39306
rect 10324 39024 10376 39030
rect 10324 38966 10376 38972
rect 10508 39024 10560 39030
rect 10508 38966 10560 38972
rect 10232 36168 10284 36174
rect 10232 36110 10284 36116
rect 10232 35624 10284 35630
rect 10232 35566 10284 35572
rect 10244 35494 10272 35566
rect 10232 35488 10284 35494
rect 10232 35430 10284 35436
rect 10140 33108 10192 33114
rect 10140 33050 10192 33056
rect 10244 31793 10272 35430
rect 10336 35290 10364 38966
rect 10416 38888 10468 38894
rect 10416 38830 10468 38836
rect 10428 37942 10456 38830
rect 10416 37936 10468 37942
rect 10416 37878 10468 37884
rect 10508 37868 10560 37874
rect 10508 37810 10560 37816
rect 10416 37800 10468 37806
rect 10416 37742 10468 37748
rect 10428 37466 10456 37742
rect 10416 37460 10468 37466
rect 10416 37402 10468 37408
rect 10324 35284 10376 35290
rect 10324 35226 10376 35232
rect 10428 35170 10456 37402
rect 10520 36922 10548 37810
rect 10508 36916 10560 36922
rect 10508 36858 10560 36864
rect 10508 36236 10560 36242
rect 10508 36178 10560 36184
rect 10336 35142 10456 35170
rect 10230 31784 10286 31793
rect 10230 31719 10286 31728
rect 9956 31680 10008 31686
rect 9956 31622 10008 31628
rect 9864 31476 9916 31482
rect 9864 31418 9916 31424
rect 10232 31476 10284 31482
rect 10232 31418 10284 31424
rect 9862 31376 9918 31385
rect 9862 31311 9918 31320
rect 10048 31340 10100 31346
rect 9876 31278 9904 31311
rect 10048 31282 10100 31288
rect 9864 31272 9916 31278
rect 9864 31214 9916 31220
rect 10060 31142 10088 31282
rect 10048 31136 10100 31142
rect 10048 31078 10100 31084
rect 10060 29238 10088 31078
rect 10244 30326 10272 31418
rect 10232 30320 10284 30326
rect 10232 30262 10284 30268
rect 10140 29504 10192 29510
rect 10140 29446 10192 29452
rect 10048 29232 10100 29238
rect 10048 29174 10100 29180
rect 9956 29096 10008 29102
rect 9956 29038 10008 29044
rect 10048 29096 10100 29102
rect 10048 29038 10100 29044
rect 9864 28960 9916 28966
rect 9864 28902 9916 28908
rect 9772 28756 9824 28762
rect 9772 28698 9824 28704
rect 9876 28218 9904 28902
rect 9968 28626 9996 29038
rect 9956 28620 10008 28626
rect 9956 28562 10008 28568
rect 9864 28212 9916 28218
rect 9864 28154 9916 28160
rect 10060 28014 10088 29038
rect 10048 28008 10100 28014
rect 10048 27950 10100 27956
rect 10048 27600 10100 27606
rect 10048 27542 10100 27548
rect 9680 26376 9732 26382
rect 9680 26318 9732 26324
rect 10060 26314 10088 27542
rect 10048 26308 10100 26314
rect 10048 26250 10100 26256
rect 10152 26194 10180 29446
rect 9968 26166 10180 26194
rect 9588 24812 9640 24818
rect 9588 24754 9640 24760
rect 9600 24138 9628 24754
rect 9772 24676 9824 24682
rect 9772 24618 9824 24624
rect 9588 24132 9640 24138
rect 9588 24074 9640 24080
rect 9600 23526 9628 24074
rect 9784 23662 9812 24618
rect 9864 24064 9916 24070
rect 9864 24006 9916 24012
rect 9772 23656 9824 23662
rect 9772 23598 9824 23604
rect 9876 23594 9904 24006
rect 9864 23588 9916 23594
rect 9864 23530 9916 23536
rect 9588 23520 9640 23526
rect 9588 23462 9640 23468
rect 9600 23186 9628 23462
rect 9588 23180 9640 23186
rect 9588 23122 9640 23128
rect 9772 23180 9824 23186
rect 9772 23122 9824 23128
rect 9588 22976 9640 22982
rect 9588 22918 9640 22924
rect 9600 22030 9628 22918
rect 9784 22094 9812 23122
rect 9876 22710 9904 23530
rect 9864 22704 9916 22710
rect 9864 22646 9916 22652
rect 9784 22066 9904 22094
rect 9588 22024 9640 22030
rect 9588 21966 9640 21972
rect 9876 20534 9904 22066
rect 9968 21622 9996 26166
rect 10244 26058 10272 30262
rect 10336 29510 10364 35142
rect 10520 35086 10548 36178
rect 10508 35080 10560 35086
rect 10508 35022 10560 35028
rect 10416 33448 10468 33454
rect 10416 33390 10468 33396
rect 10428 30122 10456 33390
rect 10612 32314 10640 43710
rect 10704 43314 10732 43726
rect 10784 43648 10836 43654
rect 10784 43590 10836 43596
rect 10796 43382 10824 43590
rect 10784 43376 10836 43382
rect 10784 43318 10836 43324
rect 10692 43308 10744 43314
rect 10692 43250 10744 43256
rect 10784 43240 10836 43246
rect 10784 43182 10836 43188
rect 10692 39500 10744 39506
rect 10692 39442 10744 39448
rect 10704 37942 10732 39442
rect 10692 37936 10744 37942
rect 10692 37878 10744 37884
rect 10704 35494 10732 37878
rect 10796 37466 10824 43182
rect 10980 42634 11008 46990
rect 11072 44470 11100 53518
rect 11256 53038 11284 56200
rect 11624 53650 11652 56200
rect 11992 54126 12020 56200
rect 12072 54188 12124 54194
rect 12072 54130 12124 54136
rect 11888 54120 11940 54126
rect 11888 54062 11940 54068
rect 11980 54120 12032 54126
rect 11980 54062 12032 54068
rect 11900 53972 11928 54062
rect 11900 53944 12020 53972
rect 11612 53644 11664 53650
rect 11612 53586 11664 53592
rect 11888 53576 11940 53582
rect 11888 53518 11940 53524
rect 11244 53032 11296 53038
rect 11244 52974 11296 52980
rect 11796 52488 11848 52494
rect 11796 52430 11848 52436
rect 11612 52012 11664 52018
rect 11612 51954 11664 51960
rect 11624 47258 11652 51954
rect 11808 48890 11836 52430
rect 11900 52154 11928 53518
rect 11888 52148 11940 52154
rect 11888 52090 11940 52096
rect 11796 48884 11848 48890
rect 11796 48826 11848 48832
rect 11704 48748 11756 48754
rect 11704 48690 11756 48696
rect 11612 47252 11664 47258
rect 11612 47194 11664 47200
rect 11520 47048 11572 47054
rect 11520 46990 11572 46996
rect 11244 44804 11296 44810
rect 11244 44746 11296 44752
rect 11060 44464 11112 44470
rect 11060 44406 11112 44412
rect 11256 44198 11284 44746
rect 11336 44328 11388 44334
rect 11336 44270 11388 44276
rect 11244 44192 11296 44198
rect 11244 44134 11296 44140
rect 11060 43240 11112 43246
rect 11060 43182 11112 43188
rect 10968 42628 11020 42634
rect 10968 42570 11020 42576
rect 11072 42566 11100 43182
rect 11244 42696 11296 42702
rect 11244 42638 11296 42644
rect 11060 42560 11112 42566
rect 11060 42502 11112 42508
rect 10968 42356 11020 42362
rect 10968 42298 11020 42304
rect 10980 41206 11008 42298
rect 11152 42152 11204 42158
rect 11152 42094 11204 42100
rect 10968 41200 11020 41206
rect 10968 41142 11020 41148
rect 10876 41064 10928 41070
rect 10876 41006 10928 41012
rect 10888 38010 10916 41006
rect 11164 40934 11192 42094
rect 11256 41682 11284 42638
rect 11244 41676 11296 41682
rect 11244 41618 11296 41624
rect 11152 40928 11204 40934
rect 11152 40870 11204 40876
rect 11256 40594 11284 41618
rect 11348 41313 11376 44270
rect 11532 42362 11560 46990
rect 11716 44538 11744 48690
rect 11992 45558 12020 53944
rect 12084 52698 12112 54130
rect 12072 52692 12124 52698
rect 12072 52634 12124 52640
rect 12360 52494 12388 56200
rect 12728 53174 12756 56200
rect 12716 53168 12768 53174
rect 12716 53110 12768 53116
rect 12820 52986 12848 56222
rect 13004 56114 13032 56222
rect 13082 56200 13138 57000
rect 13450 56200 13506 57000
rect 13818 56200 13874 57000
rect 14186 56200 14242 57000
rect 14554 56200 14610 57000
rect 14922 56200 14978 57000
rect 15290 56200 15346 57000
rect 15658 56200 15714 57000
rect 16026 56200 16082 57000
rect 16394 56200 16450 57000
rect 16762 56200 16818 57000
rect 17130 56200 17186 57000
rect 17498 56200 17554 57000
rect 17866 56200 17922 57000
rect 18234 56200 18290 57000
rect 18602 56200 18658 57000
rect 18970 56200 19026 57000
rect 19338 56200 19394 57000
rect 19706 56200 19762 57000
rect 20074 56200 20130 57000
rect 20442 56200 20498 57000
rect 20810 56200 20866 57000
rect 21178 56200 21234 57000
rect 21546 56200 21602 57000
rect 21914 56200 21970 57000
rect 22282 56200 22338 57000
rect 22650 56200 22706 57000
rect 23018 56200 23074 57000
rect 23124 56222 23336 56250
rect 13096 56114 13124 56200
rect 13004 56086 13124 56114
rect 12950 53884 13258 53893
rect 12950 53882 12956 53884
rect 13012 53882 13036 53884
rect 13092 53882 13116 53884
rect 13172 53882 13196 53884
rect 13252 53882 13258 53884
rect 13012 53830 13014 53882
rect 13194 53830 13196 53882
rect 12950 53828 12956 53830
rect 13012 53828 13036 53830
rect 13092 53828 13116 53830
rect 13172 53828 13196 53830
rect 13252 53828 13258 53830
rect 12950 53819 13258 53828
rect 13464 53106 13492 56200
rect 13832 54330 13860 56200
rect 13820 54324 13872 54330
rect 13820 54266 13872 54272
rect 13832 53582 13860 54266
rect 14200 53582 14228 56200
rect 14568 54330 14596 56200
rect 14556 54324 14608 54330
rect 14556 54266 14608 54272
rect 14936 54262 14964 56200
rect 14924 54256 14976 54262
rect 14924 54198 14976 54204
rect 14936 53786 14964 54198
rect 15304 54194 15332 56200
rect 15292 54188 15344 54194
rect 15672 54176 15700 56200
rect 16040 54262 16068 56200
rect 16028 54256 16080 54262
rect 16028 54198 16080 54204
rect 15292 54130 15344 54136
rect 15580 54148 15700 54176
rect 15844 54188 15896 54194
rect 15108 53984 15160 53990
rect 15108 53926 15160 53932
rect 14924 53780 14976 53786
rect 14924 53722 14976 53728
rect 13820 53576 13872 53582
rect 13820 53518 13872 53524
rect 14188 53576 14240 53582
rect 14188 53518 14240 53524
rect 13636 53440 13688 53446
rect 13636 53382 13688 53388
rect 13452 53100 13504 53106
rect 13452 53042 13504 53048
rect 12728 52958 12848 52986
rect 12348 52488 12400 52494
rect 12348 52430 12400 52436
rect 12360 52154 12388 52430
rect 12728 52426 12756 52958
rect 12808 52896 12860 52902
rect 12808 52838 12860 52844
rect 12716 52420 12768 52426
rect 12716 52362 12768 52368
rect 12348 52148 12400 52154
rect 12348 52090 12400 52096
rect 11980 45552 12032 45558
rect 11980 45494 12032 45500
rect 12256 45484 12308 45490
rect 12256 45426 12308 45432
rect 12268 45286 12296 45426
rect 12256 45280 12308 45286
rect 12254 45248 12256 45257
rect 12716 45280 12768 45286
rect 12308 45248 12310 45257
rect 12716 45222 12768 45228
rect 12254 45183 12310 45192
rect 12348 44736 12400 44742
rect 12348 44678 12400 44684
rect 11704 44532 11756 44538
rect 11704 44474 11756 44480
rect 12360 44334 12388 44678
rect 12624 44396 12676 44402
rect 12624 44338 12676 44344
rect 12164 44328 12216 44334
rect 12164 44270 12216 44276
rect 12348 44328 12400 44334
rect 12348 44270 12400 44276
rect 11888 44192 11940 44198
rect 11888 44134 11940 44140
rect 11796 43784 11848 43790
rect 11796 43726 11848 43732
rect 11704 43716 11756 43722
rect 11704 43658 11756 43664
rect 11520 42356 11572 42362
rect 11520 42298 11572 42304
rect 11520 42084 11572 42090
rect 11520 42026 11572 42032
rect 11428 42016 11480 42022
rect 11428 41958 11480 41964
rect 11334 41304 11390 41313
rect 11334 41239 11390 41248
rect 11336 40996 11388 41002
rect 11336 40938 11388 40944
rect 11244 40588 11296 40594
rect 11244 40530 11296 40536
rect 11348 39846 11376 40938
rect 11336 39840 11388 39846
rect 11336 39782 11388 39788
rect 11244 39296 11296 39302
rect 11244 39238 11296 39244
rect 11060 38888 11112 38894
rect 11060 38830 11112 38836
rect 11072 38350 11100 38830
rect 11060 38344 11112 38350
rect 11060 38286 11112 38292
rect 11256 38282 11284 39238
rect 11336 38752 11388 38758
rect 11336 38694 11388 38700
rect 11348 38554 11376 38694
rect 11336 38548 11388 38554
rect 11336 38490 11388 38496
rect 11244 38276 11296 38282
rect 11244 38218 11296 38224
rect 10968 38208 11020 38214
rect 10968 38150 11020 38156
rect 10876 38004 10928 38010
rect 10876 37946 10928 37952
rect 10876 37732 10928 37738
rect 10876 37674 10928 37680
rect 10784 37460 10836 37466
rect 10784 37402 10836 37408
rect 10888 37330 10916 37674
rect 10980 37670 11008 38150
rect 10968 37664 11020 37670
rect 10968 37606 11020 37612
rect 10784 37324 10836 37330
rect 10784 37266 10836 37272
rect 10876 37324 10928 37330
rect 10876 37266 10928 37272
rect 10692 35488 10744 35494
rect 10692 35430 10744 35436
rect 10796 35222 10824 37266
rect 11244 37188 11296 37194
rect 11244 37130 11296 37136
rect 10876 37120 10928 37126
rect 10876 37062 10928 37068
rect 10888 36106 10916 37062
rect 10968 36780 11020 36786
rect 10968 36722 11020 36728
rect 10876 36100 10928 36106
rect 10876 36042 10928 36048
rect 10784 35216 10836 35222
rect 10784 35158 10836 35164
rect 10692 33584 10744 33590
rect 10692 33526 10744 33532
rect 10520 32286 10640 32314
rect 10520 31482 10548 32286
rect 10600 31748 10652 31754
rect 10600 31690 10652 31696
rect 10612 31482 10640 31690
rect 10508 31476 10560 31482
rect 10508 31418 10560 31424
rect 10600 31476 10652 31482
rect 10600 31418 10652 31424
rect 10612 31362 10640 31418
rect 10520 31334 10640 31362
rect 10416 30116 10468 30122
rect 10416 30058 10468 30064
rect 10324 29504 10376 29510
rect 10324 29446 10376 29452
rect 10324 29232 10376 29238
rect 10324 29174 10376 29180
rect 10336 27606 10364 29174
rect 10416 29028 10468 29034
rect 10416 28970 10468 28976
rect 10520 28994 10548 31334
rect 10600 31272 10652 31278
rect 10600 31214 10652 31220
rect 10612 30705 10640 31214
rect 10598 30696 10654 30705
rect 10704 30666 10732 33526
rect 10796 33454 10824 35158
rect 10980 34202 11008 36722
rect 11256 36650 11284 37130
rect 11244 36644 11296 36650
rect 11244 36586 11296 36592
rect 11152 36100 11204 36106
rect 11152 36042 11204 36048
rect 11164 35630 11192 36042
rect 11152 35624 11204 35630
rect 11152 35566 11204 35572
rect 11164 34746 11192 35566
rect 11244 35488 11296 35494
rect 11244 35430 11296 35436
rect 11152 34740 11204 34746
rect 11152 34682 11204 34688
rect 10968 34196 11020 34202
rect 10968 34138 11020 34144
rect 10784 33448 10836 33454
rect 10784 33390 10836 33396
rect 11164 33130 11192 34682
rect 10980 33102 11192 33130
rect 10784 32020 10836 32026
rect 10784 31962 10836 31968
rect 10796 30938 10824 31962
rect 10980 31822 11008 33102
rect 11256 32570 11284 35430
rect 11244 32564 11296 32570
rect 11244 32506 11296 32512
rect 11256 32026 11284 32506
rect 11244 32020 11296 32026
rect 11244 31962 11296 31968
rect 10968 31816 11020 31822
rect 10874 31784 10930 31793
rect 10968 31758 11020 31764
rect 10874 31719 10930 31728
rect 10888 31278 10916 31719
rect 10876 31272 10928 31278
rect 10876 31214 10928 31220
rect 10784 30932 10836 30938
rect 10784 30874 10836 30880
rect 10980 30802 11008 31758
rect 11256 31346 11284 31962
rect 11244 31340 11296 31346
rect 11244 31282 11296 31288
rect 10968 30796 11020 30802
rect 10968 30738 11020 30744
rect 10598 30631 10654 30640
rect 10692 30660 10744 30666
rect 10692 30602 10744 30608
rect 10704 29714 10732 30602
rect 11256 30258 11284 31282
rect 11244 30252 11296 30258
rect 11244 30194 11296 30200
rect 10968 30184 11020 30190
rect 10968 30126 11020 30132
rect 10692 29708 10744 29714
rect 10692 29650 10744 29656
rect 10876 29708 10928 29714
rect 10876 29650 10928 29656
rect 10888 29306 10916 29650
rect 10980 29646 11008 30126
rect 10968 29640 11020 29646
rect 10968 29582 11020 29588
rect 10968 29504 11020 29510
rect 10968 29446 11020 29452
rect 10876 29300 10928 29306
rect 10876 29242 10928 29248
rect 10324 27600 10376 27606
rect 10324 27542 10376 27548
rect 10324 26784 10376 26790
rect 10324 26726 10376 26732
rect 10152 26030 10272 26058
rect 10336 26042 10364 26726
rect 10324 26036 10376 26042
rect 10152 22094 10180 26030
rect 10324 25978 10376 25984
rect 10428 25974 10456 28970
rect 10520 28966 10824 28994
rect 10796 28694 10824 28966
rect 10980 28744 11008 29446
rect 10888 28716 11008 28744
rect 10784 28688 10836 28694
rect 10784 28630 10836 28636
rect 10600 28008 10652 28014
rect 10520 27968 10600 27996
rect 10520 26926 10548 27968
rect 10600 27950 10652 27956
rect 10692 27872 10744 27878
rect 10692 27814 10744 27820
rect 10600 27328 10652 27334
rect 10600 27270 10652 27276
rect 10508 26920 10560 26926
rect 10508 26862 10560 26868
rect 10520 26450 10548 26862
rect 10508 26444 10560 26450
rect 10508 26386 10560 26392
rect 10612 26382 10640 27270
rect 10600 26376 10652 26382
rect 10600 26318 10652 26324
rect 10416 25968 10468 25974
rect 10416 25910 10468 25916
rect 10704 24818 10732 27814
rect 10888 27130 10916 28716
rect 10968 28620 11020 28626
rect 10968 28562 11020 28568
rect 10980 28082 11008 28562
rect 10968 28076 11020 28082
rect 10968 28018 11020 28024
rect 10968 27668 11020 27674
rect 10968 27610 11020 27616
rect 10876 27124 10928 27130
rect 10876 27066 10928 27072
rect 10692 24812 10744 24818
rect 10692 24754 10744 24760
rect 10784 24812 10836 24818
rect 10784 24754 10836 24760
rect 10796 24410 10824 24754
rect 10980 24682 11008 27610
rect 10968 24676 11020 24682
rect 10968 24618 11020 24624
rect 10980 24410 11008 24618
rect 11348 24410 11376 38490
rect 11440 37330 11468 41958
rect 11532 41682 11560 42026
rect 11520 41676 11572 41682
rect 11520 41618 11572 41624
rect 11532 38418 11560 41618
rect 11520 38412 11572 38418
rect 11520 38354 11572 38360
rect 11520 37664 11572 37670
rect 11520 37606 11572 37612
rect 11428 37324 11480 37330
rect 11428 37266 11480 37272
rect 11532 35494 11560 37606
rect 11716 36904 11744 43658
rect 11808 42702 11836 43726
rect 11900 43178 11928 44134
rect 12176 43450 12204 44270
rect 12360 43722 12388 44270
rect 12348 43716 12400 43722
rect 12348 43658 12400 43664
rect 12164 43444 12216 43450
rect 12164 43386 12216 43392
rect 11888 43172 11940 43178
rect 11888 43114 11940 43120
rect 11796 42696 11848 42702
rect 11796 42638 11848 42644
rect 11900 41070 11928 43114
rect 12532 42764 12584 42770
rect 12532 42706 12584 42712
rect 12072 42560 12124 42566
rect 12072 42502 12124 42508
rect 12440 42560 12492 42566
rect 12440 42502 12492 42508
rect 11888 41064 11940 41070
rect 11888 41006 11940 41012
rect 11888 40928 11940 40934
rect 11888 40870 11940 40876
rect 11796 39840 11848 39846
rect 11796 39782 11848 39788
rect 11808 38894 11836 39782
rect 11900 39506 11928 40870
rect 11888 39500 11940 39506
rect 11888 39442 11940 39448
rect 11796 38888 11848 38894
rect 11796 38830 11848 38836
rect 11980 38888 12032 38894
rect 11980 38830 12032 38836
rect 11716 36876 11836 36904
rect 11612 36712 11664 36718
rect 11612 36654 11664 36660
rect 11520 35488 11572 35494
rect 11520 35430 11572 35436
rect 11520 33448 11572 33454
rect 11520 33390 11572 33396
rect 11532 31754 11560 33390
rect 11624 32978 11652 36654
rect 11704 35488 11756 35494
rect 11704 35430 11756 35436
rect 11716 35154 11744 35430
rect 11704 35148 11756 35154
rect 11704 35090 11756 35096
rect 11704 34400 11756 34406
rect 11704 34342 11756 34348
rect 11716 33590 11744 34342
rect 11704 33584 11756 33590
rect 11704 33526 11756 33532
rect 11612 32972 11664 32978
rect 11612 32914 11664 32920
rect 11624 31890 11652 32914
rect 11808 32366 11836 36876
rect 11888 36644 11940 36650
rect 11888 36586 11940 36592
rect 11900 35834 11928 36586
rect 11888 35828 11940 35834
rect 11888 35770 11940 35776
rect 11992 33658 12020 38830
rect 12084 38554 12112 42502
rect 12452 42362 12480 42502
rect 12440 42356 12492 42362
rect 12440 42298 12492 42304
rect 12348 42288 12400 42294
rect 12348 42230 12400 42236
rect 12256 41268 12308 41274
rect 12256 41210 12308 41216
rect 12164 40588 12216 40594
rect 12164 40530 12216 40536
rect 12176 40050 12204 40530
rect 12164 40044 12216 40050
rect 12164 39986 12216 39992
rect 12176 39506 12204 39986
rect 12164 39500 12216 39506
rect 12164 39442 12216 39448
rect 12268 39438 12296 41210
rect 12256 39432 12308 39438
rect 12256 39374 12308 39380
rect 12360 39098 12388 42230
rect 12544 41478 12572 42706
rect 12532 41472 12584 41478
rect 12532 41414 12584 41420
rect 12636 41274 12664 44338
rect 12728 42906 12756 45222
rect 12716 42900 12768 42906
rect 12716 42842 12768 42848
rect 12624 41268 12676 41274
rect 12624 41210 12676 41216
rect 12440 39976 12492 39982
rect 12440 39918 12492 39924
rect 12348 39092 12400 39098
rect 12348 39034 12400 39040
rect 12164 38956 12216 38962
rect 12452 38944 12480 39918
rect 12624 39296 12676 39302
rect 12624 39238 12676 39244
rect 12452 38916 12572 38944
rect 12164 38898 12216 38904
rect 12072 38548 12124 38554
rect 12072 38490 12124 38496
rect 12072 38276 12124 38282
rect 12072 38218 12124 38224
rect 12084 37346 12112 38218
rect 12176 38010 12204 38898
rect 12256 38888 12308 38894
rect 12256 38830 12308 38836
rect 12268 38758 12296 38830
rect 12440 38820 12492 38826
rect 12440 38762 12492 38768
rect 12256 38752 12308 38758
rect 12256 38694 12308 38700
rect 12348 38752 12400 38758
rect 12348 38694 12400 38700
rect 12256 38208 12308 38214
rect 12256 38150 12308 38156
rect 12164 38004 12216 38010
rect 12164 37946 12216 37952
rect 12084 37330 12204 37346
rect 12072 37324 12204 37330
rect 12124 37318 12204 37324
rect 12072 37266 12124 37272
rect 12070 37224 12126 37233
rect 12070 37159 12126 37168
rect 12084 36922 12112 37159
rect 12176 36922 12204 37318
rect 12072 36916 12124 36922
rect 12072 36858 12124 36864
rect 12164 36916 12216 36922
rect 12164 36858 12216 36864
rect 12164 35760 12216 35766
rect 12164 35702 12216 35708
rect 12176 35154 12204 35702
rect 12164 35148 12216 35154
rect 12164 35090 12216 35096
rect 12164 34944 12216 34950
rect 12164 34886 12216 34892
rect 12070 33688 12126 33697
rect 11980 33652 12032 33658
rect 12070 33623 12126 33632
rect 11980 33594 12032 33600
rect 11888 33516 11940 33522
rect 11888 33458 11940 33464
rect 11796 32360 11848 32366
rect 11796 32302 11848 32308
rect 11796 32224 11848 32230
rect 11796 32166 11848 32172
rect 11612 31884 11664 31890
rect 11612 31826 11664 31832
rect 11532 31726 11652 31754
rect 11520 27328 11572 27334
rect 11520 27270 11572 27276
rect 11532 27062 11560 27270
rect 11520 27056 11572 27062
rect 11520 26998 11572 27004
rect 11520 26784 11572 26790
rect 11520 26726 11572 26732
rect 11428 24812 11480 24818
rect 11428 24754 11480 24760
rect 10784 24404 10836 24410
rect 10784 24346 10836 24352
rect 10968 24404 11020 24410
rect 10968 24346 11020 24352
rect 11336 24404 11388 24410
rect 11336 24346 11388 24352
rect 10968 24268 11020 24274
rect 10968 24210 11020 24216
rect 10876 24200 10928 24206
rect 10876 24142 10928 24148
rect 10692 23520 10744 23526
rect 10692 23462 10744 23468
rect 10232 23180 10284 23186
rect 10232 23122 10284 23128
rect 10060 22066 10180 22094
rect 9956 21616 10008 21622
rect 9956 21558 10008 21564
rect 9968 20806 9996 21558
rect 9956 20800 10008 20806
rect 9956 20742 10008 20748
rect 9864 20528 9916 20534
rect 9916 20476 9996 20482
rect 9864 20470 9996 20476
rect 9876 20454 9996 20470
rect 9864 20392 9916 20398
rect 9864 20334 9916 20340
rect 9588 19712 9640 19718
rect 9588 19654 9640 19660
rect 9600 17338 9628 19654
rect 9680 19372 9732 19378
rect 9680 19314 9732 19320
rect 9588 17332 9640 17338
rect 9588 17274 9640 17280
rect 9588 16652 9640 16658
rect 9588 16594 9640 16600
rect 9600 14618 9628 16594
rect 9692 15434 9720 19314
rect 9876 19174 9904 20334
rect 9968 20058 9996 20454
rect 9956 20052 10008 20058
rect 9956 19994 10008 20000
rect 9968 19310 9996 19994
rect 9956 19304 10008 19310
rect 9956 19246 10008 19252
rect 9864 19168 9916 19174
rect 9864 19110 9916 19116
rect 9772 18896 9824 18902
rect 9772 18838 9824 18844
rect 9784 18698 9812 18838
rect 9772 18692 9824 18698
rect 9772 18634 9824 18640
rect 9784 18290 9812 18634
rect 9772 18284 9824 18290
rect 9772 18226 9824 18232
rect 9876 16726 9904 19110
rect 9968 18902 9996 19246
rect 9956 18896 10008 18902
rect 9956 18838 10008 18844
rect 9864 16720 9916 16726
rect 9864 16662 9916 16668
rect 9680 15428 9732 15434
rect 9680 15370 9732 15376
rect 9864 14952 9916 14958
rect 9864 14894 9916 14900
rect 9588 14612 9640 14618
rect 9588 14554 9640 14560
rect 9876 14482 9904 14894
rect 9864 14476 9916 14482
rect 9864 14418 9916 14424
rect 10060 13512 10088 22066
rect 10244 21570 10272 23122
rect 10508 22772 10560 22778
rect 10508 22714 10560 22720
rect 10520 21962 10548 22714
rect 10704 22710 10732 23462
rect 10692 22704 10744 22710
rect 10692 22646 10744 22652
rect 10888 22642 10916 24142
rect 10876 22636 10928 22642
rect 10876 22578 10928 22584
rect 10508 21956 10560 21962
rect 10508 21898 10560 21904
rect 10152 21542 10272 21570
rect 10152 20330 10180 21542
rect 10232 21480 10284 21486
rect 10232 21422 10284 21428
rect 10140 20324 10192 20330
rect 10140 20266 10192 20272
rect 10244 19122 10272 21422
rect 10324 21004 10376 21010
rect 10324 20946 10376 20952
rect 10784 21004 10836 21010
rect 10784 20946 10836 20952
rect 10336 20602 10364 20946
rect 10324 20596 10376 20602
rect 10324 20538 10376 20544
rect 10336 19310 10364 20538
rect 10692 20324 10744 20330
rect 10692 20266 10744 20272
rect 10416 20256 10468 20262
rect 10416 20198 10468 20204
rect 10428 19854 10456 20198
rect 10416 19848 10468 19854
rect 10416 19790 10468 19796
rect 10600 19712 10652 19718
rect 10520 19672 10600 19700
rect 10324 19304 10376 19310
rect 10324 19246 10376 19252
rect 10244 19094 10364 19122
rect 10140 18624 10192 18630
rect 10140 18566 10192 18572
rect 9968 13484 10088 13512
rect 9588 12912 9640 12918
rect 9588 12854 9640 12860
rect 9600 12434 9628 12854
rect 9600 12406 9720 12434
rect 9692 12170 9720 12406
rect 9680 12164 9732 12170
rect 9680 12106 9732 12112
rect 9968 6914 9996 13484
rect 10152 12434 10180 18566
rect 10060 12406 10180 12434
rect 10336 12434 10364 19094
rect 10520 16522 10548 19672
rect 10600 19654 10652 19660
rect 10704 18086 10732 20266
rect 10796 19786 10824 20946
rect 10980 20398 11008 24210
rect 11348 24138 11376 24346
rect 11336 24132 11388 24138
rect 11336 24074 11388 24080
rect 11348 23662 11376 24074
rect 11336 23656 11388 23662
rect 11336 23598 11388 23604
rect 11060 22976 11112 22982
rect 11060 22918 11112 22924
rect 11072 22778 11100 22918
rect 11060 22772 11112 22778
rect 11060 22714 11112 22720
rect 11244 22636 11296 22642
rect 11244 22578 11296 22584
rect 11256 22094 11284 22578
rect 11336 22094 11388 22098
rect 11256 22092 11388 22094
rect 11256 22066 11336 22092
rect 11336 22034 11388 22040
rect 11058 21720 11114 21729
rect 11058 21655 11060 21664
rect 11112 21655 11114 21664
rect 11060 21626 11112 21632
rect 11440 21418 11468 24754
rect 11532 22506 11560 26726
rect 11624 24177 11652 31726
rect 11704 25696 11756 25702
rect 11704 25638 11756 25644
rect 11610 24168 11666 24177
rect 11610 24103 11666 24112
rect 11612 24064 11664 24070
rect 11612 24006 11664 24012
rect 11520 22500 11572 22506
rect 11520 22442 11572 22448
rect 11520 21956 11572 21962
rect 11520 21898 11572 21904
rect 11532 21690 11560 21898
rect 11520 21684 11572 21690
rect 11520 21626 11572 21632
rect 11428 21412 11480 21418
rect 11428 21354 11480 21360
rect 10968 20392 11020 20398
rect 10968 20334 11020 20340
rect 10784 19780 10836 19786
rect 10784 19722 10836 19728
rect 11428 18964 11480 18970
rect 11428 18906 11480 18912
rect 11244 18420 11296 18426
rect 11244 18362 11296 18368
rect 11152 18216 11204 18222
rect 11152 18158 11204 18164
rect 10692 18080 10744 18086
rect 10692 18022 10744 18028
rect 10600 17604 10652 17610
rect 10600 17546 10652 17552
rect 10612 16590 10640 17546
rect 10704 17134 10732 18022
rect 11164 17610 11192 18158
rect 11152 17604 11204 17610
rect 11152 17546 11204 17552
rect 10692 17128 10744 17134
rect 10692 17070 10744 17076
rect 11060 17128 11112 17134
rect 11060 17070 11112 17076
rect 10784 16652 10836 16658
rect 10784 16594 10836 16600
rect 10600 16584 10652 16590
rect 10600 16526 10652 16532
rect 10508 16516 10560 16522
rect 10508 16458 10560 16464
rect 10508 15700 10560 15706
rect 10508 15642 10560 15648
rect 10520 14618 10548 15642
rect 10612 15570 10640 16526
rect 10600 15564 10652 15570
rect 10600 15506 10652 15512
rect 10612 14958 10640 15506
rect 10600 14952 10652 14958
rect 10600 14894 10652 14900
rect 10508 14612 10560 14618
rect 10508 14554 10560 14560
rect 10796 14074 10824 16594
rect 10876 16040 10928 16046
rect 10876 15982 10928 15988
rect 10888 15162 10916 15982
rect 11072 15706 11100 17070
rect 11256 16454 11284 18362
rect 11440 16946 11468 18906
rect 11532 17746 11560 21626
rect 11624 20874 11652 24006
rect 11716 21593 11744 25638
rect 11702 21584 11758 21593
rect 11702 21519 11758 21528
rect 11704 21072 11756 21078
rect 11702 21040 11704 21049
rect 11756 21040 11758 21049
rect 11702 20975 11758 20984
rect 11612 20868 11664 20874
rect 11612 20810 11664 20816
rect 11704 20392 11756 20398
rect 11704 20334 11756 20340
rect 11716 19854 11744 20334
rect 11704 19848 11756 19854
rect 11704 19790 11756 19796
rect 11612 19440 11664 19446
rect 11612 19382 11664 19388
rect 11520 17740 11572 17746
rect 11520 17682 11572 17688
rect 11440 16918 11560 16946
rect 11428 16788 11480 16794
rect 11428 16730 11480 16736
rect 11440 16522 11468 16730
rect 11428 16516 11480 16522
rect 11428 16458 11480 16464
rect 11244 16448 11296 16454
rect 11244 16390 11296 16396
rect 11060 15700 11112 15706
rect 11060 15642 11112 15648
rect 11256 15570 11284 16390
rect 11244 15564 11296 15570
rect 11244 15506 11296 15512
rect 11256 15434 11284 15506
rect 11244 15428 11296 15434
rect 11244 15370 11296 15376
rect 10876 15156 10928 15162
rect 10876 15098 10928 15104
rect 11256 15094 11284 15370
rect 11244 15088 11296 15094
rect 11244 15030 11296 15036
rect 11060 14884 11112 14890
rect 11060 14826 11112 14832
rect 10968 14476 11020 14482
rect 10968 14418 11020 14424
rect 10784 14068 10836 14074
rect 10784 14010 10836 14016
rect 10336 12406 10456 12434
rect 10060 11642 10088 12406
rect 10060 11614 10180 11642
rect 10152 6914 10180 11614
rect 9968 6886 10088 6914
rect 10152 6886 10364 6914
rect 10060 4282 10088 6886
rect 10336 4758 10364 6886
rect 10324 4752 10376 4758
rect 10324 4694 10376 4700
rect 10048 4276 10100 4282
rect 10048 4218 10100 4224
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 9956 3528 10008 3534
rect 9956 3470 10008 3476
rect 9600 2854 9628 3470
rect 9968 2854 9996 3470
rect 10428 3126 10456 12406
rect 10692 3528 10744 3534
rect 10692 3470 10744 3476
rect 10416 3120 10468 3126
rect 10416 3062 10468 3068
rect 10324 3052 10376 3058
rect 10324 2994 10376 3000
rect 9588 2848 9640 2854
rect 9588 2790 9640 2796
rect 9956 2848 10008 2854
rect 9956 2790 10008 2796
rect 9496 2576 9548 2582
rect 9496 2518 9548 2524
rect 9600 800 9628 2790
rect 9968 800 9996 2790
rect 10336 800 10364 2994
rect 10704 800 10732 3470
rect 10796 2650 10824 14010
rect 10980 14006 11008 14418
rect 10968 14000 11020 14006
rect 10968 13942 11020 13948
rect 10968 12640 11020 12646
rect 10968 12582 11020 12588
rect 10980 12374 11008 12582
rect 10968 12368 11020 12374
rect 10968 12310 11020 12316
rect 10876 5772 10928 5778
rect 10876 5714 10928 5720
rect 10888 2990 10916 5714
rect 10968 3936 11020 3942
rect 10968 3878 11020 3884
rect 10980 3058 11008 3878
rect 10968 3052 11020 3058
rect 10968 2994 11020 3000
rect 10876 2984 10928 2990
rect 10876 2926 10928 2932
rect 10784 2644 10836 2650
rect 10784 2586 10836 2592
rect 11072 2446 11100 14826
rect 11256 14346 11284 15030
rect 11336 14612 11388 14618
rect 11336 14554 11388 14560
rect 11244 14340 11296 14346
rect 11244 14282 11296 14288
rect 11256 14006 11284 14282
rect 11244 14000 11296 14006
rect 11244 13942 11296 13948
rect 11348 12782 11376 14554
rect 11336 12776 11388 12782
rect 11336 12718 11388 12724
rect 11532 12434 11560 16918
rect 11624 14618 11652 19382
rect 11808 18630 11836 32166
rect 11900 24818 11928 33458
rect 12084 33454 12112 33623
rect 12072 33448 12124 33454
rect 12072 33390 12124 33396
rect 12176 32978 12204 34886
rect 12268 33658 12296 38150
rect 12360 37670 12388 38694
rect 12348 37664 12400 37670
rect 12348 37606 12400 37612
rect 12452 36922 12480 38762
rect 12440 36916 12492 36922
rect 12440 36858 12492 36864
rect 12348 33856 12400 33862
rect 12348 33798 12400 33804
rect 12256 33652 12308 33658
rect 12256 33594 12308 33600
rect 12164 32972 12216 32978
rect 12164 32914 12216 32920
rect 12360 32026 12388 33798
rect 12544 33454 12572 38916
rect 12636 38214 12664 39238
rect 12728 38554 12756 42842
rect 12716 38548 12768 38554
rect 12716 38490 12768 38496
rect 12624 38208 12676 38214
rect 12624 38150 12676 38156
rect 12820 37890 12848 52838
rect 12950 52796 13258 52805
rect 12950 52794 12956 52796
rect 13012 52794 13036 52796
rect 13092 52794 13116 52796
rect 13172 52794 13196 52796
rect 13252 52794 13258 52796
rect 13012 52742 13014 52794
rect 13194 52742 13196 52794
rect 12950 52740 12956 52742
rect 13012 52740 13036 52742
rect 13092 52740 13116 52742
rect 13172 52740 13196 52742
rect 13252 52740 13258 52742
rect 12950 52731 13258 52740
rect 13464 52698 13492 53042
rect 13452 52692 13504 52698
rect 13452 52634 13504 52640
rect 13360 52624 13412 52630
rect 13360 52566 13412 52572
rect 12950 51708 13258 51717
rect 12950 51706 12956 51708
rect 13012 51706 13036 51708
rect 13092 51706 13116 51708
rect 13172 51706 13196 51708
rect 13252 51706 13258 51708
rect 13012 51654 13014 51706
rect 13194 51654 13196 51706
rect 12950 51652 12956 51654
rect 13012 51652 13036 51654
rect 13092 51652 13116 51654
rect 13172 51652 13196 51654
rect 13252 51652 13258 51654
rect 12950 51643 13258 51652
rect 12950 50620 13258 50629
rect 12950 50618 12956 50620
rect 13012 50618 13036 50620
rect 13092 50618 13116 50620
rect 13172 50618 13196 50620
rect 13252 50618 13258 50620
rect 13012 50566 13014 50618
rect 13194 50566 13196 50618
rect 12950 50564 12956 50566
rect 13012 50564 13036 50566
rect 13092 50564 13116 50566
rect 13172 50564 13196 50566
rect 13252 50564 13258 50566
rect 12950 50555 13258 50564
rect 12950 49532 13258 49541
rect 12950 49530 12956 49532
rect 13012 49530 13036 49532
rect 13092 49530 13116 49532
rect 13172 49530 13196 49532
rect 13252 49530 13258 49532
rect 13012 49478 13014 49530
rect 13194 49478 13196 49530
rect 12950 49476 12956 49478
rect 13012 49476 13036 49478
rect 13092 49476 13116 49478
rect 13172 49476 13196 49478
rect 13252 49476 13258 49478
rect 12950 49467 13258 49476
rect 12950 48444 13258 48453
rect 12950 48442 12956 48444
rect 13012 48442 13036 48444
rect 13092 48442 13116 48444
rect 13172 48442 13196 48444
rect 13252 48442 13258 48444
rect 13012 48390 13014 48442
rect 13194 48390 13196 48442
rect 12950 48388 12956 48390
rect 13012 48388 13036 48390
rect 13092 48388 13116 48390
rect 13172 48388 13196 48390
rect 13252 48388 13258 48390
rect 12950 48379 13258 48388
rect 12950 47356 13258 47365
rect 12950 47354 12956 47356
rect 13012 47354 13036 47356
rect 13092 47354 13116 47356
rect 13172 47354 13196 47356
rect 13252 47354 13258 47356
rect 13012 47302 13014 47354
rect 13194 47302 13196 47354
rect 12950 47300 12956 47302
rect 13012 47300 13036 47302
rect 13092 47300 13116 47302
rect 13172 47300 13196 47302
rect 13252 47300 13258 47302
rect 12950 47291 13258 47300
rect 12950 46268 13258 46277
rect 12950 46266 12956 46268
rect 13012 46266 13036 46268
rect 13092 46266 13116 46268
rect 13172 46266 13196 46268
rect 13252 46266 13258 46268
rect 13012 46214 13014 46266
rect 13194 46214 13196 46266
rect 12950 46212 12956 46214
rect 13012 46212 13036 46214
rect 13092 46212 13116 46214
rect 13172 46212 13196 46214
rect 13252 46212 13258 46214
rect 12950 46203 13258 46212
rect 12950 45180 13258 45189
rect 12950 45178 12956 45180
rect 13012 45178 13036 45180
rect 13092 45178 13116 45180
rect 13172 45178 13196 45180
rect 13252 45178 13258 45180
rect 13012 45126 13014 45178
rect 13194 45126 13196 45178
rect 12950 45124 12956 45126
rect 13012 45124 13036 45126
rect 13092 45124 13116 45126
rect 13172 45124 13196 45126
rect 13252 45124 13258 45126
rect 12950 45115 13258 45124
rect 12950 44092 13258 44101
rect 12950 44090 12956 44092
rect 13012 44090 13036 44092
rect 13092 44090 13116 44092
rect 13172 44090 13196 44092
rect 13252 44090 13258 44092
rect 13012 44038 13014 44090
rect 13194 44038 13196 44090
rect 12950 44036 12956 44038
rect 13012 44036 13036 44038
rect 13092 44036 13116 44038
rect 13172 44036 13196 44038
rect 13252 44036 13258 44038
rect 12950 44027 13258 44036
rect 12950 43004 13258 43013
rect 12950 43002 12956 43004
rect 13012 43002 13036 43004
rect 13092 43002 13116 43004
rect 13172 43002 13196 43004
rect 13252 43002 13258 43004
rect 13012 42950 13014 43002
rect 13194 42950 13196 43002
rect 12950 42948 12956 42950
rect 13012 42948 13036 42950
rect 13092 42948 13116 42950
rect 13172 42948 13196 42950
rect 13252 42948 13258 42950
rect 12950 42939 13258 42948
rect 12950 41916 13258 41925
rect 12950 41914 12956 41916
rect 13012 41914 13036 41916
rect 13092 41914 13116 41916
rect 13172 41914 13196 41916
rect 13252 41914 13258 41916
rect 13012 41862 13014 41914
rect 13194 41862 13196 41914
rect 12950 41860 12956 41862
rect 13012 41860 13036 41862
rect 13092 41860 13116 41862
rect 13172 41860 13196 41862
rect 13252 41860 13258 41862
rect 12950 41851 13258 41860
rect 13268 41608 13320 41614
rect 13268 41550 13320 41556
rect 13280 41478 13308 41550
rect 13268 41472 13320 41478
rect 13268 41414 13320 41420
rect 13280 41274 13308 41414
rect 13268 41268 13320 41274
rect 13268 41210 13320 41216
rect 12950 40828 13258 40837
rect 12950 40826 12956 40828
rect 13012 40826 13036 40828
rect 13092 40826 13116 40828
rect 13172 40826 13196 40828
rect 13252 40826 13258 40828
rect 13012 40774 13014 40826
rect 13194 40774 13196 40826
rect 12950 40772 12956 40774
rect 13012 40772 13036 40774
rect 13092 40772 13116 40774
rect 13172 40772 13196 40774
rect 13252 40772 13258 40774
rect 12950 40763 13258 40772
rect 13372 40526 13400 52566
rect 13452 52488 13504 52494
rect 13452 52430 13504 52436
rect 13464 40769 13492 52430
rect 13544 45416 13596 45422
rect 13544 45358 13596 45364
rect 13450 40760 13506 40769
rect 13450 40695 13506 40704
rect 13452 40588 13504 40594
rect 13452 40530 13504 40536
rect 13360 40520 13412 40526
rect 13360 40462 13412 40468
rect 13360 40384 13412 40390
rect 13360 40326 13412 40332
rect 12950 39740 13258 39749
rect 12950 39738 12956 39740
rect 13012 39738 13036 39740
rect 13092 39738 13116 39740
rect 13172 39738 13196 39740
rect 13252 39738 13258 39740
rect 13012 39686 13014 39738
rect 13194 39686 13196 39738
rect 12950 39684 12956 39686
rect 13012 39684 13036 39686
rect 13092 39684 13116 39686
rect 13172 39684 13196 39686
rect 13252 39684 13258 39686
rect 12950 39675 13258 39684
rect 12900 39092 12952 39098
rect 12900 39034 12952 39040
rect 12912 38758 12940 39034
rect 12900 38752 12952 38758
rect 12900 38694 12952 38700
rect 12950 38652 13258 38661
rect 12950 38650 12956 38652
rect 13012 38650 13036 38652
rect 13092 38650 13116 38652
rect 13172 38650 13196 38652
rect 13252 38650 13258 38652
rect 13012 38598 13014 38650
rect 13194 38598 13196 38650
rect 12950 38596 12956 38598
rect 13012 38596 13036 38598
rect 13092 38596 13116 38598
rect 13172 38596 13196 38598
rect 13252 38596 13258 38598
rect 12950 38587 13258 38596
rect 12992 38548 13044 38554
rect 12992 38490 13044 38496
rect 12900 38004 12952 38010
rect 12900 37946 12952 37952
rect 12728 37862 12848 37890
rect 12624 37460 12676 37466
rect 12624 37402 12676 37408
rect 12636 37330 12664 37402
rect 12624 37324 12676 37330
rect 12624 37266 12676 37272
rect 12728 36632 12756 37862
rect 12912 37754 12940 37946
rect 13004 37806 13032 38490
rect 13372 37806 13400 40326
rect 12820 37738 12940 37754
rect 12992 37800 13044 37806
rect 12992 37742 13044 37748
rect 13360 37800 13412 37806
rect 13360 37742 13412 37748
rect 12808 37732 12940 37738
rect 12860 37726 12940 37732
rect 12808 37674 12860 37680
rect 12820 37466 12848 37674
rect 12950 37564 13258 37573
rect 12950 37562 12956 37564
rect 13012 37562 13036 37564
rect 13092 37562 13116 37564
rect 13172 37562 13196 37564
rect 13252 37562 13258 37564
rect 13012 37510 13014 37562
rect 13194 37510 13196 37562
rect 12950 37508 12956 37510
rect 13012 37508 13036 37510
rect 13092 37508 13116 37510
rect 13172 37508 13196 37510
rect 13252 37508 13258 37510
rect 12950 37499 13258 37508
rect 12808 37460 12860 37466
rect 12808 37402 12860 37408
rect 12636 36604 12756 36632
rect 12532 33448 12584 33454
rect 12532 33390 12584 33396
rect 12532 32360 12584 32366
rect 12532 32302 12584 32308
rect 12348 32020 12400 32026
rect 12348 31962 12400 31968
rect 12256 31340 12308 31346
rect 12256 31282 12308 31288
rect 12268 30666 12296 31282
rect 12544 31142 12572 32302
rect 12532 31136 12584 31142
rect 12532 31078 12584 31084
rect 12256 30660 12308 30666
rect 12256 30602 12308 30608
rect 12636 29578 12664 36604
rect 12950 36476 13258 36485
rect 12950 36474 12956 36476
rect 13012 36474 13036 36476
rect 13092 36474 13116 36476
rect 13172 36474 13196 36476
rect 13252 36474 13258 36476
rect 13012 36422 13014 36474
rect 13194 36422 13196 36474
rect 12950 36420 12956 36422
rect 13012 36420 13036 36422
rect 13092 36420 13116 36422
rect 13172 36420 13196 36422
rect 13252 36420 13258 36422
rect 12950 36411 13258 36420
rect 13360 36032 13412 36038
rect 13360 35974 13412 35980
rect 12950 35388 13258 35397
rect 12950 35386 12956 35388
rect 13012 35386 13036 35388
rect 13092 35386 13116 35388
rect 13172 35386 13196 35388
rect 13252 35386 13258 35388
rect 13012 35334 13014 35386
rect 13194 35334 13196 35386
rect 12950 35332 12956 35334
rect 13012 35332 13036 35334
rect 13092 35332 13116 35334
rect 13172 35332 13196 35334
rect 13252 35332 13258 35334
rect 12950 35323 13258 35332
rect 12714 35184 12770 35193
rect 12714 35119 12770 35128
rect 12728 32910 12756 35119
rect 13176 35012 13228 35018
rect 13176 34954 13228 34960
rect 13188 34678 13216 34954
rect 13176 34672 13228 34678
rect 13176 34614 13228 34620
rect 12808 34536 12860 34542
rect 12808 34478 12860 34484
rect 12716 32904 12768 32910
rect 12716 32846 12768 32852
rect 12728 32570 12756 32846
rect 12716 32564 12768 32570
rect 12716 32506 12768 32512
rect 12728 32230 12756 32506
rect 12716 32224 12768 32230
rect 12716 32166 12768 32172
rect 12716 31748 12768 31754
rect 12716 31690 12768 31696
rect 12348 29572 12400 29578
rect 12348 29514 12400 29520
rect 12624 29572 12676 29578
rect 12624 29514 12676 29520
rect 12164 29504 12216 29510
rect 12164 29446 12216 29452
rect 12256 29504 12308 29510
rect 12360 29481 12388 29514
rect 12256 29446 12308 29452
rect 12346 29472 12402 29481
rect 12176 29306 12204 29446
rect 12164 29300 12216 29306
rect 12164 29242 12216 29248
rect 12164 28960 12216 28966
rect 12164 28902 12216 28908
rect 12072 28008 12124 28014
rect 12072 27950 12124 27956
rect 11980 27872 12032 27878
rect 11980 27814 12032 27820
rect 11992 27674 12020 27814
rect 11980 27668 12032 27674
rect 11980 27610 12032 27616
rect 11980 26920 12032 26926
rect 11980 26862 12032 26868
rect 11992 26586 12020 26862
rect 11980 26580 12032 26586
rect 11980 26522 12032 26528
rect 11992 25974 12020 26522
rect 11980 25968 12032 25974
rect 11980 25910 12032 25916
rect 12084 25106 12112 27950
rect 11992 25078 12112 25106
rect 11888 24812 11940 24818
rect 11888 24754 11940 24760
rect 11992 23798 12020 25078
rect 11980 23792 12032 23798
rect 11980 23734 12032 23740
rect 11888 22092 11940 22098
rect 11888 22034 11940 22040
rect 11900 19514 11928 22034
rect 11992 20534 12020 23734
rect 12072 23248 12124 23254
rect 12072 23190 12124 23196
rect 12084 20874 12112 23190
rect 12176 22234 12204 28902
rect 12268 22778 12296 29446
rect 12346 29407 12402 29416
rect 12636 28762 12664 29514
rect 12624 28756 12676 28762
rect 12360 28716 12624 28744
rect 12360 28014 12388 28716
rect 12624 28698 12676 28704
rect 12532 28484 12584 28490
rect 12532 28426 12584 28432
rect 12544 28218 12572 28426
rect 12532 28212 12584 28218
rect 12532 28154 12584 28160
rect 12348 28008 12400 28014
rect 12348 27950 12400 27956
rect 12440 28008 12492 28014
rect 12440 27950 12492 27956
rect 12452 27690 12480 27950
rect 12360 27674 12480 27690
rect 12348 27668 12480 27674
rect 12400 27662 12480 27668
rect 12348 27610 12400 27616
rect 12440 27328 12492 27334
rect 12440 27270 12492 27276
rect 12452 24410 12480 27270
rect 12544 27062 12572 28154
rect 12624 28076 12676 28082
rect 12624 28018 12676 28024
rect 12532 27056 12584 27062
rect 12532 26998 12584 27004
rect 12544 26926 12572 26998
rect 12532 26920 12584 26926
rect 12532 26862 12584 26868
rect 12636 26450 12664 28018
rect 12624 26444 12676 26450
rect 12624 26386 12676 26392
rect 12624 25832 12676 25838
rect 12624 25774 12676 25780
rect 12532 25152 12584 25158
rect 12532 25094 12584 25100
rect 12544 24954 12572 25094
rect 12532 24948 12584 24954
rect 12532 24890 12584 24896
rect 12636 24818 12664 25774
rect 12624 24812 12676 24818
rect 12624 24754 12676 24760
rect 12728 24562 12756 31690
rect 12820 30938 12848 34478
rect 12950 34300 13258 34309
rect 12950 34298 12956 34300
rect 13012 34298 13036 34300
rect 13092 34298 13116 34300
rect 13172 34298 13196 34300
rect 13252 34298 13258 34300
rect 13012 34246 13014 34298
rect 13194 34246 13196 34298
rect 12950 34244 12956 34246
rect 13012 34244 13036 34246
rect 13092 34244 13116 34246
rect 13172 34244 13196 34246
rect 13252 34244 13258 34246
rect 12950 34235 13258 34244
rect 13372 33998 13400 35974
rect 13464 35630 13492 40530
rect 13556 40338 13584 45358
rect 13648 44538 13676 53382
rect 14372 52896 14424 52902
rect 14372 52838 14424 52844
rect 14384 52601 14412 52838
rect 14370 52592 14426 52601
rect 14370 52527 14426 52536
rect 13820 47252 13872 47258
rect 13820 47194 13872 47200
rect 14832 47252 14884 47258
rect 14832 47194 14884 47200
rect 13832 46714 13860 47194
rect 14556 47116 14608 47122
rect 14556 47058 14608 47064
rect 13820 46708 13872 46714
rect 13820 46650 13872 46656
rect 13728 45484 13780 45490
rect 13728 45426 13780 45432
rect 13740 44742 13768 45426
rect 14280 44872 14332 44878
rect 14280 44814 14332 44820
rect 14096 44804 14148 44810
rect 14096 44746 14148 44752
rect 13728 44736 13780 44742
rect 13728 44678 13780 44684
rect 13636 44532 13688 44538
rect 13636 44474 13688 44480
rect 13740 43654 13768 44678
rect 13636 43648 13688 43654
rect 13636 43590 13688 43596
rect 13728 43648 13780 43654
rect 13728 43590 13780 43596
rect 13648 41414 13676 43590
rect 13740 42634 13768 43590
rect 14108 43178 14136 44746
rect 14188 44192 14240 44198
rect 14188 44134 14240 44140
rect 14096 43172 14148 43178
rect 14096 43114 14148 43120
rect 13728 42628 13780 42634
rect 13728 42570 13780 42576
rect 13740 42294 13768 42570
rect 13728 42288 13780 42294
rect 13728 42230 13780 42236
rect 13740 41614 13768 42230
rect 13820 42220 13872 42226
rect 13820 42162 13872 42168
rect 13728 41608 13780 41614
rect 13728 41550 13780 41556
rect 13648 41386 13768 41414
rect 13636 40928 13688 40934
rect 13636 40870 13688 40876
rect 13648 40526 13676 40870
rect 13636 40520 13688 40526
rect 13636 40462 13688 40468
rect 13556 40310 13676 40338
rect 13648 39574 13676 40310
rect 13740 40202 13768 41386
rect 13832 40934 13860 42162
rect 13820 40928 13872 40934
rect 13820 40870 13872 40876
rect 14004 40384 14056 40390
rect 14004 40326 14056 40332
rect 13740 40174 13860 40202
rect 13728 40112 13780 40118
rect 13728 40054 13780 40060
rect 13636 39568 13688 39574
rect 13636 39510 13688 39516
rect 13740 39098 13768 40054
rect 13832 39982 13860 40174
rect 13820 39976 13872 39982
rect 13820 39918 13872 39924
rect 13912 39840 13964 39846
rect 13912 39782 13964 39788
rect 13924 39506 13952 39782
rect 13912 39500 13964 39506
rect 13912 39442 13964 39448
rect 13728 39092 13780 39098
rect 13728 39034 13780 39040
rect 13728 37800 13780 37806
rect 13728 37742 13780 37748
rect 13544 36848 13596 36854
rect 13544 36790 13596 36796
rect 13452 35624 13504 35630
rect 13452 35566 13504 35572
rect 13464 34474 13492 35566
rect 13452 34468 13504 34474
rect 13452 34410 13504 34416
rect 13360 33992 13412 33998
rect 13360 33934 13412 33940
rect 13556 33386 13584 36790
rect 13740 35290 13768 37742
rect 14016 36122 14044 40326
rect 14108 38962 14136 43114
rect 14096 38956 14148 38962
rect 14096 38898 14148 38904
rect 13924 36094 14044 36122
rect 13820 35692 13872 35698
rect 13820 35634 13872 35640
rect 13832 35494 13860 35634
rect 13820 35488 13872 35494
rect 13820 35430 13872 35436
rect 13728 35284 13780 35290
rect 13648 35244 13728 35272
rect 13544 33380 13596 33386
rect 13544 33322 13596 33328
rect 13452 33312 13504 33318
rect 13452 33254 13504 33260
rect 12950 33212 13258 33221
rect 12950 33210 12956 33212
rect 13012 33210 13036 33212
rect 13092 33210 13116 33212
rect 13172 33210 13196 33212
rect 13252 33210 13258 33212
rect 13012 33158 13014 33210
rect 13194 33158 13196 33210
rect 12950 33156 12956 33158
rect 13012 33156 13036 33158
rect 13092 33156 13116 33158
rect 13172 33156 13196 33158
rect 13252 33156 13258 33158
rect 12950 33147 13258 33156
rect 13360 32768 13412 32774
rect 13360 32710 13412 32716
rect 13372 32570 13400 32710
rect 13360 32564 13412 32570
rect 13360 32506 13412 32512
rect 12950 32124 13258 32133
rect 12950 32122 12956 32124
rect 13012 32122 13036 32124
rect 13092 32122 13116 32124
rect 13172 32122 13196 32124
rect 13252 32122 13258 32124
rect 13012 32070 13014 32122
rect 13194 32070 13196 32122
rect 12950 32068 12956 32070
rect 13012 32068 13036 32070
rect 13092 32068 13116 32070
rect 13172 32068 13196 32070
rect 13252 32068 13258 32070
rect 12950 32059 13258 32068
rect 13360 31136 13412 31142
rect 13360 31078 13412 31084
rect 12950 31036 13258 31045
rect 12950 31034 12956 31036
rect 13012 31034 13036 31036
rect 13092 31034 13116 31036
rect 13172 31034 13196 31036
rect 13252 31034 13258 31036
rect 13012 30982 13014 31034
rect 13194 30982 13196 31034
rect 12950 30980 12956 30982
rect 13012 30980 13036 30982
rect 13092 30980 13116 30982
rect 13172 30980 13196 30982
rect 13252 30980 13258 30982
rect 12950 30971 13258 30980
rect 12808 30932 12860 30938
rect 12808 30874 12860 30880
rect 13372 30666 13400 31078
rect 13360 30660 13412 30666
rect 13360 30602 13412 30608
rect 12808 30592 12860 30598
rect 12808 30534 12860 30540
rect 12820 29850 12848 30534
rect 12990 30424 13046 30433
rect 12990 30359 13046 30368
rect 13004 30326 13032 30359
rect 12992 30320 13044 30326
rect 12992 30262 13044 30268
rect 12950 29948 13258 29957
rect 12950 29946 12956 29948
rect 13012 29946 13036 29948
rect 13092 29946 13116 29948
rect 13172 29946 13196 29948
rect 13252 29946 13258 29948
rect 13012 29894 13014 29946
rect 13194 29894 13196 29946
rect 12950 29892 12956 29894
rect 13012 29892 13036 29894
rect 13092 29892 13116 29894
rect 13172 29892 13196 29894
rect 13252 29892 13258 29894
rect 12950 29883 13258 29892
rect 12808 29844 12860 29850
rect 12808 29786 12860 29792
rect 12820 28626 12848 29786
rect 13464 29714 13492 33254
rect 13648 32978 13676 35244
rect 13728 35226 13780 35232
rect 13728 35080 13780 35086
rect 13728 35022 13780 35028
rect 13740 34746 13768 35022
rect 13832 35018 13860 35430
rect 13820 35012 13872 35018
rect 13820 34954 13872 34960
rect 13728 34740 13780 34746
rect 13728 34682 13780 34688
rect 13832 34626 13860 34954
rect 13740 34598 13860 34626
rect 13740 33862 13768 34598
rect 13728 33856 13780 33862
rect 13728 33798 13780 33804
rect 13636 32972 13688 32978
rect 13636 32914 13688 32920
rect 13740 32502 13768 33798
rect 13924 33658 13952 36094
rect 14200 35834 14228 44134
rect 14292 42770 14320 44814
rect 14568 44810 14596 47058
rect 14844 45558 14872 47194
rect 14832 45552 14884 45558
rect 14832 45494 14884 45500
rect 14556 44804 14608 44810
rect 14556 44746 14608 44752
rect 14556 44260 14608 44266
rect 14556 44202 14608 44208
rect 14280 42764 14332 42770
rect 14280 42706 14332 42712
rect 14568 42022 14596 44202
rect 14924 43852 14976 43858
rect 14924 43794 14976 43800
rect 14556 42016 14608 42022
rect 14556 41958 14608 41964
rect 14568 41206 14596 41958
rect 14372 41200 14424 41206
rect 14372 41142 14424 41148
rect 14556 41200 14608 41206
rect 14556 41142 14608 41148
rect 14384 40730 14412 41142
rect 14832 41064 14884 41070
rect 14832 41006 14884 41012
rect 14464 40928 14516 40934
rect 14464 40870 14516 40876
rect 14372 40724 14424 40730
rect 14372 40666 14424 40672
rect 14280 40180 14332 40186
rect 14280 40122 14332 40128
rect 14188 35828 14240 35834
rect 14188 35770 14240 35776
rect 14002 35320 14058 35329
rect 14002 35255 14004 35264
rect 14056 35255 14058 35264
rect 14004 35226 14056 35232
rect 14096 35148 14148 35154
rect 14096 35090 14148 35096
rect 14004 34944 14056 34950
rect 14004 34886 14056 34892
rect 14016 34746 14044 34886
rect 14004 34740 14056 34746
rect 14004 34682 14056 34688
rect 13820 33652 13872 33658
rect 13820 33594 13872 33600
rect 13912 33652 13964 33658
rect 13912 33594 13964 33600
rect 13728 32496 13780 32502
rect 13728 32438 13780 32444
rect 13728 32360 13780 32366
rect 13728 32302 13780 32308
rect 13740 31754 13768 32302
rect 13728 31748 13780 31754
rect 13728 31690 13780 31696
rect 13832 30802 13860 33594
rect 13912 33516 13964 33522
rect 13912 33458 13964 33464
rect 13924 33402 13952 33458
rect 14108 33454 14136 35090
rect 14096 33448 14148 33454
rect 14002 33416 14058 33425
rect 13924 33374 14002 33402
rect 14096 33390 14148 33396
rect 14002 33351 14058 33360
rect 14016 32774 14044 33351
rect 14004 32768 14056 32774
rect 14004 32710 14056 32716
rect 14016 31754 14044 32710
rect 14016 31726 14136 31754
rect 13820 30796 13872 30802
rect 13820 30738 13872 30744
rect 13544 30592 13596 30598
rect 13544 30534 13596 30540
rect 13452 29708 13504 29714
rect 13452 29650 13504 29656
rect 13084 29504 13136 29510
rect 13084 29446 13136 29452
rect 13096 29306 13124 29446
rect 12900 29300 12952 29306
rect 12900 29242 12952 29248
rect 13084 29300 13136 29306
rect 13084 29242 13136 29248
rect 12912 29034 12940 29242
rect 13360 29232 13412 29238
rect 13360 29174 13412 29180
rect 12900 29028 12952 29034
rect 12900 28970 12952 28976
rect 13372 28966 13400 29174
rect 13360 28960 13412 28966
rect 13360 28902 13412 28908
rect 12950 28860 13258 28869
rect 12950 28858 12956 28860
rect 13012 28858 13036 28860
rect 13092 28858 13116 28860
rect 13172 28858 13196 28860
rect 13252 28858 13258 28860
rect 13012 28806 13014 28858
rect 13194 28806 13196 28858
rect 12950 28804 12956 28806
rect 13012 28804 13036 28806
rect 13092 28804 13116 28806
rect 13172 28804 13196 28806
rect 13252 28804 13258 28806
rect 12950 28795 13258 28804
rect 12808 28620 12860 28626
rect 12808 28562 12860 28568
rect 13360 28008 13412 28014
rect 13360 27950 13412 27956
rect 12950 27772 13258 27781
rect 12950 27770 12956 27772
rect 13012 27770 13036 27772
rect 13092 27770 13116 27772
rect 13172 27770 13196 27772
rect 13252 27770 13258 27772
rect 13012 27718 13014 27770
rect 13194 27718 13196 27770
rect 12950 27716 12956 27718
rect 13012 27716 13036 27718
rect 13092 27716 13116 27718
rect 13172 27716 13196 27718
rect 13252 27716 13258 27718
rect 12950 27707 13258 27716
rect 13372 27470 13400 27950
rect 13452 27940 13504 27946
rect 13452 27882 13504 27888
rect 13360 27464 13412 27470
rect 13360 27406 13412 27412
rect 13464 26994 13492 27882
rect 13452 26988 13504 26994
rect 13452 26930 13504 26936
rect 12808 26920 12860 26926
rect 12808 26862 12860 26868
rect 12820 25702 12848 26862
rect 12950 26684 13258 26693
rect 12950 26682 12956 26684
rect 13012 26682 13036 26684
rect 13092 26682 13116 26684
rect 13172 26682 13196 26684
rect 13252 26682 13258 26684
rect 13012 26630 13014 26682
rect 13194 26630 13196 26682
rect 12950 26628 12956 26630
rect 13012 26628 13036 26630
rect 13092 26628 13116 26630
rect 13172 26628 13196 26630
rect 13252 26628 13258 26630
rect 12950 26619 13258 26628
rect 13464 26058 13492 26930
rect 13556 26382 13584 30534
rect 13728 29504 13780 29510
rect 13728 29446 13780 29452
rect 13636 28620 13688 28626
rect 13636 28562 13688 28568
rect 13648 26858 13676 28562
rect 13636 26852 13688 26858
rect 13636 26794 13688 26800
rect 13544 26376 13596 26382
rect 13544 26318 13596 26324
rect 13464 26030 13584 26058
rect 13268 25968 13320 25974
rect 13268 25910 13320 25916
rect 13280 25752 13308 25910
rect 13556 25906 13584 26030
rect 13544 25900 13596 25906
rect 13544 25842 13596 25848
rect 13648 25838 13676 26794
rect 13740 26602 13768 29446
rect 13820 28416 13872 28422
rect 13820 28358 13872 28364
rect 13832 27062 13860 28358
rect 14004 27872 14056 27878
rect 14004 27814 14056 27820
rect 13820 27056 13872 27062
rect 13820 26998 13872 27004
rect 13832 26738 13860 26998
rect 13832 26710 13952 26738
rect 13740 26574 13860 26602
rect 13924 26586 13952 26710
rect 13728 26512 13780 26518
rect 13728 26454 13780 26460
rect 13636 25832 13688 25838
rect 13636 25774 13688 25780
rect 13280 25724 13400 25752
rect 12808 25696 12860 25702
rect 12808 25638 12860 25644
rect 12950 25596 13258 25605
rect 12950 25594 12956 25596
rect 13012 25594 13036 25596
rect 13092 25594 13116 25596
rect 13172 25594 13196 25596
rect 13252 25594 13258 25596
rect 13012 25542 13014 25594
rect 13194 25542 13196 25594
rect 12950 25540 12956 25542
rect 13012 25540 13036 25542
rect 13092 25540 13116 25542
rect 13172 25540 13196 25542
rect 13252 25540 13258 25542
rect 12950 25531 13258 25540
rect 12728 24534 12848 24562
rect 12440 24404 12492 24410
rect 12440 24346 12492 24352
rect 12452 24138 12480 24346
rect 12440 24132 12492 24138
rect 12360 24092 12440 24120
rect 12256 22772 12308 22778
rect 12256 22714 12308 22720
rect 12164 22228 12216 22234
rect 12164 22170 12216 22176
rect 12164 21956 12216 21962
rect 12164 21898 12216 21904
rect 12176 21622 12204 21898
rect 12164 21616 12216 21622
rect 12164 21558 12216 21564
rect 12164 21344 12216 21350
rect 12164 21286 12216 21292
rect 12072 20868 12124 20874
rect 12072 20810 12124 20816
rect 11980 20528 12032 20534
rect 11980 20470 12032 20476
rect 11980 19916 12032 19922
rect 11980 19858 12032 19864
rect 11888 19508 11940 19514
rect 11888 19450 11940 19456
rect 11796 18624 11848 18630
rect 11796 18566 11848 18572
rect 11900 18034 11928 19450
rect 11716 18006 11928 18034
rect 11716 16726 11744 18006
rect 11888 17876 11940 17882
rect 11888 17818 11940 17824
rect 11796 16992 11848 16998
rect 11796 16934 11848 16940
rect 11704 16720 11756 16726
rect 11704 16662 11756 16668
rect 11704 16108 11756 16114
rect 11704 16050 11756 16056
rect 11612 14612 11664 14618
rect 11612 14554 11664 14560
rect 11532 12406 11652 12434
rect 11244 12300 11296 12306
rect 11244 12242 11296 12248
rect 11256 11694 11284 12242
rect 11244 11688 11296 11694
rect 11244 11630 11296 11636
rect 11256 11218 11284 11630
rect 11244 11212 11296 11218
rect 11244 11154 11296 11160
rect 11624 2582 11652 12406
rect 11716 6914 11744 16050
rect 11808 12986 11836 16934
rect 11900 15706 11928 17818
rect 11992 17746 12020 19858
rect 12072 18896 12124 18902
rect 12072 18838 12124 18844
rect 11980 17740 12032 17746
rect 11980 17682 12032 17688
rect 12084 17338 12112 18838
rect 12176 17338 12204 21286
rect 12072 17332 12124 17338
rect 12072 17274 12124 17280
rect 12164 17332 12216 17338
rect 12164 17274 12216 17280
rect 11888 15700 11940 15706
rect 11888 15642 11940 15648
rect 11796 12980 11848 12986
rect 11796 12922 11848 12928
rect 11900 10962 11928 15642
rect 12070 15328 12126 15337
rect 12070 15263 12126 15272
rect 11980 12096 12032 12102
rect 11980 12038 12032 12044
rect 11992 11830 12020 12038
rect 11980 11824 12032 11830
rect 11980 11766 12032 11772
rect 11992 11354 12020 11766
rect 11980 11348 12032 11354
rect 11980 11290 12032 11296
rect 11992 11082 12020 11290
rect 11980 11076 12032 11082
rect 11980 11018 12032 11024
rect 11900 10934 12020 10962
rect 11716 6886 11928 6914
rect 11796 3936 11848 3942
rect 11796 3878 11848 3884
rect 11808 2990 11836 3878
rect 11900 3398 11928 6886
rect 11992 6390 12020 10934
rect 11980 6384 12032 6390
rect 11980 6326 12032 6332
rect 12084 4010 12112 15263
rect 12268 15094 12296 22714
rect 12360 21146 12388 24092
rect 12440 24074 12492 24080
rect 12624 23180 12676 23186
rect 12624 23122 12676 23128
rect 12532 23044 12584 23050
rect 12532 22986 12584 22992
rect 12440 22976 12492 22982
rect 12440 22918 12492 22924
rect 12348 21140 12400 21146
rect 12348 21082 12400 21088
rect 12360 20806 12388 21082
rect 12348 20800 12400 20806
rect 12348 20742 12400 20748
rect 12452 20602 12480 22918
rect 12544 22710 12572 22986
rect 12532 22704 12584 22710
rect 12530 22672 12532 22681
rect 12584 22672 12586 22681
rect 12530 22607 12586 22616
rect 12636 22574 12664 23122
rect 12624 22568 12676 22574
rect 12624 22510 12676 22516
rect 12532 22228 12584 22234
rect 12532 22170 12584 22176
rect 12440 20596 12492 20602
rect 12440 20538 12492 20544
rect 12544 20058 12572 22170
rect 12624 21616 12676 21622
rect 12624 21558 12676 21564
rect 12636 21146 12664 21558
rect 12716 21480 12768 21486
rect 12716 21422 12768 21428
rect 12728 21146 12756 21422
rect 12624 21140 12676 21146
rect 12624 21082 12676 21088
rect 12716 21140 12768 21146
rect 12716 21082 12768 21088
rect 12820 21026 12848 24534
rect 12950 24508 13258 24517
rect 12950 24506 12956 24508
rect 13012 24506 13036 24508
rect 13092 24506 13116 24508
rect 13172 24506 13196 24508
rect 13252 24506 13258 24508
rect 13012 24454 13014 24506
rect 13194 24454 13196 24506
rect 12950 24452 12956 24454
rect 13012 24452 13036 24454
rect 13092 24452 13116 24454
rect 13172 24452 13196 24454
rect 13252 24452 13258 24454
rect 12950 24443 13258 24452
rect 12950 23420 13258 23429
rect 12950 23418 12956 23420
rect 13012 23418 13036 23420
rect 13092 23418 13116 23420
rect 13172 23418 13196 23420
rect 13252 23418 13258 23420
rect 13012 23366 13014 23418
rect 13194 23366 13196 23418
rect 12950 23364 12956 23366
rect 13012 23364 13036 23366
rect 13092 23364 13116 23366
rect 13172 23364 13196 23366
rect 13252 23364 13258 23366
rect 12950 23355 13258 23364
rect 13176 23316 13228 23322
rect 13176 23258 13228 23264
rect 12992 23112 13044 23118
rect 12992 23054 13044 23060
rect 13004 22778 13032 23054
rect 13188 22982 13216 23258
rect 13176 22976 13228 22982
rect 13176 22918 13228 22924
rect 12992 22772 13044 22778
rect 12992 22714 13044 22720
rect 13372 22642 13400 25724
rect 13452 25696 13504 25702
rect 13452 25638 13504 25644
rect 13464 24274 13492 25638
rect 13636 24608 13688 24614
rect 13636 24550 13688 24556
rect 13452 24268 13504 24274
rect 13452 24210 13504 24216
rect 13648 24206 13676 24550
rect 13636 24200 13688 24206
rect 13636 24142 13688 24148
rect 13544 24064 13596 24070
rect 13544 24006 13596 24012
rect 13556 23866 13584 24006
rect 13544 23860 13596 23866
rect 13544 23802 13596 23808
rect 13648 23662 13676 24142
rect 13740 23730 13768 26454
rect 13832 25430 13860 26574
rect 13912 26580 13964 26586
rect 13912 26522 13964 26528
rect 13924 26042 13952 26522
rect 13912 26036 13964 26042
rect 13912 25978 13964 25984
rect 13912 25900 13964 25906
rect 13912 25842 13964 25848
rect 13820 25424 13872 25430
rect 13820 25366 13872 25372
rect 13820 24676 13872 24682
rect 13820 24618 13872 24624
rect 13832 24070 13860 24618
rect 13820 24064 13872 24070
rect 13820 24006 13872 24012
rect 13728 23724 13780 23730
rect 13728 23666 13780 23672
rect 13636 23656 13688 23662
rect 13636 23598 13688 23604
rect 13726 23352 13782 23361
rect 13726 23287 13728 23296
rect 13780 23287 13782 23296
rect 13728 23258 13780 23264
rect 13636 23180 13688 23186
rect 13636 23122 13688 23128
rect 13452 22772 13504 22778
rect 13452 22714 13504 22720
rect 13360 22636 13412 22642
rect 13360 22578 13412 22584
rect 13176 22568 13228 22574
rect 13174 22536 13176 22545
rect 13228 22536 13230 22545
rect 13174 22471 13230 22480
rect 12950 22332 13258 22341
rect 12950 22330 12956 22332
rect 13012 22330 13036 22332
rect 13092 22330 13116 22332
rect 13172 22330 13196 22332
rect 13252 22330 13258 22332
rect 13012 22278 13014 22330
rect 13194 22278 13196 22330
rect 12950 22276 12956 22278
rect 13012 22276 13036 22278
rect 13092 22276 13116 22278
rect 13172 22276 13196 22278
rect 13252 22276 13258 22278
rect 12950 22267 13258 22276
rect 12992 22092 13044 22098
rect 12992 22034 13044 22040
rect 13004 21894 13032 22034
rect 12992 21888 13044 21894
rect 12992 21830 13044 21836
rect 12900 21480 12952 21486
rect 12898 21448 12900 21457
rect 12952 21448 12954 21457
rect 12898 21383 12954 21392
rect 12950 21244 13258 21253
rect 12950 21242 12956 21244
rect 13012 21242 13036 21244
rect 13092 21242 13116 21244
rect 13172 21242 13196 21244
rect 13252 21242 13258 21244
rect 13012 21190 13014 21242
rect 13194 21190 13196 21242
rect 12950 21188 12956 21190
rect 13012 21188 13036 21190
rect 13092 21188 13116 21190
rect 13172 21188 13196 21190
rect 13252 21188 13258 21190
rect 12950 21179 13258 21188
rect 12636 20998 12848 21026
rect 13372 21010 13400 22578
rect 13464 21049 13492 22714
rect 13544 22704 13596 22710
rect 13544 22646 13596 22652
rect 13556 22234 13584 22646
rect 13544 22228 13596 22234
rect 13544 22170 13596 22176
rect 13556 22098 13584 22170
rect 13544 22092 13596 22098
rect 13544 22034 13596 22040
rect 13544 21548 13596 21554
rect 13544 21490 13596 21496
rect 13450 21040 13506 21049
rect 13360 21004 13412 21010
rect 12532 20052 12584 20058
rect 12532 19994 12584 20000
rect 12440 19372 12492 19378
rect 12440 19314 12492 19320
rect 12452 18426 12480 19314
rect 12544 18850 12572 19994
rect 12636 18970 12664 20998
rect 13450 20975 13506 20984
rect 13360 20946 13412 20952
rect 13556 20942 13584 21490
rect 13544 20936 13596 20942
rect 13544 20878 13596 20884
rect 13648 20618 13676 23122
rect 13728 22976 13780 22982
rect 13728 22918 13780 22924
rect 13740 22710 13768 22918
rect 13728 22704 13780 22710
rect 13728 22646 13780 22652
rect 13728 21888 13780 21894
rect 13820 21888 13872 21894
rect 13728 21830 13780 21836
rect 13818 21856 13820 21865
rect 13872 21856 13874 21865
rect 13372 20590 13676 20618
rect 12950 20156 13258 20165
rect 12950 20154 12956 20156
rect 13012 20154 13036 20156
rect 13092 20154 13116 20156
rect 13172 20154 13196 20156
rect 13252 20154 13258 20156
rect 13012 20102 13014 20154
rect 13194 20102 13196 20154
rect 12950 20100 12956 20102
rect 13012 20100 13036 20102
rect 13092 20100 13116 20102
rect 13172 20100 13196 20102
rect 13252 20100 13258 20102
rect 12950 20091 13258 20100
rect 13084 19780 13136 19786
rect 13084 19722 13136 19728
rect 13096 19514 13124 19722
rect 13084 19508 13136 19514
rect 13084 19450 13136 19456
rect 12716 19440 12768 19446
rect 13372 19394 13400 20590
rect 13452 20528 13504 20534
rect 13452 20470 13504 20476
rect 12716 19382 12768 19388
rect 12624 18964 12676 18970
rect 12624 18906 12676 18912
rect 12544 18822 12664 18850
rect 12532 18760 12584 18766
rect 12532 18702 12584 18708
rect 12440 18420 12492 18426
rect 12440 18362 12492 18368
rect 12544 18306 12572 18702
rect 12452 18290 12572 18306
rect 12440 18284 12572 18290
rect 12492 18278 12572 18284
rect 12440 18226 12492 18232
rect 12452 18154 12480 18226
rect 12440 18148 12492 18154
rect 12440 18090 12492 18096
rect 12452 16998 12480 18090
rect 12532 17536 12584 17542
rect 12532 17478 12584 17484
rect 12440 16992 12492 16998
rect 12440 16934 12492 16940
rect 12452 16130 12480 16934
rect 12544 16250 12572 17478
rect 12532 16244 12584 16250
rect 12532 16186 12584 16192
rect 12452 16102 12572 16130
rect 12256 15088 12308 15094
rect 12256 15030 12308 15036
rect 12440 15020 12492 15026
rect 12440 14962 12492 14968
rect 12256 14952 12308 14958
rect 12256 14894 12308 14900
rect 12268 14414 12296 14894
rect 12256 14408 12308 14414
rect 12256 14350 12308 14356
rect 12164 13864 12216 13870
rect 12164 13806 12216 13812
rect 12176 6914 12204 13806
rect 12268 11694 12296 14350
rect 12452 13530 12480 14962
rect 12544 13802 12572 16102
rect 12532 13796 12584 13802
rect 12532 13738 12584 13744
rect 12440 13524 12492 13530
rect 12440 13466 12492 13472
rect 12440 13388 12492 13394
rect 12440 13330 12492 13336
rect 12452 12442 12480 13330
rect 12440 12436 12492 12442
rect 12440 12378 12492 12384
rect 12256 11688 12308 11694
rect 12256 11630 12308 11636
rect 12452 11370 12480 12378
rect 12544 12050 12572 13738
rect 12636 12170 12664 18822
rect 12728 18222 12756 19382
rect 12820 19366 13400 19394
rect 12820 18834 12848 19366
rect 13360 19236 13412 19242
rect 13360 19178 13412 19184
rect 12950 19068 13258 19077
rect 12950 19066 12956 19068
rect 13012 19066 13036 19068
rect 13092 19066 13116 19068
rect 13172 19066 13196 19068
rect 13252 19066 13258 19068
rect 13012 19014 13014 19066
rect 13194 19014 13196 19066
rect 12950 19012 12956 19014
rect 13012 19012 13036 19014
rect 13092 19012 13116 19014
rect 13172 19012 13196 19014
rect 13252 19012 13258 19014
rect 12950 19003 13258 19012
rect 12808 18828 12860 18834
rect 12808 18770 12860 18776
rect 13372 18222 13400 19178
rect 12716 18216 12768 18222
rect 12716 18158 12768 18164
rect 13360 18216 13412 18222
rect 13360 18158 13412 18164
rect 12728 17338 12756 18158
rect 12950 17980 13258 17989
rect 12950 17978 12956 17980
rect 13012 17978 13036 17980
rect 13092 17978 13116 17980
rect 13172 17978 13196 17980
rect 13252 17978 13258 17980
rect 13012 17926 13014 17978
rect 13194 17926 13196 17978
rect 12950 17924 12956 17926
rect 13012 17924 13036 17926
rect 13092 17924 13116 17926
rect 13172 17924 13196 17926
rect 13252 17924 13258 17926
rect 12806 17912 12862 17921
rect 12950 17915 13258 17924
rect 12806 17847 12808 17856
rect 12860 17847 12862 17856
rect 12808 17818 12860 17824
rect 12716 17332 12768 17338
rect 12716 17274 12768 17280
rect 12716 17196 12768 17202
rect 12716 17138 12768 17144
rect 12728 14074 12756 17138
rect 12820 16114 12848 17818
rect 12950 16892 13258 16901
rect 12950 16890 12956 16892
rect 13012 16890 13036 16892
rect 13092 16890 13116 16892
rect 13172 16890 13196 16892
rect 13252 16890 13258 16892
rect 13012 16838 13014 16890
rect 13194 16838 13196 16890
rect 12950 16836 12956 16838
rect 13012 16836 13036 16838
rect 13092 16836 13116 16838
rect 13172 16836 13196 16838
rect 13252 16836 13258 16838
rect 12950 16827 13258 16836
rect 12808 16108 12860 16114
rect 12808 16050 12860 16056
rect 12806 16008 12862 16017
rect 12806 15943 12862 15952
rect 12820 15706 12848 15943
rect 12950 15804 13258 15813
rect 12950 15802 12956 15804
rect 13012 15802 13036 15804
rect 13092 15802 13116 15804
rect 13172 15802 13196 15804
rect 13252 15802 13258 15804
rect 13012 15750 13014 15802
rect 13194 15750 13196 15802
rect 12950 15748 12956 15750
rect 13012 15748 13036 15750
rect 13092 15748 13116 15750
rect 13172 15748 13196 15750
rect 13252 15748 13258 15750
rect 12950 15739 13258 15748
rect 12808 15700 12860 15706
rect 12808 15642 12860 15648
rect 12820 15094 12848 15642
rect 12808 15088 12860 15094
rect 12808 15030 12860 15036
rect 12950 14716 13258 14725
rect 12950 14714 12956 14716
rect 13012 14714 13036 14716
rect 13092 14714 13116 14716
rect 13172 14714 13196 14716
rect 13252 14714 13258 14716
rect 13012 14662 13014 14714
rect 13194 14662 13196 14714
rect 12950 14660 12956 14662
rect 13012 14660 13036 14662
rect 13092 14660 13116 14662
rect 13172 14660 13196 14662
rect 13252 14660 13258 14662
rect 12950 14651 13258 14660
rect 13372 14482 13400 18158
rect 13176 14476 13228 14482
rect 13176 14418 13228 14424
rect 13360 14476 13412 14482
rect 13360 14418 13412 14424
rect 13084 14272 13136 14278
rect 13084 14214 13136 14220
rect 13096 14074 13124 14214
rect 13188 14074 13216 14418
rect 12716 14068 12768 14074
rect 12716 14010 12768 14016
rect 13084 14068 13136 14074
rect 13084 14010 13136 14016
rect 13176 14068 13228 14074
rect 13176 14010 13228 14016
rect 13188 13870 13216 14010
rect 13176 13864 13228 13870
rect 13176 13806 13228 13812
rect 12950 13628 13258 13637
rect 12950 13626 12956 13628
rect 13012 13626 13036 13628
rect 13092 13626 13116 13628
rect 13172 13626 13196 13628
rect 13252 13626 13258 13628
rect 13012 13574 13014 13626
rect 13194 13574 13196 13626
rect 12950 13572 12956 13574
rect 13012 13572 13036 13574
rect 13092 13572 13116 13574
rect 13172 13572 13196 13574
rect 13252 13572 13258 13574
rect 12950 13563 13258 13572
rect 13464 12986 13492 20470
rect 13636 20460 13688 20466
rect 13636 20402 13688 20408
rect 13544 19304 13596 19310
rect 13544 19246 13596 19252
rect 13556 18766 13584 19246
rect 13544 18760 13596 18766
rect 13544 18702 13596 18708
rect 13544 18624 13596 18630
rect 13544 18566 13596 18572
rect 13556 14770 13584 18566
rect 13648 18426 13676 20402
rect 13740 18698 13768 21830
rect 13818 21791 13874 21800
rect 13924 19446 13952 25842
rect 14016 23798 14044 27814
rect 14004 23792 14056 23798
rect 14004 23734 14056 23740
rect 14004 21412 14056 21418
rect 14004 21354 14056 21360
rect 14016 21146 14044 21354
rect 14004 21140 14056 21146
rect 14004 21082 14056 21088
rect 13912 19440 13964 19446
rect 13912 19382 13964 19388
rect 14016 18902 14044 21082
rect 14004 18896 14056 18902
rect 14004 18838 14056 18844
rect 13728 18692 13780 18698
rect 13728 18634 13780 18640
rect 13636 18420 13688 18426
rect 13636 18362 13688 18368
rect 13912 18284 13964 18290
rect 13912 18226 13964 18232
rect 13820 18216 13872 18222
rect 13820 18158 13872 18164
rect 13832 18034 13860 18158
rect 13924 18086 13952 18226
rect 13740 18006 13860 18034
rect 13912 18080 13964 18086
rect 13912 18022 13964 18028
rect 13740 17882 13768 18006
rect 13924 17898 13952 18022
rect 13728 17876 13780 17882
rect 13728 17818 13780 17824
rect 13832 17870 13952 17898
rect 13832 17762 13860 17870
rect 13636 17740 13688 17746
rect 13636 17682 13688 17688
rect 13740 17734 13860 17762
rect 13912 17740 13964 17746
rect 13648 16454 13676 17682
rect 13740 17338 13768 17734
rect 13912 17682 13964 17688
rect 13728 17332 13780 17338
rect 13728 17274 13780 17280
rect 13924 17202 13952 17682
rect 13912 17196 13964 17202
rect 13912 17138 13964 17144
rect 13728 17128 13780 17134
rect 13780 17088 13860 17116
rect 13728 17070 13780 17076
rect 13636 16448 13688 16454
rect 13636 16390 13688 16396
rect 13648 14958 13676 16390
rect 13636 14952 13688 14958
rect 13636 14894 13688 14900
rect 13556 14742 13676 14770
rect 13544 13524 13596 13530
rect 13544 13466 13596 13472
rect 12808 12980 12860 12986
rect 12808 12922 12860 12928
rect 13452 12980 13504 12986
rect 13452 12922 13504 12928
rect 12820 12238 12848 12922
rect 13556 12850 13584 13466
rect 13452 12844 13504 12850
rect 13452 12786 13504 12792
rect 13544 12844 13596 12850
rect 13544 12786 13596 12792
rect 12950 12540 13258 12549
rect 12950 12538 12956 12540
rect 13012 12538 13036 12540
rect 13092 12538 13116 12540
rect 13172 12538 13196 12540
rect 13252 12538 13258 12540
rect 13012 12486 13014 12538
rect 13194 12486 13196 12538
rect 12950 12484 12956 12486
rect 13012 12484 13036 12486
rect 13092 12484 13116 12486
rect 13172 12484 13196 12486
rect 13252 12484 13258 12486
rect 12950 12475 13258 12484
rect 13464 12442 13492 12786
rect 13648 12730 13676 14742
rect 13556 12702 13676 12730
rect 13452 12436 13504 12442
rect 13452 12378 13504 12384
rect 12808 12232 12860 12238
rect 12808 12174 12860 12180
rect 12624 12164 12676 12170
rect 12624 12106 12676 12112
rect 13452 12164 13504 12170
rect 13452 12106 13504 12112
rect 12716 12096 12768 12102
rect 12544 12022 12664 12050
rect 12716 12038 12768 12044
rect 12452 11342 12572 11370
rect 12544 11218 12572 11342
rect 12532 11212 12584 11218
rect 12532 11154 12584 11160
rect 12348 9988 12400 9994
rect 12348 9930 12400 9936
rect 12176 6886 12296 6914
rect 12072 4004 12124 4010
rect 12072 3946 12124 3952
rect 11888 3392 11940 3398
rect 11888 3334 11940 3340
rect 12268 3058 12296 6886
rect 12256 3052 12308 3058
rect 12256 2994 12308 3000
rect 11796 2984 11848 2990
rect 11796 2926 11848 2932
rect 11612 2576 11664 2582
rect 11612 2518 11664 2524
rect 11060 2440 11112 2446
rect 11060 2382 11112 2388
rect 11428 2440 11480 2446
rect 11428 2382 11480 2388
rect 10968 2304 11020 2310
rect 11020 2264 11100 2292
rect 10968 2246 11020 2252
rect 11072 800 11100 2264
rect 11440 800 11468 2382
rect 11808 800 11836 2926
rect 12164 2508 12216 2514
rect 12164 2450 12216 2456
rect 12176 800 12204 2450
rect 12360 2446 12388 9930
rect 12636 8566 12664 12022
rect 12624 8560 12676 8566
rect 12624 8502 12676 8508
rect 12728 4146 12756 12038
rect 13360 11688 13412 11694
rect 13360 11630 13412 11636
rect 12950 11452 13258 11461
rect 12950 11450 12956 11452
rect 13012 11450 13036 11452
rect 13092 11450 13116 11452
rect 13172 11450 13196 11452
rect 13252 11450 13258 11452
rect 13012 11398 13014 11450
rect 13194 11398 13196 11450
rect 12950 11396 12956 11398
rect 13012 11396 13036 11398
rect 13092 11396 13116 11398
rect 13172 11396 13196 11398
rect 13252 11396 13258 11398
rect 12950 11387 13258 11396
rect 13372 11218 13400 11630
rect 13464 11286 13492 12106
rect 13452 11280 13504 11286
rect 13452 11222 13504 11228
rect 13360 11212 13412 11218
rect 13360 11154 13412 11160
rect 12950 10364 13258 10373
rect 12950 10362 12956 10364
rect 13012 10362 13036 10364
rect 13092 10362 13116 10364
rect 13172 10362 13196 10364
rect 13252 10362 13258 10364
rect 13012 10310 13014 10362
rect 13194 10310 13196 10362
rect 12950 10308 12956 10310
rect 13012 10308 13036 10310
rect 13092 10308 13116 10310
rect 13172 10308 13196 10310
rect 13252 10308 13258 10310
rect 12950 10299 13258 10308
rect 13556 9654 13584 12702
rect 13832 12458 13860 17088
rect 13740 12430 13860 12458
rect 13740 9674 13768 12430
rect 13820 11892 13872 11898
rect 13820 11834 13872 11840
rect 13832 10810 13860 11834
rect 13820 10804 13872 10810
rect 13820 10746 13872 10752
rect 13544 9648 13596 9654
rect 13544 9590 13596 9596
rect 13648 9646 13768 9674
rect 12950 9276 13258 9285
rect 12950 9274 12956 9276
rect 13012 9274 13036 9276
rect 13092 9274 13116 9276
rect 13172 9274 13196 9276
rect 13252 9274 13258 9276
rect 13012 9222 13014 9274
rect 13194 9222 13196 9274
rect 12950 9220 12956 9222
rect 13012 9220 13036 9222
rect 13092 9220 13116 9222
rect 13172 9220 13196 9222
rect 13252 9220 13258 9222
rect 12950 9211 13258 9220
rect 12950 8188 13258 8197
rect 12950 8186 12956 8188
rect 13012 8186 13036 8188
rect 13092 8186 13116 8188
rect 13172 8186 13196 8188
rect 13252 8186 13258 8188
rect 13012 8134 13014 8186
rect 13194 8134 13196 8186
rect 12950 8132 12956 8134
rect 13012 8132 13036 8134
rect 13092 8132 13116 8134
rect 13172 8132 13196 8134
rect 13252 8132 13258 8134
rect 12950 8123 13258 8132
rect 12950 7100 13258 7109
rect 12950 7098 12956 7100
rect 13012 7098 13036 7100
rect 13092 7098 13116 7100
rect 13172 7098 13196 7100
rect 13252 7098 13258 7100
rect 13012 7046 13014 7098
rect 13194 7046 13196 7098
rect 12950 7044 12956 7046
rect 13012 7044 13036 7046
rect 13092 7044 13116 7046
rect 13172 7044 13196 7046
rect 13252 7044 13258 7046
rect 12950 7035 13258 7044
rect 12950 6012 13258 6021
rect 12950 6010 12956 6012
rect 13012 6010 13036 6012
rect 13092 6010 13116 6012
rect 13172 6010 13196 6012
rect 13252 6010 13258 6012
rect 13012 5958 13014 6010
rect 13194 5958 13196 6010
rect 12950 5956 12956 5958
rect 13012 5956 13036 5958
rect 13092 5956 13116 5958
rect 13172 5956 13196 5958
rect 13252 5956 13258 5958
rect 12950 5947 13258 5956
rect 12950 4924 13258 4933
rect 12950 4922 12956 4924
rect 13012 4922 13036 4924
rect 13092 4922 13116 4924
rect 13172 4922 13196 4924
rect 13252 4922 13258 4924
rect 13012 4870 13014 4922
rect 13194 4870 13196 4922
rect 12950 4868 12956 4870
rect 13012 4868 13036 4870
rect 13092 4868 13116 4870
rect 13172 4868 13196 4870
rect 13252 4868 13258 4870
rect 12950 4859 13258 4868
rect 12716 4140 12768 4146
rect 12716 4082 12768 4088
rect 12808 4072 12860 4078
rect 12808 4014 12860 4020
rect 12532 3460 12584 3466
rect 12532 3402 12584 3408
rect 12348 2440 12400 2446
rect 12348 2382 12400 2388
rect 12544 800 12572 3402
rect 12820 2122 12848 4014
rect 12950 3836 13258 3845
rect 12950 3834 12956 3836
rect 13012 3834 13036 3836
rect 13092 3834 13116 3836
rect 13172 3834 13196 3836
rect 13252 3834 13258 3836
rect 13012 3782 13014 3834
rect 13194 3782 13196 3834
rect 12950 3780 12956 3782
rect 13012 3780 13036 3782
rect 13092 3780 13116 3782
rect 13172 3780 13196 3782
rect 13252 3780 13258 3782
rect 12950 3771 13258 3780
rect 13648 3738 13676 9646
rect 13924 5574 13952 17138
rect 14016 14346 14044 18838
rect 14004 14340 14056 14346
rect 14004 14282 14056 14288
rect 14108 13394 14136 31726
rect 14200 28762 14228 35770
rect 14292 34678 14320 40122
rect 14384 40118 14412 40666
rect 14372 40112 14424 40118
rect 14372 40054 14424 40060
rect 14372 39976 14424 39982
rect 14372 39918 14424 39924
rect 14384 39098 14412 39918
rect 14476 39642 14504 40870
rect 14464 39636 14516 39642
rect 14464 39578 14516 39584
rect 14648 39296 14700 39302
rect 14648 39238 14700 39244
rect 14372 39092 14424 39098
rect 14372 39034 14424 39040
rect 14464 38208 14516 38214
rect 14464 38150 14516 38156
rect 14476 36922 14504 38150
rect 14464 36916 14516 36922
rect 14464 36858 14516 36864
rect 14554 36816 14610 36825
rect 14554 36751 14610 36760
rect 14568 36038 14596 36751
rect 14556 36032 14608 36038
rect 14556 35974 14608 35980
rect 14372 35692 14424 35698
rect 14372 35634 14424 35640
rect 14280 34672 14332 34678
rect 14280 34614 14332 34620
rect 14280 30728 14332 30734
rect 14280 30670 14332 30676
rect 14188 28756 14240 28762
rect 14188 28698 14240 28704
rect 14200 25906 14228 28698
rect 14292 28626 14320 30670
rect 14384 30190 14412 35634
rect 14660 35222 14688 39238
rect 14740 39024 14792 39030
rect 14740 38966 14792 38972
rect 14752 36038 14780 38966
rect 14740 36032 14792 36038
rect 14740 35974 14792 35980
rect 14740 35624 14792 35630
rect 14740 35566 14792 35572
rect 14648 35216 14700 35222
rect 14648 35158 14700 35164
rect 14752 35086 14780 35566
rect 14844 35562 14872 41006
rect 14936 38758 14964 43794
rect 15016 42628 15068 42634
rect 15016 42570 15068 42576
rect 15028 42294 15056 42570
rect 15016 42288 15068 42294
rect 15016 42230 15068 42236
rect 14924 38752 14976 38758
rect 14924 38694 14976 38700
rect 14924 37664 14976 37670
rect 14924 37606 14976 37612
rect 14832 35556 14884 35562
rect 14832 35498 14884 35504
rect 14740 35080 14792 35086
rect 14740 35022 14792 35028
rect 14462 34504 14518 34513
rect 14462 34439 14518 34448
rect 14476 32366 14504 34439
rect 14556 34400 14608 34406
rect 14556 34342 14608 34348
rect 14568 32910 14596 34342
rect 14936 33658 14964 37606
rect 15016 36236 15068 36242
rect 15016 36178 15068 36184
rect 15028 35766 15056 36178
rect 15016 35760 15068 35766
rect 15016 35702 15068 35708
rect 14924 33652 14976 33658
rect 14924 33594 14976 33600
rect 15016 33516 15068 33522
rect 15016 33458 15068 33464
rect 15028 33114 15056 33458
rect 15016 33108 15068 33114
rect 15016 33050 15068 33056
rect 15120 32994 15148 53926
rect 15580 53786 15608 54148
rect 15844 54130 15896 54136
rect 15660 54052 15712 54058
rect 15660 53994 15712 54000
rect 15672 53961 15700 53994
rect 15658 53952 15714 53961
rect 15658 53887 15714 53896
rect 15568 53780 15620 53786
rect 15568 53722 15620 53728
rect 15580 53582 15608 53722
rect 15568 53576 15620 53582
rect 15568 53518 15620 53524
rect 15752 53440 15804 53446
rect 15752 53382 15804 53388
rect 15476 46504 15528 46510
rect 15476 46446 15528 46452
rect 15488 45490 15516 46446
rect 15476 45484 15528 45490
rect 15476 45426 15528 45432
rect 15292 45280 15344 45286
rect 15292 45222 15344 45228
rect 15304 44810 15332 45222
rect 15292 44804 15344 44810
rect 15292 44746 15344 44752
rect 15384 44260 15436 44266
rect 15384 44202 15436 44208
rect 15200 39840 15252 39846
rect 15200 39782 15252 39788
rect 15212 39438 15240 39782
rect 15200 39432 15252 39438
rect 15200 39374 15252 39380
rect 15200 38956 15252 38962
rect 15200 38898 15252 38904
rect 15212 38010 15240 38898
rect 15292 38752 15344 38758
rect 15290 38720 15292 38729
rect 15344 38720 15346 38729
rect 15290 38655 15346 38664
rect 15304 38282 15332 38655
rect 15292 38276 15344 38282
rect 15292 38218 15344 38224
rect 15396 38010 15424 44202
rect 15488 43858 15516 45426
rect 15476 43852 15528 43858
rect 15476 43794 15528 43800
rect 15488 42226 15516 43794
rect 15660 43308 15712 43314
rect 15660 43250 15712 43256
rect 15568 42560 15620 42566
rect 15568 42502 15620 42508
rect 15476 42220 15528 42226
rect 15476 42162 15528 42168
rect 15488 41682 15516 42162
rect 15580 42158 15608 42502
rect 15568 42152 15620 42158
rect 15568 42094 15620 42100
rect 15476 41676 15528 41682
rect 15476 41618 15528 41624
rect 15488 41138 15516 41618
rect 15476 41132 15528 41138
rect 15476 41074 15528 41080
rect 15476 40384 15528 40390
rect 15476 40326 15528 40332
rect 15488 39098 15516 40326
rect 15476 39092 15528 39098
rect 15476 39034 15528 39040
rect 15580 38894 15608 42094
rect 15672 40730 15700 43250
rect 15660 40724 15712 40730
rect 15660 40666 15712 40672
rect 15660 40520 15712 40526
rect 15660 40462 15712 40468
rect 15568 38888 15620 38894
rect 15568 38830 15620 38836
rect 15568 38412 15620 38418
rect 15568 38354 15620 38360
rect 15200 38004 15252 38010
rect 15200 37946 15252 37952
rect 15384 38004 15436 38010
rect 15384 37946 15436 37952
rect 15580 37942 15608 38354
rect 15568 37936 15620 37942
rect 15568 37878 15620 37884
rect 15200 37868 15252 37874
rect 15200 37810 15252 37816
rect 15212 36802 15240 37810
rect 15292 37256 15344 37262
rect 15292 37198 15344 37204
rect 15304 36922 15332 37198
rect 15476 37120 15528 37126
rect 15476 37062 15528 37068
rect 15292 36916 15344 36922
rect 15292 36858 15344 36864
rect 15384 36848 15436 36854
rect 15212 36774 15332 36802
rect 15384 36790 15436 36796
rect 15200 36644 15252 36650
rect 15200 36586 15252 36592
rect 15212 36174 15240 36586
rect 15200 36168 15252 36174
rect 15200 36110 15252 36116
rect 14660 32966 15148 32994
rect 14556 32904 14608 32910
rect 14556 32846 14608 32852
rect 14568 32366 14596 32846
rect 14464 32360 14516 32366
rect 14464 32302 14516 32308
rect 14556 32360 14608 32366
rect 14556 32302 14608 32308
rect 14556 32224 14608 32230
rect 14556 32166 14608 32172
rect 14464 31680 14516 31686
rect 14464 31622 14516 31628
rect 14476 30666 14504 31622
rect 14568 30666 14596 32166
rect 14464 30660 14516 30666
rect 14464 30602 14516 30608
rect 14556 30660 14608 30666
rect 14556 30602 14608 30608
rect 14372 30184 14424 30190
rect 14372 30126 14424 30132
rect 14476 30002 14504 30602
rect 14384 29974 14504 30002
rect 14280 28620 14332 28626
rect 14280 28562 14332 28568
rect 14280 27328 14332 27334
rect 14280 27270 14332 27276
rect 14188 25900 14240 25906
rect 14188 25842 14240 25848
rect 14188 24744 14240 24750
rect 14188 24686 14240 24692
rect 14200 19854 14228 24686
rect 14292 22030 14320 27270
rect 14280 22024 14332 22030
rect 14280 21966 14332 21972
rect 14384 21894 14412 29974
rect 14568 27538 14596 30602
rect 14660 29306 14688 32966
rect 15108 32904 15160 32910
rect 15108 32846 15160 32852
rect 14924 32564 14976 32570
rect 14924 32506 14976 32512
rect 14832 30048 14884 30054
rect 14832 29990 14884 29996
rect 14648 29300 14700 29306
rect 14648 29242 14700 29248
rect 14738 29064 14794 29073
rect 14738 28999 14794 29008
rect 14752 28014 14780 28999
rect 14740 28008 14792 28014
rect 14740 27950 14792 27956
rect 14556 27532 14608 27538
rect 14556 27474 14608 27480
rect 14464 27328 14516 27334
rect 14464 27270 14516 27276
rect 14476 26314 14504 27270
rect 14648 26784 14700 26790
rect 14648 26726 14700 26732
rect 14556 26376 14608 26382
rect 14556 26318 14608 26324
rect 14464 26308 14516 26314
rect 14464 26250 14516 26256
rect 14568 24886 14596 26318
rect 14556 24880 14608 24886
rect 14556 24822 14608 24828
rect 14660 24274 14688 26726
rect 14648 24268 14700 24274
rect 14648 24210 14700 24216
rect 14752 23508 14780 27950
rect 14844 27334 14872 29990
rect 14936 27470 14964 32506
rect 15016 30252 15068 30258
rect 15016 30194 15068 30200
rect 15028 29782 15056 30194
rect 15120 29850 15148 32846
rect 15108 29844 15160 29850
rect 15108 29786 15160 29792
rect 15016 29776 15068 29782
rect 15016 29718 15068 29724
rect 15212 29034 15240 36110
rect 15200 29028 15252 29034
rect 15200 28970 15252 28976
rect 14924 27464 14976 27470
rect 14924 27406 14976 27412
rect 14832 27328 14884 27334
rect 14832 27270 14884 27276
rect 14924 27056 14976 27062
rect 14924 26998 14976 27004
rect 14476 23480 14780 23508
rect 14832 23520 14884 23526
rect 14280 21888 14332 21894
rect 14280 21830 14332 21836
rect 14372 21888 14424 21894
rect 14372 21830 14424 21836
rect 14188 19848 14240 19854
rect 14188 19790 14240 19796
rect 14188 18624 14240 18630
rect 14188 18566 14240 18572
rect 14200 13530 14228 18566
rect 14292 17678 14320 21830
rect 14384 21486 14412 21830
rect 14372 21480 14424 21486
rect 14372 21422 14424 21428
rect 14372 20256 14424 20262
rect 14372 20198 14424 20204
rect 14280 17672 14332 17678
rect 14280 17614 14332 17620
rect 14384 17270 14412 20198
rect 14372 17264 14424 17270
rect 14372 17206 14424 17212
rect 14476 15502 14504 23480
rect 14832 23462 14884 23468
rect 14556 22772 14608 22778
rect 14556 22714 14608 22720
rect 14568 21457 14596 22714
rect 14648 21888 14700 21894
rect 14740 21888 14792 21894
rect 14648 21830 14700 21836
rect 14738 21856 14740 21865
rect 14792 21856 14794 21865
rect 14660 21486 14688 21830
rect 14738 21791 14794 21800
rect 14648 21480 14700 21486
rect 14554 21448 14610 21457
rect 14648 21422 14700 21428
rect 14554 21383 14610 21392
rect 14568 21010 14596 21383
rect 14556 21004 14608 21010
rect 14556 20946 14608 20952
rect 14660 20233 14688 21422
rect 14740 21344 14792 21350
rect 14740 21286 14792 21292
rect 14752 20602 14780 21286
rect 14740 20596 14792 20602
rect 14740 20538 14792 20544
rect 14646 20224 14702 20233
rect 14646 20159 14702 20168
rect 14844 19378 14872 23462
rect 14832 19372 14884 19378
rect 14832 19314 14884 19320
rect 14740 16992 14792 16998
rect 14740 16934 14792 16940
rect 14464 15496 14516 15502
rect 14464 15438 14516 15444
rect 14648 15360 14700 15366
rect 14648 15302 14700 15308
rect 14464 13796 14516 13802
rect 14464 13738 14516 13744
rect 14188 13524 14240 13530
rect 14188 13466 14240 13472
rect 14096 13388 14148 13394
rect 14096 13330 14148 13336
rect 14004 12912 14056 12918
rect 14004 12854 14056 12860
rect 14016 11354 14044 12854
rect 14108 12782 14136 13330
rect 14476 12918 14504 13738
rect 14556 13456 14608 13462
rect 14556 13398 14608 13404
rect 14464 12912 14516 12918
rect 14384 12860 14464 12866
rect 14384 12854 14516 12860
rect 14384 12838 14504 12854
rect 14096 12776 14148 12782
rect 14096 12718 14148 12724
rect 14280 12640 14332 12646
rect 14280 12582 14332 12588
rect 14188 12164 14240 12170
rect 14188 12106 14240 12112
rect 14004 11348 14056 11354
rect 14004 11290 14056 11296
rect 13912 5568 13964 5574
rect 13912 5510 13964 5516
rect 13728 4208 13780 4214
rect 13728 4150 13780 4156
rect 13636 3732 13688 3738
rect 13636 3674 13688 3680
rect 13740 3534 13768 4150
rect 14004 3596 14056 3602
rect 14004 3538 14056 3544
rect 13728 3528 13780 3534
rect 13728 3470 13780 3476
rect 13636 2984 13688 2990
rect 13636 2926 13688 2932
rect 12950 2748 13258 2757
rect 12950 2746 12956 2748
rect 13012 2746 13036 2748
rect 13092 2746 13116 2748
rect 13172 2746 13196 2748
rect 13252 2746 13258 2748
rect 13012 2694 13014 2746
rect 13194 2694 13196 2746
rect 12950 2692 12956 2694
rect 13012 2692 13036 2694
rect 13092 2692 13116 2694
rect 13172 2692 13196 2694
rect 13252 2692 13258 2694
rect 12950 2683 13258 2692
rect 13268 2372 13320 2378
rect 13268 2314 13320 2320
rect 12820 2094 12940 2122
rect 12912 800 12940 2094
rect 13280 800 13308 2314
rect 13648 800 13676 2926
rect 14016 800 14044 3538
rect 14200 3058 14228 12106
rect 14292 3534 14320 12582
rect 14384 11898 14412 12838
rect 14464 12436 14516 12442
rect 14464 12378 14516 12384
rect 14372 11892 14424 11898
rect 14372 11834 14424 11840
rect 14476 11830 14504 12378
rect 14464 11824 14516 11830
rect 14464 11766 14516 11772
rect 14568 11218 14596 13398
rect 14556 11212 14608 11218
rect 14556 11154 14608 11160
rect 14660 4214 14688 15302
rect 14752 14278 14780 16934
rect 14936 16794 14964 26998
rect 15016 26580 15068 26586
rect 15016 26522 15068 26528
rect 15028 24954 15056 26522
rect 15108 25152 15160 25158
rect 15108 25094 15160 25100
rect 15016 24948 15068 24954
rect 15016 24890 15068 24896
rect 15120 20602 15148 25094
rect 15212 21690 15240 28970
rect 15304 23186 15332 36774
rect 15396 35873 15424 36790
rect 15382 35864 15438 35873
rect 15382 35799 15438 35808
rect 15384 35760 15436 35766
rect 15384 35702 15436 35708
rect 15396 31482 15424 35702
rect 15384 31476 15436 31482
rect 15384 31418 15436 31424
rect 15384 30184 15436 30190
rect 15384 30126 15436 30132
rect 15396 27130 15424 30126
rect 15488 27418 15516 37062
rect 15580 33590 15608 37878
rect 15672 37738 15700 40462
rect 15660 37732 15712 37738
rect 15660 37674 15712 37680
rect 15672 36378 15700 37674
rect 15660 36372 15712 36378
rect 15660 36314 15712 36320
rect 15672 35630 15700 36314
rect 15660 35624 15712 35630
rect 15660 35566 15712 35572
rect 15764 34626 15792 53382
rect 15856 53242 15884 54130
rect 16408 53582 16436 56200
rect 16672 54256 16724 54262
rect 16672 54198 16724 54204
rect 16488 53984 16540 53990
rect 16488 53926 16540 53932
rect 16396 53576 16448 53582
rect 16396 53518 16448 53524
rect 15936 53440 15988 53446
rect 15936 53382 15988 53388
rect 15844 53236 15896 53242
rect 15844 53178 15896 53184
rect 15948 52601 15976 53382
rect 16408 53242 16436 53518
rect 16396 53236 16448 53242
rect 16396 53178 16448 53184
rect 15934 52592 15990 52601
rect 15934 52527 15990 52536
rect 16120 47456 16172 47462
rect 16120 47398 16172 47404
rect 16132 46986 16160 47398
rect 16500 47122 16528 53926
rect 16684 53242 16712 54198
rect 16776 53582 16804 56200
rect 17144 54194 17172 56200
rect 17512 54262 17540 56200
rect 17500 54256 17552 54262
rect 17500 54198 17552 54204
rect 17132 54188 17184 54194
rect 17132 54130 17184 54136
rect 16948 53984 17000 53990
rect 16948 53926 17000 53932
rect 17776 53984 17828 53990
rect 17776 53926 17828 53932
rect 16764 53576 16816 53582
rect 16764 53518 16816 53524
rect 16776 53242 16804 53518
rect 16672 53236 16724 53242
rect 16672 53178 16724 53184
rect 16764 53236 16816 53242
rect 16764 53178 16816 53184
rect 16488 47116 16540 47122
rect 16488 47058 16540 47064
rect 16856 47048 16908 47054
rect 16856 46990 16908 46996
rect 16120 46980 16172 46986
rect 16120 46922 16172 46928
rect 16580 46980 16632 46986
rect 16580 46922 16632 46928
rect 16132 46714 16160 46922
rect 16120 46708 16172 46714
rect 16120 46650 16172 46656
rect 16028 46640 16080 46646
rect 16028 46582 16080 46588
rect 15844 46028 15896 46034
rect 15844 45970 15896 45976
rect 15856 45286 15884 45970
rect 15844 45280 15896 45286
rect 15844 45222 15896 45228
rect 15856 45082 15884 45222
rect 15844 45076 15896 45082
rect 15844 45018 15896 45024
rect 16040 44742 16068 46582
rect 16132 46034 16160 46650
rect 16592 46578 16620 46922
rect 16580 46572 16632 46578
rect 16580 46514 16632 46520
rect 16592 46170 16620 46514
rect 16868 46510 16896 46990
rect 16856 46504 16908 46510
rect 16856 46446 16908 46452
rect 16580 46164 16632 46170
rect 16580 46106 16632 46112
rect 16868 46034 16896 46446
rect 16120 46028 16172 46034
rect 16120 45970 16172 45976
rect 16856 46028 16908 46034
rect 16856 45970 16908 45976
rect 16856 45280 16908 45286
rect 16856 45222 16908 45228
rect 16028 44736 16080 44742
rect 16028 44678 16080 44684
rect 15936 44328 15988 44334
rect 15936 44270 15988 44276
rect 15844 43716 15896 43722
rect 15844 43658 15896 43664
rect 15856 42838 15884 43658
rect 15844 42832 15896 42838
rect 15844 42774 15896 42780
rect 15856 38418 15884 42774
rect 15948 39386 15976 44270
rect 16040 40594 16068 44678
rect 16672 43104 16724 43110
rect 16672 43046 16724 43052
rect 16304 42560 16356 42566
rect 16304 42502 16356 42508
rect 16316 42294 16344 42502
rect 16304 42288 16356 42294
rect 16304 42230 16356 42236
rect 16316 41834 16344 42230
rect 16224 41818 16344 41834
rect 16212 41812 16344 41818
rect 16264 41806 16344 41812
rect 16212 41754 16264 41760
rect 16212 41200 16264 41206
rect 16212 41142 16264 41148
rect 16028 40588 16080 40594
rect 16028 40530 16080 40536
rect 15948 39358 16068 39386
rect 15936 39296 15988 39302
rect 15936 39238 15988 39244
rect 15844 38412 15896 38418
rect 15844 38354 15896 38360
rect 15844 37324 15896 37330
rect 15844 37266 15896 37272
rect 15856 36718 15884 37266
rect 15844 36712 15896 36718
rect 15844 36654 15896 36660
rect 15948 35290 15976 39238
rect 16040 37126 16068 39358
rect 16120 38208 16172 38214
rect 16120 38150 16172 38156
rect 16132 38010 16160 38150
rect 16120 38004 16172 38010
rect 16120 37946 16172 37952
rect 16028 37120 16080 37126
rect 16028 37062 16080 37068
rect 16224 36938 16252 41142
rect 16684 40594 16712 43046
rect 16868 42838 16896 45222
rect 16856 42832 16908 42838
rect 16856 42774 16908 42780
rect 16764 42356 16816 42362
rect 16764 42298 16816 42304
rect 16672 40588 16724 40594
rect 16672 40530 16724 40536
rect 16396 40452 16448 40458
rect 16396 40394 16448 40400
rect 16408 40118 16436 40394
rect 16672 40384 16724 40390
rect 16672 40326 16724 40332
rect 16396 40112 16448 40118
rect 16396 40054 16448 40060
rect 16304 37120 16356 37126
rect 16304 37062 16356 37068
rect 16040 36910 16252 36938
rect 16040 36242 16068 36910
rect 16316 36854 16344 37062
rect 16304 36848 16356 36854
rect 16304 36790 16356 36796
rect 16304 36712 16356 36718
rect 16304 36654 16356 36660
rect 16028 36236 16080 36242
rect 16028 36178 16080 36184
rect 16316 36174 16344 36654
rect 16304 36168 16356 36174
rect 16304 36110 16356 36116
rect 15936 35284 15988 35290
rect 15936 35226 15988 35232
rect 16028 35284 16080 35290
rect 16028 35226 16080 35232
rect 16040 34746 16068 35226
rect 16028 34740 16080 34746
rect 16028 34682 16080 34688
rect 15764 34598 16344 34626
rect 15660 33924 15712 33930
rect 15660 33866 15712 33872
rect 15568 33584 15620 33590
rect 15568 33526 15620 33532
rect 15672 30326 15700 33866
rect 16028 33312 16080 33318
rect 16028 33254 16080 33260
rect 15752 32836 15804 32842
rect 15752 32778 15804 32784
rect 15660 30320 15712 30326
rect 15660 30262 15712 30268
rect 15764 30190 15792 32778
rect 15936 32360 15988 32366
rect 15936 32302 15988 32308
rect 15948 32026 15976 32302
rect 15936 32020 15988 32026
rect 15936 31962 15988 31968
rect 16040 31754 16068 33254
rect 16120 32836 16172 32842
rect 16120 32778 16172 32784
rect 15948 31726 16068 31754
rect 15844 30388 15896 30394
rect 15844 30330 15896 30336
rect 15752 30184 15804 30190
rect 15752 30126 15804 30132
rect 15856 30054 15884 30330
rect 15844 30048 15896 30054
rect 15844 29990 15896 29996
rect 15948 28082 15976 31726
rect 16132 30818 16160 32778
rect 16212 32768 16264 32774
rect 16212 32710 16264 32716
rect 16224 31754 16252 32710
rect 16212 31748 16264 31754
rect 16212 31690 16264 31696
rect 16040 30790 16160 30818
rect 16040 30598 16068 30790
rect 16120 30660 16172 30666
rect 16224 30648 16252 31690
rect 16172 30620 16252 30648
rect 16120 30602 16172 30608
rect 16028 30592 16080 30598
rect 16028 30534 16080 30540
rect 15936 28076 15988 28082
rect 15936 28018 15988 28024
rect 15936 27940 15988 27946
rect 15936 27882 15988 27888
rect 15948 27418 15976 27882
rect 16040 27538 16068 30534
rect 16132 30394 16160 30602
rect 16316 30598 16344 34598
rect 16304 30592 16356 30598
rect 16224 30540 16304 30546
rect 16224 30534 16356 30540
rect 16224 30518 16344 30534
rect 16120 30388 16172 30394
rect 16120 30330 16172 30336
rect 16224 30054 16252 30518
rect 16304 30388 16356 30394
rect 16304 30330 16356 30336
rect 16120 30048 16172 30054
rect 16118 30016 16120 30025
rect 16212 30048 16264 30054
rect 16172 30016 16174 30025
rect 16212 29990 16264 29996
rect 16118 29951 16174 29960
rect 16224 29238 16252 29990
rect 16212 29232 16264 29238
rect 16212 29174 16264 29180
rect 16316 28098 16344 30330
rect 16132 28070 16344 28098
rect 16028 27532 16080 27538
rect 16028 27474 16080 27480
rect 15488 27390 15884 27418
rect 15948 27390 16068 27418
rect 15476 27328 15528 27334
rect 15476 27270 15528 27276
rect 15568 27328 15620 27334
rect 15568 27270 15620 27276
rect 15384 27124 15436 27130
rect 15384 27066 15436 27072
rect 15488 26976 15516 27270
rect 15396 26948 15516 26976
rect 15292 23180 15344 23186
rect 15292 23122 15344 23128
rect 15396 22982 15424 26948
rect 15476 26852 15528 26858
rect 15476 26794 15528 26800
rect 15488 24188 15516 26794
rect 15580 25362 15608 27270
rect 15750 27160 15806 27169
rect 15750 27095 15752 27104
rect 15804 27095 15806 27104
rect 15752 27066 15804 27072
rect 15568 25356 15620 25362
rect 15568 25298 15620 25304
rect 15660 25356 15712 25362
rect 15660 25298 15712 25304
rect 15488 24160 15608 24188
rect 15384 22976 15436 22982
rect 15384 22918 15436 22924
rect 15200 21684 15252 21690
rect 15200 21626 15252 21632
rect 15108 20596 15160 20602
rect 15108 20538 15160 20544
rect 15396 19334 15424 22918
rect 15580 21729 15608 24160
rect 15672 22778 15700 25298
rect 15752 23520 15804 23526
rect 15752 23462 15804 23468
rect 15660 22772 15712 22778
rect 15660 22714 15712 22720
rect 15566 21720 15622 21729
rect 15566 21655 15622 21664
rect 15474 21584 15530 21593
rect 15474 21519 15476 21528
rect 15528 21519 15530 21528
rect 15476 21490 15528 21496
rect 15304 19306 15424 19334
rect 15304 17882 15332 19306
rect 15292 17876 15344 17882
rect 15292 17818 15344 17824
rect 15476 17740 15528 17746
rect 15476 17682 15528 17688
rect 14924 16788 14976 16794
rect 14924 16730 14976 16736
rect 15384 16788 15436 16794
rect 15384 16730 15436 16736
rect 15200 16448 15252 16454
rect 15200 16390 15252 16396
rect 14832 15904 14884 15910
rect 14832 15846 14884 15852
rect 14844 15162 14872 15846
rect 14832 15156 14884 15162
rect 14832 15098 14884 15104
rect 14924 15020 14976 15026
rect 14924 14962 14976 14968
rect 15108 15020 15160 15026
rect 15108 14962 15160 14968
rect 14740 14272 14792 14278
rect 14740 14214 14792 14220
rect 14740 13524 14792 13530
rect 14740 13466 14792 13472
rect 14752 12102 14780 13466
rect 14740 12096 14792 12102
rect 14740 12038 14792 12044
rect 14648 4208 14700 4214
rect 14648 4150 14700 4156
rect 14280 3528 14332 3534
rect 14280 3470 14332 3476
rect 14752 3466 14780 12038
rect 14936 11898 14964 14962
rect 15120 14550 15148 14962
rect 15108 14544 15160 14550
rect 15108 14486 15160 14492
rect 15108 14340 15160 14346
rect 15108 14282 15160 14288
rect 15016 13184 15068 13190
rect 15016 13126 15068 13132
rect 14924 11892 14976 11898
rect 14924 11834 14976 11840
rect 15028 3534 15056 13126
rect 15120 12306 15148 14282
rect 15108 12300 15160 12306
rect 15108 12242 15160 12248
rect 15120 11218 15148 12242
rect 15212 12238 15240 16390
rect 15292 16040 15344 16046
rect 15292 15982 15344 15988
rect 15304 15162 15332 15982
rect 15292 15156 15344 15162
rect 15292 15098 15344 15104
rect 15396 12238 15424 16730
rect 15488 16726 15516 17682
rect 15476 16720 15528 16726
rect 15476 16662 15528 16668
rect 15488 16046 15516 16662
rect 15476 16040 15528 16046
rect 15476 15982 15528 15988
rect 15200 12232 15252 12238
rect 15200 12174 15252 12180
rect 15384 12232 15436 12238
rect 15384 12174 15436 12180
rect 15212 11778 15240 12174
rect 15384 11892 15436 11898
rect 15384 11834 15436 11840
rect 15212 11750 15332 11778
rect 15108 11212 15160 11218
rect 15108 11154 15160 11160
rect 15200 9444 15252 9450
rect 15200 9386 15252 9392
rect 15212 4146 15240 9386
rect 15304 6798 15332 11750
rect 15396 11694 15424 11834
rect 15488 11694 15516 15982
rect 15580 13530 15608 21655
rect 15660 20256 15712 20262
rect 15660 20198 15712 20204
rect 15672 18834 15700 20198
rect 15660 18828 15712 18834
rect 15660 18770 15712 18776
rect 15672 13954 15700 18770
rect 15764 16590 15792 23462
rect 15856 22216 15884 27390
rect 15936 27328 15988 27334
rect 15936 27270 15988 27276
rect 15948 26994 15976 27270
rect 15936 26988 15988 26994
rect 15936 26930 15988 26936
rect 16040 26586 16068 27390
rect 15936 26580 15988 26586
rect 15936 26522 15988 26528
rect 16028 26580 16080 26586
rect 16028 26522 16080 26528
rect 15948 26382 15976 26522
rect 15936 26376 15988 26382
rect 16132 26330 16160 28070
rect 16304 27124 16356 27130
rect 16304 27066 16356 27072
rect 16316 26790 16344 27066
rect 16408 26994 16436 40054
rect 16580 39296 16632 39302
rect 16580 39238 16632 39244
rect 16592 38554 16620 39238
rect 16580 38548 16632 38554
rect 16580 38490 16632 38496
rect 16488 38208 16540 38214
rect 16488 38150 16540 38156
rect 16500 36922 16528 38150
rect 16488 36916 16540 36922
rect 16488 36858 16540 36864
rect 16580 36032 16632 36038
rect 16580 35974 16632 35980
rect 16488 30864 16540 30870
rect 16488 30806 16540 30812
rect 16500 30394 16528 30806
rect 16488 30388 16540 30394
rect 16488 30330 16540 30336
rect 16592 30258 16620 35974
rect 16684 33046 16712 40326
rect 16776 38554 16804 42298
rect 16856 40928 16908 40934
rect 16856 40870 16908 40876
rect 16868 39098 16896 40870
rect 16960 40118 16988 53926
rect 17040 53440 17092 53446
rect 17040 53382 17092 53388
rect 17408 53440 17460 53446
rect 17408 53382 17460 53388
rect 17052 44538 17080 53382
rect 17316 46912 17368 46918
rect 17316 46854 17368 46860
rect 17132 46368 17184 46374
rect 17132 46310 17184 46316
rect 17040 44532 17092 44538
rect 17040 44474 17092 44480
rect 17144 43450 17172 46310
rect 17224 45484 17276 45490
rect 17224 45426 17276 45432
rect 17236 44742 17264 45426
rect 17224 44736 17276 44742
rect 17224 44678 17276 44684
rect 17132 43444 17184 43450
rect 17132 43386 17184 43392
rect 17328 41274 17356 46854
rect 17420 46714 17448 53382
rect 17788 47122 17816 53926
rect 17880 53582 17908 56200
rect 18248 54618 18276 56200
rect 18248 54590 18368 54618
rect 17950 54428 18258 54437
rect 17950 54426 17956 54428
rect 18012 54426 18036 54428
rect 18092 54426 18116 54428
rect 18172 54426 18196 54428
rect 18252 54426 18258 54428
rect 18012 54374 18014 54426
rect 18194 54374 18196 54426
rect 17950 54372 17956 54374
rect 18012 54372 18036 54374
rect 18092 54372 18116 54374
rect 18172 54372 18196 54374
rect 18252 54372 18258 54374
rect 17950 54363 18258 54372
rect 18340 53582 18368 54590
rect 18420 54256 18472 54262
rect 18420 54198 18472 54204
rect 17868 53576 17920 53582
rect 17868 53518 17920 53524
rect 18328 53576 18380 53582
rect 18328 53518 18380 53524
rect 17880 53242 17908 53518
rect 17950 53340 18258 53349
rect 17950 53338 17956 53340
rect 18012 53338 18036 53340
rect 18092 53338 18116 53340
rect 18172 53338 18196 53340
rect 18252 53338 18258 53340
rect 18012 53286 18014 53338
rect 18194 53286 18196 53338
rect 17950 53284 17956 53286
rect 18012 53284 18036 53286
rect 18092 53284 18116 53286
rect 18172 53284 18196 53286
rect 18252 53284 18258 53286
rect 17950 53275 18258 53284
rect 18340 53242 18368 53518
rect 17868 53236 17920 53242
rect 17868 53178 17920 53184
rect 18328 53236 18380 53242
rect 18328 53178 18380 53184
rect 18432 53174 18460 54198
rect 18616 54194 18644 56200
rect 18604 54188 18656 54194
rect 18604 54130 18656 54136
rect 18604 54052 18656 54058
rect 18604 53994 18656 54000
rect 18512 53440 18564 53446
rect 18512 53382 18564 53388
rect 18420 53168 18472 53174
rect 18420 53110 18472 53116
rect 17950 52252 18258 52261
rect 17950 52250 17956 52252
rect 18012 52250 18036 52252
rect 18092 52250 18116 52252
rect 18172 52250 18196 52252
rect 18252 52250 18258 52252
rect 18012 52198 18014 52250
rect 18194 52198 18196 52250
rect 17950 52196 17956 52198
rect 18012 52196 18036 52198
rect 18092 52196 18116 52198
rect 18172 52196 18196 52198
rect 18252 52196 18258 52198
rect 17950 52187 18258 52196
rect 17950 51164 18258 51173
rect 17950 51162 17956 51164
rect 18012 51162 18036 51164
rect 18092 51162 18116 51164
rect 18172 51162 18196 51164
rect 18252 51162 18258 51164
rect 18012 51110 18014 51162
rect 18194 51110 18196 51162
rect 17950 51108 17956 51110
rect 18012 51108 18036 51110
rect 18092 51108 18116 51110
rect 18172 51108 18196 51110
rect 18252 51108 18258 51110
rect 17950 51099 18258 51108
rect 17950 50076 18258 50085
rect 17950 50074 17956 50076
rect 18012 50074 18036 50076
rect 18092 50074 18116 50076
rect 18172 50074 18196 50076
rect 18252 50074 18258 50076
rect 18012 50022 18014 50074
rect 18194 50022 18196 50074
rect 17950 50020 17956 50022
rect 18012 50020 18036 50022
rect 18092 50020 18116 50022
rect 18172 50020 18196 50022
rect 18252 50020 18258 50022
rect 17950 50011 18258 50020
rect 17950 48988 18258 48997
rect 17950 48986 17956 48988
rect 18012 48986 18036 48988
rect 18092 48986 18116 48988
rect 18172 48986 18196 48988
rect 18252 48986 18258 48988
rect 18012 48934 18014 48986
rect 18194 48934 18196 48986
rect 17950 48932 17956 48934
rect 18012 48932 18036 48934
rect 18092 48932 18116 48934
rect 18172 48932 18196 48934
rect 18252 48932 18258 48934
rect 17950 48923 18258 48932
rect 17950 47900 18258 47909
rect 17950 47898 17956 47900
rect 18012 47898 18036 47900
rect 18092 47898 18116 47900
rect 18172 47898 18196 47900
rect 18252 47898 18258 47900
rect 18012 47846 18014 47898
rect 18194 47846 18196 47898
rect 17950 47844 17956 47846
rect 18012 47844 18036 47846
rect 18092 47844 18116 47846
rect 18172 47844 18196 47846
rect 18252 47844 18258 47846
rect 17950 47835 18258 47844
rect 17776 47116 17828 47122
rect 17776 47058 17828 47064
rect 17950 46812 18258 46821
rect 17950 46810 17956 46812
rect 18012 46810 18036 46812
rect 18092 46810 18116 46812
rect 18172 46810 18196 46812
rect 18252 46810 18258 46812
rect 18012 46758 18014 46810
rect 18194 46758 18196 46810
rect 17950 46756 17956 46758
rect 18012 46756 18036 46758
rect 18092 46756 18116 46758
rect 18172 46756 18196 46758
rect 18252 46756 18258 46758
rect 17950 46747 18258 46756
rect 17408 46708 17460 46714
rect 17408 46650 17460 46656
rect 18524 46578 18552 53382
rect 18616 46646 18644 53994
rect 18984 53582 19012 56200
rect 19352 54330 19380 56200
rect 19340 54324 19392 54330
rect 19340 54266 19392 54272
rect 19340 54188 19392 54194
rect 19340 54130 19392 54136
rect 18972 53576 19024 53582
rect 18972 53518 19024 53524
rect 18696 53440 18748 53446
rect 18696 53382 18748 53388
rect 18708 46714 18736 53382
rect 19352 53242 19380 54130
rect 19616 53984 19668 53990
rect 19616 53926 19668 53932
rect 19524 53440 19576 53446
rect 19524 53382 19576 53388
rect 19340 53236 19392 53242
rect 19340 53178 19392 53184
rect 18972 47048 19024 47054
rect 18972 46990 19024 46996
rect 18696 46708 18748 46714
rect 18696 46650 18748 46656
rect 18604 46640 18656 46646
rect 18656 46588 18736 46594
rect 18604 46582 18736 46588
rect 17776 46572 17828 46578
rect 17776 46514 17828 46520
rect 18512 46572 18564 46578
rect 18616 46566 18736 46582
rect 18512 46514 18564 46520
rect 17592 45892 17644 45898
rect 17592 45834 17644 45840
rect 17500 44736 17552 44742
rect 17500 44678 17552 44684
rect 17512 43722 17540 44678
rect 17500 43716 17552 43722
rect 17500 43658 17552 43664
rect 17408 42900 17460 42906
rect 17408 42842 17460 42848
rect 17316 41268 17368 41274
rect 17316 41210 17368 41216
rect 17224 41132 17276 41138
rect 17224 41074 17276 41080
rect 17236 40934 17264 41074
rect 17420 41070 17448 42842
rect 17512 41818 17540 43658
rect 17604 43654 17632 45834
rect 17592 43648 17644 43654
rect 17592 43590 17644 43596
rect 17500 41812 17552 41818
rect 17500 41754 17552 41760
rect 17408 41064 17460 41070
rect 17408 41006 17460 41012
rect 17224 40928 17276 40934
rect 17224 40870 17276 40876
rect 16948 40112 17000 40118
rect 16948 40054 17000 40060
rect 16948 39976 17000 39982
rect 16948 39918 17000 39924
rect 16856 39092 16908 39098
rect 16856 39034 16908 39040
rect 16764 38548 16816 38554
rect 16764 38490 16816 38496
rect 16764 36780 16816 36786
rect 16764 36722 16816 36728
rect 16776 34542 16804 36722
rect 16856 36576 16908 36582
rect 16856 36518 16908 36524
rect 16868 35834 16896 36518
rect 16856 35828 16908 35834
rect 16856 35770 16908 35776
rect 16960 35086 16988 39918
rect 17130 36952 17186 36961
rect 17130 36887 17186 36896
rect 17144 36310 17172 36887
rect 17236 36310 17264 40870
rect 17500 40724 17552 40730
rect 17500 40666 17552 40672
rect 17316 38820 17368 38826
rect 17316 38762 17368 38768
rect 17328 37806 17356 38762
rect 17408 38752 17460 38758
rect 17408 38694 17460 38700
rect 17316 37800 17368 37806
rect 17316 37742 17368 37748
rect 17328 36854 17356 37742
rect 17316 36848 17368 36854
rect 17316 36790 17368 36796
rect 17132 36304 17184 36310
rect 17132 36246 17184 36252
rect 17224 36304 17276 36310
rect 17224 36246 17276 36252
rect 17236 36020 17264 36246
rect 17144 35992 17264 36020
rect 16948 35080 17000 35086
rect 16948 35022 17000 35028
rect 16856 34740 16908 34746
rect 16856 34682 16908 34688
rect 16764 34536 16816 34542
rect 16764 34478 16816 34484
rect 16672 33040 16724 33046
rect 16672 32982 16724 32988
rect 16868 32978 16896 34682
rect 16948 33108 17000 33114
rect 16948 33050 17000 33056
rect 16856 32972 16908 32978
rect 16856 32914 16908 32920
rect 16868 32434 16896 32914
rect 16856 32428 16908 32434
rect 16856 32370 16908 32376
rect 16868 31872 16896 32370
rect 16960 32298 16988 33050
rect 17040 32496 17092 32502
rect 17040 32438 17092 32444
rect 16948 32292 17000 32298
rect 16948 32234 17000 32240
rect 17052 31929 17080 32438
rect 17038 31920 17094 31929
rect 16948 31884 17000 31890
rect 16868 31844 16948 31872
rect 17038 31855 17040 31864
rect 16948 31826 17000 31832
rect 17092 31855 17094 31864
rect 17040 31826 17092 31832
rect 16672 31748 16724 31754
rect 16672 31690 16724 31696
rect 16580 30252 16632 30258
rect 16580 30194 16632 30200
rect 16488 29776 16540 29782
rect 16488 29718 16540 29724
rect 16500 27946 16528 29718
rect 16684 28762 16712 31690
rect 16856 31476 16908 31482
rect 16856 31418 16908 31424
rect 16868 30190 16896 31418
rect 16948 30796 17000 30802
rect 16948 30738 17000 30744
rect 16856 30184 16908 30190
rect 16856 30126 16908 30132
rect 16764 29164 16816 29170
rect 16764 29106 16816 29112
rect 16776 29073 16804 29106
rect 16762 29064 16818 29073
rect 16762 28999 16764 29008
rect 16816 28999 16818 29008
rect 16764 28970 16816 28976
rect 16672 28756 16724 28762
rect 16672 28698 16724 28704
rect 16580 28552 16632 28558
rect 16580 28494 16632 28500
rect 16592 28218 16620 28494
rect 16580 28212 16632 28218
rect 16580 28154 16632 28160
rect 16488 27940 16540 27946
rect 16488 27882 16540 27888
rect 16500 27656 16528 27882
rect 16500 27628 16620 27656
rect 16488 27328 16540 27334
rect 16488 27270 16540 27276
rect 16396 26988 16448 26994
rect 16396 26930 16448 26936
rect 16500 26790 16528 27270
rect 16304 26784 16356 26790
rect 16488 26784 16540 26790
rect 16356 26732 16436 26738
rect 16304 26726 16436 26732
rect 16488 26726 16540 26732
rect 16316 26710 16436 26726
rect 16212 26580 16264 26586
rect 16212 26522 16264 26528
rect 15936 26318 15988 26324
rect 16040 26302 16160 26330
rect 15936 24064 15988 24070
rect 15936 24006 15988 24012
rect 15948 23866 15976 24006
rect 15936 23860 15988 23866
rect 15936 23802 15988 23808
rect 16040 23662 16068 26302
rect 16120 25696 16172 25702
rect 16118 25664 16120 25673
rect 16172 25664 16174 25673
rect 16118 25599 16174 25608
rect 16132 25498 16160 25599
rect 16120 25492 16172 25498
rect 16120 25434 16172 25440
rect 16132 25226 16160 25434
rect 16120 25220 16172 25226
rect 16120 25162 16172 25168
rect 16120 24812 16172 24818
rect 16120 24754 16172 24760
rect 16028 23656 16080 23662
rect 16028 23598 16080 23604
rect 15936 22228 15988 22234
rect 15856 22188 15936 22216
rect 15752 16584 15804 16590
rect 15752 16526 15804 16532
rect 15856 14940 15884 22188
rect 15936 22170 15988 22176
rect 16040 22094 16068 23598
rect 16132 22710 16160 24754
rect 16224 24750 16252 26522
rect 16304 26240 16356 26246
rect 16304 26182 16356 26188
rect 16316 25702 16344 26182
rect 16304 25696 16356 25702
rect 16304 25638 16356 25644
rect 16304 25152 16356 25158
rect 16304 25094 16356 25100
rect 16212 24744 16264 24750
rect 16212 24686 16264 24692
rect 16224 24206 16252 24686
rect 16316 24274 16344 25094
rect 16304 24268 16356 24274
rect 16304 24210 16356 24216
rect 16212 24200 16264 24206
rect 16212 24142 16264 24148
rect 16120 22704 16172 22710
rect 16120 22646 16172 22652
rect 15948 22066 16068 22094
rect 15948 15094 15976 22066
rect 16028 21956 16080 21962
rect 16132 21944 16160 22646
rect 16408 22094 16436 26710
rect 16500 26586 16528 26726
rect 16488 26580 16540 26586
rect 16488 26522 16540 26528
rect 16500 23508 16528 26522
rect 16592 25362 16620 27628
rect 16684 27606 16712 28698
rect 16764 28144 16816 28150
rect 16764 28086 16816 28092
rect 16672 27600 16724 27606
rect 16672 27542 16724 27548
rect 16776 27418 16804 28086
rect 16776 27390 16896 27418
rect 16764 27328 16816 27334
rect 16764 27270 16816 27276
rect 16672 26376 16724 26382
rect 16672 26318 16724 26324
rect 16684 25974 16712 26318
rect 16672 25968 16724 25974
rect 16672 25910 16724 25916
rect 16684 25498 16712 25910
rect 16672 25492 16724 25498
rect 16672 25434 16724 25440
rect 16580 25356 16632 25362
rect 16580 25298 16632 25304
rect 16684 24818 16712 25434
rect 16672 24812 16724 24818
rect 16672 24754 16724 24760
rect 16580 24744 16632 24750
rect 16580 24686 16632 24692
rect 16592 23662 16620 24686
rect 16672 24608 16724 24614
rect 16672 24550 16724 24556
rect 16580 23656 16632 23662
rect 16580 23598 16632 23604
rect 16500 23480 16620 23508
rect 16316 22066 16436 22094
rect 16212 21956 16264 21962
rect 16132 21916 16212 21944
rect 16028 21898 16080 21904
rect 16212 21898 16264 21904
rect 16040 20806 16068 21898
rect 16224 21350 16252 21898
rect 16212 21344 16264 21350
rect 16212 21286 16264 21292
rect 16224 21146 16252 21286
rect 16212 21140 16264 21146
rect 16212 21082 16264 21088
rect 16224 20874 16252 21082
rect 16212 20868 16264 20874
rect 16212 20810 16264 20816
rect 16028 20800 16080 20806
rect 16028 20742 16080 20748
rect 16040 20398 16068 20742
rect 16028 20392 16080 20398
rect 16028 20334 16080 20340
rect 16210 17640 16266 17649
rect 16210 17575 16266 17584
rect 16120 17060 16172 17066
rect 16120 17002 16172 17008
rect 16028 15972 16080 15978
rect 16028 15914 16080 15920
rect 16040 15337 16068 15914
rect 16132 15434 16160 17002
rect 16224 16794 16252 17575
rect 16212 16788 16264 16794
rect 16212 16730 16264 16736
rect 16224 16182 16252 16730
rect 16212 16176 16264 16182
rect 16212 16118 16264 16124
rect 16120 15428 16172 15434
rect 16120 15370 16172 15376
rect 16026 15328 16082 15337
rect 16026 15263 16082 15272
rect 15936 15088 15988 15094
rect 15936 15030 15988 15036
rect 15856 14912 16068 14940
rect 15936 14816 15988 14822
rect 15936 14758 15988 14764
rect 15672 13926 15884 13954
rect 15752 13864 15804 13870
rect 15752 13806 15804 13812
rect 15568 13524 15620 13530
rect 15568 13466 15620 13472
rect 15660 12776 15712 12782
rect 15660 12718 15712 12724
rect 15568 12436 15620 12442
rect 15672 12434 15700 12718
rect 15620 12406 15700 12434
rect 15568 12378 15620 12384
rect 15660 12096 15712 12102
rect 15660 12038 15712 12044
rect 15384 11688 15436 11694
rect 15384 11630 15436 11636
rect 15476 11688 15528 11694
rect 15476 11630 15528 11636
rect 15568 11688 15620 11694
rect 15568 11630 15620 11636
rect 15292 6792 15344 6798
rect 15292 6734 15344 6740
rect 15200 4140 15252 4146
rect 15200 4082 15252 4088
rect 15016 3528 15068 3534
rect 15016 3470 15068 3476
rect 14740 3460 14792 3466
rect 14740 3402 14792 3408
rect 14188 3052 14240 3058
rect 14188 2994 14240 3000
rect 14740 2984 14792 2990
rect 14740 2926 14792 2932
rect 14372 2372 14424 2378
rect 14372 2314 14424 2320
rect 14384 800 14412 2314
rect 14752 800 14780 2926
rect 15396 2650 15424 11630
rect 15580 11150 15608 11630
rect 15568 11144 15620 11150
rect 15568 11086 15620 11092
rect 15672 4706 15700 12038
rect 15764 5370 15792 13806
rect 15856 12434 15884 13926
rect 15948 13870 15976 14758
rect 16040 14006 16068 14912
rect 16132 14618 16160 15370
rect 16212 15156 16264 15162
rect 16212 15098 16264 15104
rect 16120 14612 16172 14618
rect 16120 14554 16172 14560
rect 16028 14000 16080 14006
rect 16028 13942 16080 13948
rect 15936 13864 15988 13870
rect 15936 13806 15988 13812
rect 16028 13728 16080 13734
rect 16028 13670 16080 13676
rect 15856 12406 15976 12434
rect 15844 11620 15896 11626
rect 15844 11562 15896 11568
rect 15856 11150 15884 11562
rect 15844 11144 15896 11150
rect 15844 11086 15896 11092
rect 15844 10804 15896 10810
rect 15844 10746 15896 10752
rect 15856 5778 15884 10746
rect 15948 8974 15976 12406
rect 16040 11014 16068 13670
rect 16028 11008 16080 11014
rect 16028 10950 16080 10956
rect 16040 10470 16068 10950
rect 16224 10810 16252 15098
rect 16316 15008 16344 22066
rect 16394 20632 16450 20641
rect 16394 20567 16396 20576
rect 16448 20567 16450 20576
rect 16396 20538 16448 20544
rect 16488 17604 16540 17610
rect 16488 17546 16540 17552
rect 16500 15994 16528 17546
rect 16592 16674 16620 23480
rect 16684 17338 16712 24550
rect 16776 20466 16804 27270
rect 16868 23866 16896 27390
rect 16960 26296 16988 30738
rect 17144 28558 17172 35992
rect 17328 35154 17356 36790
rect 17316 35148 17368 35154
rect 17316 35090 17368 35096
rect 17316 32292 17368 32298
rect 17316 32234 17368 32240
rect 17224 31136 17276 31142
rect 17224 31078 17276 31084
rect 17132 28552 17184 28558
rect 17132 28494 17184 28500
rect 17040 28416 17092 28422
rect 17040 28358 17092 28364
rect 17052 27470 17080 28358
rect 17040 27464 17092 27470
rect 17040 27406 17092 27412
rect 17236 27334 17264 31078
rect 17328 30802 17356 32234
rect 17420 31414 17448 38694
rect 17512 38282 17540 40666
rect 17604 39506 17632 43590
rect 17684 42560 17736 42566
rect 17684 42502 17736 42508
rect 17696 39506 17724 42502
rect 17592 39500 17644 39506
rect 17592 39442 17644 39448
rect 17684 39500 17736 39506
rect 17684 39442 17736 39448
rect 17788 39386 17816 46514
rect 18604 46504 18656 46510
rect 18604 46446 18656 46452
rect 18328 46368 18380 46374
rect 18328 46310 18380 46316
rect 17950 45724 18258 45733
rect 17950 45722 17956 45724
rect 18012 45722 18036 45724
rect 18092 45722 18116 45724
rect 18172 45722 18196 45724
rect 18252 45722 18258 45724
rect 18012 45670 18014 45722
rect 18194 45670 18196 45722
rect 17950 45668 17956 45670
rect 18012 45668 18036 45670
rect 18092 45668 18116 45670
rect 18172 45668 18196 45670
rect 18252 45668 18258 45670
rect 17950 45659 18258 45668
rect 17950 44636 18258 44645
rect 17950 44634 17956 44636
rect 18012 44634 18036 44636
rect 18092 44634 18116 44636
rect 18172 44634 18196 44636
rect 18252 44634 18258 44636
rect 18012 44582 18014 44634
rect 18194 44582 18196 44634
rect 17950 44580 17956 44582
rect 18012 44580 18036 44582
rect 18092 44580 18116 44582
rect 18172 44580 18196 44582
rect 18252 44580 18258 44582
rect 17950 44571 18258 44580
rect 18052 44396 18104 44402
rect 18052 44338 18104 44344
rect 18064 43722 18092 44338
rect 18052 43716 18104 43722
rect 18052 43658 18104 43664
rect 17950 43548 18258 43557
rect 17950 43546 17956 43548
rect 18012 43546 18036 43548
rect 18092 43546 18116 43548
rect 18172 43546 18196 43548
rect 18252 43546 18258 43548
rect 18012 43494 18014 43546
rect 18194 43494 18196 43546
rect 17950 43492 17956 43494
rect 18012 43492 18036 43494
rect 18092 43492 18116 43494
rect 18172 43492 18196 43494
rect 18252 43492 18258 43494
rect 17950 43483 18258 43492
rect 18340 42702 18368 46310
rect 18420 46164 18472 46170
rect 18420 46106 18472 46112
rect 18328 42696 18380 42702
rect 18328 42638 18380 42644
rect 17868 42560 17920 42566
rect 17868 42502 17920 42508
rect 17880 40662 17908 42502
rect 17950 42460 18258 42469
rect 17950 42458 17956 42460
rect 18012 42458 18036 42460
rect 18092 42458 18116 42460
rect 18172 42458 18196 42460
rect 18252 42458 18258 42460
rect 18012 42406 18014 42458
rect 18194 42406 18196 42458
rect 17950 42404 17956 42406
rect 18012 42404 18036 42406
rect 18092 42404 18116 42406
rect 18172 42404 18196 42406
rect 18252 42404 18258 42406
rect 17950 42395 18258 42404
rect 18432 42378 18460 46106
rect 18616 46050 18644 46446
rect 18708 46170 18736 46566
rect 18696 46164 18748 46170
rect 18696 46106 18748 46112
rect 18524 46022 18644 46050
rect 18524 45286 18552 46022
rect 18604 45892 18656 45898
rect 18604 45834 18656 45840
rect 18616 45286 18644 45834
rect 18512 45280 18564 45286
rect 18512 45222 18564 45228
rect 18604 45280 18656 45286
rect 18604 45222 18656 45228
rect 18524 44538 18552 45222
rect 18512 44532 18564 44538
rect 18512 44474 18564 44480
rect 18604 43852 18656 43858
rect 18604 43794 18656 43800
rect 18432 42350 18552 42378
rect 18420 42288 18472 42294
rect 18420 42230 18472 42236
rect 18432 41682 18460 42230
rect 18420 41676 18472 41682
rect 18420 41618 18472 41624
rect 17950 41372 18258 41381
rect 17950 41370 17956 41372
rect 18012 41370 18036 41372
rect 18092 41370 18116 41372
rect 18172 41370 18196 41372
rect 18252 41370 18258 41372
rect 18012 41318 18014 41370
rect 18194 41318 18196 41370
rect 17950 41316 17956 41318
rect 18012 41316 18036 41318
rect 18092 41316 18116 41318
rect 18172 41316 18196 41318
rect 18252 41316 18258 41318
rect 17950 41307 18258 41316
rect 18432 41138 18460 41618
rect 18420 41132 18472 41138
rect 18420 41074 18472 41080
rect 17868 40656 17920 40662
rect 17868 40598 17920 40604
rect 17696 39358 17816 39386
rect 17592 39092 17644 39098
rect 17592 39034 17644 39040
rect 17500 38276 17552 38282
rect 17500 38218 17552 38224
rect 17512 37194 17540 38218
rect 17500 37188 17552 37194
rect 17500 37130 17552 37136
rect 17604 37074 17632 39034
rect 17512 37046 17632 37074
rect 17408 31408 17460 31414
rect 17408 31350 17460 31356
rect 17408 30932 17460 30938
rect 17408 30874 17460 30880
rect 17316 30796 17368 30802
rect 17316 30738 17368 30744
rect 17316 30592 17368 30598
rect 17316 30534 17368 30540
rect 17328 28218 17356 30534
rect 17420 29034 17448 30874
rect 17512 29102 17540 37046
rect 17590 36272 17646 36281
rect 17590 36207 17646 36216
rect 17604 36174 17632 36207
rect 17592 36168 17644 36174
rect 17592 36110 17644 36116
rect 17696 33114 17724 39358
rect 17880 39098 17908 40598
rect 18328 40384 18380 40390
rect 18328 40326 18380 40332
rect 17950 40284 18258 40293
rect 17950 40282 17956 40284
rect 18012 40282 18036 40284
rect 18092 40282 18116 40284
rect 18172 40282 18196 40284
rect 18252 40282 18258 40284
rect 18012 40230 18014 40282
rect 18194 40230 18196 40282
rect 17950 40228 17956 40230
rect 18012 40228 18036 40230
rect 18092 40228 18116 40230
rect 18172 40228 18196 40230
rect 18252 40228 18258 40230
rect 17950 40219 18258 40228
rect 17950 39196 18258 39205
rect 17950 39194 17956 39196
rect 18012 39194 18036 39196
rect 18092 39194 18116 39196
rect 18172 39194 18196 39196
rect 18252 39194 18258 39196
rect 18012 39142 18014 39194
rect 18194 39142 18196 39194
rect 17950 39140 17956 39142
rect 18012 39140 18036 39142
rect 18092 39140 18116 39142
rect 18172 39140 18196 39142
rect 18252 39140 18258 39142
rect 17950 39131 18258 39140
rect 17868 39092 17920 39098
rect 17868 39034 17920 39040
rect 17950 38108 18258 38117
rect 17950 38106 17956 38108
rect 18012 38106 18036 38108
rect 18092 38106 18116 38108
rect 18172 38106 18196 38108
rect 18252 38106 18258 38108
rect 18012 38054 18014 38106
rect 18194 38054 18196 38106
rect 17950 38052 17956 38054
rect 18012 38052 18036 38054
rect 18092 38052 18116 38054
rect 18172 38052 18196 38054
rect 18252 38052 18258 38054
rect 17950 38043 18258 38052
rect 18052 37800 18104 37806
rect 18052 37742 18104 37748
rect 18064 37398 18092 37742
rect 18052 37392 18104 37398
rect 17774 37360 17830 37369
rect 18052 37334 18104 37340
rect 17830 37304 18000 37312
rect 17774 37295 17776 37304
rect 17828 37284 18000 37304
rect 17776 37266 17828 37272
rect 17972 37194 18000 37284
rect 17960 37188 18012 37194
rect 17960 37130 18012 37136
rect 17950 37020 18258 37029
rect 17950 37018 17956 37020
rect 18012 37018 18036 37020
rect 18092 37018 18116 37020
rect 18172 37018 18196 37020
rect 18252 37018 18258 37020
rect 18012 36966 18014 37018
rect 18194 36966 18196 37018
rect 17950 36964 17956 36966
rect 18012 36964 18036 36966
rect 18092 36964 18116 36966
rect 18172 36964 18196 36966
rect 18252 36964 18258 36966
rect 17950 36955 18258 36964
rect 18340 36922 18368 40326
rect 18420 39568 18472 39574
rect 18420 39510 18472 39516
rect 18432 38729 18460 39510
rect 18418 38720 18474 38729
rect 18418 38655 18474 38664
rect 18420 37664 18472 37670
rect 18420 37606 18472 37612
rect 18432 37330 18460 37606
rect 18420 37324 18472 37330
rect 18420 37266 18472 37272
rect 18236 36916 18288 36922
rect 18236 36858 18288 36864
rect 18328 36916 18380 36922
rect 18328 36858 18380 36864
rect 18248 36768 18276 36858
rect 18248 36740 18368 36768
rect 17950 35932 18258 35941
rect 17950 35930 17956 35932
rect 18012 35930 18036 35932
rect 18092 35930 18116 35932
rect 18172 35930 18196 35932
rect 18252 35930 18258 35932
rect 18012 35878 18014 35930
rect 18194 35878 18196 35930
rect 17950 35876 17956 35878
rect 18012 35876 18036 35878
rect 18092 35876 18116 35878
rect 18172 35876 18196 35878
rect 18252 35876 18258 35878
rect 17950 35867 18258 35876
rect 17950 34844 18258 34853
rect 17950 34842 17956 34844
rect 18012 34842 18036 34844
rect 18092 34842 18116 34844
rect 18172 34842 18196 34844
rect 18252 34842 18258 34844
rect 18012 34790 18014 34842
rect 18194 34790 18196 34842
rect 17950 34788 17956 34790
rect 18012 34788 18036 34790
rect 18092 34788 18116 34790
rect 18172 34788 18196 34790
rect 18252 34788 18258 34790
rect 17950 34779 18258 34788
rect 18236 34672 18288 34678
rect 18236 34614 18288 34620
rect 18248 33862 18276 34614
rect 18236 33856 18288 33862
rect 18236 33798 18288 33804
rect 17950 33756 18258 33765
rect 17950 33754 17956 33756
rect 18012 33754 18036 33756
rect 18092 33754 18116 33756
rect 18172 33754 18196 33756
rect 18252 33754 18258 33756
rect 18012 33702 18014 33754
rect 18194 33702 18196 33754
rect 17950 33700 17956 33702
rect 18012 33700 18036 33702
rect 18092 33700 18116 33702
rect 18172 33700 18196 33702
rect 18252 33700 18258 33702
rect 17950 33691 18258 33700
rect 17684 33108 17736 33114
rect 17684 33050 17736 33056
rect 17592 32224 17644 32230
rect 17592 32166 17644 32172
rect 17604 31482 17632 32166
rect 17696 32026 17724 33050
rect 18340 33046 18368 36740
rect 18432 36038 18460 37266
rect 18524 36718 18552 42350
rect 18616 40390 18644 43794
rect 18984 41414 19012 46990
rect 19536 45490 19564 53382
rect 19628 46714 19656 53926
rect 19720 53106 19748 56200
rect 20088 54262 20116 56200
rect 20076 54256 20128 54262
rect 20076 54198 20128 54204
rect 20456 53786 20484 56200
rect 20720 54256 20772 54262
rect 20720 54198 20772 54204
rect 20536 53984 20588 53990
rect 20536 53926 20588 53932
rect 20444 53780 20496 53786
rect 20444 53722 20496 53728
rect 20456 53582 20484 53722
rect 20444 53576 20496 53582
rect 20444 53518 20496 53524
rect 19708 53100 19760 53106
rect 19708 53042 19760 53048
rect 19800 52896 19852 52902
rect 19800 52838 19852 52844
rect 19616 46708 19668 46714
rect 19616 46650 19668 46656
rect 19628 45898 19656 46650
rect 19812 46034 19840 52838
rect 19892 49088 19944 49094
rect 19892 49030 19944 49036
rect 19800 46028 19852 46034
rect 19800 45970 19852 45976
rect 19616 45892 19668 45898
rect 19616 45834 19668 45840
rect 19524 45484 19576 45490
rect 19524 45426 19576 45432
rect 19432 45416 19484 45422
rect 19432 45358 19484 45364
rect 19064 45280 19116 45286
rect 19064 45222 19116 45228
rect 19076 44198 19104 45222
rect 19340 44736 19392 44742
rect 19340 44678 19392 44684
rect 19064 44192 19116 44198
rect 19064 44134 19116 44140
rect 19352 42650 19380 44678
rect 19444 44334 19472 45358
rect 19536 45286 19564 45426
rect 19524 45280 19576 45286
rect 19524 45222 19576 45228
rect 19708 45280 19760 45286
rect 19708 45222 19760 45228
rect 19432 44328 19484 44334
rect 19536 44305 19564 45222
rect 19616 44464 19668 44470
rect 19616 44406 19668 44412
rect 19432 44270 19484 44276
rect 19522 44296 19578 44305
rect 19444 43790 19472 44270
rect 19522 44231 19578 44240
rect 19432 43784 19484 43790
rect 19432 43726 19484 43732
rect 19168 42622 19380 42650
rect 19168 42158 19196 42622
rect 19340 42560 19392 42566
rect 19340 42502 19392 42508
rect 19248 42220 19300 42226
rect 19248 42162 19300 42168
rect 19156 42152 19208 42158
rect 19156 42094 19208 42100
rect 19064 41744 19116 41750
rect 19064 41686 19116 41692
rect 18892 41386 19012 41414
rect 18696 40452 18748 40458
rect 18696 40394 18748 40400
rect 18604 40384 18656 40390
rect 18604 40326 18656 40332
rect 18604 39024 18656 39030
rect 18604 38966 18656 38972
rect 18616 38894 18644 38966
rect 18604 38888 18656 38894
rect 18604 38830 18656 38836
rect 18616 38214 18644 38830
rect 18604 38208 18656 38214
rect 18604 38150 18656 38156
rect 18616 37942 18644 38150
rect 18604 37936 18656 37942
rect 18604 37878 18656 37884
rect 18512 36712 18564 36718
rect 18512 36654 18564 36660
rect 18512 36576 18564 36582
rect 18512 36518 18564 36524
rect 18420 36032 18472 36038
rect 18420 35974 18472 35980
rect 18328 33040 18380 33046
rect 18328 32982 18380 32988
rect 18156 32830 18368 32858
rect 18156 32774 18184 32830
rect 18144 32768 18196 32774
rect 18144 32710 18196 32716
rect 17950 32668 18258 32677
rect 17950 32666 17956 32668
rect 18012 32666 18036 32668
rect 18092 32666 18116 32668
rect 18172 32666 18196 32668
rect 18252 32666 18258 32668
rect 18012 32614 18014 32666
rect 18194 32614 18196 32666
rect 17950 32612 17956 32614
rect 18012 32612 18036 32614
rect 18092 32612 18116 32614
rect 18172 32612 18196 32614
rect 18252 32612 18258 32614
rect 17950 32603 18258 32612
rect 17868 32292 17920 32298
rect 17868 32234 17920 32240
rect 17684 32020 17736 32026
rect 17684 31962 17736 31968
rect 17592 31476 17644 31482
rect 17592 31418 17644 31424
rect 17696 30870 17724 31962
rect 17776 31272 17828 31278
rect 17776 31214 17828 31220
rect 17684 30864 17736 30870
rect 17684 30806 17736 30812
rect 17684 30592 17736 30598
rect 17684 30534 17736 30540
rect 17592 29708 17644 29714
rect 17592 29650 17644 29656
rect 17500 29096 17552 29102
rect 17498 29064 17500 29073
rect 17552 29064 17554 29073
rect 17408 29028 17460 29034
rect 17498 28999 17554 29008
rect 17408 28970 17460 28976
rect 17316 28212 17368 28218
rect 17316 28154 17368 28160
rect 17420 28098 17448 28970
rect 17604 28762 17632 29650
rect 17592 28756 17644 28762
rect 17592 28698 17644 28704
rect 17500 28416 17552 28422
rect 17500 28358 17552 28364
rect 17512 28218 17540 28358
rect 17500 28212 17552 28218
rect 17500 28154 17552 28160
rect 17420 28070 17540 28098
rect 17224 27328 17276 27334
rect 17224 27270 17276 27276
rect 17316 26988 17368 26994
rect 17316 26930 17368 26936
rect 17040 26308 17092 26314
rect 16960 26268 17040 26296
rect 17040 26250 17092 26256
rect 17132 26308 17184 26314
rect 17132 26250 17184 26256
rect 16948 25832 17000 25838
rect 16948 25774 17000 25780
rect 16960 24682 16988 25774
rect 17052 25362 17080 26250
rect 17040 25356 17092 25362
rect 17040 25298 17092 25304
rect 16948 24676 17000 24682
rect 16948 24618 17000 24624
rect 16856 23860 16908 23866
rect 16856 23802 16908 23808
rect 16960 23118 16988 24618
rect 17144 24070 17172 26250
rect 17224 25832 17276 25838
rect 17224 25774 17276 25780
rect 17236 24750 17264 25774
rect 17224 24744 17276 24750
rect 17224 24686 17276 24692
rect 17224 24336 17276 24342
rect 17224 24278 17276 24284
rect 17132 24064 17184 24070
rect 17132 24006 17184 24012
rect 17144 23254 17172 24006
rect 17132 23248 17184 23254
rect 17132 23190 17184 23196
rect 17040 23180 17092 23186
rect 17040 23122 17092 23128
rect 16948 23112 17000 23118
rect 16948 23054 17000 23060
rect 16960 22098 16988 23054
rect 16948 22092 17000 22098
rect 16948 22034 17000 22040
rect 16856 20800 16908 20806
rect 16856 20742 16908 20748
rect 16868 20602 16896 20742
rect 16856 20596 16908 20602
rect 16856 20538 16908 20544
rect 16764 20460 16816 20466
rect 16764 20402 16816 20408
rect 17052 19802 17080 23122
rect 17236 20874 17264 24278
rect 17328 22166 17356 26930
rect 17408 26852 17460 26858
rect 17408 26794 17460 26800
rect 17420 23186 17448 26794
rect 17512 26330 17540 28070
rect 17604 26450 17632 28698
rect 17592 26444 17644 26450
rect 17592 26386 17644 26392
rect 17512 26302 17632 26330
rect 17500 25356 17552 25362
rect 17500 25298 17552 25304
rect 17512 24410 17540 25298
rect 17604 24614 17632 26302
rect 17696 25294 17724 30534
rect 17788 28966 17816 31214
rect 17776 28960 17828 28966
rect 17776 28902 17828 28908
rect 17788 28626 17816 28902
rect 17776 28620 17828 28626
rect 17776 28562 17828 28568
rect 17880 28150 17908 32234
rect 18340 31754 18368 32830
rect 18524 32502 18552 36518
rect 18616 35204 18644 37878
rect 18708 36174 18736 40394
rect 18788 39432 18840 39438
rect 18788 39374 18840 39380
rect 18800 37806 18828 39374
rect 18788 37800 18840 37806
rect 18892 37777 18920 41386
rect 19076 39658 19104 41686
rect 19168 40594 19196 42094
rect 19260 41818 19288 42162
rect 19248 41812 19300 41818
rect 19248 41754 19300 41760
rect 19352 41750 19380 42502
rect 19444 42362 19472 43726
rect 19432 42356 19484 42362
rect 19432 42298 19484 42304
rect 19628 42022 19656 44406
rect 19616 42016 19668 42022
rect 19616 41958 19668 41964
rect 19340 41744 19392 41750
rect 19340 41686 19392 41692
rect 19352 41274 19380 41686
rect 19432 41472 19484 41478
rect 19432 41414 19484 41420
rect 19524 41472 19576 41478
rect 19524 41414 19576 41420
rect 19340 41268 19392 41274
rect 19340 41210 19392 41216
rect 19156 40588 19208 40594
rect 19156 40530 19208 40536
rect 18984 39630 19104 39658
rect 18984 38758 19012 39630
rect 19064 39024 19116 39030
rect 19064 38966 19116 38972
rect 18972 38752 19024 38758
rect 18972 38694 19024 38700
rect 18788 37742 18840 37748
rect 18878 37768 18934 37777
rect 18800 37618 18828 37742
rect 18878 37703 18934 37712
rect 18800 37590 19012 37618
rect 18696 36168 18748 36174
rect 18696 36110 18748 36116
rect 18984 35766 19012 37590
rect 19076 37194 19104 38966
rect 19168 37874 19196 40530
rect 19248 39364 19300 39370
rect 19248 39306 19300 39312
rect 19156 37868 19208 37874
rect 19156 37810 19208 37816
rect 19064 37188 19116 37194
rect 19064 37130 19116 37136
rect 19260 36922 19288 39306
rect 19444 38350 19472 41414
rect 19536 39642 19564 41414
rect 19524 39636 19576 39642
rect 19524 39578 19576 39584
rect 19628 38894 19656 41958
rect 19720 41682 19748 45222
rect 19904 43450 19932 49030
rect 20548 46714 20576 53926
rect 20732 53242 20760 54198
rect 20824 53582 20852 56200
rect 21192 54194 21220 56200
rect 21180 54188 21232 54194
rect 21180 54130 21232 54136
rect 21180 53984 21232 53990
rect 21180 53926 21232 53932
rect 20812 53576 20864 53582
rect 20812 53518 20864 53524
rect 20824 53242 20852 53518
rect 20720 53236 20772 53242
rect 20720 53178 20772 53184
rect 20812 53236 20864 53242
rect 20812 53178 20864 53184
rect 20996 51264 21048 51270
rect 20996 51206 21048 51212
rect 20720 48272 20772 48278
rect 20720 48214 20772 48220
rect 20536 46708 20588 46714
rect 20536 46650 20588 46656
rect 20548 45898 20576 46650
rect 20260 45892 20312 45898
rect 20260 45834 20312 45840
rect 20536 45892 20588 45898
rect 20536 45834 20588 45840
rect 20076 45824 20128 45830
rect 20076 45766 20128 45772
rect 19984 43716 20036 43722
rect 19984 43658 20036 43664
rect 19892 43444 19944 43450
rect 19892 43386 19944 43392
rect 19708 41676 19760 41682
rect 19708 41618 19760 41624
rect 19904 39914 19932 43386
rect 19996 40934 20024 43658
rect 19984 40928 20036 40934
rect 19984 40870 20036 40876
rect 19892 39908 19944 39914
rect 19892 39850 19944 39856
rect 19708 39840 19760 39846
rect 19708 39782 19760 39788
rect 19524 38888 19576 38894
rect 19524 38830 19576 38836
rect 19616 38888 19668 38894
rect 19616 38830 19668 38836
rect 19432 38344 19484 38350
rect 19432 38286 19484 38292
rect 19340 38208 19392 38214
rect 19340 38150 19392 38156
rect 19248 36916 19300 36922
rect 19248 36858 19300 36864
rect 19064 36780 19116 36786
rect 19064 36722 19116 36728
rect 18880 35760 18932 35766
rect 18880 35702 18932 35708
rect 18972 35760 19024 35766
rect 18972 35702 19024 35708
rect 18696 35692 18748 35698
rect 18696 35634 18748 35640
rect 18708 35494 18736 35634
rect 18696 35488 18748 35494
rect 18696 35430 18748 35436
rect 18892 35272 18920 35702
rect 18892 35244 19012 35272
rect 18788 35216 18840 35222
rect 18616 35176 18788 35204
rect 18788 35158 18840 35164
rect 18604 35080 18656 35086
rect 18604 35022 18656 35028
rect 18512 32496 18564 32502
rect 18512 32438 18564 32444
rect 18328 31748 18380 31754
rect 18328 31690 18380 31696
rect 17950 31580 18258 31589
rect 17950 31578 17956 31580
rect 18012 31578 18036 31580
rect 18092 31578 18116 31580
rect 18172 31578 18196 31580
rect 18252 31578 18258 31580
rect 18012 31526 18014 31578
rect 18194 31526 18196 31578
rect 17950 31524 17956 31526
rect 18012 31524 18036 31526
rect 18092 31524 18116 31526
rect 18172 31524 18196 31526
rect 18252 31524 18258 31526
rect 17950 31515 18258 31524
rect 18052 31272 18104 31278
rect 18052 31214 18104 31220
rect 18064 30734 18092 31214
rect 18142 30832 18198 30841
rect 18142 30767 18144 30776
rect 18196 30767 18198 30776
rect 18328 30796 18380 30802
rect 18144 30738 18196 30744
rect 18328 30738 18380 30744
rect 18052 30728 18104 30734
rect 18052 30670 18104 30676
rect 17950 30492 18258 30501
rect 17950 30490 17956 30492
rect 18012 30490 18036 30492
rect 18092 30490 18116 30492
rect 18172 30490 18196 30492
rect 18252 30490 18258 30492
rect 18012 30438 18014 30490
rect 18194 30438 18196 30490
rect 17950 30436 17956 30438
rect 18012 30436 18036 30438
rect 18092 30436 18116 30438
rect 18172 30436 18196 30438
rect 18252 30436 18258 30438
rect 17950 30427 18258 30436
rect 18234 29744 18290 29753
rect 18234 29679 18236 29688
rect 18288 29679 18290 29688
rect 18236 29650 18288 29656
rect 17950 29404 18258 29413
rect 17950 29402 17956 29404
rect 18012 29402 18036 29404
rect 18092 29402 18116 29404
rect 18172 29402 18196 29404
rect 18252 29402 18258 29404
rect 18012 29350 18014 29402
rect 18194 29350 18196 29402
rect 17950 29348 17956 29350
rect 18012 29348 18036 29350
rect 18092 29348 18116 29350
rect 18172 29348 18196 29350
rect 18252 29348 18258 29350
rect 17950 29339 18258 29348
rect 17950 28316 18258 28325
rect 17950 28314 17956 28316
rect 18012 28314 18036 28316
rect 18092 28314 18116 28316
rect 18172 28314 18196 28316
rect 18252 28314 18258 28316
rect 18012 28262 18014 28314
rect 18194 28262 18196 28314
rect 17950 28260 17956 28262
rect 18012 28260 18036 28262
rect 18092 28260 18116 28262
rect 18172 28260 18196 28262
rect 18252 28260 18258 28262
rect 17950 28251 18258 28260
rect 17868 28144 17920 28150
rect 17868 28086 17920 28092
rect 18052 28076 18104 28082
rect 18052 28018 18104 28024
rect 18064 27470 18092 28018
rect 18340 27470 18368 30738
rect 18512 30320 18564 30326
rect 18512 30262 18564 30268
rect 18420 29300 18472 29306
rect 18420 29242 18472 29248
rect 18052 27464 18104 27470
rect 17972 27424 18052 27452
rect 17972 27418 18000 27424
rect 17880 27390 18000 27418
rect 18052 27406 18104 27412
rect 18328 27464 18380 27470
rect 18328 27406 18380 27412
rect 17880 27112 17908 27390
rect 18432 27334 18460 29242
rect 18420 27328 18472 27334
rect 18420 27270 18472 27276
rect 17950 27228 18258 27237
rect 17950 27226 17956 27228
rect 18012 27226 18036 27228
rect 18092 27226 18116 27228
rect 18172 27226 18196 27228
rect 18252 27226 18258 27228
rect 18012 27174 18014 27226
rect 18194 27174 18196 27226
rect 17950 27172 17956 27174
rect 18012 27172 18036 27174
rect 18092 27172 18116 27174
rect 18172 27172 18196 27174
rect 18252 27172 18258 27174
rect 17950 27163 18258 27172
rect 18432 27130 18460 27270
rect 18420 27124 18472 27130
rect 17880 27084 18000 27112
rect 17972 26234 18000 27084
rect 18420 27066 18472 27072
rect 18328 26784 18380 26790
rect 18328 26726 18380 26732
rect 17880 26206 18000 26234
rect 17880 25922 17908 26206
rect 17950 26140 18258 26149
rect 17950 26138 17956 26140
rect 18012 26138 18036 26140
rect 18092 26138 18116 26140
rect 18172 26138 18196 26140
rect 18252 26138 18258 26140
rect 18012 26086 18014 26138
rect 18194 26086 18196 26138
rect 17950 26084 17956 26086
rect 18012 26084 18036 26086
rect 18092 26084 18116 26086
rect 18172 26084 18196 26086
rect 18252 26084 18258 26086
rect 17950 26075 18258 26084
rect 18340 26058 18368 26726
rect 18340 26030 18460 26058
rect 17880 25894 18000 25922
rect 17684 25288 17736 25294
rect 17972 25242 18000 25894
rect 17684 25230 17736 25236
rect 17880 25214 18000 25242
rect 17592 24608 17644 24614
rect 17592 24550 17644 24556
rect 17500 24404 17552 24410
rect 17500 24346 17552 24352
rect 17408 23180 17460 23186
rect 17408 23122 17460 23128
rect 17420 22234 17448 23122
rect 17512 22574 17540 24346
rect 17880 23866 17908 25214
rect 17950 25052 18258 25061
rect 17950 25050 17956 25052
rect 18012 25050 18036 25052
rect 18092 25050 18116 25052
rect 18172 25050 18196 25052
rect 18252 25050 18258 25052
rect 18012 24998 18014 25050
rect 18194 24998 18196 25050
rect 17950 24996 17956 24998
rect 18012 24996 18036 24998
rect 18092 24996 18116 24998
rect 18172 24996 18196 24998
rect 18252 24996 18258 24998
rect 17950 24987 18258 24996
rect 18432 24818 18460 26030
rect 18524 25770 18552 30262
rect 18616 28966 18644 35022
rect 18696 34944 18748 34950
rect 18696 34886 18748 34892
rect 18708 31346 18736 34886
rect 18800 33862 18828 35158
rect 18880 35148 18932 35154
rect 18880 35090 18932 35096
rect 18788 33856 18840 33862
rect 18788 33798 18840 33804
rect 18800 32774 18828 33798
rect 18788 32768 18840 32774
rect 18788 32710 18840 32716
rect 18892 32434 18920 35090
rect 18984 34746 19012 35244
rect 18972 34740 19024 34746
rect 18972 34682 19024 34688
rect 19076 34610 19104 36722
rect 19156 36712 19208 36718
rect 19156 36654 19208 36660
rect 19168 36582 19196 36654
rect 19156 36576 19208 36582
rect 19156 36518 19208 36524
rect 19064 34604 19116 34610
rect 19064 34546 19116 34552
rect 19064 34400 19116 34406
rect 19064 34342 19116 34348
rect 18972 33856 19024 33862
rect 18972 33798 19024 33804
rect 18984 33561 19012 33798
rect 18970 33552 19026 33561
rect 18970 33487 19026 33496
rect 19076 32570 19104 34342
rect 19064 32564 19116 32570
rect 19064 32506 19116 32512
rect 18880 32428 18932 32434
rect 18880 32370 18932 32376
rect 18892 31754 18920 32370
rect 18800 31726 18920 31754
rect 18696 31340 18748 31346
rect 18696 31282 18748 31288
rect 18800 29102 18828 31726
rect 18970 30696 19026 30705
rect 18970 30631 19026 30640
rect 18984 30598 19012 30631
rect 18972 30592 19024 30598
rect 18972 30534 19024 30540
rect 18880 30252 18932 30258
rect 18880 30194 18932 30200
rect 18788 29096 18840 29102
rect 18788 29038 18840 29044
rect 18604 28960 18656 28966
rect 18604 28902 18656 28908
rect 18616 28218 18644 28902
rect 18696 28416 18748 28422
rect 18696 28358 18748 28364
rect 18604 28212 18656 28218
rect 18604 28154 18656 28160
rect 18708 28098 18736 28358
rect 18616 28082 18736 28098
rect 18604 28076 18736 28082
rect 18656 28070 18736 28076
rect 18604 28018 18656 28024
rect 18800 28014 18828 29038
rect 18788 28008 18840 28014
rect 18788 27950 18840 27956
rect 18696 27328 18748 27334
rect 18696 27270 18748 27276
rect 18604 27124 18656 27130
rect 18604 27066 18656 27072
rect 18616 26994 18644 27066
rect 18604 26988 18656 26994
rect 18604 26930 18656 26936
rect 18604 26444 18656 26450
rect 18604 26386 18656 26392
rect 18616 25838 18644 26386
rect 18708 26042 18736 27270
rect 18800 26926 18828 27950
rect 18788 26920 18840 26926
rect 18788 26862 18840 26868
rect 18696 26036 18748 26042
rect 18696 25978 18748 25984
rect 18604 25832 18656 25838
rect 18604 25774 18656 25780
rect 18512 25764 18564 25770
rect 18512 25706 18564 25712
rect 18420 24812 18472 24818
rect 18420 24754 18472 24760
rect 18328 24608 18380 24614
rect 18328 24550 18380 24556
rect 17950 23964 18258 23973
rect 17950 23962 17956 23964
rect 18012 23962 18036 23964
rect 18092 23962 18116 23964
rect 18172 23962 18196 23964
rect 18252 23962 18258 23964
rect 18012 23910 18014 23962
rect 18194 23910 18196 23962
rect 17950 23908 17956 23910
rect 18012 23908 18036 23910
rect 18092 23908 18116 23910
rect 18172 23908 18196 23910
rect 18252 23908 18258 23910
rect 17950 23899 18258 23908
rect 17868 23860 17920 23866
rect 17868 23802 17920 23808
rect 17880 22710 17908 23802
rect 17950 22876 18258 22885
rect 17950 22874 17956 22876
rect 18012 22874 18036 22876
rect 18092 22874 18116 22876
rect 18172 22874 18196 22876
rect 18252 22874 18258 22876
rect 18012 22822 18014 22874
rect 18194 22822 18196 22874
rect 17950 22820 17956 22822
rect 18012 22820 18036 22822
rect 18092 22820 18116 22822
rect 18172 22820 18196 22822
rect 18252 22820 18258 22822
rect 17950 22811 18258 22820
rect 17868 22704 17920 22710
rect 17868 22646 17920 22652
rect 17500 22568 17552 22574
rect 17500 22510 17552 22516
rect 17408 22228 17460 22234
rect 17408 22170 17460 22176
rect 17316 22160 17368 22166
rect 17316 22102 17368 22108
rect 17328 21894 17356 22102
rect 17776 21956 17828 21962
rect 17776 21898 17828 21904
rect 17316 21888 17368 21894
rect 17316 21830 17368 21836
rect 17788 21690 17816 21898
rect 17950 21788 18258 21797
rect 17950 21786 17956 21788
rect 18012 21786 18036 21788
rect 18092 21786 18116 21788
rect 18172 21786 18196 21788
rect 18252 21786 18258 21788
rect 18012 21734 18014 21786
rect 18194 21734 18196 21786
rect 17950 21732 17956 21734
rect 18012 21732 18036 21734
rect 18092 21732 18116 21734
rect 18172 21732 18196 21734
rect 18252 21732 18258 21734
rect 17950 21723 18258 21732
rect 17776 21684 17828 21690
rect 17776 21626 17828 21632
rect 17224 20868 17276 20874
rect 17224 20810 17276 20816
rect 17132 20800 17184 20806
rect 17132 20742 17184 20748
rect 16960 19774 17080 19802
rect 16856 17740 16908 17746
rect 16856 17682 16908 17688
rect 16672 17332 16724 17338
rect 16672 17274 16724 17280
rect 16868 17134 16896 17682
rect 16856 17128 16908 17134
rect 16856 17070 16908 17076
rect 16592 16646 16712 16674
rect 16500 15978 16620 15994
rect 16500 15972 16632 15978
rect 16500 15966 16580 15972
rect 16500 15450 16528 15966
rect 16580 15914 16632 15920
rect 16684 15910 16712 16646
rect 16672 15904 16724 15910
rect 16672 15846 16724 15852
rect 16868 15570 16896 17070
rect 16960 16250 16988 19774
rect 17040 19712 17092 19718
rect 17040 19654 17092 19660
rect 16948 16244 17000 16250
rect 16948 16186 17000 16192
rect 17052 16130 17080 19654
rect 17144 18358 17172 20742
rect 17222 19952 17278 19961
rect 17222 19887 17278 19896
rect 17236 19854 17264 19887
rect 17224 19848 17276 19854
rect 17224 19790 17276 19796
rect 17500 19712 17552 19718
rect 17500 19654 17552 19660
rect 17408 19168 17460 19174
rect 17408 19110 17460 19116
rect 17132 18352 17184 18358
rect 17132 18294 17184 18300
rect 16960 16102 17080 16130
rect 16856 15564 16908 15570
rect 16856 15506 16908 15512
rect 16500 15434 16712 15450
rect 16500 15428 16724 15434
rect 16500 15422 16672 15428
rect 16316 14980 16528 15008
rect 16500 14890 16528 14980
rect 16396 14884 16448 14890
rect 16396 14826 16448 14832
rect 16488 14884 16540 14890
rect 16488 14826 16540 14832
rect 16304 14000 16356 14006
rect 16304 13942 16356 13948
rect 16316 12918 16344 13942
rect 16304 12912 16356 12918
rect 16304 12854 16356 12860
rect 16212 10804 16264 10810
rect 16212 10746 16264 10752
rect 16028 10464 16080 10470
rect 16028 10406 16080 10412
rect 15936 8968 15988 8974
rect 15936 8910 15988 8916
rect 16040 6914 16068 10406
rect 15948 6886 16068 6914
rect 15844 5772 15896 5778
rect 15844 5714 15896 5720
rect 15752 5364 15804 5370
rect 15752 5306 15804 5312
rect 15672 4678 15792 4706
rect 15476 3596 15528 3602
rect 15476 3538 15528 3544
rect 15384 2644 15436 2650
rect 15384 2586 15436 2592
rect 15108 2508 15160 2514
rect 15108 2450 15160 2456
rect 15120 800 15148 2450
rect 15488 800 15516 3538
rect 15658 2680 15714 2689
rect 15658 2615 15714 2624
rect 15672 2446 15700 2615
rect 15764 2446 15792 4678
rect 15844 2984 15896 2990
rect 15844 2926 15896 2932
rect 15660 2440 15712 2446
rect 15660 2382 15712 2388
rect 15752 2440 15804 2446
rect 15752 2382 15804 2388
rect 15856 800 15884 2926
rect 15948 2038 15976 6886
rect 16212 6112 16264 6118
rect 16212 6054 16264 6060
rect 16224 5302 16252 6054
rect 16212 5296 16264 5302
rect 16212 5238 16264 5244
rect 16028 5228 16080 5234
rect 16028 5170 16080 5176
rect 16040 3670 16068 5170
rect 16408 4622 16436 14826
rect 16488 14340 16540 14346
rect 16488 14282 16540 14288
rect 16500 12782 16528 14282
rect 16592 14278 16620 15422
rect 16672 15370 16724 15376
rect 16868 14414 16896 15506
rect 16856 14408 16908 14414
rect 16856 14350 16908 14356
rect 16580 14272 16632 14278
rect 16580 14214 16632 14220
rect 16592 14006 16620 14214
rect 16580 14000 16632 14006
rect 16580 13942 16632 13948
rect 16868 13870 16896 14350
rect 16856 13864 16908 13870
rect 16856 13806 16908 13812
rect 16868 12986 16896 13806
rect 16856 12980 16908 12986
rect 16856 12922 16908 12928
rect 16488 12776 16540 12782
rect 16488 12718 16540 12724
rect 16868 12306 16896 12922
rect 16856 12300 16908 12306
rect 16856 12242 16908 12248
rect 16488 9988 16540 9994
rect 16488 9930 16540 9936
rect 16396 4616 16448 4622
rect 16396 4558 16448 4564
rect 16212 4072 16264 4078
rect 16212 4014 16264 4020
rect 16028 3664 16080 3670
rect 16028 3606 16080 3612
rect 15936 2032 15988 2038
rect 15936 1974 15988 1980
rect 16224 800 16252 4014
rect 16500 3058 16528 9930
rect 16856 5364 16908 5370
rect 16856 5306 16908 5312
rect 16868 3058 16896 5306
rect 16960 5030 16988 16102
rect 17132 14952 17184 14958
rect 17132 14894 17184 14900
rect 17040 14068 17092 14074
rect 17040 14010 17092 14016
rect 17052 12986 17080 14010
rect 17144 13870 17172 14894
rect 17316 14272 17368 14278
rect 17316 14214 17368 14220
rect 17132 13864 17184 13870
rect 17132 13806 17184 13812
rect 17040 12980 17092 12986
rect 17040 12922 17092 12928
rect 17144 12442 17172 13806
rect 17224 13184 17276 13190
rect 17224 13126 17276 13132
rect 17236 12986 17264 13126
rect 17224 12980 17276 12986
rect 17224 12922 17276 12928
rect 17132 12436 17184 12442
rect 17132 12378 17184 12384
rect 17328 11830 17356 14214
rect 17316 11824 17368 11830
rect 17316 11766 17368 11772
rect 17328 6322 17356 11766
rect 17316 6316 17368 6322
rect 17316 6258 17368 6264
rect 16948 5024 17000 5030
rect 16948 4966 17000 4972
rect 16488 3052 16540 3058
rect 16488 2994 16540 3000
rect 16856 3052 16908 3058
rect 16856 2994 16908 3000
rect 16580 2916 16632 2922
rect 16580 2858 16632 2864
rect 16592 800 16620 2858
rect 17316 2848 17368 2854
rect 17316 2790 17368 2796
rect 16948 2440 17000 2446
rect 16948 2382 17000 2388
rect 16960 800 16988 2382
rect 17328 800 17356 2790
rect 17420 2378 17448 19110
rect 17512 14414 17540 19654
rect 17590 18864 17646 18873
rect 17590 18799 17592 18808
rect 17644 18799 17646 18808
rect 17592 18770 17644 18776
rect 17788 18426 17816 21626
rect 17868 21412 17920 21418
rect 17868 21354 17920 21360
rect 17776 18420 17828 18426
rect 17776 18362 17828 18368
rect 17776 18216 17828 18222
rect 17776 18158 17828 18164
rect 17788 17746 17816 18158
rect 17880 17746 17908 21354
rect 17950 20700 18258 20709
rect 17950 20698 17956 20700
rect 18012 20698 18036 20700
rect 18092 20698 18116 20700
rect 18172 20698 18196 20700
rect 18252 20698 18258 20700
rect 18012 20646 18014 20698
rect 18194 20646 18196 20698
rect 17950 20644 17956 20646
rect 18012 20644 18036 20646
rect 18092 20644 18116 20646
rect 18172 20644 18196 20646
rect 18252 20644 18258 20646
rect 17950 20635 18258 20644
rect 18236 20256 18288 20262
rect 18236 20198 18288 20204
rect 18248 19854 18276 20198
rect 18340 19922 18368 24550
rect 18524 24274 18552 25706
rect 18788 25696 18840 25702
rect 18788 25638 18840 25644
rect 18604 24744 18656 24750
rect 18604 24686 18656 24692
rect 18512 24268 18564 24274
rect 18512 24210 18564 24216
rect 18512 24064 18564 24070
rect 18512 24006 18564 24012
rect 18420 22432 18472 22438
rect 18420 22374 18472 22380
rect 18432 21690 18460 22374
rect 18420 21684 18472 21690
rect 18420 21626 18472 21632
rect 18524 21554 18552 24006
rect 18616 23322 18644 24686
rect 18800 24154 18828 25638
rect 18708 24126 18828 24154
rect 18892 24138 18920 30194
rect 18984 29730 19012 30534
rect 19064 30184 19116 30190
rect 19064 30126 19116 30132
rect 19076 29850 19104 30126
rect 19064 29844 19116 29850
rect 19064 29786 19116 29792
rect 18984 29702 19104 29730
rect 18972 27600 19024 27606
rect 18972 27542 19024 27548
rect 18984 24342 19012 27542
rect 18972 24336 19024 24342
rect 18972 24278 19024 24284
rect 18880 24132 18932 24138
rect 18604 23316 18656 23322
rect 18604 23258 18656 23264
rect 18708 23202 18736 24126
rect 18880 24074 18932 24080
rect 18788 24064 18840 24070
rect 18788 24006 18840 24012
rect 18616 23174 18736 23202
rect 18512 21548 18564 21554
rect 18512 21490 18564 21496
rect 18512 21344 18564 21350
rect 18512 21286 18564 21292
rect 18524 20942 18552 21286
rect 18616 21010 18644 23174
rect 18696 22432 18748 22438
rect 18696 22374 18748 22380
rect 18708 22098 18736 22374
rect 18696 22092 18748 22098
rect 18696 22034 18748 22040
rect 18604 21004 18656 21010
rect 18604 20946 18656 20952
rect 18512 20936 18564 20942
rect 18512 20878 18564 20884
rect 18708 20466 18736 22034
rect 18696 20460 18748 20466
rect 18696 20402 18748 20408
rect 18328 19916 18380 19922
rect 18328 19858 18380 19864
rect 18236 19848 18288 19854
rect 18236 19790 18288 19796
rect 17950 19612 18258 19621
rect 17950 19610 17956 19612
rect 18012 19610 18036 19612
rect 18092 19610 18116 19612
rect 18172 19610 18196 19612
rect 18252 19610 18258 19612
rect 18012 19558 18014 19610
rect 18194 19558 18196 19610
rect 17950 19556 17956 19558
rect 18012 19556 18036 19558
rect 18092 19556 18116 19558
rect 18172 19556 18196 19558
rect 18252 19556 18258 19558
rect 17950 19547 18258 19556
rect 18800 19378 18828 24006
rect 18880 23316 18932 23322
rect 18880 23258 18932 23264
rect 18892 20534 18920 23258
rect 18984 23186 19012 24278
rect 18972 23180 19024 23186
rect 18972 23122 19024 23128
rect 18984 22506 19012 23122
rect 18972 22500 19024 22506
rect 18972 22442 19024 22448
rect 19076 22386 19104 29702
rect 18984 22358 19104 22386
rect 18880 20528 18932 20534
rect 18880 20470 18932 20476
rect 18788 19372 18840 19378
rect 18788 19314 18840 19320
rect 18512 19236 18564 19242
rect 18512 19178 18564 19184
rect 17950 18524 18258 18533
rect 17950 18522 17956 18524
rect 18012 18522 18036 18524
rect 18092 18522 18116 18524
rect 18172 18522 18196 18524
rect 18252 18522 18258 18524
rect 18012 18470 18014 18522
rect 18194 18470 18196 18522
rect 17950 18468 17956 18470
rect 18012 18468 18036 18470
rect 18092 18468 18116 18470
rect 18172 18468 18196 18470
rect 18252 18468 18258 18470
rect 17950 18459 18258 18468
rect 18524 18329 18552 19178
rect 18788 19168 18840 19174
rect 18788 19110 18840 19116
rect 18510 18320 18566 18329
rect 18800 18290 18828 19110
rect 18510 18255 18566 18264
rect 18788 18284 18840 18290
rect 18524 18222 18552 18255
rect 18788 18226 18840 18232
rect 18512 18216 18564 18222
rect 18512 18158 18564 18164
rect 18512 18080 18564 18086
rect 18512 18022 18564 18028
rect 18328 17876 18380 17882
rect 18328 17818 18380 17824
rect 17776 17740 17828 17746
rect 17776 17682 17828 17688
rect 17868 17740 17920 17746
rect 17868 17682 17920 17688
rect 17866 17640 17922 17649
rect 18340 17610 18368 17818
rect 17866 17575 17922 17584
rect 18328 17604 18380 17610
rect 17880 17542 17908 17575
rect 18328 17546 18380 17552
rect 17868 17536 17920 17542
rect 17868 17478 17920 17484
rect 17950 17436 18258 17445
rect 17950 17434 17956 17436
rect 18012 17434 18036 17436
rect 18092 17434 18116 17436
rect 18172 17434 18196 17436
rect 18252 17434 18258 17436
rect 18012 17382 18014 17434
rect 18194 17382 18196 17434
rect 17950 17380 17956 17382
rect 18012 17380 18036 17382
rect 18092 17380 18116 17382
rect 18172 17380 18196 17382
rect 18252 17380 18258 17382
rect 17950 17371 18258 17380
rect 17592 17128 17644 17134
rect 17592 17070 17644 17076
rect 17604 15706 17632 17070
rect 18328 16992 18380 16998
rect 18328 16934 18380 16940
rect 17950 16348 18258 16357
rect 17950 16346 17956 16348
rect 18012 16346 18036 16348
rect 18092 16346 18116 16348
rect 18172 16346 18196 16348
rect 18252 16346 18258 16348
rect 18012 16294 18014 16346
rect 18194 16294 18196 16346
rect 17950 16292 17956 16294
rect 18012 16292 18036 16294
rect 18092 16292 18116 16294
rect 18172 16292 18196 16294
rect 18252 16292 18258 16294
rect 17950 16283 18258 16292
rect 17776 16244 17828 16250
rect 17776 16186 17828 16192
rect 17592 15700 17644 15706
rect 17592 15642 17644 15648
rect 17788 15502 17816 16186
rect 18340 15570 18368 16934
rect 18524 16794 18552 18022
rect 18604 17672 18656 17678
rect 18604 17614 18656 17620
rect 18512 16788 18564 16794
rect 18512 16730 18564 16736
rect 18328 15564 18380 15570
rect 18328 15506 18380 15512
rect 17776 15496 17828 15502
rect 17776 15438 17828 15444
rect 17868 15428 17920 15434
rect 17868 15370 17920 15376
rect 17500 14408 17552 14414
rect 17500 14350 17552 14356
rect 17592 14272 17644 14278
rect 17592 14214 17644 14220
rect 17604 14006 17632 14214
rect 17592 14000 17644 14006
rect 17592 13942 17644 13948
rect 17880 13734 17908 15370
rect 18512 15360 18564 15366
rect 18512 15302 18564 15308
rect 17950 15260 18258 15269
rect 17950 15258 17956 15260
rect 18012 15258 18036 15260
rect 18092 15258 18116 15260
rect 18172 15258 18196 15260
rect 18252 15258 18258 15260
rect 18012 15206 18014 15258
rect 18194 15206 18196 15258
rect 17950 15204 17956 15206
rect 18012 15204 18036 15206
rect 18092 15204 18116 15206
rect 18172 15204 18196 15206
rect 18252 15204 18258 15206
rect 17950 15195 18258 15204
rect 18524 15162 18552 15302
rect 18512 15156 18564 15162
rect 18512 15098 18564 15104
rect 18420 14884 18472 14890
rect 18420 14826 18472 14832
rect 18052 14612 18104 14618
rect 18052 14554 18104 14560
rect 18064 14414 18092 14554
rect 18052 14408 18104 14414
rect 18052 14350 18104 14356
rect 17950 14172 18258 14181
rect 17950 14170 17956 14172
rect 18012 14170 18036 14172
rect 18092 14170 18116 14172
rect 18172 14170 18196 14172
rect 18252 14170 18258 14172
rect 18012 14118 18014 14170
rect 18194 14118 18196 14170
rect 17950 14116 17956 14118
rect 18012 14116 18036 14118
rect 18092 14116 18116 14118
rect 18172 14116 18196 14118
rect 18252 14116 18258 14118
rect 17950 14107 18258 14116
rect 17868 13728 17920 13734
rect 17868 13670 17920 13676
rect 18432 13394 18460 14826
rect 18616 14074 18644 17614
rect 18696 17536 18748 17542
rect 18696 17478 18748 17484
rect 18708 17202 18736 17478
rect 18696 17196 18748 17202
rect 18696 17138 18748 17144
rect 18800 17082 18828 18226
rect 18984 17882 19012 22358
rect 19062 22264 19118 22273
rect 19062 22199 19118 22208
rect 19076 19122 19104 22199
rect 19168 19446 19196 36518
rect 19352 36378 19380 38150
rect 19536 38010 19564 38830
rect 19524 38004 19576 38010
rect 19524 37946 19576 37952
rect 19432 37800 19484 37806
rect 19432 37742 19484 37748
rect 19444 37262 19472 37742
rect 19536 37262 19564 37946
rect 19720 37738 19748 39782
rect 19800 39296 19852 39302
rect 19800 39238 19852 39244
rect 19892 39296 19944 39302
rect 19892 39238 19944 39244
rect 19708 37732 19760 37738
rect 19708 37674 19760 37680
rect 19432 37256 19484 37262
rect 19432 37198 19484 37204
rect 19524 37256 19576 37262
rect 19524 37198 19576 37204
rect 19432 36848 19484 36854
rect 19432 36790 19484 36796
rect 19340 36372 19392 36378
rect 19340 36314 19392 36320
rect 19444 36174 19472 36790
rect 19432 36168 19484 36174
rect 19432 36110 19484 36116
rect 19340 34672 19392 34678
rect 19340 34614 19392 34620
rect 19248 34604 19300 34610
rect 19248 34546 19300 34552
rect 19260 31958 19288 34546
rect 19248 31952 19300 31958
rect 19248 31894 19300 31900
rect 19248 29776 19300 29782
rect 19248 29718 19300 29724
rect 19260 28558 19288 29718
rect 19352 29238 19380 34614
rect 19444 34542 19472 36110
rect 19536 35494 19564 37198
rect 19614 36680 19670 36689
rect 19614 36615 19670 36624
rect 19628 36378 19656 36615
rect 19616 36372 19668 36378
rect 19616 36314 19668 36320
rect 19708 35828 19760 35834
rect 19708 35770 19760 35776
rect 19616 35760 19668 35766
rect 19616 35702 19668 35708
rect 19628 35494 19656 35702
rect 19524 35488 19576 35494
rect 19524 35430 19576 35436
rect 19616 35488 19668 35494
rect 19616 35430 19668 35436
rect 19536 34678 19564 35430
rect 19628 35222 19656 35430
rect 19616 35216 19668 35222
rect 19616 35158 19668 35164
rect 19524 34672 19576 34678
rect 19524 34614 19576 34620
rect 19720 34610 19748 35770
rect 19708 34604 19760 34610
rect 19708 34546 19760 34552
rect 19432 34536 19484 34542
rect 19432 34478 19484 34484
rect 19524 33924 19576 33930
rect 19524 33866 19576 33872
rect 19536 33114 19564 33866
rect 19616 33652 19668 33658
rect 19616 33594 19668 33600
rect 19524 33108 19576 33114
rect 19524 33050 19576 33056
rect 19628 31754 19656 33594
rect 19720 32570 19748 34546
rect 19708 32564 19760 32570
rect 19708 32506 19760 32512
rect 19812 32502 19840 39238
rect 19904 39001 19932 39238
rect 19890 38992 19946 39001
rect 19890 38927 19946 38936
rect 19996 38418 20024 40870
rect 20088 40594 20116 45766
rect 20076 40588 20128 40594
rect 20076 40530 20128 40536
rect 20168 40384 20220 40390
rect 20168 40326 20220 40332
rect 20076 39908 20128 39914
rect 20076 39850 20128 39856
rect 20088 39302 20116 39850
rect 20076 39296 20128 39302
rect 20076 39238 20128 39244
rect 20088 38978 20116 39238
rect 20180 39098 20208 40326
rect 20168 39092 20220 39098
rect 20168 39034 20220 39040
rect 20088 38950 20208 38978
rect 20180 38894 20208 38950
rect 20168 38888 20220 38894
rect 20168 38830 20220 38836
rect 19984 38412 20036 38418
rect 19984 38354 20036 38360
rect 19892 37868 19944 37874
rect 19892 37810 19944 37816
rect 19904 37670 19932 37810
rect 19892 37664 19944 37670
rect 19890 37632 19892 37641
rect 19944 37632 19946 37641
rect 19890 37567 19946 37576
rect 19984 35624 20036 35630
rect 20180 35578 20208 38830
rect 20272 35834 20300 45834
rect 20548 45801 20576 45834
rect 20534 45792 20590 45801
rect 20534 45727 20590 45736
rect 20536 42560 20588 42566
rect 20536 42502 20588 42508
rect 20548 42090 20576 42502
rect 20536 42084 20588 42090
rect 20536 42026 20588 42032
rect 20548 41070 20576 42026
rect 20536 41064 20588 41070
rect 20536 41006 20588 41012
rect 20536 40928 20588 40934
rect 20536 40870 20588 40876
rect 20548 40186 20576 40870
rect 20732 40594 20760 48214
rect 20904 45960 20956 45966
rect 20904 45902 20956 45908
rect 20812 45416 20864 45422
rect 20812 45358 20864 45364
rect 20824 44266 20852 45358
rect 20916 44810 20944 45902
rect 20904 44804 20956 44810
rect 20904 44746 20956 44752
rect 20812 44260 20864 44266
rect 20812 44202 20864 44208
rect 20824 43874 20852 44202
rect 20916 43994 20944 44746
rect 20904 43988 20956 43994
rect 20904 43930 20956 43936
rect 20824 43846 20944 43874
rect 20812 43784 20864 43790
rect 20812 43726 20864 43732
rect 20824 42566 20852 43726
rect 20916 42634 20944 43846
rect 20904 42628 20956 42634
rect 20904 42570 20956 42576
rect 20812 42560 20864 42566
rect 20812 42502 20864 42508
rect 20812 41676 20864 41682
rect 20812 41618 20864 41624
rect 20720 40588 20772 40594
rect 20720 40530 20772 40536
rect 20352 40180 20404 40186
rect 20352 40122 20404 40128
rect 20536 40180 20588 40186
rect 20536 40122 20588 40128
rect 20260 35828 20312 35834
rect 20260 35770 20312 35776
rect 20364 35578 20392 40122
rect 20720 39976 20772 39982
rect 20720 39918 20772 39924
rect 20444 39840 20496 39846
rect 20444 39782 20496 39788
rect 20456 37126 20484 39782
rect 20732 39386 20760 39918
rect 20824 39642 20852 41618
rect 20812 39636 20864 39642
rect 20812 39578 20864 39584
rect 20812 39500 20864 39506
rect 20916 39488 20944 42570
rect 21008 41682 21036 51206
rect 21192 44962 21220 53926
rect 21560 53582 21588 56200
rect 21824 54188 21876 54194
rect 21824 54130 21876 54136
rect 21732 54052 21784 54058
rect 21732 53994 21784 54000
rect 21548 53576 21600 53582
rect 21600 53524 21680 53530
rect 21548 53518 21680 53524
rect 21560 53502 21680 53518
rect 21272 53440 21324 53446
rect 21272 53382 21324 53388
rect 21456 53440 21508 53446
rect 21456 53382 21508 53388
rect 21548 53440 21600 53446
rect 21548 53382 21600 53388
rect 21284 45098 21312 53382
rect 21364 49972 21416 49978
rect 21364 49914 21416 49920
rect 21376 45370 21404 49914
rect 21468 45529 21496 53382
rect 21560 46034 21588 53382
rect 21652 53242 21680 53502
rect 21640 53236 21692 53242
rect 21640 53178 21692 53184
rect 21640 48544 21692 48550
rect 21640 48486 21692 48492
rect 21548 46028 21600 46034
rect 21548 45970 21600 45976
rect 21454 45520 21510 45529
rect 21454 45455 21510 45464
rect 21376 45342 21588 45370
rect 21284 45070 21404 45098
rect 21192 44934 21312 44962
rect 21180 44872 21232 44878
rect 21180 44814 21232 44820
rect 21088 44736 21140 44742
rect 21088 44678 21140 44684
rect 21100 44470 21128 44678
rect 21088 44464 21140 44470
rect 21088 44406 21140 44412
rect 21100 44198 21128 44406
rect 21088 44192 21140 44198
rect 21088 44134 21140 44140
rect 21100 43790 21128 44134
rect 21088 43784 21140 43790
rect 21088 43726 21140 43732
rect 21192 42702 21220 44814
rect 21180 42696 21232 42702
rect 21180 42638 21232 42644
rect 21192 42294 21220 42638
rect 21284 42566 21312 44934
rect 21376 44826 21404 45070
rect 21376 44798 21496 44826
rect 21468 44742 21496 44798
rect 21456 44736 21508 44742
rect 21456 44678 21508 44684
rect 21468 44334 21496 44678
rect 21456 44328 21508 44334
rect 21454 44296 21456 44305
rect 21508 44296 21510 44305
rect 21454 44231 21510 44240
rect 21272 42560 21324 42566
rect 21272 42502 21324 42508
rect 21180 42288 21232 42294
rect 21180 42230 21232 42236
rect 21088 42220 21140 42226
rect 21088 42162 21140 42168
rect 21100 42022 21128 42162
rect 21284 42106 21312 42502
rect 21192 42078 21312 42106
rect 21088 42016 21140 42022
rect 21088 41958 21140 41964
rect 20996 41676 21048 41682
rect 20996 41618 21048 41624
rect 21100 41614 21128 41958
rect 21088 41608 21140 41614
rect 21088 41550 21140 41556
rect 20996 40656 21048 40662
rect 20996 40598 21048 40604
rect 21008 40186 21036 40598
rect 20996 40180 21048 40186
rect 20996 40122 21048 40128
rect 20996 39636 21048 39642
rect 20996 39578 21048 39584
rect 20864 39460 20944 39488
rect 20812 39442 20864 39448
rect 20628 39364 20680 39370
rect 20732 39358 20944 39386
rect 20628 39306 20680 39312
rect 20640 39098 20668 39306
rect 20628 39092 20680 39098
rect 20628 39034 20680 39040
rect 20536 38752 20588 38758
rect 20536 38694 20588 38700
rect 20444 37120 20496 37126
rect 20444 37062 20496 37068
rect 20444 36372 20496 36378
rect 20444 36314 20496 36320
rect 20456 36174 20484 36314
rect 20444 36168 20496 36174
rect 20444 36110 20496 36116
rect 19984 35566 20036 35572
rect 19800 32496 19852 32502
rect 19800 32438 19852 32444
rect 19996 32434 20024 35566
rect 20088 35550 20208 35578
rect 20272 35550 20392 35578
rect 19984 32428 20036 32434
rect 19984 32370 20036 32376
rect 19984 32292 20036 32298
rect 19984 32234 20036 32240
rect 19996 32026 20024 32234
rect 19800 32020 19852 32026
rect 19800 31962 19852 31968
rect 19984 32020 20036 32026
rect 19984 31962 20036 31968
rect 19628 31726 19748 31754
rect 19616 31680 19668 31686
rect 19616 31622 19668 31628
rect 19628 31482 19656 31622
rect 19616 31476 19668 31482
rect 19616 31418 19668 31424
rect 19432 30592 19484 30598
rect 19432 30534 19484 30540
rect 19616 30592 19668 30598
rect 19616 30534 19668 30540
rect 19444 30394 19472 30534
rect 19432 30388 19484 30394
rect 19432 30330 19484 30336
rect 19444 30297 19472 30330
rect 19430 30288 19486 30297
rect 19430 30223 19486 30232
rect 19432 29504 19484 29510
rect 19432 29446 19484 29452
rect 19340 29232 19392 29238
rect 19340 29174 19392 29180
rect 19248 28552 19300 28558
rect 19248 28494 19300 28500
rect 19340 27668 19392 27674
rect 19340 27610 19392 27616
rect 19246 27568 19302 27577
rect 19246 27503 19248 27512
rect 19300 27503 19302 27512
rect 19248 27474 19300 27480
rect 19246 27160 19302 27169
rect 19246 27095 19248 27104
rect 19300 27095 19302 27104
rect 19248 27066 19300 27072
rect 19352 25226 19380 27610
rect 19340 25220 19392 25226
rect 19340 25162 19392 25168
rect 19352 24750 19380 25162
rect 19444 24954 19472 29446
rect 19524 28620 19576 28626
rect 19524 28562 19576 28568
rect 19536 27674 19564 28562
rect 19524 27668 19576 27674
rect 19524 27610 19576 27616
rect 19524 26512 19576 26518
rect 19524 26454 19576 26460
rect 19432 24948 19484 24954
rect 19432 24890 19484 24896
rect 19536 24818 19564 26454
rect 19628 25974 19656 30534
rect 19720 28694 19748 31726
rect 19812 29646 19840 31962
rect 19892 31680 19944 31686
rect 19892 31622 19944 31628
rect 19904 31482 19932 31622
rect 19892 31476 19944 31482
rect 19892 31418 19944 31424
rect 19984 30728 20036 30734
rect 19984 30670 20036 30676
rect 19996 30190 20024 30670
rect 19984 30184 20036 30190
rect 19982 30152 19984 30161
rect 20036 30152 20038 30161
rect 19982 30087 20038 30096
rect 19890 29744 19946 29753
rect 19890 29679 19892 29688
rect 19944 29679 19946 29688
rect 19984 29708 20036 29714
rect 19892 29650 19944 29656
rect 19984 29650 20036 29656
rect 19800 29640 19852 29646
rect 19800 29582 19852 29588
rect 19800 29300 19852 29306
rect 19800 29242 19852 29248
rect 19708 28688 19760 28694
rect 19708 28630 19760 28636
rect 19720 26314 19748 28630
rect 19812 27470 19840 29242
rect 19996 28506 20024 29650
rect 19904 28478 20024 28506
rect 19800 27464 19852 27470
rect 19800 27406 19852 27412
rect 19904 26858 19932 28478
rect 19984 28416 20036 28422
rect 19984 28358 20036 28364
rect 19892 26852 19944 26858
rect 19892 26794 19944 26800
rect 19708 26308 19760 26314
rect 19708 26250 19760 26256
rect 19616 25968 19668 25974
rect 19616 25910 19668 25916
rect 19524 24812 19576 24818
rect 19524 24754 19576 24760
rect 19340 24744 19392 24750
rect 19340 24686 19392 24692
rect 19892 24608 19944 24614
rect 19338 24576 19394 24585
rect 19892 24550 19944 24556
rect 19338 24511 19394 24520
rect 19352 21622 19380 24511
rect 19904 24206 19932 24550
rect 19996 24274 20024 28358
rect 20088 27878 20116 35550
rect 20168 35216 20220 35222
rect 20168 35158 20220 35164
rect 20180 35018 20208 35158
rect 20168 35012 20220 35018
rect 20168 34954 20220 34960
rect 20272 34950 20300 35550
rect 20352 35488 20404 35494
rect 20352 35430 20404 35436
rect 20260 34944 20312 34950
rect 20260 34886 20312 34892
rect 20260 34536 20312 34542
rect 20260 34478 20312 34484
rect 20168 34468 20220 34474
rect 20168 34410 20220 34416
rect 20180 33046 20208 34410
rect 20272 33998 20300 34478
rect 20260 33992 20312 33998
rect 20260 33934 20312 33940
rect 20168 33040 20220 33046
rect 20168 32982 20220 32988
rect 20180 29714 20208 32982
rect 20364 31890 20392 35430
rect 20444 35080 20496 35086
rect 20444 35022 20496 35028
rect 20456 32026 20484 35022
rect 20444 32020 20496 32026
rect 20444 31962 20496 31968
rect 20352 31884 20404 31890
rect 20352 31826 20404 31832
rect 20444 31748 20496 31754
rect 20444 31690 20496 31696
rect 20456 31482 20484 31690
rect 20444 31476 20496 31482
rect 20364 31436 20444 31464
rect 20168 29708 20220 29714
rect 20168 29650 20220 29656
rect 20076 27872 20128 27878
rect 20076 27814 20128 27820
rect 20076 27328 20128 27334
rect 20076 27270 20128 27276
rect 20088 26450 20116 27270
rect 20364 27062 20392 31436
rect 20444 31418 20496 31424
rect 20548 31346 20576 38694
rect 20720 38208 20772 38214
rect 20720 38150 20772 38156
rect 20628 37732 20680 37738
rect 20628 37674 20680 37680
rect 20640 33930 20668 37674
rect 20732 37194 20760 38150
rect 20812 37800 20864 37806
rect 20812 37742 20864 37748
rect 20720 37188 20772 37194
rect 20720 37130 20772 37136
rect 20732 36650 20760 37130
rect 20720 36644 20772 36650
rect 20720 36586 20772 36592
rect 20824 36242 20852 37742
rect 20916 37466 20944 39358
rect 21008 37890 21036 39578
rect 21100 38214 21128 41550
rect 21192 41478 21220 42078
rect 21272 41812 21324 41818
rect 21272 41754 21324 41760
rect 21180 41472 21232 41478
rect 21178 41440 21180 41449
rect 21232 41440 21234 41449
rect 21178 41375 21234 41384
rect 21088 38208 21140 38214
rect 21088 38150 21140 38156
rect 21008 37862 21128 37890
rect 20904 37460 20956 37466
rect 20904 37402 20956 37408
rect 20996 37460 21048 37466
rect 20996 37402 21048 37408
rect 20812 36236 20864 36242
rect 20812 36178 20864 36184
rect 20904 36100 20956 36106
rect 20904 36042 20956 36048
rect 20812 35828 20864 35834
rect 20812 35770 20864 35776
rect 20720 34944 20772 34950
rect 20720 34886 20772 34892
rect 20732 34202 20760 34886
rect 20720 34196 20772 34202
rect 20720 34138 20772 34144
rect 20628 33924 20680 33930
rect 20628 33866 20680 33872
rect 20720 32972 20772 32978
rect 20720 32914 20772 32920
rect 20628 32224 20680 32230
rect 20628 32166 20680 32172
rect 20536 31340 20588 31346
rect 20536 31282 20588 31288
rect 20444 30048 20496 30054
rect 20444 29990 20496 29996
rect 20456 28218 20484 29990
rect 20640 28558 20668 32166
rect 20732 32026 20760 32914
rect 20720 32020 20772 32026
rect 20720 31962 20772 31968
rect 20720 30796 20772 30802
rect 20720 30738 20772 30744
rect 20628 28552 20680 28558
rect 20628 28494 20680 28500
rect 20536 28484 20588 28490
rect 20536 28426 20588 28432
rect 20444 28212 20496 28218
rect 20444 28154 20496 28160
rect 20442 28112 20498 28121
rect 20548 28098 20576 28426
rect 20498 28070 20576 28098
rect 20442 28047 20444 28056
rect 20496 28047 20498 28056
rect 20444 28018 20496 28024
rect 20536 27872 20588 27878
rect 20536 27814 20588 27820
rect 20352 27056 20404 27062
rect 20352 26998 20404 27004
rect 20076 26444 20128 26450
rect 20076 26386 20128 26392
rect 20168 25832 20220 25838
rect 20168 25774 20220 25780
rect 20444 25832 20496 25838
rect 20444 25774 20496 25780
rect 19984 24268 20036 24274
rect 19984 24210 20036 24216
rect 19892 24200 19944 24206
rect 19892 24142 19944 24148
rect 20180 23322 20208 25774
rect 20456 24954 20484 25774
rect 20444 24948 20496 24954
rect 20444 24890 20496 24896
rect 20444 23520 20496 23526
rect 20444 23462 20496 23468
rect 20168 23316 20220 23322
rect 20168 23258 20220 23264
rect 19708 22228 19760 22234
rect 19708 22170 19760 22176
rect 19340 21616 19392 21622
rect 19340 21558 19392 21564
rect 19432 21616 19484 21622
rect 19432 21558 19484 21564
rect 19248 19508 19300 19514
rect 19248 19450 19300 19456
rect 19156 19440 19208 19446
rect 19156 19382 19208 19388
rect 19076 19094 19196 19122
rect 19064 18964 19116 18970
rect 19064 18906 19116 18912
rect 18972 17876 19024 17882
rect 18972 17818 19024 17824
rect 19076 17610 19104 18906
rect 18880 17604 18932 17610
rect 18880 17546 18932 17552
rect 19064 17604 19116 17610
rect 19064 17546 19116 17552
rect 18708 17054 18828 17082
rect 18604 14068 18656 14074
rect 18604 14010 18656 14016
rect 18616 13462 18644 14010
rect 18604 13456 18656 13462
rect 18604 13398 18656 13404
rect 18420 13388 18472 13394
rect 18420 13330 18472 13336
rect 18512 13184 18564 13190
rect 18512 13126 18564 13132
rect 17950 13084 18258 13093
rect 17950 13082 17956 13084
rect 18012 13082 18036 13084
rect 18092 13082 18116 13084
rect 18172 13082 18196 13084
rect 18252 13082 18258 13084
rect 18012 13030 18014 13082
rect 18194 13030 18196 13082
rect 17950 13028 17956 13030
rect 18012 13028 18036 13030
rect 18092 13028 18116 13030
rect 18172 13028 18196 13030
rect 18252 13028 18258 13030
rect 17950 13019 18258 13028
rect 18420 12844 18472 12850
rect 18420 12786 18472 12792
rect 17950 11996 18258 12005
rect 17950 11994 17956 11996
rect 18012 11994 18036 11996
rect 18092 11994 18116 11996
rect 18172 11994 18196 11996
rect 18252 11994 18258 11996
rect 18012 11942 18014 11994
rect 18194 11942 18196 11994
rect 17950 11940 17956 11942
rect 18012 11940 18036 11942
rect 18092 11940 18116 11942
rect 18172 11940 18196 11942
rect 18252 11940 18258 11942
rect 17950 11931 18258 11940
rect 18432 11898 18460 12786
rect 18420 11892 18472 11898
rect 18420 11834 18472 11840
rect 17950 10908 18258 10917
rect 17950 10906 17956 10908
rect 18012 10906 18036 10908
rect 18092 10906 18116 10908
rect 18172 10906 18196 10908
rect 18252 10906 18258 10908
rect 18012 10854 18014 10906
rect 18194 10854 18196 10906
rect 17950 10852 17956 10854
rect 18012 10852 18036 10854
rect 18092 10852 18116 10854
rect 18172 10852 18196 10854
rect 18252 10852 18258 10854
rect 17950 10843 18258 10852
rect 17950 9820 18258 9829
rect 17950 9818 17956 9820
rect 18012 9818 18036 9820
rect 18092 9818 18116 9820
rect 18172 9818 18196 9820
rect 18252 9818 18258 9820
rect 18012 9766 18014 9818
rect 18194 9766 18196 9818
rect 17950 9764 17956 9766
rect 18012 9764 18036 9766
rect 18092 9764 18116 9766
rect 18172 9764 18196 9766
rect 18252 9764 18258 9766
rect 17950 9755 18258 9764
rect 17776 8900 17828 8906
rect 17776 8842 17828 8848
rect 17684 3596 17736 3602
rect 17684 3538 17736 3544
rect 17408 2372 17460 2378
rect 17408 2314 17460 2320
rect 17696 800 17724 3538
rect 17788 3534 17816 8842
rect 17950 8732 18258 8741
rect 17950 8730 17956 8732
rect 18012 8730 18036 8732
rect 18092 8730 18116 8732
rect 18172 8730 18196 8732
rect 18252 8730 18258 8732
rect 18012 8678 18014 8730
rect 18194 8678 18196 8730
rect 17950 8676 17956 8678
rect 18012 8676 18036 8678
rect 18092 8676 18116 8678
rect 18172 8676 18196 8678
rect 18252 8676 18258 8678
rect 17950 8667 18258 8676
rect 17950 7644 18258 7653
rect 17950 7642 17956 7644
rect 18012 7642 18036 7644
rect 18092 7642 18116 7644
rect 18172 7642 18196 7644
rect 18252 7642 18258 7644
rect 18012 7590 18014 7642
rect 18194 7590 18196 7642
rect 17950 7588 17956 7590
rect 18012 7588 18036 7590
rect 18092 7588 18116 7590
rect 18172 7588 18196 7590
rect 18252 7588 18258 7590
rect 17950 7579 18258 7588
rect 18524 6914 18552 13126
rect 18708 12434 18736 17054
rect 18788 16788 18840 16794
rect 18788 16730 18840 16736
rect 18616 12406 18736 12434
rect 18616 8974 18644 12406
rect 18604 8968 18656 8974
rect 18604 8910 18656 8916
rect 18800 7886 18828 16730
rect 18788 7880 18840 7886
rect 18788 7822 18840 7828
rect 18524 6886 18644 6914
rect 17950 6556 18258 6565
rect 17950 6554 17956 6556
rect 18012 6554 18036 6556
rect 18092 6554 18116 6556
rect 18172 6554 18196 6556
rect 18252 6554 18258 6556
rect 18012 6502 18014 6554
rect 18194 6502 18196 6554
rect 17950 6500 17956 6502
rect 18012 6500 18036 6502
rect 18092 6500 18116 6502
rect 18172 6500 18196 6502
rect 18252 6500 18258 6502
rect 17950 6491 18258 6500
rect 17950 5468 18258 5477
rect 17950 5466 17956 5468
rect 18012 5466 18036 5468
rect 18092 5466 18116 5468
rect 18172 5466 18196 5468
rect 18252 5466 18258 5468
rect 18012 5414 18014 5466
rect 18194 5414 18196 5466
rect 17950 5412 17956 5414
rect 18012 5412 18036 5414
rect 18092 5412 18116 5414
rect 18172 5412 18196 5414
rect 18252 5412 18258 5414
rect 17950 5403 18258 5412
rect 18328 4548 18380 4554
rect 18328 4490 18380 4496
rect 17950 4380 18258 4389
rect 17950 4378 17956 4380
rect 18012 4378 18036 4380
rect 18092 4378 18116 4380
rect 18172 4378 18196 4380
rect 18252 4378 18258 4380
rect 18012 4326 18014 4378
rect 18194 4326 18196 4378
rect 17950 4324 17956 4326
rect 18012 4324 18036 4326
rect 18092 4324 18116 4326
rect 18172 4324 18196 4326
rect 18252 4324 18258 4326
rect 17950 4315 18258 4324
rect 17776 3528 17828 3534
rect 17776 3470 17828 3476
rect 17950 3292 18258 3301
rect 17950 3290 17956 3292
rect 18012 3290 18036 3292
rect 18092 3290 18116 3292
rect 18172 3290 18196 3292
rect 18252 3290 18258 3292
rect 18012 3238 18014 3290
rect 18194 3238 18196 3290
rect 17950 3236 17956 3238
rect 18012 3236 18036 3238
rect 18092 3236 18116 3238
rect 18172 3236 18196 3238
rect 18252 3236 18258 3238
rect 17950 3227 18258 3236
rect 18340 2854 18368 4490
rect 18616 4146 18644 6886
rect 18892 5778 18920 17546
rect 19076 17338 19104 17546
rect 19064 17332 19116 17338
rect 19064 17274 19116 17280
rect 19168 14618 19196 19094
rect 19260 16182 19288 19450
rect 19352 17218 19380 21558
rect 19444 21418 19472 21558
rect 19432 21412 19484 21418
rect 19432 21354 19484 21360
rect 19444 20534 19472 21354
rect 19616 21344 19668 21350
rect 19616 21286 19668 21292
rect 19628 21010 19656 21286
rect 19616 21004 19668 21010
rect 19616 20946 19668 20952
rect 19432 20528 19484 20534
rect 19432 20470 19484 20476
rect 19616 18828 19668 18834
rect 19616 18770 19668 18776
rect 19628 17338 19656 18770
rect 19616 17332 19668 17338
rect 19616 17274 19668 17280
rect 19352 17190 19656 17218
rect 19248 16176 19300 16182
rect 19248 16118 19300 16124
rect 19524 16040 19576 16046
rect 19524 15982 19576 15988
rect 19432 15904 19484 15910
rect 19432 15846 19484 15852
rect 19156 14612 19208 14618
rect 19156 14554 19208 14560
rect 18972 14340 19024 14346
rect 18972 14282 19024 14288
rect 18880 5772 18932 5778
rect 18880 5714 18932 5720
rect 18696 5024 18748 5030
rect 18696 4966 18748 4972
rect 18604 4140 18656 4146
rect 18604 4082 18656 4088
rect 18420 4072 18472 4078
rect 18420 4014 18472 4020
rect 18328 2848 18380 2854
rect 18328 2790 18380 2796
rect 17950 2204 18258 2213
rect 17950 2202 17956 2204
rect 18012 2202 18036 2204
rect 18092 2202 18116 2204
rect 18172 2202 18196 2204
rect 18252 2202 18258 2204
rect 18012 2150 18014 2202
rect 18194 2150 18196 2202
rect 17950 2148 17956 2150
rect 18012 2148 18036 2150
rect 18092 2148 18116 2150
rect 18172 2148 18196 2150
rect 18252 2148 18258 2150
rect 17950 2139 18258 2148
rect 18432 1170 18460 4014
rect 18708 3058 18736 4966
rect 18696 3052 18748 3058
rect 18696 2994 18748 3000
rect 18788 2848 18840 2854
rect 18788 2790 18840 2796
rect 18512 2372 18564 2378
rect 18512 2314 18564 2320
rect 18340 1142 18460 1170
rect 18064 870 18184 898
rect 18064 800 18092 870
rect 7852 734 8064 762
rect 8114 0 8170 800
rect 8482 0 8538 800
rect 8850 0 8906 800
rect 9218 0 9274 800
rect 9586 0 9642 800
rect 9954 0 10010 800
rect 10322 0 10378 800
rect 10690 0 10746 800
rect 11058 0 11114 800
rect 11426 0 11482 800
rect 11794 0 11850 800
rect 12162 0 12218 800
rect 12530 0 12586 800
rect 12898 0 12954 800
rect 13266 0 13322 800
rect 13634 0 13690 800
rect 14002 0 14058 800
rect 14370 0 14426 800
rect 14738 0 14794 800
rect 15106 0 15162 800
rect 15474 0 15530 800
rect 15842 0 15898 800
rect 16210 0 16266 800
rect 16578 0 16634 800
rect 16946 0 17002 800
rect 17314 0 17370 800
rect 17682 0 17738 800
rect 18050 0 18106 800
rect 18156 762 18184 870
rect 18340 762 18368 1142
rect 18524 898 18552 2314
rect 18432 870 18552 898
rect 18432 800 18460 870
rect 18800 800 18828 2790
rect 18984 2582 19012 14282
rect 19064 13864 19116 13870
rect 19064 13806 19116 13812
rect 19076 13326 19104 13806
rect 19338 13560 19394 13569
rect 19338 13495 19394 13504
rect 19352 13462 19380 13495
rect 19340 13456 19392 13462
rect 19340 13398 19392 13404
rect 19064 13320 19116 13326
rect 19064 13262 19116 13268
rect 19352 13258 19380 13398
rect 19340 13252 19392 13258
rect 19340 13194 19392 13200
rect 19444 13138 19472 15846
rect 19536 15162 19564 15982
rect 19524 15156 19576 15162
rect 19524 15098 19576 15104
rect 19628 13326 19656 17190
rect 19720 14006 19748 22170
rect 20180 22094 20208 23258
rect 20088 22066 20208 22094
rect 19800 21888 19852 21894
rect 19800 21830 19852 21836
rect 19812 21690 19840 21830
rect 19800 21684 19852 21690
rect 19800 21626 19852 21632
rect 20088 21486 20116 22066
rect 20076 21480 20128 21486
rect 20076 21422 20128 21428
rect 19800 19984 19852 19990
rect 19800 19926 19852 19932
rect 19812 16114 19840 19926
rect 20456 19786 20484 23462
rect 20444 19780 20496 19786
rect 20444 19722 20496 19728
rect 19892 19712 19944 19718
rect 19892 19654 19944 19660
rect 19800 16108 19852 16114
rect 19800 16050 19852 16056
rect 19800 15904 19852 15910
rect 19800 15846 19852 15852
rect 19812 15434 19840 15846
rect 19800 15428 19852 15434
rect 19800 15370 19852 15376
rect 19800 14476 19852 14482
rect 19800 14418 19852 14424
rect 19708 14000 19760 14006
rect 19708 13942 19760 13948
rect 19616 13320 19668 13326
rect 19616 13262 19668 13268
rect 19352 13110 19472 13138
rect 19248 12164 19300 12170
rect 19248 12106 19300 12112
rect 19064 12096 19116 12102
rect 19064 12038 19116 12044
rect 19076 11558 19104 12038
rect 19064 11552 19116 11558
rect 19064 11494 19116 11500
rect 19076 10606 19104 11494
rect 19260 11218 19288 12106
rect 19352 11830 19380 13110
rect 19432 12776 19484 12782
rect 19432 12718 19484 12724
rect 19444 12434 19472 12718
rect 19524 12640 19576 12646
rect 19708 12640 19760 12646
rect 19576 12588 19656 12594
rect 19524 12582 19656 12588
rect 19708 12582 19760 12588
rect 19536 12566 19656 12582
rect 19444 12406 19564 12434
rect 19432 12096 19484 12102
rect 19432 12038 19484 12044
rect 19340 11824 19392 11830
rect 19340 11766 19392 11772
rect 19248 11212 19300 11218
rect 19248 11154 19300 11160
rect 19260 10810 19288 11154
rect 19248 10804 19300 10810
rect 19248 10746 19300 10752
rect 19064 10600 19116 10606
rect 19064 10542 19116 10548
rect 19340 5772 19392 5778
rect 19340 5714 19392 5720
rect 19352 4622 19380 5714
rect 19444 5234 19472 12038
rect 19536 10742 19564 12406
rect 19628 11762 19656 12566
rect 19616 11756 19668 11762
rect 19616 11698 19668 11704
rect 19720 11218 19748 12582
rect 19708 11212 19760 11218
rect 19708 11154 19760 11160
rect 19524 10736 19576 10742
rect 19524 10678 19576 10684
rect 19812 6798 19840 14418
rect 19904 10062 19932 19654
rect 20548 18986 20576 27814
rect 20732 27674 20760 30738
rect 20824 30734 20852 35770
rect 20916 32570 20944 36042
rect 21008 36038 21036 37402
rect 21100 36242 21128 37862
rect 21284 36281 21312 41754
rect 21364 41064 21416 41070
rect 21364 41006 21416 41012
rect 21376 40458 21404 41006
rect 21560 41002 21588 45342
rect 21548 40996 21600 41002
rect 21548 40938 21600 40944
rect 21652 40662 21680 48486
rect 21744 45554 21772 53994
rect 21836 52698 21864 54130
rect 21928 53106 21956 56200
rect 22008 53984 22060 53990
rect 22008 53926 22060 53932
rect 21916 53100 21968 53106
rect 21916 53042 21968 53048
rect 21824 52692 21876 52698
rect 21824 52634 21876 52640
rect 22020 45558 22048 53926
rect 22296 53106 22324 56200
rect 22664 54262 22692 56200
rect 23032 56114 23060 56200
rect 23124 56114 23152 56222
rect 23032 56086 23152 56114
rect 22652 54256 22704 54262
rect 22652 54198 22704 54204
rect 22950 53884 23258 53893
rect 22950 53882 22956 53884
rect 23012 53882 23036 53884
rect 23092 53882 23116 53884
rect 23172 53882 23196 53884
rect 23252 53882 23258 53884
rect 23012 53830 23014 53882
rect 23194 53830 23196 53882
rect 22950 53828 22956 53830
rect 23012 53828 23036 53830
rect 23092 53828 23116 53830
rect 23172 53828 23196 53830
rect 23252 53828 23258 53830
rect 22950 53819 23258 53828
rect 23308 53650 23336 56222
rect 24122 56200 24178 57000
rect 24490 56200 24546 57000
rect 24858 56200 24914 57000
rect 25226 56200 25282 57000
rect 25594 56200 25650 57000
rect 25962 56200 26018 57000
rect 23940 54188 23992 54194
rect 23940 54130 23992 54136
rect 23296 53644 23348 53650
rect 23296 53586 23348 53592
rect 22284 53100 22336 53106
rect 22284 53042 22336 53048
rect 22192 52896 22244 52902
rect 22192 52838 22244 52844
rect 22744 52896 22796 52902
rect 22744 52838 22796 52844
rect 23480 52896 23532 52902
rect 23480 52838 23532 52844
rect 22204 52601 22232 52838
rect 22190 52592 22246 52601
rect 22190 52527 22246 52536
rect 22756 51270 22784 52838
rect 22950 52796 23258 52805
rect 22950 52794 22956 52796
rect 23012 52794 23036 52796
rect 23092 52794 23116 52796
rect 23172 52794 23196 52796
rect 23252 52794 23258 52796
rect 23012 52742 23014 52794
rect 23194 52742 23196 52794
rect 22950 52740 22956 52742
rect 23012 52740 23036 52742
rect 23092 52740 23116 52742
rect 23172 52740 23196 52742
rect 23252 52740 23258 52742
rect 22950 52731 23258 52740
rect 23492 52494 23520 52838
rect 23952 52698 23980 54130
rect 24136 54126 24164 56200
rect 24504 55214 24532 56200
rect 24412 55186 24532 55214
rect 24124 54120 24176 54126
rect 24124 54062 24176 54068
rect 24032 53576 24084 53582
rect 24032 53518 24084 53524
rect 23940 52692 23992 52698
rect 23940 52634 23992 52640
rect 23480 52488 23532 52494
rect 23480 52430 23532 52436
rect 23296 52352 23348 52358
rect 23296 52294 23348 52300
rect 22950 51708 23258 51717
rect 22950 51706 22956 51708
rect 23012 51706 23036 51708
rect 23092 51706 23116 51708
rect 23172 51706 23196 51708
rect 23252 51706 23258 51708
rect 23012 51654 23014 51706
rect 23194 51654 23196 51706
rect 22950 51652 22956 51654
rect 23012 51652 23036 51654
rect 23092 51652 23116 51654
rect 23172 51652 23196 51654
rect 23252 51652 23258 51654
rect 22950 51643 23258 51652
rect 22744 51264 22796 51270
rect 22744 51206 22796 51212
rect 22950 50620 23258 50629
rect 22950 50618 22956 50620
rect 23012 50618 23036 50620
rect 23092 50618 23116 50620
rect 23172 50618 23196 50620
rect 23252 50618 23258 50620
rect 23012 50566 23014 50618
rect 23194 50566 23196 50618
rect 22950 50564 22956 50566
rect 23012 50564 23036 50566
rect 23092 50564 23116 50566
rect 23172 50564 23196 50566
rect 23252 50564 23258 50566
rect 22950 50555 23258 50564
rect 22950 49532 23258 49541
rect 22950 49530 22956 49532
rect 23012 49530 23036 49532
rect 23092 49530 23116 49532
rect 23172 49530 23196 49532
rect 23252 49530 23258 49532
rect 23012 49478 23014 49530
rect 23194 49478 23196 49530
rect 22950 49476 22956 49478
rect 23012 49476 23036 49478
rect 23092 49476 23116 49478
rect 23172 49476 23196 49478
rect 23252 49476 23258 49478
rect 22950 49467 23258 49476
rect 22950 48444 23258 48453
rect 22950 48442 22956 48444
rect 23012 48442 23036 48444
rect 23092 48442 23116 48444
rect 23172 48442 23196 48444
rect 23252 48442 23258 48444
rect 23012 48390 23014 48442
rect 23194 48390 23196 48442
rect 22950 48388 22956 48390
rect 23012 48388 23036 48390
rect 23092 48388 23116 48390
rect 23172 48388 23196 48390
rect 23252 48388 23258 48390
rect 22950 48379 23258 48388
rect 22950 47356 23258 47365
rect 22950 47354 22956 47356
rect 23012 47354 23036 47356
rect 23092 47354 23116 47356
rect 23172 47354 23196 47356
rect 23252 47354 23258 47356
rect 23012 47302 23014 47354
rect 23194 47302 23196 47354
rect 22950 47300 22956 47302
rect 23012 47300 23036 47302
rect 23092 47300 23116 47302
rect 23172 47300 23196 47302
rect 23252 47300 23258 47302
rect 22950 47291 23258 47300
rect 23308 47258 23336 52294
rect 23492 52154 23520 52430
rect 23480 52148 23532 52154
rect 23480 52090 23532 52096
rect 23848 51264 23900 51270
rect 23848 51206 23900 51212
rect 23388 50176 23440 50182
rect 23388 50118 23440 50124
rect 23296 47252 23348 47258
rect 23296 47194 23348 47200
rect 23296 46368 23348 46374
rect 23296 46310 23348 46316
rect 22950 46268 23258 46277
rect 22950 46266 22956 46268
rect 23012 46266 23036 46268
rect 23092 46266 23116 46268
rect 23172 46266 23196 46268
rect 23252 46266 23258 46268
rect 23012 46214 23014 46266
rect 23194 46214 23196 46266
rect 22950 46212 22956 46214
rect 23012 46212 23036 46214
rect 23092 46212 23116 46214
rect 23172 46212 23196 46214
rect 23252 46212 23258 46214
rect 22950 46203 23258 46212
rect 22284 46096 22336 46102
rect 22284 46038 22336 46044
rect 21744 45526 21956 45554
rect 21928 44946 21956 45526
rect 22008 45552 22060 45558
rect 22008 45494 22060 45500
rect 21916 44940 21968 44946
rect 21916 44882 21968 44888
rect 22100 44328 22152 44334
rect 22100 44270 22152 44276
rect 22112 43994 22140 44270
rect 22100 43988 22152 43994
rect 22100 43930 22152 43936
rect 22008 43784 22060 43790
rect 22008 43726 22060 43732
rect 22020 43450 22048 43726
rect 22008 43444 22060 43450
rect 22008 43386 22060 43392
rect 22008 43240 22060 43246
rect 22008 43182 22060 43188
rect 22020 42702 22048 43182
rect 22008 42696 22060 42702
rect 22008 42638 22060 42644
rect 22112 41682 22140 43930
rect 22296 43382 22324 46038
rect 22650 45520 22706 45529
rect 22650 45455 22652 45464
rect 22704 45455 22706 45464
rect 22652 45426 22704 45432
rect 22664 44878 22692 45426
rect 22950 45180 23258 45189
rect 22950 45178 22956 45180
rect 23012 45178 23036 45180
rect 23092 45178 23116 45180
rect 23172 45178 23196 45180
rect 23252 45178 23258 45180
rect 23012 45126 23014 45178
rect 23194 45126 23196 45178
rect 22950 45124 22956 45126
rect 23012 45124 23036 45126
rect 23092 45124 23116 45126
rect 23172 45124 23196 45126
rect 23252 45124 23258 45126
rect 22950 45115 23258 45124
rect 22744 45008 22796 45014
rect 22744 44950 22796 44956
rect 22652 44872 22704 44878
rect 22652 44814 22704 44820
rect 22468 44736 22520 44742
rect 22468 44678 22520 44684
rect 22284 43376 22336 43382
rect 22284 43318 22336 43324
rect 22284 42696 22336 42702
rect 22284 42638 22336 42644
rect 22192 42152 22244 42158
rect 22192 42094 22244 42100
rect 22100 41676 22152 41682
rect 22100 41618 22152 41624
rect 21916 41608 21968 41614
rect 21916 41550 21968 41556
rect 21928 41414 21956 41550
rect 21836 41386 21956 41414
rect 21732 41064 21784 41070
rect 21732 41006 21784 41012
rect 21640 40656 21692 40662
rect 21640 40598 21692 40604
rect 21456 40588 21508 40594
rect 21456 40530 21508 40536
rect 21364 40452 21416 40458
rect 21364 40394 21416 40400
rect 21376 38962 21404 40394
rect 21364 38956 21416 38962
rect 21364 38898 21416 38904
rect 21270 36272 21326 36281
rect 21088 36236 21140 36242
rect 21270 36207 21326 36216
rect 21088 36178 21140 36184
rect 20996 36032 21048 36038
rect 20996 35974 21048 35980
rect 20904 32564 20956 32570
rect 20904 32506 20956 32512
rect 20904 31680 20956 31686
rect 20904 31622 20956 31628
rect 20916 31142 20944 31622
rect 21008 31482 21036 35974
rect 21100 31958 21128 36178
rect 21284 32570 21312 36207
rect 21468 36174 21496 40530
rect 21652 40474 21680 40598
rect 21560 40446 21680 40474
rect 21560 38214 21588 40446
rect 21640 40384 21692 40390
rect 21640 40326 21692 40332
rect 21652 39506 21680 40326
rect 21744 40186 21772 41006
rect 21732 40180 21784 40186
rect 21732 40122 21784 40128
rect 21836 40050 21864 41386
rect 22008 41268 22060 41274
rect 22008 41210 22060 41216
rect 21824 40044 21876 40050
rect 21824 39986 21876 39992
rect 21640 39500 21692 39506
rect 21640 39442 21692 39448
rect 21548 38208 21600 38214
rect 21548 38150 21600 38156
rect 21560 37874 21588 38150
rect 21548 37868 21600 37874
rect 21548 37810 21600 37816
rect 21652 37194 21680 39442
rect 21836 38894 21864 39986
rect 22020 39982 22048 41210
rect 22204 41070 22232 42094
rect 22192 41064 22244 41070
rect 22192 41006 22244 41012
rect 22296 40594 22324 42638
rect 22376 42220 22428 42226
rect 22376 42162 22428 42168
rect 22284 40588 22336 40594
rect 22284 40530 22336 40536
rect 22008 39976 22060 39982
rect 22008 39918 22060 39924
rect 21916 39296 21968 39302
rect 21916 39238 21968 39244
rect 21824 38888 21876 38894
rect 21824 38830 21876 38836
rect 21640 37188 21692 37194
rect 21640 37130 21692 37136
rect 21546 36816 21602 36825
rect 21546 36751 21602 36760
rect 21456 36168 21508 36174
rect 21456 36110 21508 36116
rect 21468 36038 21496 36110
rect 21456 36032 21508 36038
rect 21456 35974 21508 35980
rect 21468 32722 21496 35974
rect 21376 32694 21496 32722
rect 21272 32564 21324 32570
rect 21272 32506 21324 32512
rect 21180 32360 21232 32366
rect 21180 32302 21232 32308
rect 21088 31952 21140 31958
rect 21088 31894 21140 31900
rect 21192 31754 21220 32302
rect 21100 31726 21220 31754
rect 20996 31476 21048 31482
rect 20996 31418 21048 31424
rect 20904 31136 20956 31142
rect 20904 31078 20956 31084
rect 20812 30728 20864 30734
rect 20812 30670 20864 30676
rect 20812 30592 20864 30598
rect 20812 30534 20864 30540
rect 20824 30190 20852 30534
rect 20812 30184 20864 30190
rect 20812 30126 20864 30132
rect 20916 30002 20944 31078
rect 20824 29974 20944 30002
rect 20720 27668 20772 27674
rect 20720 27610 20772 27616
rect 20824 26518 20852 29974
rect 20996 29504 21048 29510
rect 20996 29446 21048 29452
rect 20904 28416 20956 28422
rect 20902 28384 20904 28393
rect 20956 28384 20958 28393
rect 20902 28319 20958 28328
rect 20916 28150 20944 28319
rect 20904 28144 20956 28150
rect 20904 28086 20956 28092
rect 20812 26512 20864 26518
rect 20812 26454 20864 26460
rect 20904 25492 20956 25498
rect 20904 25434 20956 25440
rect 20720 24064 20772 24070
rect 20720 24006 20772 24012
rect 20732 22030 20760 24006
rect 20812 22568 20864 22574
rect 20812 22510 20864 22516
rect 20720 22024 20772 22030
rect 20720 21966 20772 21972
rect 20720 21344 20772 21350
rect 20824 21332 20852 22510
rect 20772 21304 20852 21332
rect 20720 21286 20772 21292
rect 20720 20868 20772 20874
rect 20720 20810 20772 20816
rect 20732 20398 20760 20810
rect 20916 20806 20944 25434
rect 20904 20800 20956 20806
rect 20904 20742 20956 20748
rect 20720 20392 20772 20398
rect 20720 20334 20772 20340
rect 20628 20324 20680 20330
rect 20628 20266 20680 20272
rect 20456 18958 20576 18986
rect 19984 18896 20036 18902
rect 19984 18838 20036 18844
rect 19996 16658 20024 18838
rect 20456 18834 20484 18958
rect 20536 18896 20588 18902
rect 20536 18838 20588 18844
rect 20444 18828 20496 18834
rect 20444 18770 20496 18776
rect 20352 18624 20404 18630
rect 20352 18566 20404 18572
rect 20076 18216 20128 18222
rect 20076 18158 20128 18164
rect 19984 16652 20036 16658
rect 19984 16594 20036 16600
rect 19982 15600 20038 15609
rect 19982 15535 19984 15544
rect 20036 15535 20038 15544
rect 19984 15506 20036 15512
rect 20088 12434 20116 18158
rect 20260 16448 20312 16454
rect 20260 16390 20312 16396
rect 20272 15570 20300 16390
rect 20260 15564 20312 15570
rect 20260 15506 20312 15512
rect 20364 15162 20392 18566
rect 20548 15502 20576 18838
rect 20536 15496 20588 15502
rect 20536 15438 20588 15444
rect 20352 15156 20404 15162
rect 20352 15098 20404 15104
rect 20640 15026 20668 20266
rect 20732 19922 20760 20334
rect 20720 19916 20772 19922
rect 20720 19858 20772 19864
rect 21008 19854 21036 29446
rect 21100 28762 21128 31726
rect 21376 31686 21404 32694
rect 21180 31680 21232 31686
rect 21180 31622 21232 31628
rect 21364 31680 21416 31686
rect 21364 31622 21416 31628
rect 21192 30938 21220 31622
rect 21376 31210 21404 31622
rect 21272 31204 21324 31210
rect 21272 31146 21324 31152
rect 21364 31204 21416 31210
rect 21364 31146 21416 31152
rect 21180 30932 21232 30938
rect 21180 30874 21232 30880
rect 21180 29776 21232 29782
rect 21180 29718 21232 29724
rect 21088 28756 21140 28762
rect 21088 28698 21140 28704
rect 21100 27674 21128 28698
rect 21192 28626 21220 29718
rect 21180 28620 21232 28626
rect 21180 28562 21232 28568
rect 21088 27668 21140 27674
rect 21088 27610 21140 27616
rect 21088 25152 21140 25158
rect 21088 25094 21140 25100
rect 21100 24274 21128 25094
rect 21192 24274 21220 28562
rect 21088 24268 21140 24274
rect 21088 24210 21140 24216
rect 21180 24268 21232 24274
rect 21180 24210 21232 24216
rect 21284 24138 21312 31146
rect 21560 30734 21588 36751
rect 21652 34202 21680 37130
rect 21732 36712 21784 36718
rect 21732 36654 21784 36660
rect 21744 35154 21772 36654
rect 21824 36372 21876 36378
rect 21824 36314 21876 36320
rect 21836 36038 21864 36314
rect 21824 36032 21876 36038
rect 21824 35974 21876 35980
rect 21928 35154 21956 39238
rect 22020 39030 22048 39918
rect 22100 39296 22152 39302
rect 22388 39284 22416 42162
rect 22480 39370 22508 44678
rect 22560 43376 22612 43382
rect 22560 43318 22612 43324
rect 22572 42786 22600 43318
rect 22572 42758 22692 42786
rect 22560 42628 22612 42634
rect 22560 42570 22612 42576
rect 22572 42158 22600 42570
rect 22560 42152 22612 42158
rect 22560 42094 22612 42100
rect 22664 41970 22692 42758
rect 22756 42294 22784 44950
rect 22836 44736 22888 44742
rect 22836 44678 22888 44684
rect 22848 42362 22876 44678
rect 22950 44092 23258 44101
rect 22950 44090 22956 44092
rect 23012 44090 23036 44092
rect 23092 44090 23116 44092
rect 23172 44090 23196 44092
rect 23252 44090 23258 44092
rect 23012 44038 23014 44090
rect 23194 44038 23196 44090
rect 22950 44036 22956 44038
rect 23012 44036 23036 44038
rect 23092 44036 23116 44038
rect 23172 44036 23196 44038
rect 23252 44036 23258 44038
rect 22950 44027 23258 44036
rect 22950 43004 23258 43013
rect 22950 43002 22956 43004
rect 23012 43002 23036 43004
rect 23092 43002 23116 43004
rect 23172 43002 23196 43004
rect 23252 43002 23258 43004
rect 23012 42950 23014 43002
rect 23194 42950 23196 43002
rect 22950 42948 22956 42950
rect 23012 42948 23036 42950
rect 23092 42948 23116 42950
rect 23172 42948 23196 42950
rect 23252 42948 23258 42950
rect 22950 42939 23258 42948
rect 22836 42356 22888 42362
rect 22836 42298 22888 42304
rect 22744 42288 22796 42294
rect 22744 42230 22796 42236
rect 22572 41942 22692 41970
rect 22572 41274 22600 41942
rect 22652 41472 22704 41478
rect 22652 41414 22704 41420
rect 22756 41414 22784 42230
rect 22950 41916 23258 41925
rect 22950 41914 22956 41916
rect 23012 41914 23036 41916
rect 23092 41914 23116 41916
rect 23172 41914 23196 41916
rect 23252 41914 23258 41916
rect 23012 41862 23014 41914
rect 23194 41862 23196 41914
rect 22950 41860 22956 41862
rect 23012 41860 23036 41862
rect 23092 41860 23116 41862
rect 23172 41860 23196 41862
rect 23252 41860 23258 41862
rect 22950 41851 23258 41860
rect 23204 41744 23256 41750
rect 23204 41686 23256 41692
rect 23216 41414 23244 41686
rect 23308 41562 23336 46310
rect 23400 43432 23428 50118
rect 23860 47802 23888 51206
rect 23848 47796 23900 47802
rect 23848 47738 23900 47744
rect 24044 47734 24072 53518
rect 24216 52488 24268 52494
rect 24216 52430 24268 52436
rect 24032 47728 24084 47734
rect 24032 47670 24084 47676
rect 23848 46572 23900 46578
rect 23848 46514 23900 46520
rect 23860 46374 23888 46514
rect 23848 46368 23900 46374
rect 23848 46310 23900 46316
rect 23860 45121 23888 46310
rect 24228 45966 24256 52430
rect 24412 52018 24440 55186
rect 24492 53440 24544 53446
rect 24492 53382 24544 53388
rect 24400 52012 24452 52018
rect 24400 51954 24452 51960
rect 24400 51808 24452 51814
rect 24400 51750 24452 51756
rect 24412 47802 24440 51750
rect 24400 47796 24452 47802
rect 24400 47738 24452 47744
rect 24216 45960 24268 45966
rect 24216 45902 24268 45908
rect 24124 45824 24176 45830
rect 24124 45766 24176 45772
rect 24136 45490 24164 45766
rect 24124 45484 24176 45490
rect 24124 45426 24176 45432
rect 23846 45112 23902 45121
rect 23846 45047 23902 45056
rect 24124 44940 24176 44946
rect 24124 44882 24176 44888
rect 23572 44736 23624 44742
rect 23572 44678 23624 44684
rect 23400 43404 23520 43432
rect 23492 43194 23520 43404
rect 23400 43166 23520 43194
rect 23400 41682 23428 43166
rect 23584 41818 23612 44678
rect 23756 44328 23808 44334
rect 23756 44270 23808 44276
rect 23768 43858 23796 44270
rect 23756 43852 23808 43858
rect 23756 43794 23808 43800
rect 23756 43716 23808 43722
rect 23756 43658 23808 43664
rect 23768 43450 23796 43658
rect 23756 43444 23808 43450
rect 23756 43386 23808 43392
rect 23664 43376 23716 43382
rect 23664 43318 23716 43324
rect 23676 42702 23704 43318
rect 23664 42696 23716 42702
rect 23664 42638 23716 42644
rect 23676 42226 23704 42638
rect 23848 42356 23900 42362
rect 23848 42298 23900 42304
rect 23664 42220 23716 42226
rect 23664 42162 23716 42168
rect 23572 41812 23624 41818
rect 23572 41754 23624 41760
rect 23388 41676 23440 41682
rect 23388 41618 23440 41624
rect 23664 41676 23716 41682
rect 23664 41618 23716 41624
rect 23308 41534 23612 41562
rect 23480 41472 23532 41478
rect 23480 41414 23532 41420
rect 22560 41268 22612 41274
rect 22560 41210 22612 41216
rect 22560 41064 22612 41070
rect 22560 41006 22612 41012
rect 22468 39364 22520 39370
rect 22468 39306 22520 39312
rect 22100 39238 22152 39244
rect 22204 39256 22416 39284
rect 22008 39024 22060 39030
rect 22008 38966 22060 38972
rect 22112 38962 22140 39238
rect 22100 38956 22152 38962
rect 22100 38898 22152 38904
rect 22008 38888 22060 38894
rect 22060 38836 22140 38842
rect 22008 38830 22140 38836
rect 22020 38814 22140 38830
rect 22112 38758 22140 38814
rect 22008 38752 22060 38758
rect 22008 38694 22060 38700
rect 22100 38752 22152 38758
rect 22100 38694 22152 38700
rect 22020 36922 22048 38694
rect 22100 38412 22152 38418
rect 22100 38354 22152 38360
rect 22112 37942 22140 38354
rect 22204 38010 22232 39256
rect 22468 38888 22520 38894
rect 22468 38830 22520 38836
rect 22376 38752 22428 38758
rect 22376 38694 22428 38700
rect 22284 38344 22336 38350
rect 22284 38286 22336 38292
rect 22192 38004 22244 38010
rect 22192 37946 22244 37952
rect 22100 37936 22152 37942
rect 22100 37878 22152 37884
rect 22296 37330 22324 38286
rect 22388 38010 22416 38694
rect 22480 38282 22508 38830
rect 22468 38276 22520 38282
rect 22468 38218 22520 38224
rect 22376 38004 22428 38010
rect 22376 37946 22428 37952
rect 22480 37890 22508 38218
rect 22388 37862 22508 37890
rect 22284 37324 22336 37330
rect 22284 37266 22336 37272
rect 22008 36916 22060 36922
rect 22008 36858 22060 36864
rect 22296 36786 22324 37266
rect 22192 36780 22244 36786
rect 22192 36722 22244 36728
rect 22284 36780 22336 36786
rect 22284 36722 22336 36728
rect 22100 36032 22152 36038
rect 22100 35974 22152 35980
rect 21732 35148 21784 35154
rect 21732 35090 21784 35096
rect 21916 35148 21968 35154
rect 21916 35090 21968 35096
rect 22008 34400 22060 34406
rect 22008 34342 22060 34348
rect 21640 34196 21692 34202
rect 21640 34138 21692 34144
rect 21916 33652 21968 33658
rect 21916 33594 21968 33600
rect 21732 33108 21784 33114
rect 21732 33050 21784 33056
rect 21638 31784 21694 31793
rect 21638 31719 21694 31728
rect 21652 31142 21680 31719
rect 21640 31136 21692 31142
rect 21640 31078 21692 31084
rect 21548 30728 21600 30734
rect 21548 30670 21600 30676
rect 21744 29481 21772 33050
rect 21928 32978 21956 33594
rect 21916 32972 21968 32978
rect 21916 32914 21968 32920
rect 22020 29646 22048 34342
rect 22112 33538 22140 35974
rect 22204 34184 22232 36722
rect 22284 35080 22336 35086
rect 22284 35022 22336 35028
rect 22296 34542 22324 35022
rect 22388 34746 22416 37862
rect 22468 37732 22520 37738
rect 22468 37674 22520 37680
rect 22480 34746 22508 37674
rect 22572 36310 22600 41006
rect 22664 40186 22692 41414
rect 22756 41386 22876 41414
rect 23216 41386 23336 41414
rect 22744 41268 22796 41274
rect 22744 41210 22796 41216
rect 22652 40180 22704 40186
rect 22652 40122 22704 40128
rect 22652 39976 22704 39982
rect 22652 39918 22704 39924
rect 22664 39030 22692 39918
rect 22756 39642 22784 41210
rect 22848 40390 22876 41386
rect 22950 40828 23258 40837
rect 22950 40826 22956 40828
rect 23012 40826 23036 40828
rect 23092 40826 23116 40828
rect 23172 40826 23196 40828
rect 23252 40826 23258 40828
rect 23012 40774 23014 40826
rect 23194 40774 23196 40826
rect 22950 40772 22956 40774
rect 23012 40772 23036 40774
rect 23092 40772 23116 40774
rect 23172 40772 23196 40774
rect 23252 40772 23258 40774
rect 22950 40763 23258 40772
rect 22836 40384 22888 40390
rect 22836 40326 22888 40332
rect 22744 39636 22796 39642
rect 22744 39578 22796 39584
rect 22848 39438 22876 40326
rect 22950 39740 23258 39749
rect 22950 39738 22956 39740
rect 23012 39738 23036 39740
rect 23092 39738 23116 39740
rect 23172 39738 23196 39740
rect 23252 39738 23258 39740
rect 23012 39686 23014 39738
rect 23194 39686 23196 39738
rect 22950 39684 22956 39686
rect 23012 39684 23036 39686
rect 23092 39684 23116 39686
rect 23172 39684 23196 39686
rect 23252 39684 23258 39686
rect 22950 39675 23258 39684
rect 23204 39636 23256 39642
rect 23204 39578 23256 39584
rect 22836 39432 22888 39438
rect 22836 39374 22888 39380
rect 23216 39370 23244 39578
rect 23204 39364 23256 39370
rect 23204 39306 23256 39312
rect 22652 39024 22704 39030
rect 22652 38966 22704 38972
rect 22664 38418 22692 38966
rect 22950 38652 23258 38661
rect 22950 38650 22956 38652
rect 23012 38650 23036 38652
rect 23092 38650 23116 38652
rect 23172 38650 23196 38652
rect 23252 38650 23258 38652
rect 23012 38598 23014 38650
rect 23194 38598 23196 38650
rect 22950 38596 22956 38598
rect 23012 38596 23036 38598
rect 23092 38596 23116 38598
rect 23172 38596 23196 38598
rect 23252 38596 23258 38598
rect 22950 38587 23258 38596
rect 22744 38548 22796 38554
rect 22744 38490 22796 38496
rect 22652 38412 22704 38418
rect 22652 38354 22704 38360
rect 22652 37664 22704 37670
rect 22652 37606 22704 37612
rect 22560 36304 22612 36310
rect 22560 36246 22612 36252
rect 22376 34740 22428 34746
rect 22376 34682 22428 34688
rect 22468 34740 22520 34746
rect 22468 34682 22520 34688
rect 22284 34536 22336 34542
rect 22284 34478 22336 34484
rect 22468 34400 22520 34406
rect 22468 34342 22520 34348
rect 22204 34156 22416 34184
rect 22284 34060 22336 34066
rect 22284 34002 22336 34008
rect 22112 33510 22232 33538
rect 22100 32564 22152 32570
rect 22100 32506 22152 32512
rect 22008 29640 22060 29646
rect 22008 29582 22060 29588
rect 22112 29578 22140 32506
rect 22204 31822 22232 33510
rect 22296 32978 22324 34002
rect 22284 32972 22336 32978
rect 22284 32914 22336 32920
rect 22388 32366 22416 34156
rect 22480 33862 22508 34342
rect 22664 34082 22692 37606
rect 22756 36258 22784 38490
rect 22928 38480 22980 38486
rect 22928 38422 22980 38428
rect 22836 38208 22888 38214
rect 22836 38150 22888 38156
rect 22848 36378 22876 38150
rect 22940 37670 22968 38422
rect 23308 38418 23336 41386
rect 23388 41132 23440 41138
rect 23388 41074 23440 41080
rect 23400 40526 23428 41074
rect 23388 40520 23440 40526
rect 23388 40462 23440 40468
rect 23386 40352 23442 40361
rect 23386 40287 23442 40296
rect 23400 39642 23428 40287
rect 23388 39636 23440 39642
rect 23388 39578 23440 39584
rect 23400 39438 23428 39578
rect 23388 39432 23440 39438
rect 23388 39374 23440 39380
rect 23388 38820 23440 38826
rect 23388 38762 23440 38768
rect 23296 38412 23348 38418
rect 23296 38354 23348 38360
rect 23400 38350 23428 38762
rect 23492 38740 23520 41414
rect 23584 39982 23612 41534
rect 23676 40118 23704 41618
rect 23756 41608 23808 41614
rect 23756 41550 23808 41556
rect 23664 40112 23716 40118
rect 23664 40054 23716 40060
rect 23572 39976 23624 39982
rect 23572 39918 23624 39924
rect 23664 39976 23716 39982
rect 23664 39918 23716 39924
rect 23492 38712 23612 38740
rect 23388 38344 23440 38350
rect 23388 38286 23440 38292
rect 23400 37942 23428 38286
rect 23388 37936 23440 37942
rect 23388 37878 23440 37884
rect 22928 37664 22980 37670
rect 22928 37606 22980 37612
rect 22950 37564 23258 37573
rect 22950 37562 22956 37564
rect 23012 37562 23036 37564
rect 23092 37562 23116 37564
rect 23172 37562 23196 37564
rect 23252 37562 23258 37564
rect 23012 37510 23014 37562
rect 23194 37510 23196 37562
rect 22950 37508 22956 37510
rect 23012 37508 23036 37510
rect 23092 37508 23116 37510
rect 23172 37508 23196 37510
rect 23252 37508 23258 37510
rect 22950 37499 23258 37508
rect 23020 37120 23072 37126
rect 23020 37062 23072 37068
rect 23032 36854 23060 37062
rect 23020 36848 23072 36854
rect 23020 36790 23072 36796
rect 23032 36718 23060 36790
rect 23020 36712 23072 36718
rect 23020 36654 23072 36660
rect 23216 36638 23336 36666
rect 23216 36582 23244 36638
rect 23204 36576 23256 36582
rect 23204 36518 23256 36524
rect 22950 36476 23258 36485
rect 22950 36474 22956 36476
rect 23012 36474 23036 36476
rect 23092 36474 23116 36476
rect 23172 36474 23196 36476
rect 23252 36474 23258 36476
rect 23012 36422 23014 36474
rect 23194 36422 23196 36474
rect 22950 36420 22956 36422
rect 23012 36420 23036 36422
rect 23092 36420 23116 36422
rect 23172 36420 23196 36422
rect 23252 36420 23258 36422
rect 22950 36411 23258 36420
rect 22836 36372 22888 36378
rect 22836 36314 22888 36320
rect 22756 36230 22876 36258
rect 22744 35488 22796 35494
rect 22744 35430 22796 35436
rect 22756 35290 22784 35430
rect 22744 35284 22796 35290
rect 22744 35226 22796 35232
rect 22756 35193 22784 35226
rect 22742 35184 22798 35193
rect 22742 35119 22798 35128
rect 22744 34944 22796 34950
rect 22744 34886 22796 34892
rect 22572 34054 22692 34082
rect 22468 33856 22520 33862
rect 22468 33798 22520 33804
rect 22480 32842 22508 33798
rect 22572 33114 22600 34054
rect 22652 33924 22704 33930
rect 22652 33866 22704 33872
rect 22664 33658 22692 33866
rect 22652 33652 22704 33658
rect 22652 33594 22704 33600
rect 22560 33108 22612 33114
rect 22560 33050 22612 33056
rect 22560 32972 22612 32978
rect 22560 32914 22612 32920
rect 22468 32836 22520 32842
rect 22468 32778 22520 32784
rect 22376 32360 22428 32366
rect 22376 32302 22428 32308
rect 22284 31952 22336 31958
rect 22284 31894 22336 31900
rect 22376 31952 22428 31958
rect 22376 31894 22428 31900
rect 22192 31816 22244 31822
rect 22192 31758 22244 31764
rect 22296 30326 22324 31894
rect 22388 30326 22416 31894
rect 22468 31884 22520 31890
rect 22468 31826 22520 31832
rect 22480 30666 22508 31826
rect 22572 30802 22600 32914
rect 22652 32768 22704 32774
rect 22652 32710 22704 32716
rect 22560 30796 22612 30802
rect 22560 30738 22612 30744
rect 22468 30660 22520 30666
rect 22468 30602 22520 30608
rect 22284 30320 22336 30326
rect 22284 30262 22336 30268
rect 22376 30320 22428 30326
rect 22376 30262 22428 30268
rect 22192 30184 22244 30190
rect 22192 30126 22244 30132
rect 22100 29572 22152 29578
rect 22100 29514 22152 29520
rect 21730 29472 21786 29481
rect 22204 29458 22232 30126
rect 22572 30122 22600 30738
rect 22560 30116 22612 30122
rect 22560 30058 22612 30064
rect 22282 29744 22338 29753
rect 22282 29679 22284 29688
rect 22336 29679 22338 29688
rect 22468 29708 22520 29714
rect 22284 29650 22336 29656
rect 22468 29650 22520 29656
rect 21730 29407 21786 29416
rect 22112 29430 22232 29458
rect 22112 28626 22140 29430
rect 22192 29096 22244 29102
rect 22192 29038 22244 29044
rect 22100 28620 22152 28626
rect 22100 28562 22152 28568
rect 22204 28558 22232 29038
rect 22192 28552 22244 28558
rect 22192 28494 22244 28500
rect 21364 28416 21416 28422
rect 21364 28358 21416 28364
rect 21376 24818 21404 28358
rect 21640 27940 21692 27946
rect 21640 27882 21692 27888
rect 21456 27464 21508 27470
rect 21456 27406 21508 27412
rect 21468 26382 21496 27406
rect 21456 26376 21508 26382
rect 21456 26318 21508 26324
rect 21468 25362 21496 26318
rect 21548 25696 21600 25702
rect 21548 25638 21600 25644
rect 21456 25356 21508 25362
rect 21456 25298 21508 25304
rect 21364 24812 21416 24818
rect 21364 24754 21416 24760
rect 21456 24268 21508 24274
rect 21456 24210 21508 24216
rect 21272 24132 21324 24138
rect 21272 24074 21324 24080
rect 21088 24064 21140 24070
rect 21088 24006 21140 24012
rect 21100 23866 21128 24006
rect 21088 23860 21140 23866
rect 21088 23802 21140 23808
rect 21272 23180 21324 23186
rect 21272 23122 21324 23128
rect 21088 22772 21140 22778
rect 21088 22714 21140 22720
rect 21100 19854 21128 22714
rect 21284 22506 21312 23122
rect 21468 22778 21496 24210
rect 21456 22772 21508 22778
rect 21456 22714 21508 22720
rect 21272 22500 21324 22506
rect 21272 22442 21324 22448
rect 21272 20868 21324 20874
rect 21272 20810 21324 20816
rect 21284 20602 21312 20810
rect 21272 20596 21324 20602
rect 21272 20538 21324 20544
rect 20996 19848 21048 19854
rect 20996 19790 21048 19796
rect 21088 19848 21140 19854
rect 21088 19790 21140 19796
rect 21560 18766 21588 25638
rect 21652 22710 21680 27882
rect 22284 27464 22336 27470
rect 22284 27406 22336 27412
rect 22296 27130 22324 27406
rect 22284 27124 22336 27130
rect 22284 27066 22336 27072
rect 21732 26308 21784 26314
rect 21732 26250 21784 26256
rect 21744 25158 21772 26250
rect 22282 26072 22338 26081
rect 22282 26007 22338 26016
rect 22296 25906 22324 26007
rect 22480 25974 22508 29650
rect 22664 28218 22692 32710
rect 22756 31958 22784 34886
rect 22848 33096 22876 36230
rect 23308 36038 23336 36638
rect 23112 36032 23164 36038
rect 23112 35974 23164 35980
rect 23296 36032 23348 36038
rect 23296 35974 23348 35980
rect 23400 35986 23428 37878
rect 23480 37664 23532 37670
rect 23480 37606 23532 37612
rect 23492 36378 23520 37606
rect 23480 36372 23532 36378
rect 23480 36314 23532 36320
rect 23124 35578 23152 35974
rect 23400 35958 23520 35986
rect 23492 35834 23520 35958
rect 23480 35828 23532 35834
rect 23480 35770 23532 35776
rect 23124 35550 23336 35578
rect 22950 35388 23258 35397
rect 22950 35386 22956 35388
rect 23012 35386 23036 35388
rect 23092 35386 23116 35388
rect 23172 35386 23196 35388
rect 23252 35386 23258 35388
rect 23012 35334 23014 35386
rect 23194 35334 23196 35386
rect 22950 35332 22956 35334
rect 23012 35332 23036 35334
rect 23092 35332 23116 35334
rect 23172 35332 23196 35334
rect 23252 35332 23258 35334
rect 22950 35323 23258 35332
rect 23204 34944 23256 34950
rect 23204 34886 23256 34892
rect 23216 34746 23244 34886
rect 23204 34740 23256 34746
rect 23204 34682 23256 34688
rect 22950 34300 23258 34309
rect 22950 34298 22956 34300
rect 23012 34298 23036 34300
rect 23092 34298 23116 34300
rect 23172 34298 23196 34300
rect 23252 34298 23258 34300
rect 23012 34246 23014 34298
rect 23194 34246 23196 34298
rect 22950 34244 22956 34246
rect 23012 34244 23036 34246
rect 23092 34244 23116 34246
rect 23172 34244 23196 34246
rect 23252 34244 23258 34246
rect 22950 34235 23258 34244
rect 23308 33386 23336 35550
rect 23492 34066 23520 35770
rect 23480 34060 23532 34066
rect 23480 34002 23532 34008
rect 23492 33522 23520 34002
rect 23584 33998 23612 38712
rect 23676 37233 23704 39918
rect 23768 38298 23796 41550
rect 23860 41274 23888 42298
rect 23848 41268 23900 41274
rect 23848 41210 23900 41216
rect 24136 41070 24164 44882
rect 24228 44538 24256 45902
rect 24504 44878 24532 53382
rect 24872 53038 24900 56200
rect 24952 53100 25004 53106
rect 24952 53042 25004 53048
rect 24860 53032 24912 53038
rect 24860 52974 24912 52980
rect 24768 52624 24820 52630
rect 24674 52592 24730 52601
rect 24768 52566 24820 52572
rect 24674 52527 24730 52536
rect 24584 52352 24636 52358
rect 24584 52294 24636 52300
rect 24596 52154 24624 52294
rect 24584 52148 24636 52154
rect 24584 52090 24636 52096
rect 24688 52018 24716 52527
rect 24676 52012 24728 52018
rect 24676 51954 24728 51960
rect 24688 51610 24716 51954
rect 24676 51604 24728 51610
rect 24676 51546 24728 51552
rect 24780 51542 24808 52566
rect 24768 51536 24820 51542
rect 24768 51478 24820 51484
rect 24768 49836 24820 49842
rect 24768 49778 24820 49784
rect 24780 49201 24808 49778
rect 24766 49192 24822 49201
rect 24766 49127 24822 49136
rect 24768 48748 24820 48754
rect 24768 48690 24820 48696
rect 24780 47841 24808 48690
rect 24860 48000 24912 48006
rect 24860 47942 24912 47948
rect 24766 47832 24822 47841
rect 24766 47767 24822 47776
rect 24872 47666 24900 47942
rect 24860 47660 24912 47666
rect 24860 47602 24912 47608
rect 24964 47190 24992 53042
rect 25240 52902 25268 56200
rect 25608 53718 25636 56200
rect 25596 53712 25648 53718
rect 25596 53654 25648 53660
rect 25320 53440 25372 53446
rect 25320 53382 25372 53388
rect 25228 52896 25280 52902
rect 25228 52838 25280 52844
rect 25228 52488 25280 52494
rect 25228 52430 25280 52436
rect 25240 52018 25268 52430
rect 25228 52012 25280 52018
rect 25228 51954 25280 51960
rect 25240 51921 25268 51954
rect 25226 51912 25282 51921
rect 25226 51847 25282 51856
rect 25332 51406 25360 53382
rect 25976 52630 26004 56200
rect 25964 52624 26016 52630
rect 25964 52566 26016 52572
rect 25688 51808 25740 51814
rect 25688 51750 25740 51756
rect 25320 51400 25372 51406
rect 25320 51342 25372 51348
rect 25332 51241 25360 51342
rect 25596 51264 25648 51270
rect 25318 51232 25374 51241
rect 25596 51206 25648 51212
rect 25318 51167 25374 51176
rect 25320 50924 25372 50930
rect 25320 50866 25372 50872
rect 25136 50720 25188 50726
rect 25136 50662 25188 50668
rect 24952 47184 25004 47190
rect 24952 47126 25004 47132
rect 24952 46980 25004 46986
rect 24952 46922 25004 46928
rect 24676 46572 24728 46578
rect 24676 46514 24728 46520
rect 24584 46096 24636 46102
rect 24584 46038 24636 46044
rect 24492 44872 24544 44878
rect 24492 44814 24544 44820
rect 24216 44532 24268 44538
rect 24216 44474 24268 44480
rect 24228 43994 24256 44474
rect 24216 43988 24268 43994
rect 24216 43930 24268 43936
rect 24228 43382 24256 43930
rect 24400 43444 24452 43450
rect 24400 43386 24452 43392
rect 24216 43376 24268 43382
rect 24216 43318 24268 43324
rect 24412 41750 24440 43386
rect 24596 42566 24624 46038
rect 24688 45898 24716 46514
rect 24858 46472 24914 46481
rect 24858 46407 24860 46416
rect 24912 46407 24914 46416
rect 24860 46378 24912 46384
rect 24872 46034 24900 46378
rect 24860 46028 24912 46034
rect 24860 45970 24912 45976
rect 24964 45914 24992 46922
rect 25044 46164 25096 46170
rect 25044 46106 25096 46112
rect 24676 45892 24728 45898
rect 24676 45834 24728 45840
rect 24872 45886 24992 45914
rect 24688 43761 24716 45834
rect 24766 45792 24822 45801
rect 24766 45727 24822 45736
rect 24780 45422 24808 45727
rect 24768 45416 24820 45422
rect 24768 45358 24820 45364
rect 24766 44432 24822 44441
rect 24766 44367 24822 44376
rect 24780 43994 24808 44367
rect 24768 43988 24820 43994
rect 24768 43930 24820 43936
rect 24780 43790 24808 43930
rect 24768 43784 24820 43790
rect 24674 43752 24730 43761
rect 24768 43726 24820 43732
rect 24674 43687 24730 43696
rect 24872 42566 24900 45886
rect 25056 44010 25084 46106
rect 24964 43982 25084 44010
rect 24492 42560 24544 42566
rect 24492 42502 24544 42508
rect 24584 42560 24636 42566
rect 24584 42502 24636 42508
rect 24860 42560 24912 42566
rect 24860 42502 24912 42508
rect 24504 42294 24532 42502
rect 24492 42288 24544 42294
rect 24492 42230 24544 42236
rect 24676 42288 24728 42294
rect 24676 42230 24728 42236
rect 24400 41744 24452 41750
rect 24400 41686 24452 41692
rect 24412 41414 24440 41686
rect 24412 41386 24624 41414
rect 24216 41200 24268 41206
rect 24216 41142 24268 41148
rect 24124 41064 24176 41070
rect 24124 41006 24176 41012
rect 24032 39296 24084 39302
rect 24032 39238 24084 39244
rect 23768 38270 23980 38298
rect 23756 38208 23808 38214
rect 23756 38150 23808 38156
rect 23662 37224 23718 37233
rect 23662 37159 23718 37168
rect 23768 36242 23796 38150
rect 23848 37800 23900 37806
rect 23848 37742 23900 37748
rect 23860 37466 23888 37742
rect 23848 37460 23900 37466
rect 23848 37402 23900 37408
rect 23848 37120 23900 37126
rect 23848 37062 23900 37068
rect 23860 36922 23888 37062
rect 23848 36916 23900 36922
rect 23848 36858 23900 36864
rect 23952 36825 23980 38270
rect 23938 36816 23994 36825
rect 23938 36751 23994 36760
rect 23848 36304 23900 36310
rect 23848 36246 23900 36252
rect 23756 36236 23808 36242
rect 23756 36178 23808 36184
rect 23664 36032 23716 36038
rect 23664 35974 23716 35980
rect 23676 35290 23704 35974
rect 23860 35630 23888 36246
rect 23848 35624 23900 35630
rect 24044 35578 24072 39238
rect 24136 37806 24164 41006
rect 24228 40662 24256 41142
rect 24216 40656 24268 40662
rect 24268 40616 24348 40644
rect 24216 40598 24268 40604
rect 24216 40384 24268 40390
rect 24216 40326 24268 40332
rect 24228 39982 24256 40326
rect 24216 39976 24268 39982
rect 24216 39918 24268 39924
rect 24320 39030 24348 40616
rect 24596 40050 24624 41386
rect 24584 40044 24636 40050
rect 24584 39986 24636 39992
rect 24688 39506 24716 42230
rect 24768 41608 24820 41614
rect 24768 41550 24820 41556
rect 24780 41041 24808 41550
rect 24766 41032 24822 41041
rect 24766 40967 24822 40976
rect 24780 40662 24808 40967
rect 24768 40656 24820 40662
rect 24768 40598 24820 40604
rect 24768 40384 24820 40390
rect 24768 40326 24820 40332
rect 24676 39500 24728 39506
rect 24676 39442 24728 39448
rect 24676 39296 24728 39302
rect 24676 39238 24728 39244
rect 24308 39024 24360 39030
rect 24308 38966 24360 38972
rect 24492 38208 24544 38214
rect 24492 38150 24544 38156
rect 24124 37800 24176 37806
rect 24124 37742 24176 37748
rect 24504 37738 24532 38150
rect 24492 37732 24544 37738
rect 24492 37674 24544 37680
rect 24504 37618 24532 37674
rect 24412 37590 24532 37618
rect 24412 37330 24440 37590
rect 24400 37324 24452 37330
rect 24400 37266 24452 37272
rect 24124 37120 24176 37126
rect 24124 37062 24176 37068
rect 23848 35566 23900 35572
rect 23952 35550 24072 35578
rect 23952 35494 23980 35550
rect 23940 35488 23992 35494
rect 23940 35430 23992 35436
rect 23664 35284 23716 35290
rect 23664 35226 23716 35232
rect 24136 35222 24164 37062
rect 24412 36854 24440 37266
rect 24400 36848 24452 36854
rect 24400 36790 24452 36796
rect 24412 35766 24440 36790
rect 24492 36576 24544 36582
rect 24492 36518 24544 36524
rect 24504 36378 24532 36518
rect 24492 36372 24544 36378
rect 24492 36314 24544 36320
rect 24584 36032 24636 36038
rect 24584 35974 24636 35980
rect 24400 35760 24452 35766
rect 24400 35702 24452 35708
rect 24124 35216 24176 35222
rect 24124 35158 24176 35164
rect 24412 34950 24440 35702
rect 24400 34944 24452 34950
rect 24400 34886 24452 34892
rect 23664 34536 23716 34542
rect 23664 34478 23716 34484
rect 23572 33992 23624 33998
rect 23572 33934 23624 33940
rect 23480 33516 23532 33522
rect 23480 33458 23532 33464
rect 23296 33380 23348 33386
rect 23296 33322 23348 33328
rect 22950 33212 23258 33221
rect 22950 33210 22956 33212
rect 23012 33210 23036 33212
rect 23092 33210 23116 33212
rect 23172 33210 23196 33212
rect 23252 33210 23258 33212
rect 23012 33158 23014 33210
rect 23194 33158 23196 33210
rect 22950 33156 22956 33158
rect 23012 33156 23036 33158
rect 23092 33156 23116 33158
rect 23172 33156 23196 33158
rect 23252 33156 23258 33158
rect 22950 33147 23258 33156
rect 23112 33108 23164 33114
rect 22848 33068 22968 33096
rect 22836 32972 22888 32978
rect 22836 32914 22888 32920
rect 22744 31952 22796 31958
rect 22848 31940 22876 32914
rect 22940 32502 22968 33068
rect 23112 33050 23164 33056
rect 23124 32774 23152 33050
rect 23308 32910 23336 33322
rect 23676 33096 23704 34478
rect 24400 33856 24452 33862
rect 24400 33798 24452 33804
rect 23756 33448 23808 33454
rect 23756 33390 23808 33396
rect 23492 33068 23704 33096
rect 23296 32904 23348 32910
rect 23296 32846 23348 32852
rect 23204 32836 23256 32842
rect 23204 32778 23256 32784
rect 23112 32768 23164 32774
rect 23112 32710 23164 32716
rect 22928 32496 22980 32502
rect 22928 32438 22980 32444
rect 23216 32366 23244 32778
rect 23296 32428 23348 32434
rect 23296 32370 23348 32376
rect 23204 32360 23256 32366
rect 23204 32302 23256 32308
rect 22950 32124 23258 32133
rect 22950 32122 22956 32124
rect 23012 32122 23036 32124
rect 23092 32122 23116 32124
rect 23172 32122 23196 32124
rect 23252 32122 23258 32124
rect 23012 32070 23014 32122
rect 23194 32070 23196 32122
rect 22950 32068 22956 32070
rect 23012 32068 23036 32070
rect 23092 32068 23116 32070
rect 23172 32068 23196 32070
rect 23252 32068 23258 32070
rect 22950 32059 23258 32068
rect 22848 31912 22968 31940
rect 22744 31894 22796 31900
rect 22744 31816 22796 31822
rect 22744 31758 22796 31764
rect 22756 29714 22784 31758
rect 22940 31124 22968 31912
rect 23308 31890 23336 32370
rect 23388 31952 23440 31958
rect 23388 31894 23440 31900
rect 23296 31884 23348 31890
rect 23296 31826 23348 31832
rect 23296 31476 23348 31482
rect 23296 31418 23348 31424
rect 22848 31096 22968 31124
rect 22848 30190 22876 31096
rect 22950 31036 23258 31045
rect 22950 31034 22956 31036
rect 23012 31034 23036 31036
rect 23092 31034 23116 31036
rect 23172 31034 23196 31036
rect 23252 31034 23258 31036
rect 23012 30982 23014 31034
rect 23194 30982 23196 31034
rect 22950 30980 22956 30982
rect 23012 30980 23036 30982
rect 23092 30980 23116 30982
rect 23172 30980 23196 30982
rect 23252 30980 23258 30982
rect 22950 30971 23258 30980
rect 22836 30184 22888 30190
rect 22836 30126 22888 30132
rect 22744 29708 22796 29714
rect 22744 29650 22796 29656
rect 22744 29504 22796 29510
rect 22744 29446 22796 29452
rect 22652 28212 22704 28218
rect 22652 28154 22704 28160
rect 22468 25968 22520 25974
rect 22468 25910 22520 25916
rect 22652 25968 22704 25974
rect 22652 25910 22704 25916
rect 22284 25900 22336 25906
rect 22284 25842 22336 25848
rect 22560 25832 22612 25838
rect 22560 25774 22612 25780
rect 22284 25764 22336 25770
rect 22284 25706 22336 25712
rect 22008 25356 22060 25362
rect 22008 25298 22060 25304
rect 22020 25242 22048 25298
rect 22020 25214 22232 25242
rect 21732 25152 21784 25158
rect 21732 25094 21784 25100
rect 22100 24744 22152 24750
rect 22100 24686 22152 24692
rect 21916 23112 21968 23118
rect 21916 23054 21968 23060
rect 21640 22704 21692 22710
rect 21640 22646 21692 22652
rect 21928 22574 21956 23054
rect 21916 22568 21968 22574
rect 21916 22510 21968 22516
rect 21640 22500 21692 22506
rect 21640 22442 21692 22448
rect 21652 21622 21680 22442
rect 22112 22166 22140 24686
rect 22204 24682 22232 25214
rect 22192 24676 22244 24682
rect 22192 24618 22244 24624
rect 22192 22772 22244 22778
rect 22192 22714 22244 22720
rect 22100 22160 22152 22166
rect 22100 22102 22152 22108
rect 21640 21616 21692 21622
rect 21640 21558 21692 21564
rect 22100 21548 22152 21554
rect 22100 21490 22152 21496
rect 22112 21010 22140 21490
rect 22204 21078 22232 22714
rect 22192 21072 22244 21078
rect 22192 21014 22244 21020
rect 22100 21004 22152 21010
rect 22100 20946 22152 20952
rect 21824 20936 21876 20942
rect 21824 20878 21876 20884
rect 21836 20602 21864 20878
rect 21824 20596 21876 20602
rect 21824 20538 21876 20544
rect 21732 19712 21784 19718
rect 21732 19654 21784 19660
rect 21548 18760 21600 18766
rect 21548 18702 21600 18708
rect 21456 18624 21508 18630
rect 21456 18566 21508 18572
rect 20720 17604 20772 17610
rect 20720 17546 20772 17552
rect 20732 17270 20760 17546
rect 21180 17536 21232 17542
rect 21180 17478 21232 17484
rect 20720 17264 20772 17270
rect 20720 17206 20772 17212
rect 20732 17134 20760 17206
rect 21192 17134 21220 17478
rect 20720 17128 20772 17134
rect 20720 17070 20772 17076
rect 21180 17128 21232 17134
rect 21180 17070 21232 17076
rect 21192 16658 21220 17070
rect 21180 16652 21232 16658
rect 21180 16594 21232 16600
rect 21364 16448 21416 16454
rect 21364 16390 21416 16396
rect 20996 15360 21048 15366
rect 20996 15302 21048 15308
rect 20628 15020 20680 15026
rect 20628 14962 20680 14968
rect 20352 14816 20404 14822
rect 20352 14758 20404 14764
rect 19996 12406 20116 12434
rect 19996 12374 20024 12406
rect 19984 12368 20036 12374
rect 19984 12310 20036 12316
rect 20364 11626 20392 14758
rect 21008 14074 21036 15302
rect 21272 14816 21324 14822
rect 21272 14758 21324 14764
rect 20996 14068 21048 14074
rect 20996 14010 21048 14016
rect 20904 13796 20956 13802
rect 20904 13738 20956 13744
rect 20916 13190 20944 13738
rect 21088 13524 21140 13530
rect 21088 13466 21140 13472
rect 20904 13184 20956 13190
rect 20904 13126 20956 13132
rect 20916 12918 20944 13126
rect 20904 12912 20956 12918
rect 20904 12854 20956 12860
rect 19984 11620 20036 11626
rect 19984 11562 20036 11568
rect 20352 11620 20404 11626
rect 20352 11562 20404 11568
rect 19892 10056 19944 10062
rect 19892 9998 19944 10004
rect 19800 6792 19852 6798
rect 19800 6734 19852 6740
rect 19708 6724 19760 6730
rect 19708 6666 19760 6672
rect 19720 5234 19748 6666
rect 19996 5710 20024 11562
rect 21100 10674 21128 13466
rect 21180 13456 21232 13462
rect 21180 13398 21232 13404
rect 21088 10668 21140 10674
rect 21088 10610 21140 10616
rect 20720 8900 20772 8906
rect 20720 8842 20772 8848
rect 20260 7812 20312 7818
rect 20260 7754 20312 7760
rect 20168 6316 20220 6322
rect 20168 6258 20220 6264
rect 20180 5914 20208 6258
rect 20168 5908 20220 5914
rect 20168 5850 20220 5856
rect 20272 5846 20300 7754
rect 20260 5840 20312 5846
rect 20260 5782 20312 5788
rect 20628 5772 20680 5778
rect 20628 5714 20680 5720
rect 19984 5704 20036 5710
rect 19984 5646 20036 5652
rect 19800 5296 19852 5302
rect 19800 5238 19852 5244
rect 19432 5228 19484 5234
rect 19432 5170 19484 5176
rect 19708 5228 19760 5234
rect 19708 5170 19760 5176
rect 19524 5160 19576 5166
rect 19524 5102 19576 5108
rect 19340 4616 19392 4622
rect 19340 4558 19392 4564
rect 19156 3460 19208 3466
rect 19156 3402 19208 3408
rect 18972 2576 19024 2582
rect 18972 2518 19024 2524
rect 19168 800 19196 3402
rect 19536 800 19564 5102
rect 19812 3670 19840 5238
rect 20536 5092 20588 5098
rect 20536 5034 20588 5040
rect 19892 4684 19944 4690
rect 19892 4626 19944 4632
rect 19800 3664 19852 3670
rect 19800 3606 19852 3612
rect 19904 2854 19932 4626
rect 20260 4072 20312 4078
rect 20260 4014 20312 4020
rect 19984 2916 20036 2922
rect 19984 2858 20036 2864
rect 19892 2848 19944 2854
rect 19892 2790 19944 2796
rect 19996 2258 20024 2858
rect 19904 2230 20024 2258
rect 19904 800 19932 2230
rect 20272 800 20300 4014
rect 20548 2990 20576 5034
rect 20536 2984 20588 2990
rect 20536 2926 20588 2932
rect 20640 800 20668 5714
rect 20732 5710 20760 8842
rect 21088 7812 21140 7818
rect 21088 7754 21140 7760
rect 20996 7336 21048 7342
rect 20996 7278 21048 7284
rect 20720 5704 20772 5710
rect 20720 5646 20772 5652
rect 21008 3942 21036 7278
rect 20996 3936 21048 3942
rect 20996 3878 21048 3884
rect 21100 3534 21128 7754
rect 21192 4622 21220 13398
rect 21284 7886 21312 14758
rect 21376 13870 21404 16390
rect 21468 14414 21496 18566
rect 21548 17128 21600 17134
rect 21548 17070 21600 17076
rect 21560 16794 21588 17070
rect 21548 16788 21600 16794
rect 21548 16730 21600 16736
rect 21456 14408 21508 14414
rect 21456 14350 21508 14356
rect 21364 13864 21416 13870
rect 21364 13806 21416 13812
rect 21364 13728 21416 13734
rect 21364 13670 21416 13676
rect 21376 13190 21404 13670
rect 21560 13394 21588 16730
rect 21640 16448 21692 16454
rect 21640 16390 21692 16396
rect 21652 15609 21680 16390
rect 21638 15600 21694 15609
rect 21638 15535 21694 15544
rect 21548 13388 21600 13394
rect 21548 13330 21600 13336
rect 21364 13184 21416 13190
rect 21364 13126 21416 13132
rect 21376 12986 21404 13126
rect 21364 12980 21416 12986
rect 21364 12922 21416 12928
rect 21376 12102 21404 12922
rect 21456 12776 21508 12782
rect 21560 12764 21588 13330
rect 21652 13190 21680 15535
rect 21744 14346 21772 19654
rect 22100 19440 22152 19446
rect 22100 19382 22152 19388
rect 22112 19281 22140 19382
rect 22296 19378 22324 25706
rect 22376 23316 22428 23322
rect 22376 23258 22428 23264
rect 22388 22642 22416 23258
rect 22376 22636 22428 22642
rect 22376 22578 22428 22584
rect 22388 22234 22416 22578
rect 22376 22228 22428 22234
rect 22376 22170 22428 22176
rect 22376 21956 22428 21962
rect 22376 21898 22428 21904
rect 22388 20602 22416 21898
rect 22376 20596 22428 20602
rect 22376 20538 22428 20544
rect 22284 19372 22336 19378
rect 22284 19314 22336 19320
rect 22098 19272 22154 19281
rect 22098 19207 22154 19216
rect 22572 18970 22600 25774
rect 22664 25226 22692 25910
rect 22652 25220 22704 25226
rect 22652 25162 22704 25168
rect 22756 24954 22784 29446
rect 22848 27402 22876 30126
rect 22950 29948 23258 29957
rect 22950 29946 22956 29948
rect 23012 29946 23036 29948
rect 23092 29946 23116 29948
rect 23172 29946 23196 29948
rect 23252 29946 23258 29948
rect 23012 29894 23014 29946
rect 23194 29894 23196 29946
rect 22950 29892 22956 29894
rect 23012 29892 23036 29894
rect 23092 29892 23116 29894
rect 23172 29892 23196 29894
rect 23252 29892 23258 29894
rect 22950 29883 23258 29892
rect 22950 28860 23258 28869
rect 22950 28858 22956 28860
rect 23012 28858 23036 28860
rect 23092 28858 23116 28860
rect 23172 28858 23196 28860
rect 23252 28858 23258 28860
rect 23012 28806 23014 28858
rect 23194 28806 23196 28858
rect 22950 28804 22956 28806
rect 23012 28804 23036 28806
rect 23092 28804 23116 28806
rect 23172 28804 23196 28806
rect 23252 28804 23258 28806
rect 22950 28795 23258 28804
rect 22950 27772 23258 27781
rect 22950 27770 22956 27772
rect 23012 27770 23036 27772
rect 23092 27770 23116 27772
rect 23172 27770 23196 27772
rect 23252 27770 23258 27772
rect 23012 27718 23014 27770
rect 23194 27718 23196 27770
rect 22950 27716 22956 27718
rect 23012 27716 23036 27718
rect 23092 27716 23116 27718
rect 23172 27716 23196 27718
rect 23252 27716 23258 27718
rect 22950 27707 23258 27716
rect 23308 27418 23336 31418
rect 23400 31346 23428 31894
rect 23388 31340 23440 31346
rect 23388 31282 23440 31288
rect 23492 30598 23520 33068
rect 23664 32768 23716 32774
rect 23664 32710 23716 32716
rect 23480 30592 23532 30598
rect 23480 30534 23532 30540
rect 23572 30592 23624 30598
rect 23572 30534 23624 30540
rect 23584 30258 23612 30534
rect 23676 30326 23704 32710
rect 23664 30320 23716 30326
rect 23664 30262 23716 30268
rect 23572 30252 23624 30258
rect 23572 30194 23624 30200
rect 23388 30048 23440 30054
rect 23388 29990 23440 29996
rect 23400 29714 23428 29990
rect 23388 29708 23440 29714
rect 23388 29650 23440 29656
rect 23676 29646 23704 30262
rect 23768 30190 23796 33390
rect 23940 32224 23992 32230
rect 23940 32166 23992 32172
rect 23952 31754 23980 32166
rect 23952 31726 24072 31754
rect 23756 30184 23808 30190
rect 23756 30126 23808 30132
rect 23768 29782 23796 30126
rect 23756 29776 23808 29782
rect 23756 29718 23808 29724
rect 23664 29640 23716 29646
rect 23664 29582 23716 29588
rect 23572 29504 23624 29510
rect 23572 29446 23624 29452
rect 23940 29504 23992 29510
rect 23940 29446 23992 29452
rect 23584 28762 23612 29446
rect 23572 28756 23624 28762
rect 23572 28698 23624 28704
rect 23952 28082 23980 29446
rect 23940 28076 23992 28082
rect 23940 28018 23992 28024
rect 23940 27940 23992 27946
rect 23940 27882 23992 27888
rect 23952 27606 23980 27882
rect 23940 27600 23992 27606
rect 23860 27548 23940 27554
rect 23860 27542 23992 27548
rect 23572 27532 23624 27538
rect 23572 27474 23624 27480
rect 23860 27526 23980 27542
rect 22836 27396 22888 27402
rect 23308 27390 23428 27418
rect 22836 27338 22888 27344
rect 23296 27328 23348 27334
rect 23296 27270 23348 27276
rect 22950 26684 23258 26693
rect 22950 26682 22956 26684
rect 23012 26682 23036 26684
rect 23092 26682 23116 26684
rect 23172 26682 23196 26684
rect 23252 26682 23258 26684
rect 23012 26630 23014 26682
rect 23194 26630 23196 26682
rect 22950 26628 22956 26630
rect 23012 26628 23036 26630
rect 23092 26628 23116 26630
rect 23172 26628 23196 26630
rect 23252 26628 23258 26630
rect 22950 26619 23258 26628
rect 23308 26586 23336 27270
rect 22836 26580 22888 26586
rect 22836 26522 22888 26528
rect 23296 26580 23348 26586
rect 23296 26522 23348 26528
rect 22848 25362 22876 26522
rect 23112 26308 23164 26314
rect 23112 26250 23164 26256
rect 23124 25974 23152 26250
rect 23400 26042 23428 27390
rect 23584 27334 23612 27474
rect 23572 27328 23624 27334
rect 23572 27270 23624 27276
rect 23584 27062 23612 27270
rect 23572 27056 23624 27062
rect 23572 26998 23624 27004
rect 23584 26314 23612 26998
rect 23572 26308 23624 26314
rect 23572 26250 23624 26256
rect 23570 26208 23626 26217
rect 23570 26143 23626 26152
rect 23388 26036 23440 26042
rect 23388 25978 23440 25984
rect 23112 25968 23164 25974
rect 23112 25910 23164 25916
rect 23296 25764 23348 25770
rect 23296 25706 23348 25712
rect 22950 25596 23258 25605
rect 22950 25594 22956 25596
rect 23012 25594 23036 25596
rect 23092 25594 23116 25596
rect 23172 25594 23196 25596
rect 23252 25594 23258 25596
rect 23012 25542 23014 25594
rect 23194 25542 23196 25594
rect 22950 25540 22956 25542
rect 23012 25540 23036 25542
rect 23092 25540 23116 25542
rect 23172 25540 23196 25542
rect 23252 25540 23258 25542
rect 22950 25531 23258 25540
rect 22836 25356 22888 25362
rect 22836 25298 22888 25304
rect 22744 24948 22796 24954
rect 22744 24890 22796 24896
rect 22836 24676 22888 24682
rect 22836 24618 22888 24624
rect 22744 24608 22796 24614
rect 22744 24550 22796 24556
rect 22756 20602 22784 24550
rect 22848 22642 22876 24618
rect 22950 24508 23258 24517
rect 22950 24506 22956 24508
rect 23012 24506 23036 24508
rect 23092 24506 23116 24508
rect 23172 24506 23196 24508
rect 23252 24506 23258 24508
rect 23012 24454 23014 24506
rect 23194 24454 23196 24506
rect 22950 24452 22956 24454
rect 23012 24452 23036 24454
rect 23092 24452 23116 24454
rect 23172 24452 23196 24454
rect 23252 24452 23258 24454
rect 22950 24443 23258 24452
rect 22950 23420 23258 23429
rect 22950 23418 22956 23420
rect 23012 23418 23036 23420
rect 23092 23418 23116 23420
rect 23172 23418 23196 23420
rect 23252 23418 23258 23420
rect 23012 23366 23014 23418
rect 23194 23366 23196 23418
rect 22950 23364 22956 23366
rect 23012 23364 23036 23366
rect 23092 23364 23116 23366
rect 23172 23364 23196 23366
rect 23252 23364 23258 23366
rect 22950 23355 23258 23364
rect 22836 22636 22888 22642
rect 22836 22578 22888 22584
rect 22848 22098 22876 22578
rect 22950 22332 23258 22341
rect 22950 22330 22956 22332
rect 23012 22330 23036 22332
rect 23092 22330 23116 22332
rect 23172 22330 23196 22332
rect 23252 22330 23258 22332
rect 23012 22278 23014 22330
rect 23194 22278 23196 22330
rect 22950 22276 22956 22278
rect 23012 22276 23036 22278
rect 23092 22276 23116 22278
rect 23172 22276 23196 22278
rect 23252 22276 23258 22278
rect 22950 22267 23258 22276
rect 22836 22092 22888 22098
rect 23308 22094 23336 25706
rect 23400 25294 23428 25978
rect 23584 25974 23612 26143
rect 23572 25968 23624 25974
rect 23572 25910 23624 25916
rect 23860 25498 23888 27526
rect 23940 27396 23992 27402
rect 23940 27338 23992 27344
rect 23480 25492 23532 25498
rect 23480 25434 23532 25440
rect 23848 25492 23900 25498
rect 23848 25434 23900 25440
rect 23388 25288 23440 25294
rect 23388 25230 23440 25236
rect 23492 24750 23520 25434
rect 23480 24744 23532 24750
rect 23480 24686 23532 24692
rect 23952 23730 23980 27338
rect 24044 25974 24072 31726
rect 24308 31204 24360 31210
rect 24308 31146 24360 31152
rect 24124 29164 24176 29170
rect 24124 29106 24176 29112
rect 24136 28801 24164 29106
rect 24122 28792 24178 28801
rect 24122 28727 24178 28736
rect 24216 27940 24268 27946
rect 24216 27882 24268 27888
rect 24124 27872 24176 27878
rect 24124 27814 24176 27820
rect 24032 25968 24084 25974
rect 24032 25910 24084 25916
rect 24136 25294 24164 27814
rect 24124 25288 24176 25294
rect 24124 25230 24176 25236
rect 24124 25152 24176 25158
rect 24124 25094 24176 25100
rect 24136 23730 24164 25094
rect 23940 23724 23992 23730
rect 23940 23666 23992 23672
rect 24124 23724 24176 23730
rect 24124 23666 24176 23672
rect 23388 23656 23440 23662
rect 23388 23598 23440 23604
rect 23400 23361 23428 23598
rect 23386 23352 23442 23361
rect 23386 23287 23442 23296
rect 23940 22432 23992 22438
rect 23940 22374 23992 22380
rect 23308 22066 23428 22094
rect 22836 22034 22888 22040
rect 22848 21554 22876 22034
rect 22836 21548 22888 21554
rect 22836 21490 22888 21496
rect 22848 21350 22876 21490
rect 22836 21344 22888 21350
rect 22836 21286 22888 21292
rect 22950 21244 23258 21253
rect 22950 21242 22956 21244
rect 23012 21242 23036 21244
rect 23092 21242 23116 21244
rect 23172 21242 23196 21244
rect 23252 21242 23258 21244
rect 23012 21190 23014 21242
rect 23194 21190 23196 21242
rect 22950 21188 22956 21190
rect 23012 21188 23036 21190
rect 23092 21188 23116 21190
rect 23172 21188 23196 21190
rect 23252 21188 23258 21190
rect 22950 21179 23258 21188
rect 22744 20596 22796 20602
rect 22744 20538 22796 20544
rect 22950 20156 23258 20165
rect 22950 20154 22956 20156
rect 23012 20154 23036 20156
rect 23092 20154 23116 20156
rect 23172 20154 23196 20156
rect 23252 20154 23258 20156
rect 23012 20102 23014 20154
rect 23194 20102 23196 20154
rect 22950 20100 22956 20102
rect 23012 20100 23036 20102
rect 23092 20100 23116 20102
rect 23172 20100 23196 20102
rect 23252 20100 23258 20102
rect 22950 20091 23258 20100
rect 22652 19780 22704 19786
rect 22652 19722 22704 19728
rect 22560 18964 22612 18970
rect 22560 18906 22612 18912
rect 22560 18624 22612 18630
rect 22560 18566 22612 18572
rect 21824 18420 21876 18426
rect 21824 18362 21876 18368
rect 21836 18086 21864 18362
rect 22008 18284 22060 18290
rect 22008 18226 22060 18232
rect 21824 18080 21876 18086
rect 21824 18022 21876 18028
rect 21836 17542 21864 18022
rect 22020 17746 22048 18226
rect 22008 17740 22060 17746
rect 22008 17682 22060 17688
rect 21824 17536 21876 17542
rect 21876 17484 21956 17490
rect 21824 17478 21956 17484
rect 21836 17462 21956 17478
rect 21928 17270 21956 17462
rect 21916 17264 21968 17270
rect 21916 17206 21968 17212
rect 21928 16538 21956 17206
rect 22020 17134 22048 17682
rect 22100 17604 22152 17610
rect 22100 17546 22152 17552
rect 22008 17128 22060 17134
rect 22008 17070 22060 17076
rect 22008 16584 22060 16590
rect 21928 16532 22008 16538
rect 21928 16526 22060 16532
rect 21928 16510 22048 16526
rect 21824 16448 21876 16454
rect 21824 16390 21876 16396
rect 21836 15502 21864 16390
rect 21824 15496 21876 15502
rect 21824 15438 21876 15444
rect 21732 14340 21784 14346
rect 21732 14282 21784 14288
rect 21928 14226 21956 16510
rect 22008 15428 22060 15434
rect 22008 15370 22060 15376
rect 21744 14198 21956 14226
rect 21744 13734 21772 14198
rect 21916 14068 21968 14074
rect 21916 14010 21968 14016
rect 21824 13932 21876 13938
rect 21824 13874 21876 13880
rect 21732 13728 21784 13734
rect 21732 13670 21784 13676
rect 21640 13184 21692 13190
rect 21640 13126 21692 13132
rect 21508 12736 21588 12764
rect 21456 12718 21508 12724
rect 21364 12096 21416 12102
rect 21364 12038 21416 12044
rect 21376 10538 21404 12038
rect 21468 10606 21496 12718
rect 21456 10600 21508 10606
rect 21456 10542 21508 10548
rect 21364 10532 21416 10538
rect 21364 10474 21416 10480
rect 21272 7880 21324 7886
rect 21272 7822 21324 7828
rect 21376 6914 21404 10474
rect 21548 7404 21600 7410
rect 21548 7346 21600 7352
rect 21376 6886 21496 6914
rect 21180 4616 21232 4622
rect 21180 4558 21232 4564
rect 21364 4004 21416 4010
rect 21364 3946 21416 3952
rect 21088 3528 21140 3534
rect 21088 3470 21140 3476
rect 20996 2848 21048 2854
rect 20996 2790 21048 2796
rect 21008 800 21036 2790
rect 21376 800 21404 3946
rect 21468 3398 21496 6886
rect 21560 6458 21588 7346
rect 21548 6452 21600 6458
rect 21548 6394 21600 6400
rect 21732 4684 21784 4690
rect 21732 4626 21784 4632
rect 21456 3392 21508 3398
rect 21456 3334 21508 3340
rect 21744 2922 21772 4626
rect 21836 4214 21864 13874
rect 21928 11150 21956 14010
rect 22020 13938 22048 15370
rect 22112 15026 22140 17546
rect 22572 16658 22600 18566
rect 22560 16652 22612 16658
rect 22560 16594 22612 16600
rect 22664 15502 22692 19722
rect 23400 19378 23428 22066
rect 23756 20868 23808 20874
rect 23756 20810 23808 20816
rect 23388 19372 23440 19378
rect 23388 19314 23440 19320
rect 22950 19068 23258 19077
rect 22950 19066 22956 19068
rect 23012 19066 23036 19068
rect 23092 19066 23116 19068
rect 23172 19066 23196 19068
rect 23252 19066 23258 19068
rect 23012 19014 23014 19066
rect 23194 19014 23196 19066
rect 22950 19012 22956 19014
rect 23012 19012 23036 19014
rect 23092 19012 23116 19014
rect 23172 19012 23196 19014
rect 23252 19012 23258 19014
rect 22950 19003 23258 19012
rect 23204 18964 23256 18970
rect 23204 18906 23256 18912
rect 22836 18828 22888 18834
rect 22836 18770 22888 18776
rect 22744 18624 22796 18630
rect 22744 18566 22796 18572
rect 22756 18426 22784 18566
rect 22744 18420 22796 18426
rect 22744 18362 22796 18368
rect 22848 18358 22876 18770
rect 23216 18426 23244 18906
rect 23664 18692 23716 18698
rect 23664 18634 23716 18640
rect 23386 18592 23442 18601
rect 23386 18527 23442 18536
rect 22928 18420 22980 18426
rect 22928 18362 22980 18368
rect 23204 18420 23256 18426
rect 23204 18362 23256 18368
rect 22836 18352 22888 18358
rect 22836 18294 22888 18300
rect 22940 18170 22968 18362
rect 22848 18142 22968 18170
rect 23296 18216 23348 18222
rect 23296 18158 23348 18164
rect 22652 15496 22704 15502
rect 22652 15438 22704 15444
rect 22100 15020 22152 15026
rect 22100 14962 22152 14968
rect 22848 14958 22876 18142
rect 22950 17980 23258 17989
rect 22950 17978 22956 17980
rect 23012 17978 23036 17980
rect 23092 17978 23116 17980
rect 23172 17978 23196 17980
rect 23252 17978 23258 17980
rect 23012 17926 23014 17978
rect 23194 17926 23196 17978
rect 22950 17924 22956 17926
rect 23012 17924 23036 17926
rect 23092 17924 23116 17926
rect 23172 17924 23196 17926
rect 23252 17924 23258 17926
rect 22950 17915 23258 17924
rect 23308 17338 23336 18158
rect 23400 17746 23428 18527
rect 23388 17740 23440 17746
rect 23388 17682 23440 17688
rect 23296 17332 23348 17338
rect 23296 17274 23348 17280
rect 22950 16892 23258 16901
rect 22950 16890 22956 16892
rect 23012 16890 23036 16892
rect 23092 16890 23116 16892
rect 23172 16890 23196 16892
rect 23252 16890 23258 16892
rect 23012 16838 23014 16890
rect 23194 16838 23196 16890
rect 22950 16836 22956 16838
rect 23012 16836 23036 16838
rect 23092 16836 23116 16838
rect 23172 16836 23196 16838
rect 23252 16836 23258 16838
rect 22950 16827 23258 16836
rect 22950 15804 23258 15813
rect 22950 15802 22956 15804
rect 23012 15802 23036 15804
rect 23092 15802 23116 15804
rect 23172 15802 23196 15804
rect 23252 15802 23258 15804
rect 23012 15750 23014 15802
rect 23194 15750 23196 15802
rect 22950 15748 22956 15750
rect 23012 15748 23036 15750
rect 23092 15748 23116 15750
rect 23172 15748 23196 15750
rect 23252 15748 23258 15750
rect 22950 15739 23258 15748
rect 23308 15570 23336 17274
rect 23676 16114 23704 18634
rect 23664 16108 23716 16114
rect 23664 16050 23716 16056
rect 23664 15904 23716 15910
rect 23664 15846 23716 15852
rect 23296 15564 23348 15570
rect 23296 15506 23348 15512
rect 23296 15360 23348 15366
rect 23296 15302 23348 15308
rect 22836 14952 22888 14958
rect 22836 14894 22888 14900
rect 22950 14716 23258 14725
rect 22950 14714 22956 14716
rect 23012 14714 23036 14716
rect 23092 14714 23116 14716
rect 23172 14714 23196 14716
rect 23252 14714 23258 14716
rect 23012 14662 23014 14714
rect 23194 14662 23196 14714
rect 22950 14660 22956 14662
rect 23012 14660 23036 14662
rect 23092 14660 23116 14662
rect 23172 14660 23196 14662
rect 23252 14660 23258 14662
rect 22950 14651 23258 14660
rect 22928 14340 22980 14346
rect 22928 14282 22980 14288
rect 22560 14272 22612 14278
rect 22560 14214 22612 14220
rect 22008 13932 22060 13938
rect 22008 13874 22060 13880
rect 22100 12844 22152 12850
rect 22100 12786 22152 12792
rect 22112 12442 22140 12786
rect 22100 12436 22152 12442
rect 22100 12378 22152 12384
rect 22468 11756 22520 11762
rect 22468 11698 22520 11704
rect 22480 11354 22508 11698
rect 22468 11348 22520 11354
rect 22468 11290 22520 11296
rect 22008 11280 22060 11286
rect 22008 11222 22060 11228
rect 21916 11144 21968 11150
rect 21916 11086 21968 11092
rect 22020 9586 22048 11222
rect 22572 11218 22600 14214
rect 22744 14068 22796 14074
rect 22744 14010 22796 14016
rect 22756 12238 22784 14010
rect 22836 14000 22888 14006
rect 22836 13942 22888 13948
rect 22848 13394 22876 13942
rect 22940 13938 22968 14282
rect 22928 13932 22980 13938
rect 22928 13874 22980 13880
rect 22950 13628 23258 13637
rect 22950 13626 22956 13628
rect 23012 13626 23036 13628
rect 23092 13626 23116 13628
rect 23172 13626 23196 13628
rect 23252 13626 23258 13628
rect 23012 13574 23014 13626
rect 23194 13574 23196 13626
rect 22950 13572 22956 13574
rect 23012 13572 23036 13574
rect 23092 13572 23116 13574
rect 23172 13572 23196 13574
rect 23252 13572 23258 13574
rect 22950 13563 23258 13572
rect 22836 13388 22888 13394
rect 22836 13330 22888 13336
rect 23308 13326 23336 15302
rect 23388 13864 23440 13870
rect 23388 13806 23440 13812
rect 23296 13320 23348 13326
rect 23296 13262 23348 13268
rect 22950 12540 23258 12549
rect 22950 12538 22956 12540
rect 23012 12538 23036 12540
rect 23092 12538 23116 12540
rect 23172 12538 23196 12540
rect 23252 12538 23258 12540
rect 23012 12486 23014 12538
rect 23194 12486 23196 12538
rect 22950 12484 22956 12486
rect 23012 12484 23036 12486
rect 23092 12484 23116 12486
rect 23172 12484 23196 12486
rect 23252 12484 23258 12486
rect 22950 12475 23258 12484
rect 22652 12232 22704 12238
rect 22652 12174 22704 12180
rect 22744 12232 22796 12238
rect 22744 12174 22796 12180
rect 22664 11898 22692 12174
rect 22652 11892 22704 11898
rect 22652 11834 22704 11840
rect 22950 11452 23258 11461
rect 22950 11450 22956 11452
rect 23012 11450 23036 11452
rect 23092 11450 23116 11452
rect 23172 11450 23196 11452
rect 23252 11450 23258 11452
rect 23012 11398 23014 11450
rect 23194 11398 23196 11450
rect 22950 11396 22956 11398
rect 23012 11396 23036 11398
rect 23092 11396 23116 11398
rect 23172 11396 23196 11398
rect 23252 11396 23258 11398
rect 22950 11387 23258 11396
rect 22836 11280 22888 11286
rect 22836 11222 22888 11228
rect 22560 11212 22612 11218
rect 22560 11154 22612 11160
rect 22008 9580 22060 9586
rect 22008 9522 22060 9528
rect 22848 8974 22876 11222
rect 23400 11150 23428 13806
rect 23676 11762 23704 15846
rect 23768 15026 23796 20810
rect 23952 16114 23980 22374
rect 24228 22030 24256 27882
rect 24320 27470 24348 31146
rect 24412 28150 24440 33798
rect 24492 32224 24544 32230
rect 24492 32166 24544 32172
rect 24400 28144 24452 28150
rect 24400 28086 24452 28092
rect 24308 27464 24360 27470
rect 24308 27406 24360 27412
rect 24400 27328 24452 27334
rect 24400 27270 24452 27276
rect 24308 26852 24360 26858
rect 24308 26794 24360 26800
rect 24320 23118 24348 26794
rect 24412 26790 24440 27270
rect 24400 26784 24452 26790
rect 24400 26726 24452 26732
rect 24412 26518 24440 26726
rect 24400 26512 24452 26518
rect 24400 26454 24452 26460
rect 24504 26382 24532 32166
rect 24596 30734 24624 35974
rect 24688 33998 24716 39238
rect 24780 38321 24808 40326
rect 24766 38312 24822 38321
rect 24766 38247 24822 38256
rect 24768 38208 24820 38214
rect 24768 38150 24820 38156
rect 24780 36786 24808 38150
rect 24768 36780 24820 36786
rect 24768 36722 24820 36728
rect 24780 35601 24808 36722
rect 24872 36530 24900 42502
rect 24964 41478 24992 43982
rect 25044 43852 25096 43858
rect 25044 43794 25096 43800
rect 25056 42158 25084 43794
rect 25148 42838 25176 50662
rect 25332 50561 25360 50866
rect 25318 50552 25374 50561
rect 25318 50487 25374 50496
rect 25320 50312 25372 50318
rect 25320 50254 25372 50260
rect 25332 49881 25360 50254
rect 25318 49872 25374 49881
rect 25318 49807 25374 49816
rect 25320 49224 25372 49230
rect 25320 49166 25372 49172
rect 25332 48521 25360 49166
rect 25318 48512 25374 48521
rect 25318 48447 25374 48456
rect 25504 48136 25556 48142
rect 25504 48078 25556 48084
rect 25516 47462 25544 48078
rect 25504 47456 25556 47462
rect 25504 47398 25556 47404
rect 25516 47161 25544 47398
rect 25502 47152 25558 47161
rect 25502 47087 25558 47096
rect 25320 44872 25372 44878
rect 25320 44814 25372 44820
rect 25228 43104 25280 43110
rect 25228 43046 25280 43052
rect 25136 42832 25188 42838
rect 25136 42774 25188 42780
rect 25044 42152 25096 42158
rect 25044 42094 25096 42100
rect 24952 41472 25004 41478
rect 24952 41414 25004 41420
rect 24952 41064 25004 41070
rect 25056 41052 25084 42094
rect 25136 42016 25188 42022
rect 25136 41958 25188 41964
rect 25004 41024 25084 41052
rect 24952 41006 25004 41012
rect 24964 40594 24992 41006
rect 24952 40588 25004 40594
rect 24952 40530 25004 40536
rect 24952 39976 25004 39982
rect 24952 39918 25004 39924
rect 25044 39976 25096 39982
rect 25044 39918 25096 39924
rect 24964 39681 24992 39918
rect 24950 39672 25006 39681
rect 24950 39607 25006 39616
rect 25056 39574 25084 39918
rect 25044 39568 25096 39574
rect 25044 39510 25096 39516
rect 25148 39370 25176 41958
rect 25136 39364 25188 39370
rect 25136 39306 25188 39312
rect 25044 39024 25096 39030
rect 25044 38966 25096 38972
rect 24952 37188 25004 37194
rect 24952 37130 25004 37136
rect 24964 36961 24992 37130
rect 24950 36952 25006 36961
rect 24950 36887 25006 36896
rect 24872 36502 24992 36530
rect 24766 35592 24822 35601
rect 24766 35527 24822 35536
rect 24768 34944 24820 34950
rect 24768 34886 24820 34892
rect 24780 34490 24808 34886
rect 24780 34462 24900 34490
rect 24676 33992 24728 33998
rect 24676 33934 24728 33940
rect 24872 33930 24900 34462
rect 24860 33924 24912 33930
rect 24860 33866 24912 33872
rect 24676 33856 24728 33862
rect 24676 33798 24728 33804
rect 24584 30728 24636 30734
rect 24584 30670 24636 30676
rect 24584 30592 24636 30598
rect 24584 30534 24636 30540
rect 24596 30190 24624 30534
rect 24584 30184 24636 30190
rect 24584 30126 24636 30132
rect 24688 29238 24716 33798
rect 24872 33522 24900 33866
rect 24860 33516 24912 33522
rect 24860 33458 24912 33464
rect 24872 31482 24900 33458
rect 24860 31476 24912 31482
rect 24860 31418 24912 31424
rect 24872 30938 24900 31418
rect 24860 30932 24912 30938
rect 24860 30874 24912 30880
rect 24872 30666 24900 30874
rect 24860 30660 24912 30666
rect 24860 30602 24912 30608
rect 24768 30592 24820 30598
rect 24768 30534 24820 30540
rect 24676 29232 24728 29238
rect 24676 29174 24728 29180
rect 24584 29028 24636 29034
rect 24584 28970 24636 28976
rect 24492 26376 24544 26382
rect 24492 26318 24544 26324
rect 24596 24970 24624 28970
rect 24676 28620 24728 28626
rect 24676 28562 24728 28568
rect 24688 28014 24716 28562
rect 24676 28008 24728 28014
rect 24676 27950 24728 27956
rect 24688 26761 24716 27950
rect 24780 27062 24808 30534
rect 24872 30394 24900 30602
rect 24860 30388 24912 30394
rect 24860 30330 24912 30336
rect 24860 28416 24912 28422
rect 24860 28358 24912 28364
rect 24872 28121 24900 28358
rect 24858 28112 24914 28121
rect 24858 28047 24914 28056
rect 24768 27056 24820 27062
rect 24768 26998 24820 27004
rect 24860 26920 24912 26926
rect 24860 26862 24912 26868
rect 24674 26752 24730 26761
rect 24674 26687 24730 26696
rect 24676 26512 24728 26518
rect 24676 26454 24728 26460
rect 24504 24942 24624 24970
rect 24400 24404 24452 24410
rect 24400 24346 24452 24352
rect 24412 23322 24440 24346
rect 24504 24206 24532 24942
rect 24688 24834 24716 26454
rect 24768 25764 24820 25770
rect 24768 25706 24820 25712
rect 24596 24818 24716 24834
rect 24584 24812 24716 24818
rect 24636 24806 24716 24812
rect 24584 24754 24636 24760
rect 24596 24410 24624 24754
rect 24584 24404 24636 24410
rect 24584 24346 24636 24352
rect 24492 24200 24544 24206
rect 24492 24142 24544 24148
rect 24492 24064 24544 24070
rect 24492 24006 24544 24012
rect 24676 24064 24728 24070
rect 24676 24006 24728 24012
rect 24400 23316 24452 23322
rect 24400 23258 24452 23264
rect 24308 23112 24360 23118
rect 24308 23054 24360 23060
rect 24412 22658 24440 23258
rect 24504 22778 24532 24006
rect 24584 22976 24636 22982
rect 24584 22918 24636 22924
rect 24492 22772 24544 22778
rect 24492 22714 24544 22720
rect 24412 22642 24532 22658
rect 24412 22636 24544 22642
rect 24412 22630 24492 22636
rect 24492 22578 24544 22584
rect 24308 22432 24360 22438
rect 24308 22374 24360 22380
rect 24320 22166 24348 22374
rect 24504 22166 24532 22578
rect 24308 22160 24360 22166
rect 24308 22102 24360 22108
rect 24492 22160 24544 22166
rect 24492 22102 24544 22108
rect 24216 22024 24268 22030
rect 24216 21966 24268 21972
rect 24320 21842 24348 22102
rect 24228 21814 24348 21842
rect 24228 20398 24256 21814
rect 24400 21480 24452 21486
rect 24400 21422 24452 21428
rect 24308 21140 24360 21146
rect 24308 21082 24360 21088
rect 24216 20392 24268 20398
rect 24216 20334 24268 20340
rect 24216 20052 24268 20058
rect 24216 19994 24268 20000
rect 24228 18970 24256 19994
rect 24216 18964 24268 18970
rect 24216 18906 24268 18912
rect 24228 18630 24256 18906
rect 24320 18766 24348 21082
rect 24412 20602 24440 21422
rect 24490 21312 24546 21321
rect 24490 21247 24546 21256
rect 24400 20596 24452 20602
rect 24400 20538 24452 20544
rect 24504 19378 24532 21247
rect 24492 19372 24544 19378
rect 24492 19314 24544 19320
rect 24308 18760 24360 18766
rect 24308 18702 24360 18708
rect 24216 18624 24268 18630
rect 24216 18566 24268 18572
rect 24228 18358 24256 18566
rect 24216 18352 24268 18358
rect 24216 18294 24268 18300
rect 24228 17338 24256 18294
rect 24216 17332 24268 17338
rect 24216 17274 24268 17280
rect 24228 16794 24256 17274
rect 24216 16788 24268 16794
rect 24216 16730 24268 16736
rect 23940 16108 23992 16114
rect 23940 16050 23992 16056
rect 23940 15972 23992 15978
rect 23940 15914 23992 15920
rect 23756 15020 23808 15026
rect 23756 14962 23808 14968
rect 23848 13184 23900 13190
rect 23848 13126 23900 13132
rect 23664 11756 23716 11762
rect 23664 11698 23716 11704
rect 23480 11620 23532 11626
rect 23480 11562 23532 11568
rect 23388 11144 23440 11150
rect 23388 11086 23440 11092
rect 22950 10364 23258 10373
rect 22950 10362 22956 10364
rect 23012 10362 23036 10364
rect 23092 10362 23116 10364
rect 23172 10362 23196 10364
rect 23252 10362 23258 10364
rect 23012 10310 23014 10362
rect 23194 10310 23196 10362
rect 22950 10308 22956 10310
rect 23012 10308 23036 10310
rect 23092 10308 23116 10310
rect 23172 10308 23196 10310
rect 23252 10308 23258 10310
rect 22950 10299 23258 10308
rect 22950 9276 23258 9285
rect 22950 9274 22956 9276
rect 23012 9274 23036 9276
rect 23092 9274 23116 9276
rect 23172 9274 23196 9276
rect 23252 9274 23258 9276
rect 23012 9222 23014 9274
rect 23194 9222 23196 9274
rect 22950 9220 22956 9222
rect 23012 9220 23036 9222
rect 23092 9220 23116 9222
rect 23172 9220 23196 9222
rect 23252 9220 23258 9222
rect 22950 9211 23258 9220
rect 22836 8968 22888 8974
rect 22836 8910 22888 8916
rect 22744 8900 22796 8906
rect 22744 8842 22796 8848
rect 22756 7478 22784 8842
rect 23296 8832 23348 8838
rect 23296 8774 23348 8780
rect 22950 8188 23258 8197
rect 22950 8186 22956 8188
rect 23012 8186 23036 8188
rect 23092 8186 23116 8188
rect 23172 8186 23196 8188
rect 23252 8186 23258 8188
rect 23012 8134 23014 8186
rect 23194 8134 23196 8186
rect 22950 8132 22956 8134
rect 23012 8132 23036 8134
rect 23092 8132 23116 8134
rect 23172 8132 23196 8134
rect 23252 8132 23258 8134
rect 22950 8123 23258 8132
rect 22744 7472 22796 7478
rect 22744 7414 22796 7420
rect 22468 7336 22520 7342
rect 22468 7278 22520 7284
rect 22008 6724 22060 6730
rect 22008 6666 22060 6672
rect 21916 5636 21968 5642
rect 21916 5578 21968 5584
rect 21824 4208 21876 4214
rect 21824 4150 21876 4156
rect 21732 2916 21784 2922
rect 21732 2858 21784 2864
rect 21928 2802 21956 5578
rect 22020 3058 22048 6666
rect 22100 6180 22152 6186
rect 22100 6122 22152 6128
rect 22008 3052 22060 3058
rect 22008 2994 22060 3000
rect 21744 2774 21956 2802
rect 21744 800 21772 2774
rect 22112 800 22140 6122
rect 22284 5160 22336 5166
rect 22284 5102 22336 5108
rect 22296 2854 22324 5102
rect 22284 2848 22336 2854
rect 22284 2790 22336 2796
rect 22480 800 22508 7278
rect 22950 7100 23258 7109
rect 22950 7098 22956 7100
rect 23012 7098 23036 7100
rect 23092 7098 23116 7100
rect 23172 7098 23196 7100
rect 23252 7098 23258 7100
rect 23012 7046 23014 7098
rect 23194 7046 23196 7098
rect 22950 7044 22956 7046
rect 23012 7044 23036 7046
rect 23092 7044 23116 7046
rect 23172 7044 23196 7046
rect 23252 7044 23258 7046
rect 22950 7035 23258 7044
rect 23308 6322 23336 8774
rect 23388 6384 23440 6390
rect 23388 6326 23440 6332
rect 23296 6316 23348 6322
rect 23296 6258 23348 6264
rect 22950 6012 23258 6021
rect 22950 6010 22956 6012
rect 23012 6010 23036 6012
rect 23092 6010 23116 6012
rect 23172 6010 23196 6012
rect 23252 6010 23258 6012
rect 23012 5958 23014 6010
rect 23194 5958 23196 6010
rect 22950 5956 22956 5958
rect 23012 5956 23036 5958
rect 23092 5956 23116 5958
rect 23172 5956 23196 5958
rect 23252 5956 23258 5958
rect 22950 5947 23258 5956
rect 22950 4924 23258 4933
rect 22950 4922 22956 4924
rect 23012 4922 23036 4924
rect 23092 4922 23116 4924
rect 23172 4922 23196 4924
rect 23252 4922 23258 4924
rect 23012 4870 23014 4922
rect 23194 4870 23196 4922
rect 22950 4868 22956 4870
rect 23012 4868 23036 4870
rect 23092 4868 23116 4870
rect 23172 4868 23196 4870
rect 23252 4868 23258 4870
rect 22950 4859 23258 4868
rect 23400 4321 23428 6326
rect 23386 4312 23442 4321
rect 23386 4247 23442 4256
rect 23492 4146 23520 11562
rect 23860 9994 23888 13126
rect 23952 12850 23980 15914
rect 24596 15162 24624 22918
rect 24688 17678 24716 24006
rect 24780 19854 24808 25706
rect 24872 24750 24900 26862
rect 24860 24744 24912 24750
rect 24860 24686 24912 24692
rect 24860 24268 24912 24274
rect 24860 24210 24912 24216
rect 24872 24041 24900 24210
rect 24858 24032 24914 24041
rect 24858 23967 24914 23976
rect 24860 23180 24912 23186
rect 24860 23122 24912 23128
rect 24872 22681 24900 23122
rect 24858 22672 24914 22681
rect 24858 22607 24914 22616
rect 24860 22092 24912 22098
rect 24860 22034 24912 22040
rect 24872 22001 24900 22034
rect 24858 21992 24914 22001
rect 24858 21927 24914 21936
rect 24860 21616 24912 21622
rect 24860 21558 24912 21564
rect 24872 21078 24900 21558
rect 24860 21072 24912 21078
rect 24860 21014 24912 21020
rect 24872 20602 24900 21014
rect 24860 20596 24912 20602
rect 24860 20538 24912 20544
rect 24872 20058 24900 20538
rect 24860 20052 24912 20058
rect 24860 19994 24912 20000
rect 24858 19952 24914 19961
rect 24858 19887 24914 19896
rect 24768 19848 24820 19854
rect 24768 19790 24820 19796
rect 24872 19446 24900 19887
rect 24860 19440 24912 19446
rect 24860 19382 24912 19388
rect 24766 17912 24822 17921
rect 24766 17847 24822 17856
rect 24676 17672 24728 17678
rect 24676 17614 24728 17620
rect 24674 17232 24730 17241
rect 24674 17167 24730 17176
rect 24584 15156 24636 15162
rect 24584 15098 24636 15104
rect 24688 14958 24716 17167
rect 24780 16046 24808 17847
rect 24858 16552 24914 16561
rect 24858 16487 24914 16496
rect 24872 16114 24900 16487
rect 24860 16108 24912 16114
rect 24860 16050 24912 16056
rect 24768 16040 24820 16046
rect 24768 15982 24820 15988
rect 24858 15872 24914 15881
rect 24858 15807 24914 15816
rect 24872 15570 24900 15807
rect 24860 15564 24912 15570
rect 24860 15506 24912 15512
rect 24860 15088 24912 15094
rect 24860 15030 24912 15036
rect 24676 14952 24728 14958
rect 24676 14894 24728 14900
rect 24872 14521 24900 15030
rect 24858 14512 24914 14521
rect 24858 14447 24914 14456
rect 24766 13832 24822 13841
rect 24766 13767 24822 13776
rect 24674 13152 24730 13161
rect 24674 13087 24730 13096
rect 23940 12844 23992 12850
rect 23940 12786 23992 12792
rect 24584 12096 24636 12102
rect 24584 12038 24636 12044
rect 23940 11552 23992 11558
rect 23940 11494 23992 11500
rect 23952 10674 23980 11494
rect 24216 11076 24268 11082
rect 24216 11018 24268 11024
rect 24032 11008 24084 11014
rect 24032 10950 24084 10956
rect 23940 10668 23992 10674
rect 23940 10610 23992 10616
rect 23848 9988 23900 9994
rect 23848 9930 23900 9936
rect 23940 9580 23992 9586
rect 23940 9522 23992 9528
rect 23952 6118 23980 9522
rect 24044 8498 24072 10950
rect 24124 9920 24176 9926
rect 24124 9862 24176 9868
rect 24032 8492 24084 8498
rect 24032 8434 24084 8440
rect 24136 7410 24164 9862
rect 24228 7886 24256 11018
rect 24308 10464 24360 10470
rect 24308 10406 24360 10412
rect 24320 7886 24348 10406
rect 24596 10062 24624 12038
rect 24688 11694 24716 13087
rect 24780 12782 24808 13767
rect 24860 12912 24912 12918
rect 24860 12854 24912 12860
rect 24768 12776 24820 12782
rect 24768 12718 24820 12724
rect 24872 12481 24900 12854
rect 24858 12472 24914 12481
rect 24858 12407 24914 12416
rect 24964 12434 24992 36502
rect 25056 36310 25084 38966
rect 25136 38480 25188 38486
rect 25136 38422 25188 38428
rect 25148 37670 25176 38422
rect 25136 37664 25188 37670
rect 25136 37606 25188 37612
rect 25044 36304 25096 36310
rect 25044 36246 25096 36252
rect 25148 36122 25176 37606
rect 25056 36094 25176 36122
rect 25056 35630 25084 36094
rect 25044 35624 25096 35630
rect 25044 35566 25096 35572
rect 25056 35154 25084 35566
rect 25240 35494 25268 43046
rect 25332 42401 25360 44814
rect 25504 44328 25556 44334
rect 25504 44270 25556 44276
rect 25516 43654 25544 44270
rect 25504 43648 25556 43654
rect 25504 43590 25556 43596
rect 25412 43308 25464 43314
rect 25412 43250 25464 43256
rect 25424 42922 25452 43250
rect 25516 43081 25544 43590
rect 25502 43072 25558 43081
rect 25502 43007 25558 43016
rect 25424 42894 25544 42922
rect 25412 42832 25464 42838
rect 25412 42774 25464 42780
rect 25318 42392 25374 42401
rect 25318 42327 25374 42336
rect 25320 40928 25372 40934
rect 25320 40870 25372 40876
rect 25332 39982 25360 40870
rect 25320 39976 25372 39982
rect 25320 39918 25372 39924
rect 25332 39001 25360 39918
rect 25424 39438 25452 42774
rect 25516 42566 25544 42894
rect 25504 42560 25556 42566
rect 25504 42502 25556 42508
rect 25516 41721 25544 42502
rect 25502 41712 25558 41721
rect 25502 41647 25558 41656
rect 25412 39432 25464 39438
rect 25412 39374 25464 39380
rect 25318 38992 25374 39001
rect 25318 38927 25374 38936
rect 25412 38344 25464 38350
rect 25412 38286 25464 38292
rect 25320 37664 25372 37670
rect 25424 37641 25452 38286
rect 25320 37606 25372 37612
rect 25410 37632 25466 37641
rect 25332 37262 25360 37606
rect 25410 37567 25466 37576
rect 25504 37460 25556 37466
rect 25504 37402 25556 37408
rect 25320 37256 25372 37262
rect 25320 37198 25372 37204
rect 25332 36281 25360 37198
rect 25318 36272 25374 36281
rect 25318 36207 25374 36216
rect 25320 36168 25372 36174
rect 25320 36110 25372 36116
rect 25228 35488 25280 35494
rect 25228 35430 25280 35436
rect 25044 35148 25096 35154
rect 25044 35090 25096 35096
rect 25332 34921 25360 36110
rect 25412 35080 25464 35086
rect 25412 35022 25464 35028
rect 25318 34912 25374 34921
rect 25318 34847 25374 34856
rect 25228 34604 25280 34610
rect 25228 34546 25280 34552
rect 25320 34604 25372 34610
rect 25320 34546 25372 34552
rect 25136 32564 25188 32570
rect 25136 32506 25188 32512
rect 25044 31136 25096 31142
rect 25044 31078 25096 31084
rect 25056 25974 25084 31078
rect 25148 29850 25176 32506
rect 25136 29844 25188 29850
rect 25136 29786 25188 29792
rect 25240 28762 25268 34546
rect 25332 33862 25360 34546
rect 25424 34241 25452 35022
rect 25410 34232 25466 34241
rect 25410 34167 25466 34176
rect 25320 33856 25372 33862
rect 25320 33798 25372 33804
rect 25332 33561 25360 33798
rect 25516 33658 25544 37402
rect 25504 33652 25556 33658
rect 25504 33594 25556 33600
rect 25318 33552 25374 33561
rect 25318 33487 25374 33496
rect 25320 32904 25372 32910
rect 25318 32872 25320 32881
rect 25372 32872 25374 32881
rect 25318 32807 25374 32816
rect 25320 32428 25372 32434
rect 25320 32370 25372 32376
rect 25332 32201 25360 32370
rect 25318 32192 25374 32201
rect 25318 32127 25374 32136
rect 25608 31958 25636 51206
rect 25700 37398 25728 51750
rect 25872 47524 25924 47530
rect 25872 47466 25924 47472
rect 25688 37392 25740 37398
rect 25688 37334 25740 37340
rect 25596 31952 25648 31958
rect 25596 31894 25648 31900
rect 25412 31816 25464 31822
rect 25412 31758 25464 31764
rect 25318 31512 25374 31521
rect 25318 31447 25374 31456
rect 25332 31346 25360 31447
rect 25320 31340 25372 31346
rect 25320 31282 25372 31288
rect 25332 30938 25360 31282
rect 25320 30932 25372 30938
rect 25320 30874 25372 30880
rect 25424 30841 25452 31758
rect 25410 30832 25466 30841
rect 25410 30767 25466 30776
rect 25318 30152 25374 30161
rect 25318 30087 25374 30096
rect 25332 29646 25360 30087
rect 25320 29640 25372 29646
rect 25320 29582 25372 29588
rect 25332 29306 25360 29582
rect 25410 29472 25466 29481
rect 25410 29407 25466 29416
rect 25320 29300 25372 29306
rect 25320 29242 25372 29248
rect 25228 28756 25280 28762
rect 25228 28698 25280 28704
rect 25424 28558 25452 29407
rect 25412 28552 25464 28558
rect 25412 28494 25464 28500
rect 25424 28218 25452 28494
rect 25412 28212 25464 28218
rect 25412 28154 25464 28160
rect 25504 28144 25556 28150
rect 25504 28086 25556 28092
rect 25410 27432 25466 27441
rect 25410 27367 25466 27376
rect 25424 27130 25452 27367
rect 25412 27124 25464 27130
rect 25412 27066 25464 27072
rect 25424 26450 25452 27066
rect 25412 26444 25464 26450
rect 25412 26386 25464 26392
rect 25228 26308 25280 26314
rect 25228 26250 25280 26256
rect 25044 25968 25096 25974
rect 25044 25910 25096 25916
rect 25044 25424 25096 25430
rect 25044 25366 25096 25372
rect 25056 23118 25084 25366
rect 25134 24712 25190 24721
rect 25134 24647 25190 24656
rect 25148 23798 25176 24647
rect 25136 23792 25188 23798
rect 25136 23734 25188 23740
rect 25044 23112 25096 23118
rect 25044 23054 25096 23060
rect 25044 22092 25096 22098
rect 25044 22034 25096 22040
rect 25056 21690 25084 22034
rect 25044 21684 25096 21690
rect 25044 21626 25096 21632
rect 25044 21480 25096 21486
rect 25044 21422 25096 21428
rect 25056 20466 25084 21422
rect 25134 20632 25190 20641
rect 25134 20567 25190 20576
rect 25044 20460 25096 20466
rect 25044 20402 25096 20408
rect 25148 19922 25176 20567
rect 25136 19916 25188 19922
rect 25136 19858 25188 19864
rect 25240 19378 25268 26250
rect 25318 25392 25374 25401
rect 25318 25327 25374 25336
rect 25332 22642 25360 25327
rect 25412 24744 25464 24750
rect 25412 24686 25464 24692
rect 25424 23186 25452 24686
rect 25412 23180 25464 23186
rect 25412 23122 25464 23128
rect 25516 22982 25544 28086
rect 25504 22976 25556 22982
rect 25504 22918 25556 22924
rect 25320 22636 25372 22642
rect 25320 22578 25372 22584
rect 25332 22234 25360 22578
rect 25320 22228 25372 22234
rect 25320 22170 25372 22176
rect 25884 22094 25912 47466
rect 26056 46504 26108 46510
rect 26056 46446 26108 46452
rect 25964 44396 26016 44402
rect 25964 44338 26016 44344
rect 25976 38554 26004 44338
rect 26068 41002 26096 46446
rect 26056 40996 26108 41002
rect 26056 40938 26108 40944
rect 25964 38548 26016 38554
rect 25964 38490 26016 38496
rect 25516 22066 25912 22094
rect 25228 19372 25280 19378
rect 25228 19314 25280 19320
rect 25134 15192 25190 15201
rect 25134 15127 25190 15136
rect 25148 14006 25176 15127
rect 25136 14000 25188 14006
rect 25136 13942 25188 13948
rect 24964 12406 25084 12434
rect 24952 12164 25004 12170
rect 24952 12106 25004 12112
rect 24964 11801 24992 12106
rect 24950 11792 25006 11801
rect 24950 11727 25006 11736
rect 24676 11688 24728 11694
rect 24676 11630 24728 11636
rect 24766 11112 24822 11121
rect 24766 11047 24822 11056
rect 24780 10606 24808 11047
rect 24768 10600 24820 10606
rect 24768 10542 24820 10548
rect 24766 10432 24822 10441
rect 24766 10367 24822 10376
rect 24584 10056 24636 10062
rect 24584 9998 24636 10004
rect 24780 9518 24808 10367
rect 24860 10124 24912 10130
rect 24860 10066 24912 10072
rect 24872 9761 24900 10066
rect 24858 9752 24914 9761
rect 24858 9687 24914 9696
rect 24768 9512 24820 9518
rect 24768 9454 24820 9460
rect 24492 9376 24544 9382
rect 24492 9318 24544 9324
rect 24216 7880 24268 7886
rect 24216 7822 24268 7828
rect 24308 7880 24360 7886
rect 24308 7822 24360 7828
rect 24124 7404 24176 7410
rect 24124 7346 24176 7352
rect 24504 6798 24532 9318
rect 25056 8974 25084 12406
rect 25134 9072 25190 9081
rect 25134 9007 25190 9016
rect 24860 8968 24912 8974
rect 24860 8910 24912 8916
rect 25044 8968 25096 8974
rect 25044 8910 25096 8916
rect 24676 8832 24728 8838
rect 24676 8774 24728 8780
rect 24688 8566 24716 8774
rect 24676 8560 24728 8566
rect 24676 8502 24728 8508
rect 24584 8424 24636 8430
rect 24584 8366 24636 8372
rect 24766 8392 24822 8401
rect 24492 6792 24544 6798
rect 24492 6734 24544 6740
rect 23940 6112 23992 6118
rect 23940 6054 23992 6060
rect 23480 4140 23532 4146
rect 23480 4082 23532 4088
rect 22950 3836 23258 3845
rect 22950 3834 22956 3836
rect 23012 3834 23036 3836
rect 23092 3834 23116 3836
rect 23172 3834 23196 3836
rect 23252 3834 23258 3836
rect 23012 3782 23014 3834
rect 23194 3782 23196 3834
rect 22950 3780 22956 3782
rect 23012 3780 23036 3782
rect 23092 3780 23116 3782
rect 23172 3780 23196 3782
rect 23252 3780 23258 3782
rect 22950 3771 23258 3780
rect 23848 3528 23900 3534
rect 23294 3496 23350 3505
rect 23848 3470 23900 3476
rect 23294 3431 23350 3440
rect 22836 3052 22888 3058
rect 22836 2994 22888 3000
rect 22848 800 22876 2994
rect 22950 2748 23258 2757
rect 22950 2746 22956 2748
rect 23012 2746 23036 2748
rect 23092 2746 23116 2748
rect 23172 2746 23196 2748
rect 23252 2746 23258 2748
rect 23012 2694 23014 2746
rect 23194 2694 23196 2746
rect 22950 2692 22956 2694
rect 23012 2692 23036 2694
rect 23092 2692 23116 2694
rect 23172 2692 23196 2694
rect 23252 2692 23258 2694
rect 22950 2683 23258 2692
rect 23308 2530 23336 3431
rect 23860 3194 23888 3470
rect 23848 3188 23900 3194
rect 23848 3130 23900 3136
rect 23940 2984 23992 2990
rect 23940 2926 23992 2932
rect 23572 2916 23624 2922
rect 23572 2858 23624 2864
rect 23216 2502 23336 2530
rect 23216 800 23244 2502
rect 23584 800 23612 2858
rect 23952 800 23980 2926
rect 24596 2774 24624 8366
rect 24766 8327 24822 8336
rect 24676 7744 24728 7750
rect 24676 7686 24728 7692
rect 24688 5234 24716 7686
rect 24780 7342 24808 8327
rect 24872 7562 24900 8910
rect 25148 8566 25176 9007
rect 25516 8906 25544 22066
rect 25504 8900 25556 8906
rect 25504 8842 25556 8848
rect 25228 8832 25280 8838
rect 25228 8774 25280 8780
rect 25136 8560 25188 8566
rect 25136 8502 25188 8508
rect 24952 7948 25004 7954
rect 24952 7890 25004 7896
rect 24964 7721 24992 7890
rect 24950 7712 25006 7721
rect 24950 7647 25006 7656
rect 24872 7534 24992 7562
rect 24768 7336 24820 7342
rect 24768 7278 24820 7284
rect 24766 7032 24822 7041
rect 24766 6967 24822 6976
rect 24780 6254 24808 6967
rect 24860 6860 24912 6866
rect 24860 6802 24912 6808
rect 24872 6361 24900 6802
rect 24858 6352 24914 6361
rect 24858 6287 24914 6296
rect 24768 6248 24820 6254
rect 24768 6190 24820 6196
rect 24766 5672 24822 5681
rect 24766 5607 24822 5616
rect 24676 5228 24728 5234
rect 24676 5170 24728 5176
rect 24780 5166 24808 5607
rect 24768 5160 24820 5166
rect 24768 5102 24820 5108
rect 24596 2746 24716 2774
rect 24308 2440 24360 2446
rect 24308 2382 24360 2388
rect 24320 800 24348 2382
rect 24688 800 24716 2746
rect 24964 2650 24992 7534
rect 25240 3738 25268 8774
rect 25318 4992 25374 5001
rect 25318 4927 25374 4936
rect 25332 4826 25360 4927
rect 25320 4820 25372 4826
rect 25320 4762 25372 4768
rect 25320 3936 25372 3942
rect 25320 3878 25372 3884
rect 25228 3732 25280 3738
rect 25228 3674 25280 3680
rect 25044 3528 25096 3534
rect 25044 3470 25096 3476
rect 24952 2644 25004 2650
rect 24952 2586 25004 2592
rect 25056 800 25084 3470
rect 25332 2530 25360 3878
rect 25412 2916 25464 2922
rect 25412 2858 25464 2864
rect 25424 2650 25452 2858
rect 25412 2644 25464 2650
rect 25412 2586 25464 2592
rect 25332 2502 25452 2530
rect 25424 800 25452 2502
rect 18156 734 18368 762
rect 18418 0 18474 800
rect 18786 0 18842 800
rect 19154 0 19210 800
rect 19522 0 19578 800
rect 19890 0 19946 800
rect 20258 0 20314 800
rect 20626 0 20682 800
rect 20994 0 21050 800
rect 21362 0 21418 800
rect 21730 0 21786 800
rect 22098 0 22154 800
rect 22466 0 22522 800
rect 22834 0 22890 800
rect 23202 0 23258 800
rect 23570 0 23626 800
rect 23938 0 23994 800
rect 24306 0 24362 800
rect 24674 0 24730 800
rect 25042 0 25098 800
rect 25410 0 25466 800
<< via2 >>
rect 1214 52672 1270 52728
rect 1122 50396 1124 50416
rect 1124 50396 1176 50416
rect 1176 50396 1178 50416
rect 1122 50360 1178 50396
rect 2778 54984 2834 55040
rect 2956 53882 3012 53884
rect 3036 53882 3092 53884
rect 3116 53882 3172 53884
rect 3196 53882 3252 53884
rect 2956 53830 3002 53882
rect 3002 53830 3012 53882
rect 3036 53830 3066 53882
rect 3066 53830 3078 53882
rect 3078 53830 3092 53882
rect 3116 53830 3130 53882
rect 3130 53830 3142 53882
rect 3142 53830 3172 53882
rect 3196 53830 3206 53882
rect 3206 53830 3252 53882
rect 2956 53828 3012 53830
rect 3036 53828 3092 53830
rect 3116 53828 3172 53830
rect 3196 53828 3252 53830
rect 2956 52794 3012 52796
rect 3036 52794 3092 52796
rect 3116 52794 3172 52796
rect 3196 52794 3252 52796
rect 2956 52742 3002 52794
rect 3002 52742 3012 52794
rect 3036 52742 3066 52794
rect 3066 52742 3078 52794
rect 3078 52742 3092 52794
rect 3116 52742 3130 52794
rect 3130 52742 3142 52794
rect 3142 52742 3172 52794
rect 3196 52742 3206 52794
rect 3206 52742 3252 52794
rect 2956 52740 3012 52742
rect 3036 52740 3092 52742
rect 3116 52740 3172 52742
rect 3196 52740 3252 52742
rect 2956 51706 3012 51708
rect 3036 51706 3092 51708
rect 3116 51706 3172 51708
rect 3196 51706 3252 51708
rect 2956 51654 3002 51706
rect 3002 51654 3012 51706
rect 3036 51654 3066 51706
rect 3066 51654 3078 51706
rect 3078 51654 3092 51706
rect 3116 51654 3130 51706
rect 3130 51654 3142 51706
rect 3142 51654 3172 51706
rect 3196 51654 3206 51706
rect 3206 51654 3252 51706
rect 2956 51652 3012 51654
rect 3036 51652 3092 51654
rect 3116 51652 3172 51654
rect 3196 51652 3252 51654
rect 2956 50618 3012 50620
rect 3036 50618 3092 50620
rect 3116 50618 3172 50620
rect 3196 50618 3252 50620
rect 2956 50566 3002 50618
rect 3002 50566 3012 50618
rect 3036 50566 3066 50618
rect 3066 50566 3078 50618
rect 3078 50566 3092 50618
rect 3116 50566 3130 50618
rect 3130 50566 3142 50618
rect 3142 50566 3172 50618
rect 3196 50566 3206 50618
rect 3206 50566 3252 50618
rect 2956 50564 3012 50566
rect 3036 50564 3092 50566
rect 3116 50564 3172 50566
rect 3196 50564 3252 50566
rect 2956 49530 3012 49532
rect 3036 49530 3092 49532
rect 3116 49530 3172 49532
rect 3196 49530 3252 49532
rect 2956 49478 3002 49530
rect 3002 49478 3012 49530
rect 3036 49478 3066 49530
rect 3066 49478 3078 49530
rect 3078 49478 3092 49530
rect 3116 49478 3130 49530
rect 3130 49478 3142 49530
rect 3142 49478 3172 49530
rect 3196 49478 3206 49530
rect 3206 49478 3252 49530
rect 2956 49476 3012 49478
rect 3036 49476 3092 49478
rect 3116 49476 3172 49478
rect 3196 49476 3252 49478
rect 2956 48442 3012 48444
rect 3036 48442 3092 48444
rect 3116 48442 3172 48444
rect 3196 48442 3252 48444
rect 2956 48390 3002 48442
rect 3002 48390 3012 48442
rect 3036 48390 3066 48442
rect 3066 48390 3078 48442
rect 3078 48390 3092 48442
rect 3116 48390 3130 48442
rect 3130 48390 3142 48442
rect 3142 48390 3172 48442
rect 3196 48390 3206 48442
rect 3206 48390 3252 48442
rect 2956 48388 3012 48390
rect 3036 48388 3092 48390
rect 3116 48388 3172 48390
rect 3196 48388 3252 48390
rect 1306 48068 1362 48104
rect 1306 48048 1308 48068
rect 1308 48048 1360 48068
rect 1360 48048 1362 48068
rect 2956 47354 3012 47356
rect 3036 47354 3092 47356
rect 3116 47354 3172 47356
rect 3196 47354 3252 47356
rect 2956 47302 3002 47354
rect 3002 47302 3012 47354
rect 3036 47302 3066 47354
rect 3066 47302 3078 47354
rect 3078 47302 3092 47354
rect 3116 47302 3130 47354
rect 3130 47302 3142 47354
rect 3142 47302 3172 47354
rect 3196 47302 3206 47354
rect 3206 47302 3252 47354
rect 2956 47300 3012 47302
rect 3036 47300 3092 47302
rect 3116 47300 3172 47302
rect 3196 47300 3252 47302
rect 2956 46266 3012 46268
rect 3036 46266 3092 46268
rect 3116 46266 3172 46268
rect 3196 46266 3252 46268
rect 2956 46214 3002 46266
rect 3002 46214 3012 46266
rect 3036 46214 3066 46266
rect 3066 46214 3078 46266
rect 3078 46214 3092 46266
rect 3116 46214 3130 46266
rect 3130 46214 3142 46266
rect 3142 46214 3172 46266
rect 3196 46214 3206 46266
rect 3206 46214 3252 46266
rect 2956 46212 3012 46214
rect 3036 46212 3092 46214
rect 3116 46212 3172 46214
rect 3196 46212 3252 46214
rect 1214 45736 1270 45792
rect 2956 45178 3012 45180
rect 3036 45178 3092 45180
rect 3116 45178 3172 45180
rect 3196 45178 3252 45180
rect 2956 45126 3002 45178
rect 3002 45126 3012 45178
rect 3036 45126 3066 45178
rect 3066 45126 3078 45178
rect 3078 45126 3092 45178
rect 3116 45126 3130 45178
rect 3130 45126 3142 45178
rect 3142 45126 3172 45178
rect 3196 45126 3206 45178
rect 3206 45126 3252 45178
rect 2956 45124 3012 45126
rect 3036 45124 3092 45126
rect 3116 45124 3172 45126
rect 3196 45124 3252 45126
rect 2956 44090 3012 44092
rect 3036 44090 3092 44092
rect 3116 44090 3172 44092
rect 3196 44090 3252 44092
rect 2956 44038 3002 44090
rect 3002 44038 3012 44090
rect 3036 44038 3066 44090
rect 3066 44038 3078 44090
rect 3078 44038 3092 44090
rect 3116 44038 3130 44090
rect 3130 44038 3142 44090
rect 3142 44038 3172 44090
rect 3196 44038 3206 44090
rect 3206 44038 3252 44090
rect 2956 44036 3012 44038
rect 3036 44036 3092 44038
rect 3116 44036 3172 44038
rect 3196 44036 3252 44038
rect 1306 43424 1362 43480
rect 2956 43002 3012 43004
rect 3036 43002 3092 43004
rect 3116 43002 3172 43004
rect 3196 43002 3252 43004
rect 2956 42950 3002 43002
rect 3002 42950 3012 43002
rect 3036 42950 3066 43002
rect 3066 42950 3078 43002
rect 3078 42950 3092 43002
rect 3116 42950 3130 43002
rect 3130 42950 3142 43002
rect 3142 42950 3172 43002
rect 3196 42950 3206 43002
rect 3206 42950 3252 43002
rect 2956 42948 3012 42950
rect 3036 42948 3092 42950
rect 3116 42948 3172 42950
rect 3196 42948 3252 42950
rect 2956 41914 3012 41916
rect 3036 41914 3092 41916
rect 3116 41914 3172 41916
rect 3196 41914 3252 41916
rect 2956 41862 3002 41914
rect 3002 41862 3012 41914
rect 3036 41862 3066 41914
rect 3066 41862 3078 41914
rect 3078 41862 3092 41914
rect 3116 41862 3130 41914
rect 3130 41862 3142 41914
rect 3142 41862 3172 41914
rect 3196 41862 3206 41914
rect 3206 41862 3252 41914
rect 2956 41860 3012 41862
rect 3036 41860 3092 41862
rect 3116 41860 3172 41862
rect 3196 41860 3252 41862
rect 1674 41112 1730 41168
rect 2956 40826 3012 40828
rect 3036 40826 3092 40828
rect 3116 40826 3172 40828
rect 3196 40826 3252 40828
rect 2956 40774 3002 40826
rect 3002 40774 3012 40826
rect 3036 40774 3066 40826
rect 3066 40774 3078 40826
rect 3078 40774 3092 40826
rect 3116 40774 3130 40826
rect 3130 40774 3142 40826
rect 3142 40774 3172 40826
rect 3196 40774 3206 40826
rect 3206 40774 3252 40826
rect 2956 40772 3012 40774
rect 3036 40772 3092 40774
rect 3116 40772 3172 40774
rect 3196 40772 3252 40774
rect 2956 39738 3012 39740
rect 3036 39738 3092 39740
rect 3116 39738 3172 39740
rect 3196 39738 3252 39740
rect 2956 39686 3002 39738
rect 3002 39686 3012 39738
rect 3036 39686 3066 39738
rect 3066 39686 3078 39738
rect 3078 39686 3092 39738
rect 3116 39686 3130 39738
rect 3130 39686 3142 39738
rect 3142 39686 3172 39738
rect 3196 39686 3206 39738
rect 3206 39686 3252 39738
rect 2956 39684 3012 39686
rect 3036 39684 3092 39686
rect 3116 39684 3172 39686
rect 3196 39684 3252 39686
rect 1214 38800 1270 38856
rect 2956 38650 3012 38652
rect 3036 38650 3092 38652
rect 3116 38650 3172 38652
rect 3196 38650 3252 38652
rect 2956 38598 3002 38650
rect 3002 38598 3012 38650
rect 3036 38598 3066 38650
rect 3066 38598 3078 38650
rect 3078 38598 3092 38650
rect 3116 38598 3130 38650
rect 3130 38598 3142 38650
rect 3142 38598 3172 38650
rect 3196 38598 3206 38650
rect 3206 38598 3252 38650
rect 2956 38596 3012 38598
rect 3036 38596 3092 38598
rect 3116 38596 3172 38598
rect 3196 38596 3252 38598
rect 2956 37562 3012 37564
rect 3036 37562 3092 37564
rect 3116 37562 3172 37564
rect 3196 37562 3252 37564
rect 2956 37510 3002 37562
rect 3002 37510 3012 37562
rect 3036 37510 3066 37562
rect 3066 37510 3078 37562
rect 3078 37510 3092 37562
rect 3116 37510 3130 37562
rect 3130 37510 3142 37562
rect 3142 37510 3172 37562
rect 3196 37510 3206 37562
rect 3206 37510 3252 37562
rect 2956 37508 3012 37510
rect 3036 37508 3092 37510
rect 3116 37508 3172 37510
rect 3196 37508 3252 37510
rect 1306 36488 1362 36544
rect 1582 34176 1638 34232
rect 1306 31864 1362 31920
rect 1306 29552 1362 29608
rect 1306 27240 1362 27296
rect 2956 36474 3012 36476
rect 3036 36474 3092 36476
rect 3116 36474 3172 36476
rect 3196 36474 3252 36476
rect 2956 36422 3002 36474
rect 3002 36422 3012 36474
rect 3036 36422 3066 36474
rect 3066 36422 3078 36474
rect 3078 36422 3092 36474
rect 3116 36422 3130 36474
rect 3130 36422 3142 36474
rect 3142 36422 3172 36474
rect 3196 36422 3206 36474
rect 3206 36422 3252 36474
rect 2956 36420 3012 36422
rect 3036 36420 3092 36422
rect 3116 36420 3172 36422
rect 3196 36420 3252 36422
rect 2956 35386 3012 35388
rect 3036 35386 3092 35388
rect 3116 35386 3172 35388
rect 3196 35386 3252 35388
rect 2956 35334 3002 35386
rect 3002 35334 3012 35386
rect 3036 35334 3066 35386
rect 3066 35334 3078 35386
rect 3078 35334 3092 35386
rect 3116 35334 3130 35386
rect 3130 35334 3142 35386
rect 3142 35334 3172 35386
rect 3196 35334 3206 35386
rect 3206 35334 3252 35386
rect 2956 35332 3012 35334
rect 3036 35332 3092 35334
rect 3116 35332 3172 35334
rect 3196 35332 3252 35334
rect 1306 24928 1362 24984
rect 2956 34298 3012 34300
rect 3036 34298 3092 34300
rect 3116 34298 3172 34300
rect 3196 34298 3252 34300
rect 2956 34246 3002 34298
rect 3002 34246 3012 34298
rect 3036 34246 3066 34298
rect 3066 34246 3078 34298
rect 3078 34246 3092 34298
rect 3116 34246 3130 34298
rect 3130 34246 3142 34298
rect 3142 34246 3172 34298
rect 3196 34246 3206 34298
rect 3206 34246 3252 34298
rect 2956 34244 3012 34246
rect 3036 34244 3092 34246
rect 3116 34244 3172 34246
rect 3196 34244 3252 34246
rect 2956 33210 3012 33212
rect 3036 33210 3092 33212
rect 3116 33210 3172 33212
rect 3196 33210 3252 33212
rect 2956 33158 3002 33210
rect 3002 33158 3012 33210
rect 3036 33158 3066 33210
rect 3066 33158 3078 33210
rect 3078 33158 3092 33210
rect 3116 33158 3130 33210
rect 3130 33158 3142 33210
rect 3142 33158 3172 33210
rect 3196 33158 3206 33210
rect 3206 33158 3252 33210
rect 2956 33156 3012 33158
rect 3036 33156 3092 33158
rect 3116 33156 3172 33158
rect 3196 33156 3252 33158
rect 2956 32122 3012 32124
rect 3036 32122 3092 32124
rect 3116 32122 3172 32124
rect 3196 32122 3252 32124
rect 2956 32070 3002 32122
rect 3002 32070 3012 32122
rect 3036 32070 3066 32122
rect 3066 32070 3078 32122
rect 3078 32070 3092 32122
rect 3116 32070 3130 32122
rect 3130 32070 3142 32122
rect 3142 32070 3172 32122
rect 3196 32070 3206 32122
rect 3206 32070 3252 32122
rect 2956 32068 3012 32070
rect 3036 32068 3092 32070
rect 3116 32068 3172 32070
rect 3196 32068 3252 32070
rect 2956 31034 3012 31036
rect 3036 31034 3092 31036
rect 3116 31034 3172 31036
rect 3196 31034 3252 31036
rect 2956 30982 3002 31034
rect 3002 30982 3012 31034
rect 3036 30982 3066 31034
rect 3066 30982 3078 31034
rect 3078 30982 3092 31034
rect 3116 30982 3130 31034
rect 3130 30982 3142 31034
rect 3142 30982 3172 31034
rect 3196 30982 3206 31034
rect 3206 30982 3252 31034
rect 2956 30980 3012 30982
rect 3036 30980 3092 30982
rect 3116 30980 3172 30982
rect 3196 30980 3252 30982
rect 2956 29946 3012 29948
rect 3036 29946 3092 29948
rect 3116 29946 3172 29948
rect 3196 29946 3252 29948
rect 2956 29894 3002 29946
rect 3002 29894 3012 29946
rect 3036 29894 3066 29946
rect 3066 29894 3078 29946
rect 3078 29894 3092 29946
rect 3116 29894 3130 29946
rect 3130 29894 3142 29946
rect 3142 29894 3172 29946
rect 3196 29894 3206 29946
rect 3206 29894 3252 29946
rect 2956 29892 3012 29894
rect 3036 29892 3092 29894
rect 3116 29892 3172 29894
rect 3196 29892 3252 29894
rect 2956 28858 3012 28860
rect 3036 28858 3092 28860
rect 3116 28858 3172 28860
rect 3196 28858 3252 28860
rect 2956 28806 3002 28858
rect 3002 28806 3012 28858
rect 3036 28806 3066 28858
rect 3066 28806 3078 28858
rect 3078 28806 3092 28858
rect 3116 28806 3130 28858
rect 3130 28806 3142 28858
rect 3142 28806 3172 28858
rect 3196 28806 3206 28858
rect 3206 28806 3252 28858
rect 2956 28804 3012 28806
rect 3036 28804 3092 28806
rect 3116 28804 3172 28806
rect 3196 28804 3252 28806
rect 2956 27770 3012 27772
rect 3036 27770 3092 27772
rect 3116 27770 3172 27772
rect 3196 27770 3252 27772
rect 2956 27718 3002 27770
rect 3002 27718 3012 27770
rect 3036 27718 3066 27770
rect 3066 27718 3078 27770
rect 3078 27718 3092 27770
rect 3116 27718 3130 27770
rect 3130 27718 3142 27770
rect 3142 27718 3172 27770
rect 3196 27718 3206 27770
rect 3206 27718 3252 27770
rect 2956 27716 3012 27718
rect 3036 27716 3092 27718
rect 3116 27716 3172 27718
rect 3196 27716 3252 27718
rect 2956 26682 3012 26684
rect 3036 26682 3092 26684
rect 3116 26682 3172 26684
rect 3196 26682 3252 26684
rect 2956 26630 3002 26682
rect 3002 26630 3012 26682
rect 3036 26630 3066 26682
rect 3066 26630 3078 26682
rect 3078 26630 3092 26682
rect 3116 26630 3130 26682
rect 3130 26630 3142 26682
rect 3142 26630 3172 26682
rect 3196 26630 3206 26682
rect 3206 26630 3252 26682
rect 2956 26628 3012 26630
rect 3036 26628 3092 26630
rect 3116 26628 3172 26630
rect 3196 26628 3252 26630
rect 2956 25594 3012 25596
rect 3036 25594 3092 25596
rect 3116 25594 3172 25596
rect 3196 25594 3252 25596
rect 2956 25542 3002 25594
rect 3002 25542 3012 25594
rect 3036 25542 3066 25594
rect 3066 25542 3078 25594
rect 3078 25542 3092 25594
rect 3116 25542 3130 25594
rect 3130 25542 3142 25594
rect 3142 25542 3172 25594
rect 3196 25542 3206 25594
rect 3206 25542 3252 25594
rect 2956 25540 3012 25542
rect 3036 25540 3092 25542
rect 3116 25540 3172 25542
rect 3196 25540 3252 25542
rect 2956 24506 3012 24508
rect 3036 24506 3092 24508
rect 3116 24506 3172 24508
rect 3196 24506 3252 24508
rect 2956 24454 3002 24506
rect 3002 24454 3012 24506
rect 3036 24454 3066 24506
rect 3066 24454 3078 24506
rect 3078 24454 3092 24506
rect 3116 24454 3130 24506
rect 3130 24454 3142 24506
rect 3142 24454 3172 24506
rect 3196 24454 3206 24506
rect 3206 24454 3252 24506
rect 2956 24452 3012 24454
rect 3036 24452 3092 24454
rect 3116 24452 3172 24454
rect 3196 24452 3252 24454
rect 938 22616 994 22672
rect 2956 23418 3012 23420
rect 3036 23418 3092 23420
rect 3116 23418 3172 23420
rect 3196 23418 3252 23420
rect 2956 23366 3002 23418
rect 3002 23366 3012 23418
rect 3036 23366 3066 23418
rect 3066 23366 3078 23418
rect 3078 23366 3092 23418
rect 3116 23366 3130 23418
rect 3130 23366 3142 23418
rect 3142 23366 3172 23418
rect 3196 23366 3206 23418
rect 3206 23366 3252 23418
rect 2956 23364 3012 23366
rect 3036 23364 3092 23366
rect 3116 23364 3172 23366
rect 3196 23364 3252 23366
rect 2956 22330 3012 22332
rect 3036 22330 3092 22332
rect 3116 22330 3172 22332
rect 3196 22330 3252 22332
rect 2956 22278 3002 22330
rect 3002 22278 3012 22330
rect 3036 22278 3066 22330
rect 3066 22278 3078 22330
rect 3078 22278 3092 22330
rect 3116 22278 3130 22330
rect 3130 22278 3142 22330
rect 3142 22278 3172 22330
rect 3196 22278 3206 22330
rect 3206 22278 3252 22330
rect 2956 22276 3012 22278
rect 3036 22276 3092 22278
rect 3116 22276 3172 22278
rect 3196 22276 3252 22278
rect 1306 20340 1308 20360
rect 1308 20340 1360 20360
rect 1360 20340 1362 20360
rect 1306 20304 1362 20340
rect 1306 17992 1362 18048
rect 2956 21242 3012 21244
rect 3036 21242 3092 21244
rect 3116 21242 3172 21244
rect 3196 21242 3252 21244
rect 2956 21190 3002 21242
rect 3002 21190 3012 21242
rect 3036 21190 3066 21242
rect 3066 21190 3078 21242
rect 3078 21190 3092 21242
rect 3116 21190 3130 21242
rect 3130 21190 3142 21242
rect 3142 21190 3172 21242
rect 3196 21190 3206 21242
rect 3206 21190 3252 21242
rect 2956 21188 3012 21190
rect 3036 21188 3092 21190
rect 3116 21188 3172 21190
rect 3196 21188 3252 21190
rect 2956 20154 3012 20156
rect 3036 20154 3092 20156
rect 3116 20154 3172 20156
rect 3196 20154 3252 20156
rect 2956 20102 3002 20154
rect 3002 20102 3012 20154
rect 3036 20102 3066 20154
rect 3066 20102 3078 20154
rect 3078 20102 3092 20154
rect 3116 20102 3130 20154
rect 3130 20102 3142 20154
rect 3142 20102 3172 20154
rect 3196 20102 3206 20154
rect 3206 20102 3252 20154
rect 2956 20100 3012 20102
rect 3036 20100 3092 20102
rect 3116 20100 3172 20102
rect 3196 20100 3252 20102
rect 2956 19066 3012 19068
rect 3036 19066 3092 19068
rect 3116 19066 3172 19068
rect 3196 19066 3252 19068
rect 2956 19014 3002 19066
rect 3002 19014 3012 19066
rect 3036 19014 3066 19066
rect 3066 19014 3078 19066
rect 3078 19014 3092 19066
rect 3116 19014 3130 19066
rect 3130 19014 3142 19066
rect 3142 19014 3172 19066
rect 3196 19014 3206 19066
rect 3206 19014 3252 19066
rect 2956 19012 3012 19014
rect 3036 19012 3092 19014
rect 3116 19012 3172 19014
rect 3196 19012 3252 19014
rect 1306 15680 1362 15736
rect 1766 13368 1822 13424
rect 2956 17978 3012 17980
rect 3036 17978 3092 17980
rect 3116 17978 3172 17980
rect 3196 17978 3252 17980
rect 2956 17926 3002 17978
rect 3002 17926 3012 17978
rect 3036 17926 3066 17978
rect 3066 17926 3078 17978
rect 3078 17926 3092 17978
rect 3116 17926 3130 17978
rect 3130 17926 3142 17978
rect 3142 17926 3172 17978
rect 3196 17926 3206 17978
rect 3206 17926 3252 17978
rect 2956 17924 3012 17926
rect 3036 17924 3092 17926
rect 3116 17924 3172 17926
rect 3196 17924 3252 17926
rect 2956 16890 3012 16892
rect 3036 16890 3092 16892
rect 3116 16890 3172 16892
rect 3196 16890 3252 16892
rect 2956 16838 3002 16890
rect 3002 16838 3012 16890
rect 3036 16838 3066 16890
rect 3066 16838 3078 16890
rect 3078 16838 3092 16890
rect 3116 16838 3130 16890
rect 3130 16838 3142 16890
rect 3142 16838 3172 16890
rect 3196 16838 3206 16890
rect 3206 16838 3252 16890
rect 2956 16836 3012 16838
rect 3036 16836 3092 16838
rect 3116 16836 3172 16838
rect 3196 16836 3252 16838
rect 2956 15802 3012 15804
rect 3036 15802 3092 15804
rect 3116 15802 3172 15804
rect 3196 15802 3252 15804
rect 2956 15750 3002 15802
rect 3002 15750 3012 15802
rect 3036 15750 3066 15802
rect 3066 15750 3078 15802
rect 3078 15750 3092 15802
rect 3116 15750 3130 15802
rect 3130 15750 3142 15802
rect 3142 15750 3172 15802
rect 3196 15750 3206 15802
rect 3206 15750 3252 15802
rect 2956 15748 3012 15750
rect 3036 15748 3092 15750
rect 3116 15748 3172 15750
rect 3196 15748 3252 15750
rect 2956 14714 3012 14716
rect 3036 14714 3092 14716
rect 3116 14714 3172 14716
rect 3196 14714 3252 14716
rect 2956 14662 3002 14714
rect 3002 14662 3012 14714
rect 3036 14662 3066 14714
rect 3066 14662 3078 14714
rect 3078 14662 3092 14714
rect 3116 14662 3130 14714
rect 3130 14662 3142 14714
rect 3142 14662 3172 14714
rect 3196 14662 3206 14714
rect 3206 14662 3252 14714
rect 2956 14660 3012 14662
rect 3036 14660 3092 14662
rect 3116 14660 3172 14662
rect 3196 14660 3252 14662
rect 2956 13626 3012 13628
rect 3036 13626 3092 13628
rect 3116 13626 3172 13628
rect 3196 13626 3252 13628
rect 2956 13574 3002 13626
rect 3002 13574 3012 13626
rect 3036 13574 3066 13626
rect 3066 13574 3078 13626
rect 3078 13574 3092 13626
rect 3116 13574 3130 13626
rect 3130 13574 3142 13626
rect 3142 13574 3172 13626
rect 3196 13574 3206 13626
rect 3206 13574 3252 13626
rect 2956 13572 3012 13574
rect 3036 13572 3092 13574
rect 3116 13572 3172 13574
rect 3196 13572 3252 13574
rect 2956 12538 3012 12540
rect 3036 12538 3092 12540
rect 3116 12538 3172 12540
rect 3196 12538 3252 12540
rect 2956 12486 3002 12538
rect 3002 12486 3012 12538
rect 3036 12486 3066 12538
rect 3066 12486 3078 12538
rect 3078 12486 3092 12538
rect 3116 12486 3130 12538
rect 3130 12486 3142 12538
rect 3142 12486 3172 12538
rect 3196 12486 3206 12538
rect 3206 12486 3252 12538
rect 2956 12484 3012 12486
rect 3036 12484 3092 12486
rect 3116 12484 3172 12486
rect 3196 12484 3252 12486
rect 2956 11450 3012 11452
rect 3036 11450 3092 11452
rect 3116 11450 3172 11452
rect 3196 11450 3252 11452
rect 2956 11398 3002 11450
rect 3002 11398 3012 11450
rect 3036 11398 3066 11450
rect 3066 11398 3078 11450
rect 3078 11398 3092 11450
rect 3116 11398 3130 11450
rect 3130 11398 3142 11450
rect 3142 11398 3172 11450
rect 3196 11398 3206 11450
rect 3206 11398 3252 11450
rect 2956 11396 3012 11398
rect 3036 11396 3092 11398
rect 3116 11396 3172 11398
rect 3196 11396 3252 11398
rect 3330 11056 3386 11112
rect 2956 10362 3012 10364
rect 3036 10362 3092 10364
rect 3116 10362 3172 10364
rect 3196 10362 3252 10364
rect 2956 10310 3002 10362
rect 3002 10310 3012 10362
rect 3036 10310 3066 10362
rect 3066 10310 3078 10362
rect 3078 10310 3092 10362
rect 3116 10310 3130 10362
rect 3130 10310 3142 10362
rect 3142 10310 3172 10362
rect 3196 10310 3206 10362
rect 3206 10310 3252 10362
rect 2956 10308 3012 10310
rect 3036 10308 3092 10310
rect 3116 10308 3172 10310
rect 3196 10308 3252 10310
rect 2956 9274 3012 9276
rect 3036 9274 3092 9276
rect 3116 9274 3172 9276
rect 3196 9274 3252 9276
rect 2956 9222 3002 9274
rect 3002 9222 3012 9274
rect 3036 9222 3066 9274
rect 3066 9222 3078 9274
rect 3078 9222 3092 9274
rect 3116 9222 3130 9274
rect 3130 9222 3142 9274
rect 3142 9222 3172 9274
rect 3196 9222 3206 9274
rect 3206 9222 3252 9274
rect 2956 9220 3012 9222
rect 3036 9220 3092 9222
rect 3116 9220 3172 9222
rect 3196 9220 3252 9222
rect 2870 8744 2926 8800
rect 2956 8186 3012 8188
rect 3036 8186 3092 8188
rect 3116 8186 3172 8188
rect 3196 8186 3252 8188
rect 2956 8134 3002 8186
rect 3002 8134 3012 8186
rect 3036 8134 3066 8186
rect 3066 8134 3078 8186
rect 3078 8134 3092 8186
rect 3116 8134 3130 8186
rect 3130 8134 3142 8186
rect 3142 8134 3172 8186
rect 3196 8134 3206 8186
rect 3206 8134 3252 8186
rect 2956 8132 3012 8134
rect 3036 8132 3092 8134
rect 3116 8132 3172 8134
rect 3196 8132 3252 8134
rect 2956 7098 3012 7100
rect 3036 7098 3092 7100
rect 3116 7098 3172 7100
rect 3196 7098 3252 7100
rect 2956 7046 3002 7098
rect 3002 7046 3012 7098
rect 3036 7046 3066 7098
rect 3066 7046 3078 7098
rect 3078 7046 3092 7098
rect 3116 7046 3130 7098
rect 3130 7046 3142 7098
rect 3142 7046 3172 7098
rect 3196 7046 3206 7098
rect 3206 7046 3252 7098
rect 2956 7044 3012 7046
rect 3036 7044 3092 7046
rect 3116 7044 3172 7046
rect 3196 7044 3252 7046
rect 3146 6432 3202 6488
rect 2956 6010 3012 6012
rect 3036 6010 3092 6012
rect 3116 6010 3172 6012
rect 3196 6010 3252 6012
rect 2956 5958 3002 6010
rect 3002 5958 3012 6010
rect 3036 5958 3066 6010
rect 3066 5958 3078 6010
rect 3078 5958 3092 6010
rect 3116 5958 3130 6010
rect 3130 5958 3142 6010
rect 3142 5958 3172 6010
rect 3196 5958 3206 6010
rect 3206 5958 3252 6010
rect 2956 5956 3012 5958
rect 3036 5956 3092 5958
rect 3116 5956 3172 5958
rect 3196 5956 3252 5958
rect 2956 4922 3012 4924
rect 3036 4922 3092 4924
rect 3116 4922 3172 4924
rect 3196 4922 3252 4924
rect 2956 4870 3002 4922
rect 3002 4870 3012 4922
rect 3036 4870 3066 4922
rect 3066 4870 3078 4922
rect 3078 4870 3092 4922
rect 3116 4870 3130 4922
rect 3130 4870 3142 4922
rect 3142 4870 3172 4922
rect 3196 4870 3206 4922
rect 3206 4870 3252 4922
rect 2956 4868 3012 4870
rect 3036 4868 3092 4870
rect 3116 4868 3172 4870
rect 3196 4868 3252 4870
rect 3238 4120 3294 4176
rect 2956 3834 3012 3836
rect 3036 3834 3092 3836
rect 3116 3834 3172 3836
rect 3196 3834 3252 3836
rect 2956 3782 3002 3834
rect 3002 3782 3012 3834
rect 3036 3782 3066 3834
rect 3066 3782 3078 3834
rect 3078 3782 3092 3834
rect 3116 3782 3130 3834
rect 3130 3782 3142 3834
rect 3142 3782 3172 3834
rect 3196 3782 3206 3834
rect 3206 3782 3252 3834
rect 2956 3780 3012 3782
rect 3036 3780 3092 3782
rect 3116 3780 3172 3782
rect 3196 3780 3252 3782
rect 2956 2746 3012 2748
rect 3036 2746 3092 2748
rect 3116 2746 3172 2748
rect 3196 2746 3252 2748
rect 2956 2694 3002 2746
rect 3002 2694 3012 2746
rect 3036 2694 3066 2746
rect 3066 2694 3078 2746
rect 3078 2694 3092 2746
rect 3116 2694 3130 2746
rect 3130 2694 3142 2746
rect 3142 2694 3172 2746
rect 3196 2694 3206 2746
rect 3206 2694 3252 2746
rect 2956 2692 3012 2694
rect 3036 2692 3092 2694
rect 3116 2692 3172 2694
rect 3196 2692 3252 2694
rect 2778 1808 2834 1864
rect 7956 54426 8012 54428
rect 8036 54426 8092 54428
rect 8116 54426 8172 54428
rect 8196 54426 8252 54428
rect 7956 54374 8002 54426
rect 8002 54374 8012 54426
rect 8036 54374 8066 54426
rect 8066 54374 8078 54426
rect 8078 54374 8092 54426
rect 8116 54374 8130 54426
rect 8130 54374 8142 54426
rect 8142 54374 8172 54426
rect 8196 54374 8206 54426
rect 8206 54374 8252 54426
rect 7956 54372 8012 54374
rect 8036 54372 8092 54374
rect 8116 54372 8172 54374
rect 8196 54372 8252 54374
rect 7956 53338 8012 53340
rect 8036 53338 8092 53340
rect 8116 53338 8172 53340
rect 8196 53338 8252 53340
rect 7956 53286 8002 53338
rect 8002 53286 8012 53338
rect 8036 53286 8066 53338
rect 8066 53286 8078 53338
rect 8078 53286 8092 53338
rect 8116 53286 8130 53338
rect 8130 53286 8142 53338
rect 8142 53286 8172 53338
rect 8196 53286 8206 53338
rect 8206 53286 8252 53338
rect 7956 53284 8012 53286
rect 8036 53284 8092 53286
rect 8116 53284 8172 53286
rect 8196 53284 8252 53286
rect 7956 52250 8012 52252
rect 8036 52250 8092 52252
rect 8116 52250 8172 52252
rect 8196 52250 8252 52252
rect 7956 52198 8002 52250
rect 8002 52198 8012 52250
rect 8036 52198 8066 52250
rect 8066 52198 8078 52250
rect 8078 52198 8092 52250
rect 8116 52198 8130 52250
rect 8130 52198 8142 52250
rect 8142 52198 8172 52250
rect 8196 52198 8206 52250
rect 8206 52198 8252 52250
rect 7956 52196 8012 52198
rect 8036 52196 8092 52198
rect 8116 52196 8172 52198
rect 8196 52196 8252 52198
rect 7956 51162 8012 51164
rect 8036 51162 8092 51164
rect 8116 51162 8172 51164
rect 8196 51162 8252 51164
rect 7956 51110 8002 51162
rect 8002 51110 8012 51162
rect 8036 51110 8066 51162
rect 8066 51110 8078 51162
rect 8078 51110 8092 51162
rect 8116 51110 8130 51162
rect 8130 51110 8142 51162
rect 8142 51110 8172 51162
rect 8196 51110 8206 51162
rect 8206 51110 8252 51162
rect 7956 51108 8012 51110
rect 8036 51108 8092 51110
rect 8116 51108 8172 51110
rect 8196 51108 8252 51110
rect 7956 50074 8012 50076
rect 8036 50074 8092 50076
rect 8116 50074 8172 50076
rect 8196 50074 8252 50076
rect 7956 50022 8002 50074
rect 8002 50022 8012 50074
rect 8036 50022 8066 50074
rect 8066 50022 8078 50074
rect 8078 50022 8092 50074
rect 8116 50022 8130 50074
rect 8130 50022 8142 50074
rect 8142 50022 8172 50074
rect 8196 50022 8206 50074
rect 8206 50022 8252 50074
rect 7956 50020 8012 50022
rect 8036 50020 8092 50022
rect 8116 50020 8172 50022
rect 8196 50020 8252 50022
rect 7956 48986 8012 48988
rect 8036 48986 8092 48988
rect 8116 48986 8172 48988
rect 8196 48986 8252 48988
rect 7956 48934 8002 48986
rect 8002 48934 8012 48986
rect 8036 48934 8066 48986
rect 8066 48934 8078 48986
rect 8078 48934 8092 48986
rect 8116 48934 8130 48986
rect 8130 48934 8142 48986
rect 8142 48934 8172 48986
rect 8196 48934 8206 48986
rect 8206 48934 8252 48986
rect 7956 48932 8012 48934
rect 8036 48932 8092 48934
rect 8116 48932 8172 48934
rect 8196 48932 8252 48934
rect 7956 47898 8012 47900
rect 8036 47898 8092 47900
rect 8116 47898 8172 47900
rect 8196 47898 8252 47900
rect 7956 47846 8002 47898
rect 8002 47846 8012 47898
rect 8036 47846 8066 47898
rect 8066 47846 8078 47898
rect 8078 47846 8092 47898
rect 8116 47846 8130 47898
rect 8130 47846 8142 47898
rect 8142 47846 8172 47898
rect 8196 47846 8206 47898
rect 8206 47846 8252 47898
rect 7956 47844 8012 47846
rect 8036 47844 8092 47846
rect 8116 47844 8172 47846
rect 8196 47844 8252 47846
rect 7956 46810 8012 46812
rect 8036 46810 8092 46812
rect 8116 46810 8172 46812
rect 8196 46810 8252 46812
rect 7956 46758 8002 46810
rect 8002 46758 8012 46810
rect 8036 46758 8066 46810
rect 8066 46758 8078 46810
rect 8078 46758 8092 46810
rect 8116 46758 8130 46810
rect 8130 46758 8142 46810
rect 8142 46758 8172 46810
rect 8196 46758 8206 46810
rect 8206 46758 8252 46810
rect 7956 46756 8012 46758
rect 8036 46756 8092 46758
rect 8116 46756 8172 46758
rect 8196 46756 8252 46758
rect 7956 45722 8012 45724
rect 8036 45722 8092 45724
rect 8116 45722 8172 45724
rect 8196 45722 8252 45724
rect 7956 45670 8002 45722
rect 8002 45670 8012 45722
rect 8036 45670 8066 45722
rect 8066 45670 8078 45722
rect 8078 45670 8092 45722
rect 8116 45670 8130 45722
rect 8130 45670 8142 45722
rect 8142 45670 8172 45722
rect 8196 45670 8206 45722
rect 8206 45670 8252 45722
rect 7956 45668 8012 45670
rect 8036 45668 8092 45670
rect 8116 45668 8172 45670
rect 8196 45668 8252 45670
rect 7956 44634 8012 44636
rect 8036 44634 8092 44636
rect 8116 44634 8172 44636
rect 8196 44634 8252 44636
rect 7956 44582 8002 44634
rect 8002 44582 8012 44634
rect 8036 44582 8066 44634
rect 8066 44582 8078 44634
rect 8078 44582 8092 44634
rect 8116 44582 8130 44634
rect 8130 44582 8142 44634
rect 8142 44582 8172 44634
rect 8196 44582 8206 44634
rect 8206 44582 8252 44634
rect 7956 44580 8012 44582
rect 8036 44580 8092 44582
rect 8116 44580 8172 44582
rect 8196 44580 8252 44582
rect 7956 43546 8012 43548
rect 8036 43546 8092 43548
rect 8116 43546 8172 43548
rect 8196 43546 8252 43548
rect 7956 43494 8002 43546
rect 8002 43494 8012 43546
rect 8036 43494 8066 43546
rect 8066 43494 8078 43546
rect 8078 43494 8092 43546
rect 8116 43494 8130 43546
rect 8130 43494 8142 43546
rect 8142 43494 8172 43546
rect 8196 43494 8206 43546
rect 8206 43494 8252 43546
rect 7956 43492 8012 43494
rect 8036 43492 8092 43494
rect 8116 43492 8172 43494
rect 8196 43492 8252 43494
rect 7956 42458 8012 42460
rect 8036 42458 8092 42460
rect 8116 42458 8172 42460
rect 8196 42458 8252 42460
rect 7956 42406 8002 42458
rect 8002 42406 8012 42458
rect 8036 42406 8066 42458
rect 8066 42406 8078 42458
rect 8078 42406 8092 42458
rect 8116 42406 8130 42458
rect 8130 42406 8142 42458
rect 8142 42406 8172 42458
rect 8196 42406 8206 42458
rect 8206 42406 8252 42458
rect 7956 42404 8012 42406
rect 8036 42404 8092 42406
rect 8116 42404 8172 42406
rect 8196 42404 8252 42406
rect 7956 41370 8012 41372
rect 8036 41370 8092 41372
rect 8116 41370 8172 41372
rect 8196 41370 8252 41372
rect 7956 41318 8002 41370
rect 8002 41318 8012 41370
rect 8036 41318 8066 41370
rect 8066 41318 8078 41370
rect 8078 41318 8092 41370
rect 8116 41318 8130 41370
rect 8130 41318 8142 41370
rect 8142 41318 8172 41370
rect 8196 41318 8206 41370
rect 8206 41318 8252 41370
rect 7956 41316 8012 41318
rect 8036 41316 8092 41318
rect 8116 41316 8172 41318
rect 8196 41316 8252 41318
rect 7956 40282 8012 40284
rect 8036 40282 8092 40284
rect 8116 40282 8172 40284
rect 8196 40282 8252 40284
rect 7956 40230 8002 40282
rect 8002 40230 8012 40282
rect 8036 40230 8066 40282
rect 8066 40230 8078 40282
rect 8078 40230 8092 40282
rect 8116 40230 8130 40282
rect 8130 40230 8142 40282
rect 8142 40230 8172 40282
rect 8196 40230 8206 40282
rect 8206 40230 8252 40282
rect 7956 40228 8012 40230
rect 8036 40228 8092 40230
rect 8116 40228 8172 40230
rect 8196 40228 8252 40230
rect 7956 39194 8012 39196
rect 8036 39194 8092 39196
rect 8116 39194 8172 39196
rect 8196 39194 8252 39196
rect 7956 39142 8002 39194
rect 8002 39142 8012 39194
rect 8036 39142 8066 39194
rect 8066 39142 8078 39194
rect 8078 39142 8092 39194
rect 8116 39142 8130 39194
rect 8130 39142 8142 39194
rect 8142 39142 8172 39194
rect 8196 39142 8206 39194
rect 8206 39142 8252 39194
rect 7956 39140 8012 39142
rect 8036 39140 8092 39142
rect 8116 39140 8172 39142
rect 8196 39140 8252 39142
rect 7956 38106 8012 38108
rect 8036 38106 8092 38108
rect 8116 38106 8172 38108
rect 8196 38106 8252 38108
rect 7956 38054 8002 38106
rect 8002 38054 8012 38106
rect 8036 38054 8066 38106
rect 8066 38054 8078 38106
rect 8078 38054 8092 38106
rect 8116 38054 8130 38106
rect 8130 38054 8142 38106
rect 8142 38054 8172 38106
rect 8196 38054 8206 38106
rect 8206 38054 8252 38106
rect 7956 38052 8012 38054
rect 8036 38052 8092 38054
rect 8116 38052 8172 38054
rect 8196 38052 8252 38054
rect 7956 37018 8012 37020
rect 8036 37018 8092 37020
rect 8116 37018 8172 37020
rect 8196 37018 8252 37020
rect 7956 36966 8002 37018
rect 8002 36966 8012 37018
rect 8036 36966 8066 37018
rect 8066 36966 8078 37018
rect 8078 36966 8092 37018
rect 8116 36966 8130 37018
rect 8130 36966 8142 37018
rect 8142 36966 8172 37018
rect 8196 36966 8206 37018
rect 8206 36966 8252 37018
rect 7956 36964 8012 36966
rect 8036 36964 8092 36966
rect 8116 36964 8172 36966
rect 8196 36964 8252 36966
rect 7956 35930 8012 35932
rect 8036 35930 8092 35932
rect 8116 35930 8172 35932
rect 8196 35930 8252 35932
rect 7956 35878 8002 35930
rect 8002 35878 8012 35930
rect 8036 35878 8066 35930
rect 8066 35878 8078 35930
rect 8078 35878 8092 35930
rect 8116 35878 8130 35930
rect 8130 35878 8142 35930
rect 8142 35878 8172 35930
rect 8196 35878 8206 35930
rect 8206 35878 8252 35930
rect 7956 35876 8012 35878
rect 8036 35876 8092 35878
rect 8116 35876 8172 35878
rect 8196 35876 8252 35878
rect 7194 31728 7250 31784
rect 7378 31728 7434 31784
rect 7956 34842 8012 34844
rect 8036 34842 8092 34844
rect 8116 34842 8172 34844
rect 8196 34842 8252 34844
rect 7956 34790 8002 34842
rect 8002 34790 8012 34842
rect 8036 34790 8066 34842
rect 8066 34790 8078 34842
rect 8078 34790 8092 34842
rect 8116 34790 8130 34842
rect 8130 34790 8142 34842
rect 8142 34790 8172 34842
rect 8196 34790 8206 34842
rect 8206 34790 8252 34842
rect 7956 34788 8012 34790
rect 8036 34788 8092 34790
rect 8116 34788 8172 34790
rect 8196 34788 8252 34790
rect 9678 44684 9680 44704
rect 9680 44684 9732 44704
rect 9732 44684 9734 44704
rect 9678 44648 9734 44684
rect 9862 36896 9918 36952
rect 8758 35808 8814 35864
rect 7956 33754 8012 33756
rect 8036 33754 8092 33756
rect 8116 33754 8172 33756
rect 8196 33754 8252 33756
rect 7956 33702 8002 33754
rect 8002 33702 8012 33754
rect 8036 33702 8066 33754
rect 8066 33702 8078 33754
rect 8078 33702 8092 33754
rect 8116 33702 8130 33754
rect 8130 33702 8142 33754
rect 8142 33702 8172 33754
rect 8196 33702 8206 33754
rect 8206 33702 8252 33754
rect 7956 33700 8012 33702
rect 8036 33700 8092 33702
rect 8116 33700 8172 33702
rect 8196 33700 8252 33702
rect 7956 32666 8012 32668
rect 8036 32666 8092 32668
rect 8116 32666 8172 32668
rect 8196 32666 8252 32668
rect 7956 32614 8002 32666
rect 8002 32614 8012 32666
rect 8036 32614 8066 32666
rect 8066 32614 8078 32666
rect 8078 32614 8092 32666
rect 8116 32614 8130 32666
rect 8130 32614 8142 32666
rect 8142 32614 8172 32666
rect 8196 32614 8206 32666
rect 8206 32614 8252 32666
rect 7956 32612 8012 32614
rect 8036 32612 8092 32614
rect 8116 32612 8172 32614
rect 8196 32612 8252 32614
rect 7956 31578 8012 31580
rect 8036 31578 8092 31580
rect 8116 31578 8172 31580
rect 8196 31578 8252 31580
rect 7956 31526 8002 31578
rect 8002 31526 8012 31578
rect 8036 31526 8066 31578
rect 8066 31526 8078 31578
rect 8078 31526 8092 31578
rect 8116 31526 8130 31578
rect 8130 31526 8142 31578
rect 8142 31526 8172 31578
rect 8196 31526 8206 31578
rect 8206 31526 8252 31578
rect 7956 31524 8012 31526
rect 8036 31524 8092 31526
rect 8116 31524 8172 31526
rect 8196 31524 8252 31526
rect 7956 30490 8012 30492
rect 8036 30490 8092 30492
rect 8116 30490 8172 30492
rect 8196 30490 8252 30492
rect 7956 30438 8002 30490
rect 8002 30438 8012 30490
rect 8036 30438 8066 30490
rect 8066 30438 8078 30490
rect 8078 30438 8092 30490
rect 8116 30438 8130 30490
rect 8130 30438 8142 30490
rect 8142 30438 8172 30490
rect 8196 30438 8206 30490
rect 8206 30438 8252 30490
rect 7956 30436 8012 30438
rect 8036 30436 8092 30438
rect 8116 30436 8172 30438
rect 8196 30436 8252 30438
rect 7956 29402 8012 29404
rect 8036 29402 8092 29404
rect 8116 29402 8172 29404
rect 8196 29402 8252 29404
rect 7956 29350 8002 29402
rect 8002 29350 8012 29402
rect 8036 29350 8066 29402
rect 8066 29350 8078 29402
rect 8078 29350 8092 29402
rect 8116 29350 8130 29402
rect 8130 29350 8142 29402
rect 8142 29350 8172 29402
rect 8196 29350 8206 29402
rect 8206 29350 8252 29402
rect 7956 29348 8012 29350
rect 8036 29348 8092 29350
rect 8116 29348 8172 29350
rect 8196 29348 8252 29350
rect 7956 28314 8012 28316
rect 8036 28314 8092 28316
rect 8116 28314 8172 28316
rect 8196 28314 8252 28316
rect 7956 28262 8002 28314
rect 8002 28262 8012 28314
rect 8036 28262 8066 28314
rect 8066 28262 8078 28314
rect 8078 28262 8092 28314
rect 8116 28262 8130 28314
rect 8130 28262 8142 28314
rect 8142 28262 8172 28314
rect 8196 28262 8206 28314
rect 8206 28262 8252 28314
rect 7956 28260 8012 28262
rect 8036 28260 8092 28262
rect 8116 28260 8172 28262
rect 8196 28260 8252 28262
rect 7956 27226 8012 27228
rect 8036 27226 8092 27228
rect 8116 27226 8172 27228
rect 8196 27226 8252 27228
rect 7956 27174 8002 27226
rect 8002 27174 8012 27226
rect 8036 27174 8066 27226
rect 8066 27174 8078 27226
rect 8078 27174 8092 27226
rect 8116 27174 8130 27226
rect 8130 27174 8142 27226
rect 8142 27174 8172 27226
rect 8196 27174 8206 27226
rect 8206 27174 8252 27226
rect 7956 27172 8012 27174
rect 8036 27172 8092 27174
rect 8116 27172 8172 27174
rect 8196 27172 8252 27174
rect 7956 26138 8012 26140
rect 8036 26138 8092 26140
rect 8116 26138 8172 26140
rect 8196 26138 8252 26140
rect 7956 26086 8002 26138
rect 8002 26086 8012 26138
rect 8036 26086 8066 26138
rect 8066 26086 8078 26138
rect 8078 26086 8092 26138
rect 8116 26086 8130 26138
rect 8130 26086 8142 26138
rect 8142 26086 8172 26138
rect 8196 26086 8206 26138
rect 8206 26086 8252 26138
rect 7956 26084 8012 26086
rect 8036 26084 8092 26086
rect 8116 26084 8172 26086
rect 8196 26084 8252 26086
rect 7956 25050 8012 25052
rect 8036 25050 8092 25052
rect 8116 25050 8172 25052
rect 8196 25050 8252 25052
rect 7956 24998 8002 25050
rect 8002 24998 8012 25050
rect 8036 24998 8066 25050
rect 8066 24998 8078 25050
rect 8078 24998 8092 25050
rect 8116 24998 8130 25050
rect 8130 24998 8142 25050
rect 8142 24998 8172 25050
rect 8196 24998 8206 25050
rect 8206 24998 8252 25050
rect 7956 24996 8012 24998
rect 8036 24996 8092 24998
rect 8116 24996 8172 24998
rect 8196 24996 8252 24998
rect 7956 23962 8012 23964
rect 8036 23962 8092 23964
rect 8116 23962 8172 23964
rect 8196 23962 8252 23964
rect 7956 23910 8002 23962
rect 8002 23910 8012 23962
rect 8036 23910 8066 23962
rect 8066 23910 8078 23962
rect 8078 23910 8092 23962
rect 8116 23910 8130 23962
rect 8130 23910 8142 23962
rect 8142 23910 8172 23962
rect 8196 23910 8206 23962
rect 8206 23910 8252 23962
rect 7956 23908 8012 23910
rect 8036 23908 8092 23910
rect 8116 23908 8172 23910
rect 8196 23908 8252 23910
rect 7956 22874 8012 22876
rect 8036 22874 8092 22876
rect 8116 22874 8172 22876
rect 8196 22874 8252 22876
rect 7956 22822 8002 22874
rect 8002 22822 8012 22874
rect 8036 22822 8066 22874
rect 8066 22822 8078 22874
rect 8078 22822 8092 22874
rect 8116 22822 8130 22874
rect 8130 22822 8142 22874
rect 8142 22822 8172 22874
rect 8196 22822 8206 22874
rect 8206 22822 8252 22874
rect 7956 22820 8012 22822
rect 8036 22820 8092 22822
rect 8116 22820 8172 22822
rect 8196 22820 8252 22822
rect 7956 21786 8012 21788
rect 8036 21786 8092 21788
rect 8116 21786 8172 21788
rect 8196 21786 8252 21788
rect 7956 21734 8002 21786
rect 8002 21734 8012 21786
rect 8036 21734 8066 21786
rect 8066 21734 8078 21786
rect 8078 21734 8092 21786
rect 8116 21734 8130 21786
rect 8130 21734 8142 21786
rect 8142 21734 8172 21786
rect 8196 21734 8206 21786
rect 8206 21734 8252 21786
rect 7956 21732 8012 21734
rect 8036 21732 8092 21734
rect 8116 21732 8172 21734
rect 8196 21732 8252 21734
rect 7956 20698 8012 20700
rect 8036 20698 8092 20700
rect 8116 20698 8172 20700
rect 8196 20698 8252 20700
rect 7956 20646 8002 20698
rect 8002 20646 8012 20698
rect 8036 20646 8066 20698
rect 8066 20646 8078 20698
rect 8078 20646 8092 20698
rect 8116 20646 8130 20698
rect 8130 20646 8142 20698
rect 8142 20646 8172 20698
rect 8196 20646 8206 20698
rect 8206 20646 8252 20698
rect 7956 20644 8012 20646
rect 8036 20644 8092 20646
rect 8116 20644 8172 20646
rect 8196 20644 8252 20646
rect 7956 19610 8012 19612
rect 8036 19610 8092 19612
rect 8116 19610 8172 19612
rect 8196 19610 8252 19612
rect 7956 19558 8002 19610
rect 8002 19558 8012 19610
rect 8036 19558 8066 19610
rect 8066 19558 8078 19610
rect 8078 19558 8092 19610
rect 8116 19558 8130 19610
rect 8130 19558 8142 19610
rect 8142 19558 8172 19610
rect 8196 19558 8206 19610
rect 8206 19558 8252 19610
rect 7956 19556 8012 19558
rect 8036 19556 8092 19558
rect 8116 19556 8172 19558
rect 8196 19556 8252 19558
rect 7956 18522 8012 18524
rect 8036 18522 8092 18524
rect 8116 18522 8172 18524
rect 8196 18522 8252 18524
rect 7956 18470 8002 18522
rect 8002 18470 8012 18522
rect 8036 18470 8066 18522
rect 8066 18470 8078 18522
rect 8078 18470 8092 18522
rect 8116 18470 8130 18522
rect 8130 18470 8142 18522
rect 8142 18470 8172 18522
rect 8196 18470 8206 18522
rect 8206 18470 8252 18522
rect 7956 18468 8012 18470
rect 8036 18468 8092 18470
rect 8116 18468 8172 18470
rect 8196 18468 8252 18470
rect 7956 17434 8012 17436
rect 8036 17434 8092 17436
rect 8116 17434 8172 17436
rect 8196 17434 8252 17436
rect 7956 17382 8002 17434
rect 8002 17382 8012 17434
rect 8036 17382 8066 17434
rect 8066 17382 8078 17434
rect 8078 17382 8092 17434
rect 8116 17382 8130 17434
rect 8130 17382 8142 17434
rect 8142 17382 8172 17434
rect 8196 17382 8206 17434
rect 8206 17382 8252 17434
rect 7956 17380 8012 17382
rect 8036 17380 8092 17382
rect 8116 17380 8172 17382
rect 8196 17380 8252 17382
rect 7956 16346 8012 16348
rect 8036 16346 8092 16348
rect 8116 16346 8172 16348
rect 8196 16346 8252 16348
rect 7956 16294 8002 16346
rect 8002 16294 8012 16346
rect 8036 16294 8066 16346
rect 8066 16294 8078 16346
rect 8078 16294 8092 16346
rect 8116 16294 8130 16346
rect 8130 16294 8142 16346
rect 8142 16294 8172 16346
rect 8196 16294 8206 16346
rect 8206 16294 8252 16346
rect 7956 16292 8012 16294
rect 8036 16292 8092 16294
rect 8116 16292 8172 16294
rect 8196 16292 8252 16294
rect 7956 15258 8012 15260
rect 8036 15258 8092 15260
rect 8116 15258 8172 15260
rect 8196 15258 8252 15260
rect 7956 15206 8002 15258
rect 8002 15206 8012 15258
rect 8036 15206 8066 15258
rect 8066 15206 8078 15258
rect 8078 15206 8092 15258
rect 8116 15206 8130 15258
rect 8130 15206 8142 15258
rect 8142 15206 8172 15258
rect 8196 15206 8206 15258
rect 8206 15206 8252 15258
rect 7956 15204 8012 15206
rect 8036 15204 8092 15206
rect 8116 15204 8172 15206
rect 8196 15204 8252 15206
rect 7956 14170 8012 14172
rect 8036 14170 8092 14172
rect 8116 14170 8172 14172
rect 8196 14170 8252 14172
rect 7956 14118 8002 14170
rect 8002 14118 8012 14170
rect 8036 14118 8066 14170
rect 8066 14118 8078 14170
rect 8078 14118 8092 14170
rect 8116 14118 8130 14170
rect 8130 14118 8142 14170
rect 8142 14118 8172 14170
rect 8196 14118 8206 14170
rect 8206 14118 8252 14170
rect 7956 14116 8012 14118
rect 8036 14116 8092 14118
rect 8116 14116 8172 14118
rect 8196 14116 8252 14118
rect 7956 13082 8012 13084
rect 8036 13082 8092 13084
rect 8116 13082 8172 13084
rect 8196 13082 8252 13084
rect 7956 13030 8002 13082
rect 8002 13030 8012 13082
rect 8036 13030 8066 13082
rect 8066 13030 8078 13082
rect 8078 13030 8092 13082
rect 8116 13030 8130 13082
rect 8130 13030 8142 13082
rect 8142 13030 8172 13082
rect 8196 13030 8206 13082
rect 8206 13030 8252 13082
rect 7956 13028 8012 13030
rect 8036 13028 8092 13030
rect 8116 13028 8172 13030
rect 8196 13028 8252 13030
rect 7956 11994 8012 11996
rect 8036 11994 8092 11996
rect 8116 11994 8172 11996
rect 8196 11994 8252 11996
rect 7956 11942 8002 11994
rect 8002 11942 8012 11994
rect 8036 11942 8066 11994
rect 8066 11942 8078 11994
rect 8078 11942 8092 11994
rect 8116 11942 8130 11994
rect 8130 11942 8142 11994
rect 8142 11942 8172 11994
rect 8196 11942 8206 11994
rect 8206 11942 8252 11994
rect 7956 11940 8012 11942
rect 8036 11940 8092 11942
rect 8116 11940 8172 11942
rect 8196 11940 8252 11942
rect 7956 10906 8012 10908
rect 8036 10906 8092 10908
rect 8116 10906 8172 10908
rect 8196 10906 8252 10908
rect 7956 10854 8002 10906
rect 8002 10854 8012 10906
rect 8036 10854 8066 10906
rect 8066 10854 8078 10906
rect 8078 10854 8092 10906
rect 8116 10854 8130 10906
rect 8130 10854 8142 10906
rect 8142 10854 8172 10906
rect 8196 10854 8206 10906
rect 8206 10854 8252 10906
rect 7956 10852 8012 10854
rect 8036 10852 8092 10854
rect 8116 10852 8172 10854
rect 8196 10852 8252 10854
rect 7956 9818 8012 9820
rect 8036 9818 8092 9820
rect 8116 9818 8172 9820
rect 8196 9818 8252 9820
rect 7956 9766 8002 9818
rect 8002 9766 8012 9818
rect 8036 9766 8066 9818
rect 8066 9766 8078 9818
rect 8078 9766 8092 9818
rect 8116 9766 8130 9818
rect 8130 9766 8142 9818
rect 8142 9766 8172 9818
rect 8196 9766 8206 9818
rect 8206 9766 8252 9818
rect 7956 9764 8012 9766
rect 8036 9764 8092 9766
rect 8116 9764 8172 9766
rect 8196 9764 8252 9766
rect 7956 8730 8012 8732
rect 8036 8730 8092 8732
rect 8116 8730 8172 8732
rect 8196 8730 8252 8732
rect 7956 8678 8002 8730
rect 8002 8678 8012 8730
rect 8036 8678 8066 8730
rect 8066 8678 8078 8730
rect 8078 8678 8092 8730
rect 8116 8678 8130 8730
rect 8130 8678 8142 8730
rect 8142 8678 8172 8730
rect 8196 8678 8206 8730
rect 8206 8678 8252 8730
rect 7956 8676 8012 8678
rect 8036 8676 8092 8678
rect 8116 8676 8172 8678
rect 8196 8676 8252 8678
rect 7956 7642 8012 7644
rect 8036 7642 8092 7644
rect 8116 7642 8172 7644
rect 8196 7642 8252 7644
rect 7956 7590 8002 7642
rect 8002 7590 8012 7642
rect 8036 7590 8066 7642
rect 8066 7590 8078 7642
rect 8078 7590 8092 7642
rect 8116 7590 8130 7642
rect 8130 7590 8142 7642
rect 8142 7590 8172 7642
rect 8196 7590 8206 7642
rect 8206 7590 8252 7642
rect 7956 7588 8012 7590
rect 8036 7588 8092 7590
rect 8116 7588 8172 7590
rect 8196 7588 8252 7590
rect 7956 6554 8012 6556
rect 8036 6554 8092 6556
rect 8116 6554 8172 6556
rect 8196 6554 8252 6556
rect 7956 6502 8002 6554
rect 8002 6502 8012 6554
rect 8036 6502 8066 6554
rect 8066 6502 8078 6554
rect 8078 6502 8092 6554
rect 8116 6502 8130 6554
rect 8130 6502 8142 6554
rect 8142 6502 8172 6554
rect 8196 6502 8206 6554
rect 8206 6502 8252 6554
rect 7956 6500 8012 6502
rect 8036 6500 8092 6502
rect 8116 6500 8172 6502
rect 8196 6500 8252 6502
rect 7838 5752 7894 5808
rect 7746 5616 7802 5672
rect 7956 5466 8012 5468
rect 8036 5466 8092 5468
rect 8116 5466 8172 5468
rect 8196 5466 8252 5468
rect 7956 5414 8002 5466
rect 8002 5414 8012 5466
rect 8036 5414 8066 5466
rect 8066 5414 8078 5466
rect 8078 5414 8092 5466
rect 8116 5414 8130 5466
rect 8130 5414 8142 5466
rect 8142 5414 8172 5466
rect 8196 5414 8206 5466
rect 8206 5414 8252 5466
rect 7956 5412 8012 5414
rect 8036 5412 8092 5414
rect 8116 5412 8172 5414
rect 8196 5412 8252 5414
rect 7956 4378 8012 4380
rect 8036 4378 8092 4380
rect 8116 4378 8172 4380
rect 8196 4378 8252 4380
rect 7956 4326 8002 4378
rect 8002 4326 8012 4378
rect 8036 4326 8066 4378
rect 8066 4326 8078 4378
rect 8078 4326 8092 4378
rect 8116 4326 8130 4378
rect 8130 4326 8142 4378
rect 8142 4326 8172 4378
rect 8196 4326 8206 4378
rect 8206 4326 8252 4378
rect 7956 4324 8012 4326
rect 8036 4324 8092 4326
rect 8116 4324 8172 4326
rect 8196 4324 8252 4326
rect 7956 3290 8012 3292
rect 8036 3290 8092 3292
rect 8116 3290 8172 3292
rect 8196 3290 8252 3292
rect 7956 3238 8002 3290
rect 8002 3238 8012 3290
rect 8036 3238 8066 3290
rect 8066 3238 8078 3290
rect 8078 3238 8092 3290
rect 8116 3238 8130 3290
rect 8130 3238 8142 3290
rect 8142 3238 8172 3290
rect 8196 3238 8206 3290
rect 8206 3238 8252 3290
rect 7956 3236 8012 3238
rect 8036 3236 8092 3238
rect 8116 3236 8172 3238
rect 8196 3236 8252 3238
rect 7956 2202 8012 2204
rect 8036 2202 8092 2204
rect 8116 2202 8172 2204
rect 8196 2202 8252 2204
rect 7956 2150 8002 2202
rect 8002 2150 8012 2202
rect 8036 2150 8066 2202
rect 8066 2150 8078 2202
rect 8078 2150 8092 2202
rect 8116 2150 8130 2202
rect 8130 2150 8142 2202
rect 8142 2150 8172 2202
rect 8196 2150 8206 2202
rect 8206 2150 8252 2202
rect 7956 2148 8012 2150
rect 8036 2148 8092 2150
rect 8116 2148 8172 2150
rect 8196 2148 8252 2150
rect 10230 31728 10286 31784
rect 9862 31320 9918 31376
rect 12956 53882 13012 53884
rect 13036 53882 13092 53884
rect 13116 53882 13172 53884
rect 13196 53882 13252 53884
rect 12956 53830 13002 53882
rect 13002 53830 13012 53882
rect 13036 53830 13066 53882
rect 13066 53830 13078 53882
rect 13078 53830 13092 53882
rect 13116 53830 13130 53882
rect 13130 53830 13142 53882
rect 13142 53830 13172 53882
rect 13196 53830 13206 53882
rect 13206 53830 13252 53882
rect 12956 53828 13012 53830
rect 13036 53828 13092 53830
rect 13116 53828 13172 53830
rect 13196 53828 13252 53830
rect 12254 45228 12256 45248
rect 12256 45228 12308 45248
rect 12308 45228 12310 45248
rect 12254 45192 12310 45228
rect 11334 41248 11390 41304
rect 10598 30640 10654 30696
rect 10874 31728 10930 31784
rect 12070 37168 12126 37224
rect 12070 33632 12126 33688
rect 11058 21684 11114 21720
rect 11058 21664 11060 21684
rect 11060 21664 11112 21684
rect 11112 21664 11114 21684
rect 11610 24112 11666 24168
rect 11702 21528 11758 21584
rect 11702 21020 11704 21040
rect 11704 21020 11756 21040
rect 11756 21020 11758 21040
rect 11702 20984 11758 21020
rect 12956 52794 13012 52796
rect 13036 52794 13092 52796
rect 13116 52794 13172 52796
rect 13196 52794 13252 52796
rect 12956 52742 13002 52794
rect 13002 52742 13012 52794
rect 13036 52742 13066 52794
rect 13066 52742 13078 52794
rect 13078 52742 13092 52794
rect 13116 52742 13130 52794
rect 13130 52742 13142 52794
rect 13142 52742 13172 52794
rect 13196 52742 13206 52794
rect 13206 52742 13252 52794
rect 12956 52740 13012 52742
rect 13036 52740 13092 52742
rect 13116 52740 13172 52742
rect 13196 52740 13252 52742
rect 12956 51706 13012 51708
rect 13036 51706 13092 51708
rect 13116 51706 13172 51708
rect 13196 51706 13252 51708
rect 12956 51654 13002 51706
rect 13002 51654 13012 51706
rect 13036 51654 13066 51706
rect 13066 51654 13078 51706
rect 13078 51654 13092 51706
rect 13116 51654 13130 51706
rect 13130 51654 13142 51706
rect 13142 51654 13172 51706
rect 13196 51654 13206 51706
rect 13206 51654 13252 51706
rect 12956 51652 13012 51654
rect 13036 51652 13092 51654
rect 13116 51652 13172 51654
rect 13196 51652 13252 51654
rect 12956 50618 13012 50620
rect 13036 50618 13092 50620
rect 13116 50618 13172 50620
rect 13196 50618 13252 50620
rect 12956 50566 13002 50618
rect 13002 50566 13012 50618
rect 13036 50566 13066 50618
rect 13066 50566 13078 50618
rect 13078 50566 13092 50618
rect 13116 50566 13130 50618
rect 13130 50566 13142 50618
rect 13142 50566 13172 50618
rect 13196 50566 13206 50618
rect 13206 50566 13252 50618
rect 12956 50564 13012 50566
rect 13036 50564 13092 50566
rect 13116 50564 13172 50566
rect 13196 50564 13252 50566
rect 12956 49530 13012 49532
rect 13036 49530 13092 49532
rect 13116 49530 13172 49532
rect 13196 49530 13252 49532
rect 12956 49478 13002 49530
rect 13002 49478 13012 49530
rect 13036 49478 13066 49530
rect 13066 49478 13078 49530
rect 13078 49478 13092 49530
rect 13116 49478 13130 49530
rect 13130 49478 13142 49530
rect 13142 49478 13172 49530
rect 13196 49478 13206 49530
rect 13206 49478 13252 49530
rect 12956 49476 13012 49478
rect 13036 49476 13092 49478
rect 13116 49476 13172 49478
rect 13196 49476 13252 49478
rect 12956 48442 13012 48444
rect 13036 48442 13092 48444
rect 13116 48442 13172 48444
rect 13196 48442 13252 48444
rect 12956 48390 13002 48442
rect 13002 48390 13012 48442
rect 13036 48390 13066 48442
rect 13066 48390 13078 48442
rect 13078 48390 13092 48442
rect 13116 48390 13130 48442
rect 13130 48390 13142 48442
rect 13142 48390 13172 48442
rect 13196 48390 13206 48442
rect 13206 48390 13252 48442
rect 12956 48388 13012 48390
rect 13036 48388 13092 48390
rect 13116 48388 13172 48390
rect 13196 48388 13252 48390
rect 12956 47354 13012 47356
rect 13036 47354 13092 47356
rect 13116 47354 13172 47356
rect 13196 47354 13252 47356
rect 12956 47302 13002 47354
rect 13002 47302 13012 47354
rect 13036 47302 13066 47354
rect 13066 47302 13078 47354
rect 13078 47302 13092 47354
rect 13116 47302 13130 47354
rect 13130 47302 13142 47354
rect 13142 47302 13172 47354
rect 13196 47302 13206 47354
rect 13206 47302 13252 47354
rect 12956 47300 13012 47302
rect 13036 47300 13092 47302
rect 13116 47300 13172 47302
rect 13196 47300 13252 47302
rect 12956 46266 13012 46268
rect 13036 46266 13092 46268
rect 13116 46266 13172 46268
rect 13196 46266 13252 46268
rect 12956 46214 13002 46266
rect 13002 46214 13012 46266
rect 13036 46214 13066 46266
rect 13066 46214 13078 46266
rect 13078 46214 13092 46266
rect 13116 46214 13130 46266
rect 13130 46214 13142 46266
rect 13142 46214 13172 46266
rect 13196 46214 13206 46266
rect 13206 46214 13252 46266
rect 12956 46212 13012 46214
rect 13036 46212 13092 46214
rect 13116 46212 13172 46214
rect 13196 46212 13252 46214
rect 12956 45178 13012 45180
rect 13036 45178 13092 45180
rect 13116 45178 13172 45180
rect 13196 45178 13252 45180
rect 12956 45126 13002 45178
rect 13002 45126 13012 45178
rect 13036 45126 13066 45178
rect 13066 45126 13078 45178
rect 13078 45126 13092 45178
rect 13116 45126 13130 45178
rect 13130 45126 13142 45178
rect 13142 45126 13172 45178
rect 13196 45126 13206 45178
rect 13206 45126 13252 45178
rect 12956 45124 13012 45126
rect 13036 45124 13092 45126
rect 13116 45124 13172 45126
rect 13196 45124 13252 45126
rect 12956 44090 13012 44092
rect 13036 44090 13092 44092
rect 13116 44090 13172 44092
rect 13196 44090 13252 44092
rect 12956 44038 13002 44090
rect 13002 44038 13012 44090
rect 13036 44038 13066 44090
rect 13066 44038 13078 44090
rect 13078 44038 13092 44090
rect 13116 44038 13130 44090
rect 13130 44038 13142 44090
rect 13142 44038 13172 44090
rect 13196 44038 13206 44090
rect 13206 44038 13252 44090
rect 12956 44036 13012 44038
rect 13036 44036 13092 44038
rect 13116 44036 13172 44038
rect 13196 44036 13252 44038
rect 12956 43002 13012 43004
rect 13036 43002 13092 43004
rect 13116 43002 13172 43004
rect 13196 43002 13252 43004
rect 12956 42950 13002 43002
rect 13002 42950 13012 43002
rect 13036 42950 13066 43002
rect 13066 42950 13078 43002
rect 13078 42950 13092 43002
rect 13116 42950 13130 43002
rect 13130 42950 13142 43002
rect 13142 42950 13172 43002
rect 13196 42950 13206 43002
rect 13206 42950 13252 43002
rect 12956 42948 13012 42950
rect 13036 42948 13092 42950
rect 13116 42948 13172 42950
rect 13196 42948 13252 42950
rect 12956 41914 13012 41916
rect 13036 41914 13092 41916
rect 13116 41914 13172 41916
rect 13196 41914 13252 41916
rect 12956 41862 13002 41914
rect 13002 41862 13012 41914
rect 13036 41862 13066 41914
rect 13066 41862 13078 41914
rect 13078 41862 13092 41914
rect 13116 41862 13130 41914
rect 13130 41862 13142 41914
rect 13142 41862 13172 41914
rect 13196 41862 13206 41914
rect 13206 41862 13252 41914
rect 12956 41860 13012 41862
rect 13036 41860 13092 41862
rect 13116 41860 13172 41862
rect 13196 41860 13252 41862
rect 12956 40826 13012 40828
rect 13036 40826 13092 40828
rect 13116 40826 13172 40828
rect 13196 40826 13252 40828
rect 12956 40774 13002 40826
rect 13002 40774 13012 40826
rect 13036 40774 13066 40826
rect 13066 40774 13078 40826
rect 13078 40774 13092 40826
rect 13116 40774 13130 40826
rect 13130 40774 13142 40826
rect 13142 40774 13172 40826
rect 13196 40774 13206 40826
rect 13206 40774 13252 40826
rect 12956 40772 13012 40774
rect 13036 40772 13092 40774
rect 13116 40772 13172 40774
rect 13196 40772 13252 40774
rect 13450 40704 13506 40760
rect 12956 39738 13012 39740
rect 13036 39738 13092 39740
rect 13116 39738 13172 39740
rect 13196 39738 13252 39740
rect 12956 39686 13002 39738
rect 13002 39686 13012 39738
rect 13036 39686 13066 39738
rect 13066 39686 13078 39738
rect 13078 39686 13092 39738
rect 13116 39686 13130 39738
rect 13130 39686 13142 39738
rect 13142 39686 13172 39738
rect 13196 39686 13206 39738
rect 13206 39686 13252 39738
rect 12956 39684 13012 39686
rect 13036 39684 13092 39686
rect 13116 39684 13172 39686
rect 13196 39684 13252 39686
rect 12956 38650 13012 38652
rect 13036 38650 13092 38652
rect 13116 38650 13172 38652
rect 13196 38650 13252 38652
rect 12956 38598 13002 38650
rect 13002 38598 13012 38650
rect 13036 38598 13066 38650
rect 13066 38598 13078 38650
rect 13078 38598 13092 38650
rect 13116 38598 13130 38650
rect 13130 38598 13142 38650
rect 13142 38598 13172 38650
rect 13196 38598 13206 38650
rect 13206 38598 13252 38650
rect 12956 38596 13012 38598
rect 13036 38596 13092 38598
rect 13116 38596 13172 38598
rect 13196 38596 13252 38598
rect 12956 37562 13012 37564
rect 13036 37562 13092 37564
rect 13116 37562 13172 37564
rect 13196 37562 13252 37564
rect 12956 37510 13002 37562
rect 13002 37510 13012 37562
rect 13036 37510 13066 37562
rect 13066 37510 13078 37562
rect 13078 37510 13092 37562
rect 13116 37510 13130 37562
rect 13130 37510 13142 37562
rect 13142 37510 13172 37562
rect 13196 37510 13206 37562
rect 13206 37510 13252 37562
rect 12956 37508 13012 37510
rect 13036 37508 13092 37510
rect 13116 37508 13172 37510
rect 13196 37508 13252 37510
rect 12956 36474 13012 36476
rect 13036 36474 13092 36476
rect 13116 36474 13172 36476
rect 13196 36474 13252 36476
rect 12956 36422 13002 36474
rect 13002 36422 13012 36474
rect 13036 36422 13066 36474
rect 13066 36422 13078 36474
rect 13078 36422 13092 36474
rect 13116 36422 13130 36474
rect 13130 36422 13142 36474
rect 13142 36422 13172 36474
rect 13196 36422 13206 36474
rect 13206 36422 13252 36474
rect 12956 36420 13012 36422
rect 13036 36420 13092 36422
rect 13116 36420 13172 36422
rect 13196 36420 13252 36422
rect 12956 35386 13012 35388
rect 13036 35386 13092 35388
rect 13116 35386 13172 35388
rect 13196 35386 13252 35388
rect 12956 35334 13002 35386
rect 13002 35334 13012 35386
rect 13036 35334 13066 35386
rect 13066 35334 13078 35386
rect 13078 35334 13092 35386
rect 13116 35334 13130 35386
rect 13130 35334 13142 35386
rect 13142 35334 13172 35386
rect 13196 35334 13206 35386
rect 13206 35334 13252 35386
rect 12956 35332 13012 35334
rect 13036 35332 13092 35334
rect 13116 35332 13172 35334
rect 13196 35332 13252 35334
rect 12714 35128 12770 35184
rect 12346 29416 12402 29472
rect 12956 34298 13012 34300
rect 13036 34298 13092 34300
rect 13116 34298 13172 34300
rect 13196 34298 13252 34300
rect 12956 34246 13002 34298
rect 13002 34246 13012 34298
rect 13036 34246 13066 34298
rect 13066 34246 13078 34298
rect 13078 34246 13092 34298
rect 13116 34246 13130 34298
rect 13130 34246 13142 34298
rect 13142 34246 13172 34298
rect 13196 34246 13206 34298
rect 13206 34246 13252 34298
rect 12956 34244 13012 34246
rect 13036 34244 13092 34246
rect 13116 34244 13172 34246
rect 13196 34244 13252 34246
rect 14370 52536 14426 52592
rect 12956 33210 13012 33212
rect 13036 33210 13092 33212
rect 13116 33210 13172 33212
rect 13196 33210 13252 33212
rect 12956 33158 13002 33210
rect 13002 33158 13012 33210
rect 13036 33158 13066 33210
rect 13066 33158 13078 33210
rect 13078 33158 13092 33210
rect 13116 33158 13130 33210
rect 13130 33158 13142 33210
rect 13142 33158 13172 33210
rect 13196 33158 13206 33210
rect 13206 33158 13252 33210
rect 12956 33156 13012 33158
rect 13036 33156 13092 33158
rect 13116 33156 13172 33158
rect 13196 33156 13252 33158
rect 12956 32122 13012 32124
rect 13036 32122 13092 32124
rect 13116 32122 13172 32124
rect 13196 32122 13252 32124
rect 12956 32070 13002 32122
rect 13002 32070 13012 32122
rect 13036 32070 13066 32122
rect 13066 32070 13078 32122
rect 13078 32070 13092 32122
rect 13116 32070 13130 32122
rect 13130 32070 13142 32122
rect 13142 32070 13172 32122
rect 13196 32070 13206 32122
rect 13206 32070 13252 32122
rect 12956 32068 13012 32070
rect 13036 32068 13092 32070
rect 13116 32068 13172 32070
rect 13196 32068 13252 32070
rect 12956 31034 13012 31036
rect 13036 31034 13092 31036
rect 13116 31034 13172 31036
rect 13196 31034 13252 31036
rect 12956 30982 13002 31034
rect 13002 30982 13012 31034
rect 13036 30982 13066 31034
rect 13066 30982 13078 31034
rect 13078 30982 13092 31034
rect 13116 30982 13130 31034
rect 13130 30982 13142 31034
rect 13142 30982 13172 31034
rect 13196 30982 13206 31034
rect 13206 30982 13252 31034
rect 12956 30980 13012 30982
rect 13036 30980 13092 30982
rect 13116 30980 13172 30982
rect 13196 30980 13252 30982
rect 12990 30368 13046 30424
rect 12956 29946 13012 29948
rect 13036 29946 13092 29948
rect 13116 29946 13172 29948
rect 13196 29946 13252 29948
rect 12956 29894 13002 29946
rect 13002 29894 13012 29946
rect 13036 29894 13066 29946
rect 13066 29894 13078 29946
rect 13078 29894 13092 29946
rect 13116 29894 13130 29946
rect 13130 29894 13142 29946
rect 13142 29894 13172 29946
rect 13196 29894 13206 29946
rect 13206 29894 13252 29946
rect 12956 29892 13012 29894
rect 13036 29892 13092 29894
rect 13116 29892 13172 29894
rect 13196 29892 13252 29894
rect 14002 35284 14058 35320
rect 14002 35264 14004 35284
rect 14004 35264 14056 35284
rect 14056 35264 14058 35284
rect 14002 33360 14058 33416
rect 12956 28858 13012 28860
rect 13036 28858 13092 28860
rect 13116 28858 13172 28860
rect 13196 28858 13252 28860
rect 12956 28806 13002 28858
rect 13002 28806 13012 28858
rect 13036 28806 13066 28858
rect 13066 28806 13078 28858
rect 13078 28806 13092 28858
rect 13116 28806 13130 28858
rect 13130 28806 13142 28858
rect 13142 28806 13172 28858
rect 13196 28806 13206 28858
rect 13206 28806 13252 28858
rect 12956 28804 13012 28806
rect 13036 28804 13092 28806
rect 13116 28804 13172 28806
rect 13196 28804 13252 28806
rect 12956 27770 13012 27772
rect 13036 27770 13092 27772
rect 13116 27770 13172 27772
rect 13196 27770 13252 27772
rect 12956 27718 13002 27770
rect 13002 27718 13012 27770
rect 13036 27718 13066 27770
rect 13066 27718 13078 27770
rect 13078 27718 13092 27770
rect 13116 27718 13130 27770
rect 13130 27718 13142 27770
rect 13142 27718 13172 27770
rect 13196 27718 13206 27770
rect 13206 27718 13252 27770
rect 12956 27716 13012 27718
rect 13036 27716 13092 27718
rect 13116 27716 13172 27718
rect 13196 27716 13252 27718
rect 12956 26682 13012 26684
rect 13036 26682 13092 26684
rect 13116 26682 13172 26684
rect 13196 26682 13252 26684
rect 12956 26630 13002 26682
rect 13002 26630 13012 26682
rect 13036 26630 13066 26682
rect 13066 26630 13078 26682
rect 13078 26630 13092 26682
rect 13116 26630 13130 26682
rect 13130 26630 13142 26682
rect 13142 26630 13172 26682
rect 13196 26630 13206 26682
rect 13206 26630 13252 26682
rect 12956 26628 13012 26630
rect 13036 26628 13092 26630
rect 13116 26628 13172 26630
rect 13196 26628 13252 26630
rect 12956 25594 13012 25596
rect 13036 25594 13092 25596
rect 13116 25594 13172 25596
rect 13196 25594 13252 25596
rect 12956 25542 13002 25594
rect 13002 25542 13012 25594
rect 13036 25542 13066 25594
rect 13066 25542 13078 25594
rect 13078 25542 13092 25594
rect 13116 25542 13130 25594
rect 13130 25542 13142 25594
rect 13142 25542 13172 25594
rect 13196 25542 13206 25594
rect 13206 25542 13252 25594
rect 12956 25540 13012 25542
rect 13036 25540 13092 25542
rect 13116 25540 13172 25542
rect 13196 25540 13252 25542
rect 12070 15272 12126 15328
rect 12530 22652 12532 22672
rect 12532 22652 12584 22672
rect 12584 22652 12586 22672
rect 12530 22616 12586 22652
rect 12956 24506 13012 24508
rect 13036 24506 13092 24508
rect 13116 24506 13172 24508
rect 13196 24506 13252 24508
rect 12956 24454 13002 24506
rect 13002 24454 13012 24506
rect 13036 24454 13066 24506
rect 13066 24454 13078 24506
rect 13078 24454 13092 24506
rect 13116 24454 13130 24506
rect 13130 24454 13142 24506
rect 13142 24454 13172 24506
rect 13196 24454 13206 24506
rect 13206 24454 13252 24506
rect 12956 24452 13012 24454
rect 13036 24452 13092 24454
rect 13116 24452 13172 24454
rect 13196 24452 13252 24454
rect 12956 23418 13012 23420
rect 13036 23418 13092 23420
rect 13116 23418 13172 23420
rect 13196 23418 13252 23420
rect 12956 23366 13002 23418
rect 13002 23366 13012 23418
rect 13036 23366 13066 23418
rect 13066 23366 13078 23418
rect 13078 23366 13092 23418
rect 13116 23366 13130 23418
rect 13130 23366 13142 23418
rect 13142 23366 13172 23418
rect 13196 23366 13206 23418
rect 13206 23366 13252 23418
rect 12956 23364 13012 23366
rect 13036 23364 13092 23366
rect 13116 23364 13172 23366
rect 13196 23364 13252 23366
rect 13726 23316 13782 23352
rect 13726 23296 13728 23316
rect 13728 23296 13780 23316
rect 13780 23296 13782 23316
rect 13174 22516 13176 22536
rect 13176 22516 13228 22536
rect 13228 22516 13230 22536
rect 13174 22480 13230 22516
rect 12956 22330 13012 22332
rect 13036 22330 13092 22332
rect 13116 22330 13172 22332
rect 13196 22330 13252 22332
rect 12956 22278 13002 22330
rect 13002 22278 13012 22330
rect 13036 22278 13066 22330
rect 13066 22278 13078 22330
rect 13078 22278 13092 22330
rect 13116 22278 13130 22330
rect 13130 22278 13142 22330
rect 13142 22278 13172 22330
rect 13196 22278 13206 22330
rect 13206 22278 13252 22330
rect 12956 22276 13012 22278
rect 13036 22276 13092 22278
rect 13116 22276 13172 22278
rect 13196 22276 13252 22278
rect 12898 21428 12900 21448
rect 12900 21428 12952 21448
rect 12952 21428 12954 21448
rect 12898 21392 12954 21428
rect 12956 21242 13012 21244
rect 13036 21242 13092 21244
rect 13116 21242 13172 21244
rect 13196 21242 13252 21244
rect 12956 21190 13002 21242
rect 13002 21190 13012 21242
rect 13036 21190 13066 21242
rect 13066 21190 13078 21242
rect 13078 21190 13092 21242
rect 13116 21190 13130 21242
rect 13130 21190 13142 21242
rect 13142 21190 13172 21242
rect 13196 21190 13206 21242
rect 13206 21190 13252 21242
rect 12956 21188 13012 21190
rect 13036 21188 13092 21190
rect 13116 21188 13172 21190
rect 13196 21188 13252 21190
rect 13450 20984 13506 21040
rect 13818 21836 13820 21856
rect 13820 21836 13872 21856
rect 13872 21836 13874 21856
rect 12956 20154 13012 20156
rect 13036 20154 13092 20156
rect 13116 20154 13172 20156
rect 13196 20154 13252 20156
rect 12956 20102 13002 20154
rect 13002 20102 13012 20154
rect 13036 20102 13066 20154
rect 13066 20102 13078 20154
rect 13078 20102 13092 20154
rect 13116 20102 13130 20154
rect 13130 20102 13142 20154
rect 13142 20102 13172 20154
rect 13196 20102 13206 20154
rect 13206 20102 13252 20154
rect 12956 20100 13012 20102
rect 13036 20100 13092 20102
rect 13116 20100 13172 20102
rect 13196 20100 13252 20102
rect 12956 19066 13012 19068
rect 13036 19066 13092 19068
rect 13116 19066 13172 19068
rect 13196 19066 13252 19068
rect 12956 19014 13002 19066
rect 13002 19014 13012 19066
rect 13036 19014 13066 19066
rect 13066 19014 13078 19066
rect 13078 19014 13092 19066
rect 13116 19014 13130 19066
rect 13130 19014 13142 19066
rect 13142 19014 13172 19066
rect 13196 19014 13206 19066
rect 13206 19014 13252 19066
rect 12956 19012 13012 19014
rect 13036 19012 13092 19014
rect 13116 19012 13172 19014
rect 13196 19012 13252 19014
rect 12956 17978 13012 17980
rect 13036 17978 13092 17980
rect 13116 17978 13172 17980
rect 13196 17978 13252 17980
rect 12956 17926 13002 17978
rect 13002 17926 13012 17978
rect 13036 17926 13066 17978
rect 13066 17926 13078 17978
rect 13078 17926 13092 17978
rect 13116 17926 13130 17978
rect 13130 17926 13142 17978
rect 13142 17926 13172 17978
rect 13196 17926 13206 17978
rect 13206 17926 13252 17978
rect 12956 17924 13012 17926
rect 13036 17924 13092 17926
rect 13116 17924 13172 17926
rect 13196 17924 13252 17926
rect 12806 17876 12862 17912
rect 12806 17856 12808 17876
rect 12808 17856 12860 17876
rect 12860 17856 12862 17876
rect 12956 16890 13012 16892
rect 13036 16890 13092 16892
rect 13116 16890 13172 16892
rect 13196 16890 13252 16892
rect 12956 16838 13002 16890
rect 13002 16838 13012 16890
rect 13036 16838 13066 16890
rect 13066 16838 13078 16890
rect 13078 16838 13092 16890
rect 13116 16838 13130 16890
rect 13130 16838 13142 16890
rect 13142 16838 13172 16890
rect 13196 16838 13206 16890
rect 13206 16838 13252 16890
rect 12956 16836 13012 16838
rect 13036 16836 13092 16838
rect 13116 16836 13172 16838
rect 13196 16836 13252 16838
rect 12806 15952 12862 16008
rect 12956 15802 13012 15804
rect 13036 15802 13092 15804
rect 13116 15802 13172 15804
rect 13196 15802 13252 15804
rect 12956 15750 13002 15802
rect 13002 15750 13012 15802
rect 13036 15750 13066 15802
rect 13066 15750 13078 15802
rect 13078 15750 13092 15802
rect 13116 15750 13130 15802
rect 13130 15750 13142 15802
rect 13142 15750 13172 15802
rect 13196 15750 13206 15802
rect 13206 15750 13252 15802
rect 12956 15748 13012 15750
rect 13036 15748 13092 15750
rect 13116 15748 13172 15750
rect 13196 15748 13252 15750
rect 12956 14714 13012 14716
rect 13036 14714 13092 14716
rect 13116 14714 13172 14716
rect 13196 14714 13252 14716
rect 12956 14662 13002 14714
rect 13002 14662 13012 14714
rect 13036 14662 13066 14714
rect 13066 14662 13078 14714
rect 13078 14662 13092 14714
rect 13116 14662 13130 14714
rect 13130 14662 13142 14714
rect 13142 14662 13172 14714
rect 13196 14662 13206 14714
rect 13206 14662 13252 14714
rect 12956 14660 13012 14662
rect 13036 14660 13092 14662
rect 13116 14660 13172 14662
rect 13196 14660 13252 14662
rect 12956 13626 13012 13628
rect 13036 13626 13092 13628
rect 13116 13626 13172 13628
rect 13196 13626 13252 13628
rect 12956 13574 13002 13626
rect 13002 13574 13012 13626
rect 13036 13574 13066 13626
rect 13066 13574 13078 13626
rect 13078 13574 13092 13626
rect 13116 13574 13130 13626
rect 13130 13574 13142 13626
rect 13142 13574 13172 13626
rect 13196 13574 13206 13626
rect 13206 13574 13252 13626
rect 12956 13572 13012 13574
rect 13036 13572 13092 13574
rect 13116 13572 13172 13574
rect 13196 13572 13252 13574
rect 13818 21800 13874 21836
rect 12956 12538 13012 12540
rect 13036 12538 13092 12540
rect 13116 12538 13172 12540
rect 13196 12538 13252 12540
rect 12956 12486 13002 12538
rect 13002 12486 13012 12538
rect 13036 12486 13066 12538
rect 13066 12486 13078 12538
rect 13078 12486 13092 12538
rect 13116 12486 13130 12538
rect 13130 12486 13142 12538
rect 13142 12486 13172 12538
rect 13196 12486 13206 12538
rect 13206 12486 13252 12538
rect 12956 12484 13012 12486
rect 13036 12484 13092 12486
rect 13116 12484 13172 12486
rect 13196 12484 13252 12486
rect 12956 11450 13012 11452
rect 13036 11450 13092 11452
rect 13116 11450 13172 11452
rect 13196 11450 13252 11452
rect 12956 11398 13002 11450
rect 13002 11398 13012 11450
rect 13036 11398 13066 11450
rect 13066 11398 13078 11450
rect 13078 11398 13092 11450
rect 13116 11398 13130 11450
rect 13130 11398 13142 11450
rect 13142 11398 13172 11450
rect 13196 11398 13206 11450
rect 13206 11398 13252 11450
rect 12956 11396 13012 11398
rect 13036 11396 13092 11398
rect 13116 11396 13172 11398
rect 13196 11396 13252 11398
rect 12956 10362 13012 10364
rect 13036 10362 13092 10364
rect 13116 10362 13172 10364
rect 13196 10362 13252 10364
rect 12956 10310 13002 10362
rect 13002 10310 13012 10362
rect 13036 10310 13066 10362
rect 13066 10310 13078 10362
rect 13078 10310 13092 10362
rect 13116 10310 13130 10362
rect 13130 10310 13142 10362
rect 13142 10310 13172 10362
rect 13196 10310 13206 10362
rect 13206 10310 13252 10362
rect 12956 10308 13012 10310
rect 13036 10308 13092 10310
rect 13116 10308 13172 10310
rect 13196 10308 13252 10310
rect 12956 9274 13012 9276
rect 13036 9274 13092 9276
rect 13116 9274 13172 9276
rect 13196 9274 13252 9276
rect 12956 9222 13002 9274
rect 13002 9222 13012 9274
rect 13036 9222 13066 9274
rect 13066 9222 13078 9274
rect 13078 9222 13092 9274
rect 13116 9222 13130 9274
rect 13130 9222 13142 9274
rect 13142 9222 13172 9274
rect 13196 9222 13206 9274
rect 13206 9222 13252 9274
rect 12956 9220 13012 9222
rect 13036 9220 13092 9222
rect 13116 9220 13172 9222
rect 13196 9220 13252 9222
rect 12956 8186 13012 8188
rect 13036 8186 13092 8188
rect 13116 8186 13172 8188
rect 13196 8186 13252 8188
rect 12956 8134 13002 8186
rect 13002 8134 13012 8186
rect 13036 8134 13066 8186
rect 13066 8134 13078 8186
rect 13078 8134 13092 8186
rect 13116 8134 13130 8186
rect 13130 8134 13142 8186
rect 13142 8134 13172 8186
rect 13196 8134 13206 8186
rect 13206 8134 13252 8186
rect 12956 8132 13012 8134
rect 13036 8132 13092 8134
rect 13116 8132 13172 8134
rect 13196 8132 13252 8134
rect 12956 7098 13012 7100
rect 13036 7098 13092 7100
rect 13116 7098 13172 7100
rect 13196 7098 13252 7100
rect 12956 7046 13002 7098
rect 13002 7046 13012 7098
rect 13036 7046 13066 7098
rect 13066 7046 13078 7098
rect 13078 7046 13092 7098
rect 13116 7046 13130 7098
rect 13130 7046 13142 7098
rect 13142 7046 13172 7098
rect 13196 7046 13206 7098
rect 13206 7046 13252 7098
rect 12956 7044 13012 7046
rect 13036 7044 13092 7046
rect 13116 7044 13172 7046
rect 13196 7044 13252 7046
rect 12956 6010 13012 6012
rect 13036 6010 13092 6012
rect 13116 6010 13172 6012
rect 13196 6010 13252 6012
rect 12956 5958 13002 6010
rect 13002 5958 13012 6010
rect 13036 5958 13066 6010
rect 13066 5958 13078 6010
rect 13078 5958 13092 6010
rect 13116 5958 13130 6010
rect 13130 5958 13142 6010
rect 13142 5958 13172 6010
rect 13196 5958 13206 6010
rect 13206 5958 13252 6010
rect 12956 5956 13012 5958
rect 13036 5956 13092 5958
rect 13116 5956 13172 5958
rect 13196 5956 13252 5958
rect 12956 4922 13012 4924
rect 13036 4922 13092 4924
rect 13116 4922 13172 4924
rect 13196 4922 13252 4924
rect 12956 4870 13002 4922
rect 13002 4870 13012 4922
rect 13036 4870 13066 4922
rect 13066 4870 13078 4922
rect 13078 4870 13092 4922
rect 13116 4870 13130 4922
rect 13130 4870 13142 4922
rect 13142 4870 13172 4922
rect 13196 4870 13206 4922
rect 13206 4870 13252 4922
rect 12956 4868 13012 4870
rect 13036 4868 13092 4870
rect 13116 4868 13172 4870
rect 13196 4868 13252 4870
rect 12956 3834 13012 3836
rect 13036 3834 13092 3836
rect 13116 3834 13172 3836
rect 13196 3834 13252 3836
rect 12956 3782 13002 3834
rect 13002 3782 13012 3834
rect 13036 3782 13066 3834
rect 13066 3782 13078 3834
rect 13078 3782 13092 3834
rect 13116 3782 13130 3834
rect 13130 3782 13142 3834
rect 13142 3782 13172 3834
rect 13196 3782 13206 3834
rect 13206 3782 13252 3834
rect 12956 3780 13012 3782
rect 13036 3780 13092 3782
rect 13116 3780 13172 3782
rect 13196 3780 13252 3782
rect 14554 36760 14610 36816
rect 14462 34448 14518 34504
rect 15658 53896 15714 53952
rect 15290 38700 15292 38720
rect 15292 38700 15344 38720
rect 15344 38700 15346 38720
rect 15290 38664 15346 38700
rect 14738 29008 14794 29064
rect 14738 21836 14740 21856
rect 14740 21836 14792 21856
rect 14792 21836 14794 21856
rect 14738 21800 14794 21836
rect 14554 21392 14610 21448
rect 14646 20168 14702 20224
rect 12956 2746 13012 2748
rect 13036 2746 13092 2748
rect 13116 2746 13172 2748
rect 13196 2746 13252 2748
rect 12956 2694 13002 2746
rect 13002 2694 13012 2746
rect 13036 2694 13066 2746
rect 13066 2694 13078 2746
rect 13078 2694 13092 2746
rect 13116 2694 13130 2746
rect 13130 2694 13142 2746
rect 13142 2694 13172 2746
rect 13196 2694 13206 2746
rect 13206 2694 13252 2746
rect 12956 2692 13012 2694
rect 13036 2692 13092 2694
rect 13116 2692 13172 2694
rect 13196 2692 13252 2694
rect 15382 35808 15438 35864
rect 15934 52536 15990 52592
rect 16118 29996 16120 30016
rect 16120 29996 16172 30016
rect 16172 29996 16174 30016
rect 16118 29960 16174 29996
rect 15750 27124 15806 27160
rect 15750 27104 15752 27124
rect 15752 27104 15804 27124
rect 15804 27104 15806 27124
rect 15566 21664 15622 21720
rect 15474 21548 15530 21584
rect 15474 21528 15476 21548
rect 15476 21528 15528 21548
rect 15528 21528 15530 21548
rect 17956 54426 18012 54428
rect 18036 54426 18092 54428
rect 18116 54426 18172 54428
rect 18196 54426 18252 54428
rect 17956 54374 18002 54426
rect 18002 54374 18012 54426
rect 18036 54374 18066 54426
rect 18066 54374 18078 54426
rect 18078 54374 18092 54426
rect 18116 54374 18130 54426
rect 18130 54374 18142 54426
rect 18142 54374 18172 54426
rect 18196 54374 18206 54426
rect 18206 54374 18252 54426
rect 17956 54372 18012 54374
rect 18036 54372 18092 54374
rect 18116 54372 18172 54374
rect 18196 54372 18252 54374
rect 17956 53338 18012 53340
rect 18036 53338 18092 53340
rect 18116 53338 18172 53340
rect 18196 53338 18252 53340
rect 17956 53286 18002 53338
rect 18002 53286 18012 53338
rect 18036 53286 18066 53338
rect 18066 53286 18078 53338
rect 18078 53286 18092 53338
rect 18116 53286 18130 53338
rect 18130 53286 18142 53338
rect 18142 53286 18172 53338
rect 18196 53286 18206 53338
rect 18206 53286 18252 53338
rect 17956 53284 18012 53286
rect 18036 53284 18092 53286
rect 18116 53284 18172 53286
rect 18196 53284 18252 53286
rect 17956 52250 18012 52252
rect 18036 52250 18092 52252
rect 18116 52250 18172 52252
rect 18196 52250 18252 52252
rect 17956 52198 18002 52250
rect 18002 52198 18012 52250
rect 18036 52198 18066 52250
rect 18066 52198 18078 52250
rect 18078 52198 18092 52250
rect 18116 52198 18130 52250
rect 18130 52198 18142 52250
rect 18142 52198 18172 52250
rect 18196 52198 18206 52250
rect 18206 52198 18252 52250
rect 17956 52196 18012 52198
rect 18036 52196 18092 52198
rect 18116 52196 18172 52198
rect 18196 52196 18252 52198
rect 17956 51162 18012 51164
rect 18036 51162 18092 51164
rect 18116 51162 18172 51164
rect 18196 51162 18252 51164
rect 17956 51110 18002 51162
rect 18002 51110 18012 51162
rect 18036 51110 18066 51162
rect 18066 51110 18078 51162
rect 18078 51110 18092 51162
rect 18116 51110 18130 51162
rect 18130 51110 18142 51162
rect 18142 51110 18172 51162
rect 18196 51110 18206 51162
rect 18206 51110 18252 51162
rect 17956 51108 18012 51110
rect 18036 51108 18092 51110
rect 18116 51108 18172 51110
rect 18196 51108 18252 51110
rect 17956 50074 18012 50076
rect 18036 50074 18092 50076
rect 18116 50074 18172 50076
rect 18196 50074 18252 50076
rect 17956 50022 18002 50074
rect 18002 50022 18012 50074
rect 18036 50022 18066 50074
rect 18066 50022 18078 50074
rect 18078 50022 18092 50074
rect 18116 50022 18130 50074
rect 18130 50022 18142 50074
rect 18142 50022 18172 50074
rect 18196 50022 18206 50074
rect 18206 50022 18252 50074
rect 17956 50020 18012 50022
rect 18036 50020 18092 50022
rect 18116 50020 18172 50022
rect 18196 50020 18252 50022
rect 17956 48986 18012 48988
rect 18036 48986 18092 48988
rect 18116 48986 18172 48988
rect 18196 48986 18252 48988
rect 17956 48934 18002 48986
rect 18002 48934 18012 48986
rect 18036 48934 18066 48986
rect 18066 48934 18078 48986
rect 18078 48934 18092 48986
rect 18116 48934 18130 48986
rect 18130 48934 18142 48986
rect 18142 48934 18172 48986
rect 18196 48934 18206 48986
rect 18206 48934 18252 48986
rect 17956 48932 18012 48934
rect 18036 48932 18092 48934
rect 18116 48932 18172 48934
rect 18196 48932 18252 48934
rect 17956 47898 18012 47900
rect 18036 47898 18092 47900
rect 18116 47898 18172 47900
rect 18196 47898 18252 47900
rect 17956 47846 18002 47898
rect 18002 47846 18012 47898
rect 18036 47846 18066 47898
rect 18066 47846 18078 47898
rect 18078 47846 18092 47898
rect 18116 47846 18130 47898
rect 18130 47846 18142 47898
rect 18142 47846 18172 47898
rect 18196 47846 18206 47898
rect 18206 47846 18252 47898
rect 17956 47844 18012 47846
rect 18036 47844 18092 47846
rect 18116 47844 18172 47846
rect 18196 47844 18252 47846
rect 17956 46810 18012 46812
rect 18036 46810 18092 46812
rect 18116 46810 18172 46812
rect 18196 46810 18252 46812
rect 17956 46758 18002 46810
rect 18002 46758 18012 46810
rect 18036 46758 18066 46810
rect 18066 46758 18078 46810
rect 18078 46758 18092 46810
rect 18116 46758 18130 46810
rect 18130 46758 18142 46810
rect 18142 46758 18172 46810
rect 18196 46758 18206 46810
rect 18206 46758 18252 46810
rect 17956 46756 18012 46758
rect 18036 46756 18092 46758
rect 18116 46756 18172 46758
rect 18196 46756 18252 46758
rect 17130 36896 17186 36952
rect 17038 31884 17094 31920
rect 17038 31864 17040 31884
rect 17040 31864 17092 31884
rect 17092 31864 17094 31884
rect 16762 29028 16818 29064
rect 16762 29008 16764 29028
rect 16764 29008 16816 29028
rect 16816 29008 16818 29028
rect 16118 25644 16120 25664
rect 16120 25644 16172 25664
rect 16172 25644 16174 25664
rect 16118 25608 16174 25644
rect 16210 17584 16266 17640
rect 16026 15272 16082 15328
rect 16394 20596 16450 20632
rect 16394 20576 16396 20596
rect 16396 20576 16448 20596
rect 16448 20576 16450 20596
rect 17956 45722 18012 45724
rect 18036 45722 18092 45724
rect 18116 45722 18172 45724
rect 18196 45722 18252 45724
rect 17956 45670 18002 45722
rect 18002 45670 18012 45722
rect 18036 45670 18066 45722
rect 18066 45670 18078 45722
rect 18078 45670 18092 45722
rect 18116 45670 18130 45722
rect 18130 45670 18142 45722
rect 18142 45670 18172 45722
rect 18196 45670 18206 45722
rect 18206 45670 18252 45722
rect 17956 45668 18012 45670
rect 18036 45668 18092 45670
rect 18116 45668 18172 45670
rect 18196 45668 18252 45670
rect 17956 44634 18012 44636
rect 18036 44634 18092 44636
rect 18116 44634 18172 44636
rect 18196 44634 18252 44636
rect 17956 44582 18002 44634
rect 18002 44582 18012 44634
rect 18036 44582 18066 44634
rect 18066 44582 18078 44634
rect 18078 44582 18092 44634
rect 18116 44582 18130 44634
rect 18130 44582 18142 44634
rect 18142 44582 18172 44634
rect 18196 44582 18206 44634
rect 18206 44582 18252 44634
rect 17956 44580 18012 44582
rect 18036 44580 18092 44582
rect 18116 44580 18172 44582
rect 18196 44580 18252 44582
rect 17956 43546 18012 43548
rect 18036 43546 18092 43548
rect 18116 43546 18172 43548
rect 18196 43546 18252 43548
rect 17956 43494 18002 43546
rect 18002 43494 18012 43546
rect 18036 43494 18066 43546
rect 18066 43494 18078 43546
rect 18078 43494 18092 43546
rect 18116 43494 18130 43546
rect 18130 43494 18142 43546
rect 18142 43494 18172 43546
rect 18196 43494 18206 43546
rect 18206 43494 18252 43546
rect 17956 43492 18012 43494
rect 18036 43492 18092 43494
rect 18116 43492 18172 43494
rect 18196 43492 18252 43494
rect 17956 42458 18012 42460
rect 18036 42458 18092 42460
rect 18116 42458 18172 42460
rect 18196 42458 18252 42460
rect 17956 42406 18002 42458
rect 18002 42406 18012 42458
rect 18036 42406 18066 42458
rect 18066 42406 18078 42458
rect 18078 42406 18092 42458
rect 18116 42406 18130 42458
rect 18130 42406 18142 42458
rect 18142 42406 18172 42458
rect 18196 42406 18206 42458
rect 18206 42406 18252 42458
rect 17956 42404 18012 42406
rect 18036 42404 18092 42406
rect 18116 42404 18172 42406
rect 18196 42404 18252 42406
rect 17956 41370 18012 41372
rect 18036 41370 18092 41372
rect 18116 41370 18172 41372
rect 18196 41370 18252 41372
rect 17956 41318 18002 41370
rect 18002 41318 18012 41370
rect 18036 41318 18066 41370
rect 18066 41318 18078 41370
rect 18078 41318 18092 41370
rect 18116 41318 18130 41370
rect 18130 41318 18142 41370
rect 18142 41318 18172 41370
rect 18196 41318 18206 41370
rect 18206 41318 18252 41370
rect 17956 41316 18012 41318
rect 18036 41316 18092 41318
rect 18116 41316 18172 41318
rect 18196 41316 18252 41318
rect 17590 36216 17646 36272
rect 17956 40282 18012 40284
rect 18036 40282 18092 40284
rect 18116 40282 18172 40284
rect 18196 40282 18252 40284
rect 17956 40230 18002 40282
rect 18002 40230 18012 40282
rect 18036 40230 18066 40282
rect 18066 40230 18078 40282
rect 18078 40230 18092 40282
rect 18116 40230 18130 40282
rect 18130 40230 18142 40282
rect 18142 40230 18172 40282
rect 18196 40230 18206 40282
rect 18206 40230 18252 40282
rect 17956 40228 18012 40230
rect 18036 40228 18092 40230
rect 18116 40228 18172 40230
rect 18196 40228 18252 40230
rect 17956 39194 18012 39196
rect 18036 39194 18092 39196
rect 18116 39194 18172 39196
rect 18196 39194 18252 39196
rect 17956 39142 18002 39194
rect 18002 39142 18012 39194
rect 18036 39142 18066 39194
rect 18066 39142 18078 39194
rect 18078 39142 18092 39194
rect 18116 39142 18130 39194
rect 18130 39142 18142 39194
rect 18142 39142 18172 39194
rect 18196 39142 18206 39194
rect 18206 39142 18252 39194
rect 17956 39140 18012 39142
rect 18036 39140 18092 39142
rect 18116 39140 18172 39142
rect 18196 39140 18252 39142
rect 17956 38106 18012 38108
rect 18036 38106 18092 38108
rect 18116 38106 18172 38108
rect 18196 38106 18252 38108
rect 17956 38054 18002 38106
rect 18002 38054 18012 38106
rect 18036 38054 18066 38106
rect 18066 38054 18078 38106
rect 18078 38054 18092 38106
rect 18116 38054 18130 38106
rect 18130 38054 18142 38106
rect 18142 38054 18172 38106
rect 18196 38054 18206 38106
rect 18206 38054 18252 38106
rect 17956 38052 18012 38054
rect 18036 38052 18092 38054
rect 18116 38052 18172 38054
rect 18196 38052 18252 38054
rect 17774 37324 17830 37360
rect 17774 37304 17776 37324
rect 17776 37304 17828 37324
rect 17828 37304 17830 37324
rect 17956 37018 18012 37020
rect 18036 37018 18092 37020
rect 18116 37018 18172 37020
rect 18196 37018 18252 37020
rect 17956 36966 18002 37018
rect 18002 36966 18012 37018
rect 18036 36966 18066 37018
rect 18066 36966 18078 37018
rect 18078 36966 18092 37018
rect 18116 36966 18130 37018
rect 18130 36966 18142 37018
rect 18142 36966 18172 37018
rect 18196 36966 18206 37018
rect 18206 36966 18252 37018
rect 17956 36964 18012 36966
rect 18036 36964 18092 36966
rect 18116 36964 18172 36966
rect 18196 36964 18252 36966
rect 18418 38664 18474 38720
rect 17956 35930 18012 35932
rect 18036 35930 18092 35932
rect 18116 35930 18172 35932
rect 18196 35930 18252 35932
rect 17956 35878 18002 35930
rect 18002 35878 18012 35930
rect 18036 35878 18066 35930
rect 18066 35878 18078 35930
rect 18078 35878 18092 35930
rect 18116 35878 18130 35930
rect 18130 35878 18142 35930
rect 18142 35878 18172 35930
rect 18196 35878 18206 35930
rect 18206 35878 18252 35930
rect 17956 35876 18012 35878
rect 18036 35876 18092 35878
rect 18116 35876 18172 35878
rect 18196 35876 18252 35878
rect 17956 34842 18012 34844
rect 18036 34842 18092 34844
rect 18116 34842 18172 34844
rect 18196 34842 18252 34844
rect 17956 34790 18002 34842
rect 18002 34790 18012 34842
rect 18036 34790 18066 34842
rect 18066 34790 18078 34842
rect 18078 34790 18092 34842
rect 18116 34790 18130 34842
rect 18130 34790 18142 34842
rect 18142 34790 18172 34842
rect 18196 34790 18206 34842
rect 18206 34790 18252 34842
rect 17956 34788 18012 34790
rect 18036 34788 18092 34790
rect 18116 34788 18172 34790
rect 18196 34788 18252 34790
rect 17956 33754 18012 33756
rect 18036 33754 18092 33756
rect 18116 33754 18172 33756
rect 18196 33754 18252 33756
rect 17956 33702 18002 33754
rect 18002 33702 18012 33754
rect 18036 33702 18066 33754
rect 18066 33702 18078 33754
rect 18078 33702 18092 33754
rect 18116 33702 18130 33754
rect 18130 33702 18142 33754
rect 18142 33702 18172 33754
rect 18196 33702 18206 33754
rect 18206 33702 18252 33754
rect 17956 33700 18012 33702
rect 18036 33700 18092 33702
rect 18116 33700 18172 33702
rect 18196 33700 18252 33702
rect 19522 44240 19578 44296
rect 17956 32666 18012 32668
rect 18036 32666 18092 32668
rect 18116 32666 18172 32668
rect 18196 32666 18252 32668
rect 17956 32614 18002 32666
rect 18002 32614 18012 32666
rect 18036 32614 18066 32666
rect 18066 32614 18078 32666
rect 18078 32614 18092 32666
rect 18116 32614 18130 32666
rect 18130 32614 18142 32666
rect 18142 32614 18172 32666
rect 18196 32614 18206 32666
rect 18206 32614 18252 32666
rect 17956 32612 18012 32614
rect 18036 32612 18092 32614
rect 18116 32612 18172 32614
rect 18196 32612 18252 32614
rect 17498 29044 17500 29064
rect 17500 29044 17552 29064
rect 17552 29044 17554 29064
rect 17498 29008 17554 29044
rect 18878 37712 18934 37768
rect 17956 31578 18012 31580
rect 18036 31578 18092 31580
rect 18116 31578 18172 31580
rect 18196 31578 18252 31580
rect 17956 31526 18002 31578
rect 18002 31526 18012 31578
rect 18036 31526 18066 31578
rect 18066 31526 18078 31578
rect 18078 31526 18092 31578
rect 18116 31526 18130 31578
rect 18130 31526 18142 31578
rect 18142 31526 18172 31578
rect 18196 31526 18206 31578
rect 18206 31526 18252 31578
rect 17956 31524 18012 31526
rect 18036 31524 18092 31526
rect 18116 31524 18172 31526
rect 18196 31524 18252 31526
rect 18142 30796 18198 30832
rect 18142 30776 18144 30796
rect 18144 30776 18196 30796
rect 18196 30776 18198 30796
rect 17956 30490 18012 30492
rect 18036 30490 18092 30492
rect 18116 30490 18172 30492
rect 18196 30490 18252 30492
rect 17956 30438 18002 30490
rect 18002 30438 18012 30490
rect 18036 30438 18066 30490
rect 18066 30438 18078 30490
rect 18078 30438 18092 30490
rect 18116 30438 18130 30490
rect 18130 30438 18142 30490
rect 18142 30438 18172 30490
rect 18196 30438 18206 30490
rect 18206 30438 18252 30490
rect 17956 30436 18012 30438
rect 18036 30436 18092 30438
rect 18116 30436 18172 30438
rect 18196 30436 18252 30438
rect 18234 29708 18290 29744
rect 18234 29688 18236 29708
rect 18236 29688 18288 29708
rect 18288 29688 18290 29708
rect 17956 29402 18012 29404
rect 18036 29402 18092 29404
rect 18116 29402 18172 29404
rect 18196 29402 18252 29404
rect 17956 29350 18002 29402
rect 18002 29350 18012 29402
rect 18036 29350 18066 29402
rect 18066 29350 18078 29402
rect 18078 29350 18092 29402
rect 18116 29350 18130 29402
rect 18130 29350 18142 29402
rect 18142 29350 18172 29402
rect 18196 29350 18206 29402
rect 18206 29350 18252 29402
rect 17956 29348 18012 29350
rect 18036 29348 18092 29350
rect 18116 29348 18172 29350
rect 18196 29348 18252 29350
rect 17956 28314 18012 28316
rect 18036 28314 18092 28316
rect 18116 28314 18172 28316
rect 18196 28314 18252 28316
rect 17956 28262 18002 28314
rect 18002 28262 18012 28314
rect 18036 28262 18066 28314
rect 18066 28262 18078 28314
rect 18078 28262 18092 28314
rect 18116 28262 18130 28314
rect 18130 28262 18142 28314
rect 18142 28262 18172 28314
rect 18196 28262 18206 28314
rect 18206 28262 18252 28314
rect 17956 28260 18012 28262
rect 18036 28260 18092 28262
rect 18116 28260 18172 28262
rect 18196 28260 18252 28262
rect 17956 27226 18012 27228
rect 18036 27226 18092 27228
rect 18116 27226 18172 27228
rect 18196 27226 18252 27228
rect 17956 27174 18002 27226
rect 18002 27174 18012 27226
rect 18036 27174 18066 27226
rect 18066 27174 18078 27226
rect 18078 27174 18092 27226
rect 18116 27174 18130 27226
rect 18130 27174 18142 27226
rect 18142 27174 18172 27226
rect 18196 27174 18206 27226
rect 18206 27174 18252 27226
rect 17956 27172 18012 27174
rect 18036 27172 18092 27174
rect 18116 27172 18172 27174
rect 18196 27172 18252 27174
rect 17956 26138 18012 26140
rect 18036 26138 18092 26140
rect 18116 26138 18172 26140
rect 18196 26138 18252 26140
rect 17956 26086 18002 26138
rect 18002 26086 18012 26138
rect 18036 26086 18066 26138
rect 18066 26086 18078 26138
rect 18078 26086 18092 26138
rect 18116 26086 18130 26138
rect 18130 26086 18142 26138
rect 18142 26086 18172 26138
rect 18196 26086 18206 26138
rect 18206 26086 18252 26138
rect 17956 26084 18012 26086
rect 18036 26084 18092 26086
rect 18116 26084 18172 26086
rect 18196 26084 18252 26086
rect 17956 25050 18012 25052
rect 18036 25050 18092 25052
rect 18116 25050 18172 25052
rect 18196 25050 18252 25052
rect 17956 24998 18002 25050
rect 18002 24998 18012 25050
rect 18036 24998 18066 25050
rect 18066 24998 18078 25050
rect 18078 24998 18092 25050
rect 18116 24998 18130 25050
rect 18130 24998 18142 25050
rect 18142 24998 18172 25050
rect 18196 24998 18206 25050
rect 18206 24998 18252 25050
rect 17956 24996 18012 24998
rect 18036 24996 18092 24998
rect 18116 24996 18172 24998
rect 18196 24996 18252 24998
rect 18970 33496 19026 33552
rect 18970 30640 19026 30696
rect 17956 23962 18012 23964
rect 18036 23962 18092 23964
rect 18116 23962 18172 23964
rect 18196 23962 18252 23964
rect 17956 23910 18002 23962
rect 18002 23910 18012 23962
rect 18036 23910 18066 23962
rect 18066 23910 18078 23962
rect 18078 23910 18092 23962
rect 18116 23910 18130 23962
rect 18130 23910 18142 23962
rect 18142 23910 18172 23962
rect 18196 23910 18206 23962
rect 18206 23910 18252 23962
rect 17956 23908 18012 23910
rect 18036 23908 18092 23910
rect 18116 23908 18172 23910
rect 18196 23908 18252 23910
rect 17956 22874 18012 22876
rect 18036 22874 18092 22876
rect 18116 22874 18172 22876
rect 18196 22874 18252 22876
rect 17956 22822 18002 22874
rect 18002 22822 18012 22874
rect 18036 22822 18066 22874
rect 18066 22822 18078 22874
rect 18078 22822 18092 22874
rect 18116 22822 18130 22874
rect 18130 22822 18142 22874
rect 18142 22822 18172 22874
rect 18196 22822 18206 22874
rect 18206 22822 18252 22874
rect 17956 22820 18012 22822
rect 18036 22820 18092 22822
rect 18116 22820 18172 22822
rect 18196 22820 18252 22822
rect 17956 21786 18012 21788
rect 18036 21786 18092 21788
rect 18116 21786 18172 21788
rect 18196 21786 18252 21788
rect 17956 21734 18002 21786
rect 18002 21734 18012 21786
rect 18036 21734 18066 21786
rect 18066 21734 18078 21786
rect 18078 21734 18092 21786
rect 18116 21734 18130 21786
rect 18130 21734 18142 21786
rect 18142 21734 18172 21786
rect 18196 21734 18206 21786
rect 18206 21734 18252 21786
rect 17956 21732 18012 21734
rect 18036 21732 18092 21734
rect 18116 21732 18172 21734
rect 18196 21732 18252 21734
rect 17222 19896 17278 19952
rect 15658 2624 15714 2680
rect 17590 18828 17646 18864
rect 17590 18808 17592 18828
rect 17592 18808 17644 18828
rect 17644 18808 17646 18828
rect 17956 20698 18012 20700
rect 18036 20698 18092 20700
rect 18116 20698 18172 20700
rect 18196 20698 18252 20700
rect 17956 20646 18002 20698
rect 18002 20646 18012 20698
rect 18036 20646 18066 20698
rect 18066 20646 18078 20698
rect 18078 20646 18092 20698
rect 18116 20646 18130 20698
rect 18130 20646 18142 20698
rect 18142 20646 18172 20698
rect 18196 20646 18206 20698
rect 18206 20646 18252 20698
rect 17956 20644 18012 20646
rect 18036 20644 18092 20646
rect 18116 20644 18172 20646
rect 18196 20644 18252 20646
rect 17956 19610 18012 19612
rect 18036 19610 18092 19612
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 17956 19558 18002 19610
rect 18002 19558 18012 19610
rect 18036 19558 18066 19610
rect 18066 19558 18078 19610
rect 18078 19558 18092 19610
rect 18116 19558 18130 19610
rect 18130 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 17956 19556 18012 19558
rect 18036 19556 18092 19558
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 17956 18522 18012 18524
rect 18036 18522 18092 18524
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 17956 18470 18002 18522
rect 18002 18470 18012 18522
rect 18036 18470 18066 18522
rect 18066 18470 18078 18522
rect 18078 18470 18092 18522
rect 18116 18470 18130 18522
rect 18130 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 17956 18468 18012 18470
rect 18036 18468 18092 18470
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 18510 18264 18566 18320
rect 17866 17584 17922 17640
rect 17956 17434 18012 17436
rect 18036 17434 18092 17436
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 17956 17382 18002 17434
rect 18002 17382 18012 17434
rect 18036 17382 18066 17434
rect 18066 17382 18078 17434
rect 18078 17382 18092 17434
rect 18116 17382 18130 17434
rect 18130 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 17956 17380 18012 17382
rect 18036 17380 18092 17382
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 17956 16346 18012 16348
rect 18036 16346 18092 16348
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 17956 16294 18002 16346
rect 18002 16294 18012 16346
rect 18036 16294 18066 16346
rect 18066 16294 18078 16346
rect 18078 16294 18092 16346
rect 18116 16294 18130 16346
rect 18130 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 17956 16292 18012 16294
rect 18036 16292 18092 16294
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 17956 15258 18012 15260
rect 18036 15258 18092 15260
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 17956 15206 18002 15258
rect 18002 15206 18012 15258
rect 18036 15206 18066 15258
rect 18066 15206 18078 15258
rect 18078 15206 18092 15258
rect 18116 15206 18130 15258
rect 18130 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 17956 15204 18012 15206
rect 18036 15204 18092 15206
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 17956 14170 18012 14172
rect 18036 14170 18092 14172
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 17956 14118 18002 14170
rect 18002 14118 18012 14170
rect 18036 14118 18066 14170
rect 18066 14118 18078 14170
rect 18078 14118 18092 14170
rect 18116 14118 18130 14170
rect 18130 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 17956 14116 18012 14118
rect 18036 14116 18092 14118
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 19062 22208 19118 22264
rect 19614 36624 19670 36680
rect 19890 38936 19946 38992
rect 19890 37612 19892 37632
rect 19892 37612 19944 37632
rect 19944 37612 19946 37632
rect 19890 37576 19946 37612
rect 20534 45736 20590 45792
rect 21454 45464 21510 45520
rect 21454 44276 21456 44296
rect 21456 44276 21508 44296
rect 21508 44276 21510 44296
rect 21454 44240 21510 44276
rect 19430 30232 19486 30288
rect 19246 27532 19302 27568
rect 19246 27512 19248 27532
rect 19248 27512 19300 27532
rect 19300 27512 19302 27532
rect 19246 27124 19302 27160
rect 19246 27104 19248 27124
rect 19248 27104 19300 27124
rect 19300 27104 19302 27124
rect 19982 30132 19984 30152
rect 19984 30132 20036 30152
rect 20036 30132 20038 30152
rect 19982 30096 20038 30132
rect 19890 29708 19946 29744
rect 19890 29688 19892 29708
rect 19892 29688 19944 29708
rect 19944 29688 19946 29708
rect 19338 24520 19394 24576
rect 21178 41420 21180 41440
rect 21180 41420 21232 41440
rect 21232 41420 21234 41440
rect 21178 41384 21234 41420
rect 20442 28076 20498 28112
rect 20442 28056 20444 28076
rect 20444 28056 20496 28076
rect 20496 28056 20498 28076
rect 17956 13082 18012 13084
rect 18036 13082 18092 13084
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 17956 13030 18002 13082
rect 18002 13030 18012 13082
rect 18036 13030 18066 13082
rect 18066 13030 18078 13082
rect 18078 13030 18092 13082
rect 18116 13030 18130 13082
rect 18130 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 17956 13028 18012 13030
rect 18036 13028 18092 13030
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 17956 11994 18012 11996
rect 18036 11994 18092 11996
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 17956 11942 18002 11994
rect 18002 11942 18012 11994
rect 18036 11942 18066 11994
rect 18066 11942 18078 11994
rect 18078 11942 18092 11994
rect 18116 11942 18130 11994
rect 18130 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 17956 11940 18012 11942
rect 18036 11940 18092 11942
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 17956 10906 18012 10908
rect 18036 10906 18092 10908
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 17956 10854 18002 10906
rect 18002 10854 18012 10906
rect 18036 10854 18066 10906
rect 18066 10854 18078 10906
rect 18078 10854 18092 10906
rect 18116 10854 18130 10906
rect 18130 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 17956 10852 18012 10854
rect 18036 10852 18092 10854
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 17956 9818 18012 9820
rect 18036 9818 18092 9820
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 17956 9766 18002 9818
rect 18002 9766 18012 9818
rect 18036 9766 18066 9818
rect 18066 9766 18078 9818
rect 18078 9766 18092 9818
rect 18116 9766 18130 9818
rect 18130 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 17956 9764 18012 9766
rect 18036 9764 18092 9766
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 17956 8730 18012 8732
rect 18036 8730 18092 8732
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 17956 8678 18002 8730
rect 18002 8678 18012 8730
rect 18036 8678 18066 8730
rect 18066 8678 18078 8730
rect 18078 8678 18092 8730
rect 18116 8678 18130 8730
rect 18130 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 17956 8676 18012 8678
rect 18036 8676 18092 8678
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 17956 7642 18012 7644
rect 18036 7642 18092 7644
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 17956 7590 18002 7642
rect 18002 7590 18012 7642
rect 18036 7590 18066 7642
rect 18066 7590 18078 7642
rect 18078 7590 18092 7642
rect 18116 7590 18130 7642
rect 18130 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 17956 7588 18012 7590
rect 18036 7588 18092 7590
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 17956 6554 18012 6556
rect 18036 6554 18092 6556
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 17956 6502 18002 6554
rect 18002 6502 18012 6554
rect 18036 6502 18066 6554
rect 18066 6502 18078 6554
rect 18078 6502 18092 6554
rect 18116 6502 18130 6554
rect 18130 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 17956 6500 18012 6502
rect 18036 6500 18092 6502
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 17956 5466 18012 5468
rect 18036 5466 18092 5468
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 17956 5414 18002 5466
rect 18002 5414 18012 5466
rect 18036 5414 18066 5466
rect 18066 5414 18078 5466
rect 18078 5414 18092 5466
rect 18116 5414 18130 5466
rect 18130 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 17956 5412 18012 5414
rect 18036 5412 18092 5414
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 17956 4378 18012 4380
rect 18036 4378 18092 4380
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 17956 4326 18002 4378
rect 18002 4326 18012 4378
rect 18036 4326 18066 4378
rect 18066 4326 18078 4378
rect 18078 4326 18092 4378
rect 18116 4326 18130 4378
rect 18130 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 17956 4324 18012 4326
rect 18036 4324 18092 4326
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 17956 3290 18012 3292
rect 18036 3290 18092 3292
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 17956 3238 18002 3290
rect 18002 3238 18012 3290
rect 18036 3238 18066 3290
rect 18066 3238 18078 3290
rect 18078 3238 18092 3290
rect 18116 3238 18130 3290
rect 18130 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 17956 3236 18012 3238
rect 18036 3236 18092 3238
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 17956 2202 18012 2204
rect 18036 2202 18092 2204
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 17956 2150 18002 2202
rect 18002 2150 18012 2202
rect 18036 2150 18066 2202
rect 18066 2150 18078 2202
rect 18078 2150 18092 2202
rect 18116 2150 18130 2202
rect 18130 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 17956 2148 18012 2150
rect 18036 2148 18092 2150
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 19338 13504 19394 13560
rect 22956 53882 23012 53884
rect 23036 53882 23092 53884
rect 23116 53882 23172 53884
rect 23196 53882 23252 53884
rect 22956 53830 23002 53882
rect 23002 53830 23012 53882
rect 23036 53830 23066 53882
rect 23066 53830 23078 53882
rect 23078 53830 23092 53882
rect 23116 53830 23130 53882
rect 23130 53830 23142 53882
rect 23142 53830 23172 53882
rect 23196 53830 23206 53882
rect 23206 53830 23252 53882
rect 22956 53828 23012 53830
rect 23036 53828 23092 53830
rect 23116 53828 23172 53830
rect 23196 53828 23252 53830
rect 22190 52536 22246 52592
rect 22956 52794 23012 52796
rect 23036 52794 23092 52796
rect 23116 52794 23172 52796
rect 23196 52794 23252 52796
rect 22956 52742 23002 52794
rect 23002 52742 23012 52794
rect 23036 52742 23066 52794
rect 23066 52742 23078 52794
rect 23078 52742 23092 52794
rect 23116 52742 23130 52794
rect 23130 52742 23142 52794
rect 23142 52742 23172 52794
rect 23196 52742 23206 52794
rect 23206 52742 23252 52794
rect 22956 52740 23012 52742
rect 23036 52740 23092 52742
rect 23116 52740 23172 52742
rect 23196 52740 23252 52742
rect 22956 51706 23012 51708
rect 23036 51706 23092 51708
rect 23116 51706 23172 51708
rect 23196 51706 23252 51708
rect 22956 51654 23002 51706
rect 23002 51654 23012 51706
rect 23036 51654 23066 51706
rect 23066 51654 23078 51706
rect 23078 51654 23092 51706
rect 23116 51654 23130 51706
rect 23130 51654 23142 51706
rect 23142 51654 23172 51706
rect 23196 51654 23206 51706
rect 23206 51654 23252 51706
rect 22956 51652 23012 51654
rect 23036 51652 23092 51654
rect 23116 51652 23172 51654
rect 23196 51652 23252 51654
rect 22956 50618 23012 50620
rect 23036 50618 23092 50620
rect 23116 50618 23172 50620
rect 23196 50618 23252 50620
rect 22956 50566 23002 50618
rect 23002 50566 23012 50618
rect 23036 50566 23066 50618
rect 23066 50566 23078 50618
rect 23078 50566 23092 50618
rect 23116 50566 23130 50618
rect 23130 50566 23142 50618
rect 23142 50566 23172 50618
rect 23196 50566 23206 50618
rect 23206 50566 23252 50618
rect 22956 50564 23012 50566
rect 23036 50564 23092 50566
rect 23116 50564 23172 50566
rect 23196 50564 23252 50566
rect 22956 49530 23012 49532
rect 23036 49530 23092 49532
rect 23116 49530 23172 49532
rect 23196 49530 23252 49532
rect 22956 49478 23002 49530
rect 23002 49478 23012 49530
rect 23036 49478 23066 49530
rect 23066 49478 23078 49530
rect 23078 49478 23092 49530
rect 23116 49478 23130 49530
rect 23130 49478 23142 49530
rect 23142 49478 23172 49530
rect 23196 49478 23206 49530
rect 23206 49478 23252 49530
rect 22956 49476 23012 49478
rect 23036 49476 23092 49478
rect 23116 49476 23172 49478
rect 23196 49476 23252 49478
rect 22956 48442 23012 48444
rect 23036 48442 23092 48444
rect 23116 48442 23172 48444
rect 23196 48442 23252 48444
rect 22956 48390 23002 48442
rect 23002 48390 23012 48442
rect 23036 48390 23066 48442
rect 23066 48390 23078 48442
rect 23078 48390 23092 48442
rect 23116 48390 23130 48442
rect 23130 48390 23142 48442
rect 23142 48390 23172 48442
rect 23196 48390 23206 48442
rect 23206 48390 23252 48442
rect 22956 48388 23012 48390
rect 23036 48388 23092 48390
rect 23116 48388 23172 48390
rect 23196 48388 23252 48390
rect 22956 47354 23012 47356
rect 23036 47354 23092 47356
rect 23116 47354 23172 47356
rect 23196 47354 23252 47356
rect 22956 47302 23002 47354
rect 23002 47302 23012 47354
rect 23036 47302 23066 47354
rect 23066 47302 23078 47354
rect 23078 47302 23092 47354
rect 23116 47302 23130 47354
rect 23130 47302 23142 47354
rect 23142 47302 23172 47354
rect 23196 47302 23206 47354
rect 23206 47302 23252 47354
rect 22956 47300 23012 47302
rect 23036 47300 23092 47302
rect 23116 47300 23172 47302
rect 23196 47300 23252 47302
rect 22956 46266 23012 46268
rect 23036 46266 23092 46268
rect 23116 46266 23172 46268
rect 23196 46266 23252 46268
rect 22956 46214 23002 46266
rect 23002 46214 23012 46266
rect 23036 46214 23066 46266
rect 23066 46214 23078 46266
rect 23078 46214 23092 46266
rect 23116 46214 23130 46266
rect 23130 46214 23142 46266
rect 23142 46214 23172 46266
rect 23196 46214 23206 46266
rect 23206 46214 23252 46266
rect 22956 46212 23012 46214
rect 23036 46212 23092 46214
rect 23116 46212 23172 46214
rect 23196 46212 23252 46214
rect 22650 45484 22706 45520
rect 22650 45464 22652 45484
rect 22652 45464 22704 45484
rect 22704 45464 22706 45484
rect 22956 45178 23012 45180
rect 23036 45178 23092 45180
rect 23116 45178 23172 45180
rect 23196 45178 23252 45180
rect 22956 45126 23002 45178
rect 23002 45126 23012 45178
rect 23036 45126 23066 45178
rect 23066 45126 23078 45178
rect 23078 45126 23092 45178
rect 23116 45126 23130 45178
rect 23130 45126 23142 45178
rect 23142 45126 23172 45178
rect 23196 45126 23206 45178
rect 23206 45126 23252 45178
rect 22956 45124 23012 45126
rect 23036 45124 23092 45126
rect 23116 45124 23172 45126
rect 23196 45124 23252 45126
rect 21270 36216 21326 36272
rect 21546 36760 21602 36816
rect 20902 28364 20904 28384
rect 20904 28364 20956 28384
rect 20956 28364 20958 28384
rect 20902 28328 20958 28364
rect 19982 15564 20038 15600
rect 19982 15544 19984 15564
rect 19984 15544 20036 15564
rect 20036 15544 20038 15564
rect 22956 44090 23012 44092
rect 23036 44090 23092 44092
rect 23116 44090 23172 44092
rect 23196 44090 23252 44092
rect 22956 44038 23002 44090
rect 23002 44038 23012 44090
rect 23036 44038 23066 44090
rect 23066 44038 23078 44090
rect 23078 44038 23092 44090
rect 23116 44038 23130 44090
rect 23130 44038 23142 44090
rect 23142 44038 23172 44090
rect 23196 44038 23206 44090
rect 23206 44038 23252 44090
rect 22956 44036 23012 44038
rect 23036 44036 23092 44038
rect 23116 44036 23172 44038
rect 23196 44036 23252 44038
rect 22956 43002 23012 43004
rect 23036 43002 23092 43004
rect 23116 43002 23172 43004
rect 23196 43002 23252 43004
rect 22956 42950 23002 43002
rect 23002 42950 23012 43002
rect 23036 42950 23066 43002
rect 23066 42950 23078 43002
rect 23078 42950 23092 43002
rect 23116 42950 23130 43002
rect 23130 42950 23142 43002
rect 23142 42950 23172 43002
rect 23196 42950 23206 43002
rect 23206 42950 23252 43002
rect 22956 42948 23012 42950
rect 23036 42948 23092 42950
rect 23116 42948 23172 42950
rect 23196 42948 23252 42950
rect 22956 41914 23012 41916
rect 23036 41914 23092 41916
rect 23116 41914 23172 41916
rect 23196 41914 23252 41916
rect 22956 41862 23002 41914
rect 23002 41862 23012 41914
rect 23036 41862 23066 41914
rect 23066 41862 23078 41914
rect 23078 41862 23092 41914
rect 23116 41862 23130 41914
rect 23130 41862 23142 41914
rect 23142 41862 23172 41914
rect 23196 41862 23206 41914
rect 23206 41862 23252 41914
rect 22956 41860 23012 41862
rect 23036 41860 23092 41862
rect 23116 41860 23172 41862
rect 23196 41860 23252 41862
rect 23846 45056 23902 45112
rect 21638 31728 21694 31784
rect 22956 40826 23012 40828
rect 23036 40826 23092 40828
rect 23116 40826 23172 40828
rect 23196 40826 23252 40828
rect 22956 40774 23002 40826
rect 23002 40774 23012 40826
rect 23036 40774 23066 40826
rect 23066 40774 23078 40826
rect 23078 40774 23092 40826
rect 23116 40774 23130 40826
rect 23130 40774 23142 40826
rect 23142 40774 23172 40826
rect 23196 40774 23206 40826
rect 23206 40774 23252 40826
rect 22956 40772 23012 40774
rect 23036 40772 23092 40774
rect 23116 40772 23172 40774
rect 23196 40772 23252 40774
rect 22956 39738 23012 39740
rect 23036 39738 23092 39740
rect 23116 39738 23172 39740
rect 23196 39738 23252 39740
rect 22956 39686 23002 39738
rect 23002 39686 23012 39738
rect 23036 39686 23066 39738
rect 23066 39686 23078 39738
rect 23078 39686 23092 39738
rect 23116 39686 23130 39738
rect 23130 39686 23142 39738
rect 23142 39686 23172 39738
rect 23196 39686 23206 39738
rect 23206 39686 23252 39738
rect 22956 39684 23012 39686
rect 23036 39684 23092 39686
rect 23116 39684 23172 39686
rect 23196 39684 23252 39686
rect 22956 38650 23012 38652
rect 23036 38650 23092 38652
rect 23116 38650 23172 38652
rect 23196 38650 23252 38652
rect 22956 38598 23002 38650
rect 23002 38598 23012 38650
rect 23036 38598 23066 38650
rect 23066 38598 23078 38650
rect 23078 38598 23092 38650
rect 23116 38598 23130 38650
rect 23130 38598 23142 38650
rect 23142 38598 23172 38650
rect 23196 38598 23206 38650
rect 23206 38598 23252 38650
rect 22956 38596 23012 38598
rect 23036 38596 23092 38598
rect 23116 38596 23172 38598
rect 23196 38596 23252 38598
rect 23386 40296 23442 40352
rect 22956 37562 23012 37564
rect 23036 37562 23092 37564
rect 23116 37562 23172 37564
rect 23196 37562 23252 37564
rect 22956 37510 23002 37562
rect 23002 37510 23012 37562
rect 23036 37510 23066 37562
rect 23066 37510 23078 37562
rect 23078 37510 23092 37562
rect 23116 37510 23130 37562
rect 23130 37510 23142 37562
rect 23142 37510 23172 37562
rect 23196 37510 23206 37562
rect 23206 37510 23252 37562
rect 22956 37508 23012 37510
rect 23036 37508 23092 37510
rect 23116 37508 23172 37510
rect 23196 37508 23252 37510
rect 22956 36474 23012 36476
rect 23036 36474 23092 36476
rect 23116 36474 23172 36476
rect 23196 36474 23252 36476
rect 22956 36422 23002 36474
rect 23002 36422 23012 36474
rect 23036 36422 23066 36474
rect 23066 36422 23078 36474
rect 23078 36422 23092 36474
rect 23116 36422 23130 36474
rect 23130 36422 23142 36474
rect 23142 36422 23172 36474
rect 23196 36422 23206 36474
rect 23206 36422 23252 36474
rect 22956 36420 23012 36422
rect 23036 36420 23092 36422
rect 23116 36420 23172 36422
rect 23196 36420 23252 36422
rect 22742 35128 22798 35184
rect 21730 29416 21786 29472
rect 22282 29708 22338 29744
rect 22282 29688 22284 29708
rect 22284 29688 22336 29708
rect 22336 29688 22338 29708
rect 22282 26016 22338 26072
rect 22956 35386 23012 35388
rect 23036 35386 23092 35388
rect 23116 35386 23172 35388
rect 23196 35386 23252 35388
rect 22956 35334 23002 35386
rect 23002 35334 23012 35386
rect 23036 35334 23066 35386
rect 23066 35334 23078 35386
rect 23078 35334 23092 35386
rect 23116 35334 23130 35386
rect 23130 35334 23142 35386
rect 23142 35334 23172 35386
rect 23196 35334 23206 35386
rect 23206 35334 23252 35386
rect 22956 35332 23012 35334
rect 23036 35332 23092 35334
rect 23116 35332 23172 35334
rect 23196 35332 23252 35334
rect 22956 34298 23012 34300
rect 23036 34298 23092 34300
rect 23116 34298 23172 34300
rect 23196 34298 23252 34300
rect 22956 34246 23002 34298
rect 23002 34246 23012 34298
rect 23036 34246 23066 34298
rect 23066 34246 23078 34298
rect 23078 34246 23092 34298
rect 23116 34246 23130 34298
rect 23130 34246 23142 34298
rect 23142 34246 23172 34298
rect 23196 34246 23206 34298
rect 23206 34246 23252 34298
rect 22956 34244 23012 34246
rect 23036 34244 23092 34246
rect 23116 34244 23172 34246
rect 23196 34244 23252 34246
rect 24674 52536 24730 52592
rect 24766 49136 24822 49192
rect 24766 47776 24822 47832
rect 25226 51856 25282 51912
rect 25318 51176 25374 51232
rect 24858 46436 24914 46472
rect 24858 46416 24860 46436
rect 24860 46416 24912 46436
rect 24912 46416 24914 46436
rect 24766 45736 24822 45792
rect 24766 44376 24822 44432
rect 24674 43696 24730 43752
rect 23662 37168 23718 37224
rect 23938 36760 23994 36816
rect 24766 40976 24822 41032
rect 22956 33210 23012 33212
rect 23036 33210 23092 33212
rect 23116 33210 23172 33212
rect 23196 33210 23252 33212
rect 22956 33158 23002 33210
rect 23002 33158 23012 33210
rect 23036 33158 23066 33210
rect 23066 33158 23078 33210
rect 23078 33158 23092 33210
rect 23116 33158 23130 33210
rect 23130 33158 23142 33210
rect 23142 33158 23172 33210
rect 23196 33158 23206 33210
rect 23206 33158 23252 33210
rect 22956 33156 23012 33158
rect 23036 33156 23092 33158
rect 23116 33156 23172 33158
rect 23196 33156 23252 33158
rect 22956 32122 23012 32124
rect 23036 32122 23092 32124
rect 23116 32122 23172 32124
rect 23196 32122 23252 32124
rect 22956 32070 23002 32122
rect 23002 32070 23012 32122
rect 23036 32070 23066 32122
rect 23066 32070 23078 32122
rect 23078 32070 23092 32122
rect 23116 32070 23130 32122
rect 23130 32070 23142 32122
rect 23142 32070 23172 32122
rect 23196 32070 23206 32122
rect 23206 32070 23252 32122
rect 22956 32068 23012 32070
rect 23036 32068 23092 32070
rect 23116 32068 23172 32070
rect 23196 32068 23252 32070
rect 22956 31034 23012 31036
rect 23036 31034 23092 31036
rect 23116 31034 23172 31036
rect 23196 31034 23252 31036
rect 22956 30982 23002 31034
rect 23002 30982 23012 31034
rect 23036 30982 23066 31034
rect 23066 30982 23078 31034
rect 23078 30982 23092 31034
rect 23116 30982 23130 31034
rect 23130 30982 23142 31034
rect 23142 30982 23172 31034
rect 23196 30982 23206 31034
rect 23206 30982 23252 31034
rect 22956 30980 23012 30982
rect 23036 30980 23092 30982
rect 23116 30980 23172 30982
rect 23196 30980 23252 30982
rect 21638 15544 21694 15600
rect 22098 19216 22154 19272
rect 22956 29946 23012 29948
rect 23036 29946 23092 29948
rect 23116 29946 23172 29948
rect 23196 29946 23252 29948
rect 22956 29894 23002 29946
rect 23002 29894 23012 29946
rect 23036 29894 23066 29946
rect 23066 29894 23078 29946
rect 23078 29894 23092 29946
rect 23116 29894 23130 29946
rect 23130 29894 23142 29946
rect 23142 29894 23172 29946
rect 23196 29894 23206 29946
rect 23206 29894 23252 29946
rect 22956 29892 23012 29894
rect 23036 29892 23092 29894
rect 23116 29892 23172 29894
rect 23196 29892 23252 29894
rect 22956 28858 23012 28860
rect 23036 28858 23092 28860
rect 23116 28858 23172 28860
rect 23196 28858 23252 28860
rect 22956 28806 23002 28858
rect 23002 28806 23012 28858
rect 23036 28806 23066 28858
rect 23066 28806 23078 28858
rect 23078 28806 23092 28858
rect 23116 28806 23130 28858
rect 23130 28806 23142 28858
rect 23142 28806 23172 28858
rect 23196 28806 23206 28858
rect 23206 28806 23252 28858
rect 22956 28804 23012 28806
rect 23036 28804 23092 28806
rect 23116 28804 23172 28806
rect 23196 28804 23252 28806
rect 22956 27770 23012 27772
rect 23036 27770 23092 27772
rect 23116 27770 23172 27772
rect 23196 27770 23252 27772
rect 22956 27718 23002 27770
rect 23002 27718 23012 27770
rect 23036 27718 23066 27770
rect 23066 27718 23078 27770
rect 23078 27718 23092 27770
rect 23116 27718 23130 27770
rect 23130 27718 23142 27770
rect 23142 27718 23172 27770
rect 23196 27718 23206 27770
rect 23206 27718 23252 27770
rect 22956 27716 23012 27718
rect 23036 27716 23092 27718
rect 23116 27716 23172 27718
rect 23196 27716 23252 27718
rect 22956 26682 23012 26684
rect 23036 26682 23092 26684
rect 23116 26682 23172 26684
rect 23196 26682 23252 26684
rect 22956 26630 23002 26682
rect 23002 26630 23012 26682
rect 23036 26630 23066 26682
rect 23066 26630 23078 26682
rect 23078 26630 23092 26682
rect 23116 26630 23130 26682
rect 23130 26630 23142 26682
rect 23142 26630 23172 26682
rect 23196 26630 23206 26682
rect 23206 26630 23252 26682
rect 22956 26628 23012 26630
rect 23036 26628 23092 26630
rect 23116 26628 23172 26630
rect 23196 26628 23252 26630
rect 23570 26152 23626 26208
rect 22956 25594 23012 25596
rect 23036 25594 23092 25596
rect 23116 25594 23172 25596
rect 23196 25594 23252 25596
rect 22956 25542 23002 25594
rect 23002 25542 23012 25594
rect 23036 25542 23066 25594
rect 23066 25542 23078 25594
rect 23078 25542 23092 25594
rect 23116 25542 23130 25594
rect 23130 25542 23142 25594
rect 23142 25542 23172 25594
rect 23196 25542 23206 25594
rect 23206 25542 23252 25594
rect 22956 25540 23012 25542
rect 23036 25540 23092 25542
rect 23116 25540 23172 25542
rect 23196 25540 23252 25542
rect 22956 24506 23012 24508
rect 23036 24506 23092 24508
rect 23116 24506 23172 24508
rect 23196 24506 23252 24508
rect 22956 24454 23002 24506
rect 23002 24454 23012 24506
rect 23036 24454 23066 24506
rect 23066 24454 23078 24506
rect 23078 24454 23092 24506
rect 23116 24454 23130 24506
rect 23130 24454 23142 24506
rect 23142 24454 23172 24506
rect 23196 24454 23206 24506
rect 23206 24454 23252 24506
rect 22956 24452 23012 24454
rect 23036 24452 23092 24454
rect 23116 24452 23172 24454
rect 23196 24452 23252 24454
rect 22956 23418 23012 23420
rect 23036 23418 23092 23420
rect 23116 23418 23172 23420
rect 23196 23418 23252 23420
rect 22956 23366 23002 23418
rect 23002 23366 23012 23418
rect 23036 23366 23066 23418
rect 23066 23366 23078 23418
rect 23078 23366 23092 23418
rect 23116 23366 23130 23418
rect 23130 23366 23142 23418
rect 23142 23366 23172 23418
rect 23196 23366 23206 23418
rect 23206 23366 23252 23418
rect 22956 23364 23012 23366
rect 23036 23364 23092 23366
rect 23116 23364 23172 23366
rect 23196 23364 23252 23366
rect 22956 22330 23012 22332
rect 23036 22330 23092 22332
rect 23116 22330 23172 22332
rect 23196 22330 23252 22332
rect 22956 22278 23002 22330
rect 23002 22278 23012 22330
rect 23036 22278 23066 22330
rect 23066 22278 23078 22330
rect 23078 22278 23092 22330
rect 23116 22278 23130 22330
rect 23130 22278 23142 22330
rect 23142 22278 23172 22330
rect 23196 22278 23206 22330
rect 23206 22278 23252 22330
rect 22956 22276 23012 22278
rect 23036 22276 23092 22278
rect 23116 22276 23172 22278
rect 23196 22276 23252 22278
rect 24122 28736 24178 28792
rect 23386 23296 23442 23352
rect 22956 21242 23012 21244
rect 23036 21242 23092 21244
rect 23116 21242 23172 21244
rect 23196 21242 23252 21244
rect 22956 21190 23002 21242
rect 23002 21190 23012 21242
rect 23036 21190 23066 21242
rect 23066 21190 23078 21242
rect 23078 21190 23092 21242
rect 23116 21190 23130 21242
rect 23130 21190 23142 21242
rect 23142 21190 23172 21242
rect 23196 21190 23206 21242
rect 23206 21190 23252 21242
rect 22956 21188 23012 21190
rect 23036 21188 23092 21190
rect 23116 21188 23172 21190
rect 23196 21188 23252 21190
rect 22956 20154 23012 20156
rect 23036 20154 23092 20156
rect 23116 20154 23172 20156
rect 23196 20154 23252 20156
rect 22956 20102 23002 20154
rect 23002 20102 23012 20154
rect 23036 20102 23066 20154
rect 23066 20102 23078 20154
rect 23078 20102 23092 20154
rect 23116 20102 23130 20154
rect 23130 20102 23142 20154
rect 23142 20102 23172 20154
rect 23196 20102 23206 20154
rect 23206 20102 23252 20154
rect 22956 20100 23012 20102
rect 23036 20100 23092 20102
rect 23116 20100 23172 20102
rect 23196 20100 23252 20102
rect 22956 19066 23012 19068
rect 23036 19066 23092 19068
rect 23116 19066 23172 19068
rect 23196 19066 23252 19068
rect 22956 19014 23002 19066
rect 23002 19014 23012 19066
rect 23036 19014 23066 19066
rect 23066 19014 23078 19066
rect 23078 19014 23092 19066
rect 23116 19014 23130 19066
rect 23130 19014 23142 19066
rect 23142 19014 23172 19066
rect 23196 19014 23206 19066
rect 23206 19014 23252 19066
rect 22956 19012 23012 19014
rect 23036 19012 23092 19014
rect 23116 19012 23172 19014
rect 23196 19012 23252 19014
rect 23386 18536 23442 18592
rect 22956 17978 23012 17980
rect 23036 17978 23092 17980
rect 23116 17978 23172 17980
rect 23196 17978 23252 17980
rect 22956 17926 23002 17978
rect 23002 17926 23012 17978
rect 23036 17926 23066 17978
rect 23066 17926 23078 17978
rect 23078 17926 23092 17978
rect 23116 17926 23130 17978
rect 23130 17926 23142 17978
rect 23142 17926 23172 17978
rect 23196 17926 23206 17978
rect 23206 17926 23252 17978
rect 22956 17924 23012 17926
rect 23036 17924 23092 17926
rect 23116 17924 23172 17926
rect 23196 17924 23252 17926
rect 22956 16890 23012 16892
rect 23036 16890 23092 16892
rect 23116 16890 23172 16892
rect 23196 16890 23252 16892
rect 22956 16838 23002 16890
rect 23002 16838 23012 16890
rect 23036 16838 23066 16890
rect 23066 16838 23078 16890
rect 23078 16838 23092 16890
rect 23116 16838 23130 16890
rect 23130 16838 23142 16890
rect 23142 16838 23172 16890
rect 23196 16838 23206 16890
rect 23206 16838 23252 16890
rect 22956 16836 23012 16838
rect 23036 16836 23092 16838
rect 23116 16836 23172 16838
rect 23196 16836 23252 16838
rect 22956 15802 23012 15804
rect 23036 15802 23092 15804
rect 23116 15802 23172 15804
rect 23196 15802 23252 15804
rect 22956 15750 23002 15802
rect 23002 15750 23012 15802
rect 23036 15750 23066 15802
rect 23066 15750 23078 15802
rect 23078 15750 23092 15802
rect 23116 15750 23130 15802
rect 23130 15750 23142 15802
rect 23142 15750 23172 15802
rect 23196 15750 23206 15802
rect 23206 15750 23252 15802
rect 22956 15748 23012 15750
rect 23036 15748 23092 15750
rect 23116 15748 23172 15750
rect 23196 15748 23252 15750
rect 22956 14714 23012 14716
rect 23036 14714 23092 14716
rect 23116 14714 23172 14716
rect 23196 14714 23252 14716
rect 22956 14662 23002 14714
rect 23002 14662 23012 14714
rect 23036 14662 23066 14714
rect 23066 14662 23078 14714
rect 23078 14662 23092 14714
rect 23116 14662 23130 14714
rect 23130 14662 23142 14714
rect 23142 14662 23172 14714
rect 23196 14662 23206 14714
rect 23206 14662 23252 14714
rect 22956 14660 23012 14662
rect 23036 14660 23092 14662
rect 23116 14660 23172 14662
rect 23196 14660 23252 14662
rect 22956 13626 23012 13628
rect 23036 13626 23092 13628
rect 23116 13626 23172 13628
rect 23196 13626 23252 13628
rect 22956 13574 23002 13626
rect 23002 13574 23012 13626
rect 23036 13574 23066 13626
rect 23066 13574 23078 13626
rect 23078 13574 23092 13626
rect 23116 13574 23130 13626
rect 23130 13574 23142 13626
rect 23142 13574 23172 13626
rect 23196 13574 23206 13626
rect 23206 13574 23252 13626
rect 22956 13572 23012 13574
rect 23036 13572 23092 13574
rect 23116 13572 23172 13574
rect 23196 13572 23252 13574
rect 22956 12538 23012 12540
rect 23036 12538 23092 12540
rect 23116 12538 23172 12540
rect 23196 12538 23252 12540
rect 22956 12486 23002 12538
rect 23002 12486 23012 12538
rect 23036 12486 23066 12538
rect 23066 12486 23078 12538
rect 23078 12486 23092 12538
rect 23116 12486 23130 12538
rect 23130 12486 23142 12538
rect 23142 12486 23172 12538
rect 23196 12486 23206 12538
rect 23206 12486 23252 12538
rect 22956 12484 23012 12486
rect 23036 12484 23092 12486
rect 23116 12484 23172 12486
rect 23196 12484 23252 12486
rect 22956 11450 23012 11452
rect 23036 11450 23092 11452
rect 23116 11450 23172 11452
rect 23196 11450 23252 11452
rect 22956 11398 23002 11450
rect 23002 11398 23012 11450
rect 23036 11398 23066 11450
rect 23066 11398 23078 11450
rect 23078 11398 23092 11450
rect 23116 11398 23130 11450
rect 23130 11398 23142 11450
rect 23142 11398 23172 11450
rect 23196 11398 23206 11450
rect 23206 11398 23252 11450
rect 22956 11396 23012 11398
rect 23036 11396 23092 11398
rect 23116 11396 23172 11398
rect 23196 11396 23252 11398
rect 24766 38256 24822 38312
rect 25318 50496 25374 50552
rect 25318 49816 25374 49872
rect 25318 48456 25374 48512
rect 25502 47096 25558 47152
rect 24950 39616 25006 39672
rect 24950 36896 25006 36952
rect 24766 35536 24822 35592
rect 24858 28056 24914 28112
rect 24674 26696 24730 26752
rect 24490 21256 24546 21312
rect 22956 10362 23012 10364
rect 23036 10362 23092 10364
rect 23116 10362 23172 10364
rect 23196 10362 23252 10364
rect 22956 10310 23002 10362
rect 23002 10310 23012 10362
rect 23036 10310 23066 10362
rect 23066 10310 23078 10362
rect 23078 10310 23092 10362
rect 23116 10310 23130 10362
rect 23130 10310 23142 10362
rect 23142 10310 23172 10362
rect 23196 10310 23206 10362
rect 23206 10310 23252 10362
rect 22956 10308 23012 10310
rect 23036 10308 23092 10310
rect 23116 10308 23172 10310
rect 23196 10308 23252 10310
rect 22956 9274 23012 9276
rect 23036 9274 23092 9276
rect 23116 9274 23172 9276
rect 23196 9274 23252 9276
rect 22956 9222 23002 9274
rect 23002 9222 23012 9274
rect 23036 9222 23066 9274
rect 23066 9222 23078 9274
rect 23078 9222 23092 9274
rect 23116 9222 23130 9274
rect 23130 9222 23142 9274
rect 23142 9222 23172 9274
rect 23196 9222 23206 9274
rect 23206 9222 23252 9274
rect 22956 9220 23012 9222
rect 23036 9220 23092 9222
rect 23116 9220 23172 9222
rect 23196 9220 23252 9222
rect 22956 8186 23012 8188
rect 23036 8186 23092 8188
rect 23116 8186 23172 8188
rect 23196 8186 23252 8188
rect 22956 8134 23002 8186
rect 23002 8134 23012 8186
rect 23036 8134 23066 8186
rect 23066 8134 23078 8186
rect 23078 8134 23092 8186
rect 23116 8134 23130 8186
rect 23130 8134 23142 8186
rect 23142 8134 23172 8186
rect 23196 8134 23206 8186
rect 23206 8134 23252 8186
rect 22956 8132 23012 8134
rect 23036 8132 23092 8134
rect 23116 8132 23172 8134
rect 23196 8132 23252 8134
rect 22956 7098 23012 7100
rect 23036 7098 23092 7100
rect 23116 7098 23172 7100
rect 23196 7098 23252 7100
rect 22956 7046 23002 7098
rect 23002 7046 23012 7098
rect 23036 7046 23066 7098
rect 23066 7046 23078 7098
rect 23078 7046 23092 7098
rect 23116 7046 23130 7098
rect 23130 7046 23142 7098
rect 23142 7046 23172 7098
rect 23196 7046 23206 7098
rect 23206 7046 23252 7098
rect 22956 7044 23012 7046
rect 23036 7044 23092 7046
rect 23116 7044 23172 7046
rect 23196 7044 23252 7046
rect 22956 6010 23012 6012
rect 23036 6010 23092 6012
rect 23116 6010 23172 6012
rect 23196 6010 23252 6012
rect 22956 5958 23002 6010
rect 23002 5958 23012 6010
rect 23036 5958 23066 6010
rect 23066 5958 23078 6010
rect 23078 5958 23092 6010
rect 23116 5958 23130 6010
rect 23130 5958 23142 6010
rect 23142 5958 23172 6010
rect 23196 5958 23206 6010
rect 23206 5958 23252 6010
rect 22956 5956 23012 5958
rect 23036 5956 23092 5958
rect 23116 5956 23172 5958
rect 23196 5956 23252 5958
rect 22956 4922 23012 4924
rect 23036 4922 23092 4924
rect 23116 4922 23172 4924
rect 23196 4922 23252 4924
rect 22956 4870 23002 4922
rect 23002 4870 23012 4922
rect 23036 4870 23066 4922
rect 23066 4870 23078 4922
rect 23078 4870 23092 4922
rect 23116 4870 23130 4922
rect 23130 4870 23142 4922
rect 23142 4870 23172 4922
rect 23196 4870 23206 4922
rect 23206 4870 23252 4922
rect 22956 4868 23012 4870
rect 23036 4868 23092 4870
rect 23116 4868 23172 4870
rect 23196 4868 23252 4870
rect 23386 4256 23442 4312
rect 24858 23976 24914 24032
rect 24858 22616 24914 22672
rect 24858 21936 24914 21992
rect 24858 19896 24914 19952
rect 24766 17856 24822 17912
rect 24674 17176 24730 17232
rect 24858 16496 24914 16552
rect 24858 15816 24914 15872
rect 24858 14456 24914 14512
rect 24766 13776 24822 13832
rect 24674 13096 24730 13152
rect 24858 12416 24914 12472
rect 25502 43016 25558 43072
rect 25318 42336 25374 42392
rect 25502 41656 25558 41712
rect 25318 38936 25374 38992
rect 25410 37576 25466 37632
rect 25318 36216 25374 36272
rect 25318 34856 25374 34912
rect 25410 34176 25466 34232
rect 25318 33496 25374 33552
rect 25318 32852 25320 32872
rect 25320 32852 25372 32872
rect 25372 32852 25374 32872
rect 25318 32816 25374 32852
rect 25318 32136 25374 32192
rect 25318 31456 25374 31512
rect 25410 30776 25466 30832
rect 25318 30096 25374 30152
rect 25410 29416 25466 29472
rect 25410 27376 25466 27432
rect 25134 24656 25190 24712
rect 25134 20576 25190 20632
rect 25318 25336 25374 25392
rect 25134 15136 25190 15192
rect 24950 11736 25006 11792
rect 24766 11056 24822 11112
rect 24766 10376 24822 10432
rect 24858 9696 24914 9752
rect 25134 9016 25190 9072
rect 22956 3834 23012 3836
rect 23036 3834 23092 3836
rect 23116 3834 23172 3836
rect 23196 3834 23252 3836
rect 22956 3782 23002 3834
rect 23002 3782 23012 3834
rect 23036 3782 23066 3834
rect 23066 3782 23078 3834
rect 23078 3782 23092 3834
rect 23116 3782 23130 3834
rect 23130 3782 23142 3834
rect 23142 3782 23172 3834
rect 23196 3782 23206 3834
rect 23206 3782 23252 3834
rect 22956 3780 23012 3782
rect 23036 3780 23092 3782
rect 23116 3780 23172 3782
rect 23196 3780 23252 3782
rect 23294 3440 23350 3496
rect 22956 2746 23012 2748
rect 23036 2746 23092 2748
rect 23116 2746 23172 2748
rect 23196 2746 23252 2748
rect 22956 2694 23002 2746
rect 23002 2694 23012 2746
rect 23036 2694 23066 2746
rect 23066 2694 23078 2746
rect 23078 2694 23092 2746
rect 23116 2694 23130 2746
rect 23130 2694 23142 2746
rect 23142 2694 23172 2746
rect 23196 2694 23206 2746
rect 23206 2694 23252 2746
rect 22956 2692 23012 2694
rect 23036 2692 23092 2694
rect 23116 2692 23172 2694
rect 23196 2692 23252 2694
rect 24766 8336 24822 8392
rect 24950 7656 25006 7712
rect 24766 6976 24822 7032
rect 24858 6296 24914 6352
rect 24766 5616 24822 5672
rect 25318 4936 25374 4992
<< metal3 >>
rect 0 55042 800 55072
rect 2773 55042 2839 55045
rect 0 55040 2839 55042
rect 0 54984 2778 55040
rect 2834 54984 2839 55040
rect 0 54982 2839 54984
rect 0 54952 800 54982
rect 2773 54979 2839 54982
rect 7946 54432 8262 54433
rect 7946 54368 7952 54432
rect 8016 54368 8032 54432
rect 8096 54368 8112 54432
rect 8176 54368 8192 54432
rect 8256 54368 8262 54432
rect 7946 54367 8262 54368
rect 17946 54432 18262 54433
rect 17946 54368 17952 54432
rect 18016 54368 18032 54432
rect 18096 54368 18112 54432
rect 18176 54368 18192 54432
rect 18256 54368 18262 54432
rect 17946 54367 18262 54368
rect 15653 53954 15719 53957
rect 15878 53954 15884 53956
rect 15653 53952 15884 53954
rect 15653 53896 15658 53952
rect 15714 53896 15884 53952
rect 15653 53894 15884 53896
rect 15653 53891 15719 53894
rect 15878 53892 15884 53894
rect 15948 53892 15954 53956
rect 2946 53888 3262 53889
rect 2946 53824 2952 53888
rect 3016 53824 3032 53888
rect 3096 53824 3112 53888
rect 3176 53824 3192 53888
rect 3256 53824 3262 53888
rect 2946 53823 3262 53824
rect 12946 53888 13262 53889
rect 12946 53824 12952 53888
rect 13016 53824 13032 53888
rect 13096 53824 13112 53888
rect 13176 53824 13192 53888
rect 13256 53824 13262 53888
rect 12946 53823 13262 53824
rect 22946 53888 23262 53889
rect 22946 53824 22952 53888
rect 23016 53824 23032 53888
rect 23096 53824 23112 53888
rect 23176 53824 23192 53888
rect 23256 53824 23262 53888
rect 22946 53823 23262 53824
rect 7946 53344 8262 53345
rect 7946 53280 7952 53344
rect 8016 53280 8032 53344
rect 8096 53280 8112 53344
rect 8176 53280 8192 53344
rect 8256 53280 8262 53344
rect 7946 53279 8262 53280
rect 17946 53344 18262 53345
rect 17946 53280 17952 53344
rect 18016 53280 18032 53344
rect 18096 53280 18112 53344
rect 18176 53280 18192 53344
rect 18256 53280 18262 53344
rect 17946 53279 18262 53280
rect 2946 52800 3262 52801
rect 0 52730 800 52760
rect 2946 52736 2952 52800
rect 3016 52736 3032 52800
rect 3096 52736 3112 52800
rect 3176 52736 3192 52800
rect 3256 52736 3262 52800
rect 2946 52735 3262 52736
rect 12946 52800 13262 52801
rect 12946 52736 12952 52800
rect 13016 52736 13032 52800
rect 13096 52736 13112 52800
rect 13176 52736 13192 52800
rect 13256 52736 13262 52800
rect 12946 52735 13262 52736
rect 22946 52800 23262 52801
rect 22946 52736 22952 52800
rect 23016 52736 23032 52800
rect 23096 52736 23112 52800
rect 23176 52736 23192 52800
rect 23256 52736 23262 52800
rect 22946 52735 23262 52736
rect 1209 52730 1275 52733
rect 0 52728 1275 52730
rect 0 52672 1214 52728
rect 1270 52672 1275 52728
rect 0 52670 1275 52672
rect 0 52640 800 52670
rect 1209 52667 1275 52670
rect 14365 52596 14431 52597
rect 14365 52592 14412 52596
rect 14476 52594 14482 52596
rect 14365 52536 14370 52592
rect 14365 52532 14412 52536
rect 14476 52534 14522 52594
rect 14476 52532 14482 52534
rect 15694 52532 15700 52596
rect 15764 52594 15770 52596
rect 15929 52594 15995 52597
rect 15764 52592 15995 52594
rect 15764 52536 15934 52592
rect 15990 52536 15995 52592
rect 15764 52534 15995 52536
rect 15764 52532 15770 52534
rect 14365 52531 14431 52532
rect 15929 52531 15995 52534
rect 22185 52594 22251 52597
rect 22318 52594 22324 52596
rect 22185 52592 22324 52594
rect 22185 52536 22190 52592
rect 22246 52536 22324 52592
rect 22185 52534 22324 52536
rect 22185 52531 22251 52534
rect 22318 52532 22324 52534
rect 22388 52532 22394 52596
rect 24669 52594 24735 52597
rect 26200 52594 27000 52624
rect 24669 52592 27000 52594
rect 24669 52536 24674 52592
rect 24730 52536 27000 52592
rect 24669 52534 27000 52536
rect 24669 52531 24735 52534
rect 26200 52504 27000 52534
rect 7946 52256 8262 52257
rect 7946 52192 7952 52256
rect 8016 52192 8032 52256
rect 8096 52192 8112 52256
rect 8176 52192 8192 52256
rect 8256 52192 8262 52256
rect 7946 52191 8262 52192
rect 17946 52256 18262 52257
rect 17946 52192 17952 52256
rect 18016 52192 18032 52256
rect 18096 52192 18112 52256
rect 18176 52192 18192 52256
rect 18256 52192 18262 52256
rect 17946 52191 18262 52192
rect 25221 51914 25287 51917
rect 26200 51914 27000 51944
rect 25221 51912 27000 51914
rect 25221 51856 25226 51912
rect 25282 51856 27000 51912
rect 25221 51854 27000 51856
rect 25221 51851 25287 51854
rect 26200 51824 27000 51854
rect 2946 51712 3262 51713
rect 2946 51648 2952 51712
rect 3016 51648 3032 51712
rect 3096 51648 3112 51712
rect 3176 51648 3192 51712
rect 3256 51648 3262 51712
rect 2946 51647 3262 51648
rect 12946 51712 13262 51713
rect 12946 51648 12952 51712
rect 13016 51648 13032 51712
rect 13096 51648 13112 51712
rect 13176 51648 13192 51712
rect 13256 51648 13262 51712
rect 12946 51647 13262 51648
rect 22946 51712 23262 51713
rect 22946 51648 22952 51712
rect 23016 51648 23032 51712
rect 23096 51648 23112 51712
rect 23176 51648 23192 51712
rect 23256 51648 23262 51712
rect 22946 51647 23262 51648
rect 25313 51234 25379 51237
rect 26200 51234 27000 51264
rect 25313 51232 27000 51234
rect 25313 51176 25318 51232
rect 25374 51176 27000 51232
rect 25313 51174 27000 51176
rect 25313 51171 25379 51174
rect 7946 51168 8262 51169
rect 7946 51104 7952 51168
rect 8016 51104 8032 51168
rect 8096 51104 8112 51168
rect 8176 51104 8192 51168
rect 8256 51104 8262 51168
rect 7946 51103 8262 51104
rect 17946 51168 18262 51169
rect 17946 51104 17952 51168
rect 18016 51104 18032 51168
rect 18096 51104 18112 51168
rect 18176 51104 18192 51168
rect 18256 51104 18262 51168
rect 26200 51144 27000 51174
rect 17946 51103 18262 51104
rect 2946 50624 3262 50625
rect 2946 50560 2952 50624
rect 3016 50560 3032 50624
rect 3096 50560 3112 50624
rect 3176 50560 3192 50624
rect 3256 50560 3262 50624
rect 2946 50559 3262 50560
rect 12946 50624 13262 50625
rect 12946 50560 12952 50624
rect 13016 50560 13032 50624
rect 13096 50560 13112 50624
rect 13176 50560 13192 50624
rect 13256 50560 13262 50624
rect 12946 50559 13262 50560
rect 22946 50624 23262 50625
rect 22946 50560 22952 50624
rect 23016 50560 23032 50624
rect 23096 50560 23112 50624
rect 23176 50560 23192 50624
rect 23256 50560 23262 50624
rect 22946 50559 23262 50560
rect 25313 50554 25379 50557
rect 26200 50554 27000 50584
rect 25313 50552 27000 50554
rect 25313 50496 25318 50552
rect 25374 50496 27000 50552
rect 25313 50494 27000 50496
rect 25313 50491 25379 50494
rect 26200 50464 27000 50494
rect 0 50418 800 50448
rect 1117 50418 1183 50421
rect 0 50416 1183 50418
rect 0 50360 1122 50416
rect 1178 50360 1183 50416
rect 0 50358 1183 50360
rect 0 50328 800 50358
rect 1117 50355 1183 50358
rect 7946 50080 8262 50081
rect 7946 50016 7952 50080
rect 8016 50016 8032 50080
rect 8096 50016 8112 50080
rect 8176 50016 8192 50080
rect 8256 50016 8262 50080
rect 7946 50015 8262 50016
rect 17946 50080 18262 50081
rect 17946 50016 17952 50080
rect 18016 50016 18032 50080
rect 18096 50016 18112 50080
rect 18176 50016 18192 50080
rect 18256 50016 18262 50080
rect 17946 50015 18262 50016
rect 25313 49874 25379 49877
rect 26200 49874 27000 49904
rect 25313 49872 27000 49874
rect 25313 49816 25318 49872
rect 25374 49816 27000 49872
rect 25313 49814 27000 49816
rect 25313 49811 25379 49814
rect 26200 49784 27000 49814
rect 2946 49536 3262 49537
rect 2946 49472 2952 49536
rect 3016 49472 3032 49536
rect 3096 49472 3112 49536
rect 3176 49472 3192 49536
rect 3256 49472 3262 49536
rect 2946 49471 3262 49472
rect 12946 49536 13262 49537
rect 12946 49472 12952 49536
rect 13016 49472 13032 49536
rect 13096 49472 13112 49536
rect 13176 49472 13192 49536
rect 13256 49472 13262 49536
rect 12946 49471 13262 49472
rect 22946 49536 23262 49537
rect 22946 49472 22952 49536
rect 23016 49472 23032 49536
rect 23096 49472 23112 49536
rect 23176 49472 23192 49536
rect 23256 49472 23262 49536
rect 22946 49471 23262 49472
rect 24761 49194 24827 49197
rect 26200 49194 27000 49224
rect 24761 49192 27000 49194
rect 24761 49136 24766 49192
rect 24822 49136 27000 49192
rect 24761 49134 27000 49136
rect 24761 49131 24827 49134
rect 26200 49104 27000 49134
rect 7946 48992 8262 48993
rect 7946 48928 7952 48992
rect 8016 48928 8032 48992
rect 8096 48928 8112 48992
rect 8176 48928 8192 48992
rect 8256 48928 8262 48992
rect 7946 48927 8262 48928
rect 17946 48992 18262 48993
rect 17946 48928 17952 48992
rect 18016 48928 18032 48992
rect 18096 48928 18112 48992
rect 18176 48928 18192 48992
rect 18256 48928 18262 48992
rect 17946 48927 18262 48928
rect 25313 48514 25379 48517
rect 26200 48514 27000 48544
rect 25313 48512 27000 48514
rect 25313 48456 25318 48512
rect 25374 48456 27000 48512
rect 25313 48454 27000 48456
rect 25313 48451 25379 48454
rect 2946 48448 3262 48449
rect 2946 48384 2952 48448
rect 3016 48384 3032 48448
rect 3096 48384 3112 48448
rect 3176 48384 3192 48448
rect 3256 48384 3262 48448
rect 2946 48383 3262 48384
rect 12946 48448 13262 48449
rect 12946 48384 12952 48448
rect 13016 48384 13032 48448
rect 13096 48384 13112 48448
rect 13176 48384 13192 48448
rect 13256 48384 13262 48448
rect 12946 48383 13262 48384
rect 22946 48448 23262 48449
rect 22946 48384 22952 48448
rect 23016 48384 23032 48448
rect 23096 48384 23112 48448
rect 23176 48384 23192 48448
rect 23256 48384 23262 48448
rect 26200 48424 27000 48454
rect 22946 48383 23262 48384
rect 0 48106 800 48136
rect 1301 48106 1367 48109
rect 0 48104 1367 48106
rect 0 48048 1306 48104
rect 1362 48048 1367 48104
rect 0 48046 1367 48048
rect 0 48016 800 48046
rect 1301 48043 1367 48046
rect 7946 47904 8262 47905
rect 7946 47840 7952 47904
rect 8016 47840 8032 47904
rect 8096 47840 8112 47904
rect 8176 47840 8192 47904
rect 8256 47840 8262 47904
rect 7946 47839 8262 47840
rect 17946 47904 18262 47905
rect 17946 47840 17952 47904
rect 18016 47840 18032 47904
rect 18096 47840 18112 47904
rect 18176 47840 18192 47904
rect 18256 47840 18262 47904
rect 17946 47839 18262 47840
rect 24761 47834 24827 47837
rect 26200 47834 27000 47864
rect 24761 47832 27000 47834
rect 24761 47776 24766 47832
rect 24822 47776 27000 47832
rect 24761 47774 27000 47776
rect 24761 47771 24827 47774
rect 26200 47744 27000 47774
rect 2946 47360 3262 47361
rect 2946 47296 2952 47360
rect 3016 47296 3032 47360
rect 3096 47296 3112 47360
rect 3176 47296 3192 47360
rect 3256 47296 3262 47360
rect 2946 47295 3262 47296
rect 12946 47360 13262 47361
rect 12946 47296 12952 47360
rect 13016 47296 13032 47360
rect 13096 47296 13112 47360
rect 13176 47296 13192 47360
rect 13256 47296 13262 47360
rect 12946 47295 13262 47296
rect 22946 47360 23262 47361
rect 22946 47296 22952 47360
rect 23016 47296 23032 47360
rect 23096 47296 23112 47360
rect 23176 47296 23192 47360
rect 23256 47296 23262 47360
rect 22946 47295 23262 47296
rect 25497 47154 25563 47157
rect 26200 47154 27000 47184
rect 25497 47152 27000 47154
rect 25497 47096 25502 47152
rect 25558 47096 27000 47152
rect 25497 47094 27000 47096
rect 25497 47091 25563 47094
rect 26200 47064 27000 47094
rect 7946 46816 8262 46817
rect 7946 46752 7952 46816
rect 8016 46752 8032 46816
rect 8096 46752 8112 46816
rect 8176 46752 8192 46816
rect 8256 46752 8262 46816
rect 7946 46751 8262 46752
rect 17946 46816 18262 46817
rect 17946 46752 17952 46816
rect 18016 46752 18032 46816
rect 18096 46752 18112 46816
rect 18176 46752 18192 46816
rect 18256 46752 18262 46816
rect 17946 46751 18262 46752
rect 24853 46474 24919 46477
rect 26200 46474 27000 46504
rect 24853 46472 27000 46474
rect 24853 46416 24858 46472
rect 24914 46416 27000 46472
rect 24853 46414 27000 46416
rect 24853 46411 24919 46414
rect 26200 46384 27000 46414
rect 2946 46272 3262 46273
rect 2946 46208 2952 46272
rect 3016 46208 3032 46272
rect 3096 46208 3112 46272
rect 3176 46208 3192 46272
rect 3256 46208 3262 46272
rect 2946 46207 3262 46208
rect 12946 46272 13262 46273
rect 12946 46208 12952 46272
rect 13016 46208 13032 46272
rect 13096 46208 13112 46272
rect 13176 46208 13192 46272
rect 13256 46208 13262 46272
rect 12946 46207 13262 46208
rect 22946 46272 23262 46273
rect 22946 46208 22952 46272
rect 23016 46208 23032 46272
rect 23096 46208 23112 46272
rect 23176 46208 23192 46272
rect 23256 46208 23262 46272
rect 22946 46207 23262 46208
rect 0 45794 800 45824
rect 1209 45794 1275 45797
rect 20529 45796 20595 45797
rect 20478 45794 20484 45796
rect 0 45792 1275 45794
rect 0 45736 1214 45792
rect 1270 45736 1275 45792
rect 0 45734 1275 45736
rect 20438 45734 20484 45794
rect 20548 45792 20595 45796
rect 20590 45736 20595 45792
rect 0 45704 800 45734
rect 1209 45731 1275 45734
rect 20478 45732 20484 45734
rect 20548 45732 20595 45736
rect 20529 45731 20595 45732
rect 24761 45794 24827 45797
rect 26200 45794 27000 45824
rect 24761 45792 27000 45794
rect 24761 45736 24766 45792
rect 24822 45736 27000 45792
rect 24761 45734 27000 45736
rect 24761 45731 24827 45734
rect 7946 45728 8262 45729
rect 7946 45664 7952 45728
rect 8016 45664 8032 45728
rect 8096 45664 8112 45728
rect 8176 45664 8192 45728
rect 8256 45664 8262 45728
rect 7946 45663 8262 45664
rect 17946 45728 18262 45729
rect 17946 45664 17952 45728
rect 18016 45664 18032 45728
rect 18096 45664 18112 45728
rect 18176 45664 18192 45728
rect 18256 45664 18262 45728
rect 26200 45704 27000 45734
rect 17946 45663 18262 45664
rect 21449 45524 21515 45525
rect 21398 45460 21404 45524
rect 21468 45522 21515 45524
rect 22645 45522 22711 45525
rect 21468 45520 22711 45522
rect 21510 45464 22650 45520
rect 22706 45464 22711 45520
rect 21468 45462 22711 45464
rect 21468 45460 21515 45462
rect 21449 45459 21515 45460
rect 22645 45459 22711 45462
rect 12014 45188 12020 45252
rect 12084 45250 12090 45252
rect 12249 45250 12315 45253
rect 12084 45248 12315 45250
rect 12084 45192 12254 45248
rect 12310 45192 12315 45248
rect 12084 45190 12315 45192
rect 12084 45188 12090 45190
rect 12249 45187 12315 45190
rect 2946 45184 3262 45185
rect 2946 45120 2952 45184
rect 3016 45120 3032 45184
rect 3096 45120 3112 45184
rect 3176 45120 3192 45184
rect 3256 45120 3262 45184
rect 2946 45119 3262 45120
rect 12946 45184 13262 45185
rect 12946 45120 12952 45184
rect 13016 45120 13032 45184
rect 13096 45120 13112 45184
rect 13176 45120 13192 45184
rect 13256 45120 13262 45184
rect 12946 45119 13262 45120
rect 22946 45184 23262 45185
rect 22946 45120 22952 45184
rect 23016 45120 23032 45184
rect 23096 45120 23112 45184
rect 23176 45120 23192 45184
rect 23256 45120 23262 45184
rect 22946 45119 23262 45120
rect 23841 45114 23907 45117
rect 26200 45114 27000 45144
rect 23841 45112 27000 45114
rect 23841 45056 23846 45112
rect 23902 45056 27000 45112
rect 23841 45054 27000 45056
rect 23841 45051 23907 45054
rect 26200 45024 27000 45054
rect 9673 44706 9739 44709
rect 9806 44706 9812 44708
rect 9673 44704 9812 44706
rect 9673 44648 9678 44704
rect 9734 44648 9812 44704
rect 9673 44646 9812 44648
rect 9673 44643 9739 44646
rect 9806 44644 9812 44646
rect 9876 44644 9882 44708
rect 7946 44640 8262 44641
rect 7946 44576 7952 44640
rect 8016 44576 8032 44640
rect 8096 44576 8112 44640
rect 8176 44576 8192 44640
rect 8256 44576 8262 44640
rect 7946 44575 8262 44576
rect 17946 44640 18262 44641
rect 17946 44576 17952 44640
rect 18016 44576 18032 44640
rect 18096 44576 18112 44640
rect 18176 44576 18192 44640
rect 18256 44576 18262 44640
rect 17946 44575 18262 44576
rect 24761 44434 24827 44437
rect 26200 44434 27000 44464
rect 24761 44432 27000 44434
rect 24761 44376 24766 44432
rect 24822 44376 27000 44432
rect 24761 44374 27000 44376
rect 24761 44371 24827 44374
rect 26200 44344 27000 44374
rect 19374 44236 19380 44300
rect 19444 44298 19450 44300
rect 19517 44298 19583 44301
rect 19444 44296 19583 44298
rect 19444 44240 19522 44296
rect 19578 44240 19583 44296
rect 19444 44238 19583 44240
rect 19444 44236 19450 44238
rect 19517 44235 19583 44238
rect 21030 44236 21036 44300
rect 21100 44298 21106 44300
rect 21449 44298 21515 44301
rect 21100 44296 21515 44298
rect 21100 44240 21454 44296
rect 21510 44240 21515 44296
rect 21100 44238 21515 44240
rect 21100 44236 21106 44238
rect 21449 44235 21515 44238
rect 2946 44096 3262 44097
rect 2946 44032 2952 44096
rect 3016 44032 3032 44096
rect 3096 44032 3112 44096
rect 3176 44032 3192 44096
rect 3256 44032 3262 44096
rect 2946 44031 3262 44032
rect 12946 44096 13262 44097
rect 12946 44032 12952 44096
rect 13016 44032 13032 44096
rect 13096 44032 13112 44096
rect 13176 44032 13192 44096
rect 13256 44032 13262 44096
rect 12946 44031 13262 44032
rect 22946 44096 23262 44097
rect 22946 44032 22952 44096
rect 23016 44032 23032 44096
rect 23096 44032 23112 44096
rect 23176 44032 23192 44096
rect 23256 44032 23262 44096
rect 22946 44031 23262 44032
rect 24669 43754 24735 43757
rect 26200 43754 27000 43784
rect 24669 43752 27000 43754
rect 24669 43696 24674 43752
rect 24730 43696 27000 43752
rect 24669 43694 27000 43696
rect 24669 43691 24735 43694
rect 26200 43664 27000 43694
rect 7946 43552 8262 43553
rect 0 43482 800 43512
rect 7946 43488 7952 43552
rect 8016 43488 8032 43552
rect 8096 43488 8112 43552
rect 8176 43488 8192 43552
rect 8256 43488 8262 43552
rect 7946 43487 8262 43488
rect 17946 43552 18262 43553
rect 17946 43488 17952 43552
rect 18016 43488 18032 43552
rect 18096 43488 18112 43552
rect 18176 43488 18192 43552
rect 18256 43488 18262 43552
rect 17946 43487 18262 43488
rect 1301 43482 1367 43485
rect 0 43480 1367 43482
rect 0 43424 1306 43480
rect 1362 43424 1367 43480
rect 0 43422 1367 43424
rect 0 43392 800 43422
rect 1301 43419 1367 43422
rect 25497 43074 25563 43077
rect 26200 43074 27000 43104
rect 25497 43072 27000 43074
rect 25497 43016 25502 43072
rect 25558 43016 27000 43072
rect 25497 43014 27000 43016
rect 25497 43011 25563 43014
rect 2946 43008 3262 43009
rect 2946 42944 2952 43008
rect 3016 42944 3032 43008
rect 3096 42944 3112 43008
rect 3176 42944 3192 43008
rect 3256 42944 3262 43008
rect 2946 42943 3262 42944
rect 12946 43008 13262 43009
rect 12946 42944 12952 43008
rect 13016 42944 13032 43008
rect 13096 42944 13112 43008
rect 13176 42944 13192 43008
rect 13256 42944 13262 43008
rect 12946 42943 13262 42944
rect 22946 43008 23262 43009
rect 22946 42944 22952 43008
rect 23016 42944 23032 43008
rect 23096 42944 23112 43008
rect 23176 42944 23192 43008
rect 23256 42944 23262 43008
rect 26200 42984 27000 43014
rect 22946 42943 23262 42944
rect 7946 42464 8262 42465
rect 7946 42400 7952 42464
rect 8016 42400 8032 42464
rect 8096 42400 8112 42464
rect 8176 42400 8192 42464
rect 8256 42400 8262 42464
rect 7946 42399 8262 42400
rect 17946 42464 18262 42465
rect 17946 42400 17952 42464
rect 18016 42400 18032 42464
rect 18096 42400 18112 42464
rect 18176 42400 18192 42464
rect 18256 42400 18262 42464
rect 17946 42399 18262 42400
rect 25313 42394 25379 42397
rect 26200 42394 27000 42424
rect 25313 42392 27000 42394
rect 25313 42336 25318 42392
rect 25374 42336 27000 42392
rect 25313 42334 27000 42336
rect 25313 42331 25379 42334
rect 26200 42304 27000 42334
rect 2946 41920 3262 41921
rect 2946 41856 2952 41920
rect 3016 41856 3032 41920
rect 3096 41856 3112 41920
rect 3176 41856 3192 41920
rect 3256 41856 3262 41920
rect 2946 41855 3262 41856
rect 12946 41920 13262 41921
rect 12946 41856 12952 41920
rect 13016 41856 13032 41920
rect 13096 41856 13112 41920
rect 13176 41856 13192 41920
rect 13256 41856 13262 41920
rect 12946 41855 13262 41856
rect 22946 41920 23262 41921
rect 22946 41856 22952 41920
rect 23016 41856 23032 41920
rect 23096 41856 23112 41920
rect 23176 41856 23192 41920
rect 23256 41856 23262 41920
rect 22946 41855 23262 41856
rect 25497 41714 25563 41717
rect 26200 41714 27000 41744
rect 25497 41712 27000 41714
rect 25497 41656 25502 41712
rect 25558 41656 27000 41712
rect 25497 41654 27000 41656
rect 25497 41651 25563 41654
rect 26200 41624 27000 41654
rect 21173 41444 21239 41445
rect 21173 41442 21220 41444
rect 21128 41440 21220 41442
rect 21128 41384 21178 41440
rect 21128 41382 21220 41384
rect 21173 41380 21220 41382
rect 21284 41380 21290 41444
rect 21173 41379 21239 41380
rect 7946 41376 8262 41377
rect 7946 41312 7952 41376
rect 8016 41312 8032 41376
rect 8096 41312 8112 41376
rect 8176 41312 8192 41376
rect 8256 41312 8262 41376
rect 7946 41311 8262 41312
rect 17946 41376 18262 41377
rect 17946 41312 17952 41376
rect 18016 41312 18032 41376
rect 18096 41312 18112 41376
rect 18176 41312 18192 41376
rect 18256 41312 18262 41376
rect 17946 41311 18262 41312
rect 11329 41306 11395 41309
rect 13670 41306 13676 41308
rect 11329 41304 13676 41306
rect 11329 41248 11334 41304
rect 11390 41248 13676 41304
rect 11329 41246 13676 41248
rect 11329 41243 11395 41246
rect 13670 41244 13676 41246
rect 13740 41244 13746 41308
rect 0 41170 800 41200
rect 1669 41170 1735 41173
rect 0 41168 1735 41170
rect 0 41112 1674 41168
rect 1730 41112 1735 41168
rect 0 41110 1735 41112
rect 0 41080 800 41110
rect 1669 41107 1735 41110
rect 24761 41034 24827 41037
rect 26200 41034 27000 41064
rect 24761 41032 27000 41034
rect 24761 40976 24766 41032
rect 24822 40976 27000 41032
rect 24761 40974 27000 40976
rect 24761 40971 24827 40974
rect 26200 40944 27000 40974
rect 2946 40832 3262 40833
rect 2946 40768 2952 40832
rect 3016 40768 3032 40832
rect 3096 40768 3112 40832
rect 3176 40768 3192 40832
rect 3256 40768 3262 40832
rect 2946 40767 3262 40768
rect 12946 40832 13262 40833
rect 12946 40768 12952 40832
rect 13016 40768 13032 40832
rect 13096 40768 13112 40832
rect 13176 40768 13192 40832
rect 13256 40768 13262 40832
rect 12946 40767 13262 40768
rect 22946 40832 23262 40833
rect 22946 40768 22952 40832
rect 23016 40768 23032 40832
rect 23096 40768 23112 40832
rect 23176 40768 23192 40832
rect 23256 40768 23262 40832
rect 22946 40767 23262 40768
rect 13445 40762 13511 40765
rect 14590 40762 14596 40764
rect 13445 40760 14596 40762
rect 13445 40704 13450 40760
rect 13506 40704 14596 40760
rect 13445 40702 14596 40704
rect 13445 40699 13511 40702
rect 14590 40700 14596 40702
rect 14660 40700 14666 40764
rect 23381 40354 23447 40357
rect 26200 40354 27000 40384
rect 23381 40352 27000 40354
rect 23381 40296 23386 40352
rect 23442 40296 27000 40352
rect 23381 40294 27000 40296
rect 23381 40291 23447 40294
rect 7946 40288 8262 40289
rect 7946 40224 7952 40288
rect 8016 40224 8032 40288
rect 8096 40224 8112 40288
rect 8176 40224 8192 40288
rect 8256 40224 8262 40288
rect 7946 40223 8262 40224
rect 17946 40288 18262 40289
rect 17946 40224 17952 40288
rect 18016 40224 18032 40288
rect 18096 40224 18112 40288
rect 18176 40224 18192 40288
rect 18256 40224 18262 40288
rect 26200 40264 27000 40294
rect 17946 40223 18262 40224
rect 2946 39744 3262 39745
rect 2946 39680 2952 39744
rect 3016 39680 3032 39744
rect 3096 39680 3112 39744
rect 3176 39680 3192 39744
rect 3256 39680 3262 39744
rect 2946 39679 3262 39680
rect 12946 39744 13262 39745
rect 12946 39680 12952 39744
rect 13016 39680 13032 39744
rect 13096 39680 13112 39744
rect 13176 39680 13192 39744
rect 13256 39680 13262 39744
rect 12946 39679 13262 39680
rect 22946 39744 23262 39745
rect 22946 39680 22952 39744
rect 23016 39680 23032 39744
rect 23096 39680 23112 39744
rect 23176 39680 23192 39744
rect 23256 39680 23262 39744
rect 22946 39679 23262 39680
rect 24945 39674 25011 39677
rect 26200 39674 27000 39704
rect 24945 39672 27000 39674
rect 24945 39616 24950 39672
rect 25006 39616 27000 39672
rect 24945 39614 27000 39616
rect 24945 39611 25011 39614
rect 26200 39584 27000 39614
rect 7946 39200 8262 39201
rect 7946 39136 7952 39200
rect 8016 39136 8032 39200
rect 8096 39136 8112 39200
rect 8176 39136 8192 39200
rect 8256 39136 8262 39200
rect 7946 39135 8262 39136
rect 17946 39200 18262 39201
rect 17946 39136 17952 39200
rect 18016 39136 18032 39200
rect 18096 39136 18112 39200
rect 18176 39136 18192 39200
rect 18256 39136 18262 39200
rect 17946 39135 18262 39136
rect 17534 38932 17540 38996
rect 17604 38994 17610 38996
rect 19885 38994 19951 38997
rect 17604 38992 19951 38994
rect 17604 38936 19890 38992
rect 19946 38936 19951 38992
rect 17604 38934 19951 38936
rect 17604 38932 17610 38934
rect 19885 38931 19951 38934
rect 25313 38994 25379 38997
rect 26200 38994 27000 39024
rect 25313 38992 27000 38994
rect 25313 38936 25318 38992
rect 25374 38936 27000 38992
rect 25313 38934 27000 38936
rect 25313 38931 25379 38934
rect 26200 38904 27000 38934
rect 0 38858 800 38888
rect 1209 38858 1275 38861
rect 0 38856 1275 38858
rect 0 38800 1214 38856
rect 1270 38800 1275 38856
rect 0 38798 1275 38800
rect 0 38768 800 38798
rect 1209 38795 1275 38798
rect 15142 38660 15148 38724
rect 15212 38722 15218 38724
rect 15285 38722 15351 38725
rect 15212 38720 15351 38722
rect 15212 38664 15290 38720
rect 15346 38664 15351 38720
rect 15212 38662 15351 38664
rect 15212 38660 15218 38662
rect 15285 38659 15351 38662
rect 18413 38724 18479 38725
rect 18413 38720 18460 38724
rect 18524 38722 18530 38724
rect 18413 38664 18418 38720
rect 18413 38660 18460 38664
rect 18524 38662 18570 38722
rect 18524 38660 18530 38662
rect 18413 38659 18479 38660
rect 2946 38656 3262 38657
rect 2946 38592 2952 38656
rect 3016 38592 3032 38656
rect 3096 38592 3112 38656
rect 3176 38592 3192 38656
rect 3256 38592 3262 38656
rect 2946 38591 3262 38592
rect 12946 38656 13262 38657
rect 12946 38592 12952 38656
rect 13016 38592 13032 38656
rect 13096 38592 13112 38656
rect 13176 38592 13192 38656
rect 13256 38592 13262 38656
rect 12946 38591 13262 38592
rect 22946 38656 23262 38657
rect 22946 38592 22952 38656
rect 23016 38592 23032 38656
rect 23096 38592 23112 38656
rect 23176 38592 23192 38656
rect 23256 38592 23262 38656
rect 22946 38591 23262 38592
rect 24761 38314 24827 38317
rect 26200 38314 27000 38344
rect 24761 38312 27000 38314
rect 24761 38256 24766 38312
rect 24822 38256 27000 38312
rect 24761 38254 27000 38256
rect 24761 38251 24827 38254
rect 26200 38224 27000 38254
rect 7946 38112 8262 38113
rect 7946 38048 7952 38112
rect 8016 38048 8032 38112
rect 8096 38048 8112 38112
rect 8176 38048 8192 38112
rect 8256 38048 8262 38112
rect 7946 38047 8262 38048
rect 17946 38112 18262 38113
rect 17946 38048 17952 38112
rect 18016 38048 18032 38112
rect 18096 38048 18112 38112
rect 18176 38048 18192 38112
rect 18256 38048 18262 38112
rect 17946 38047 18262 38048
rect 18873 37770 18939 37773
rect 18830 37768 18939 37770
rect 18830 37712 18878 37768
rect 18934 37712 18939 37768
rect 18830 37707 18939 37712
rect 18638 37572 18644 37636
rect 18708 37634 18714 37636
rect 18830 37634 18890 37707
rect 19885 37634 19951 37637
rect 18708 37632 19951 37634
rect 18708 37576 19890 37632
rect 19946 37576 19951 37632
rect 18708 37574 19951 37576
rect 18708 37572 18714 37574
rect 19885 37571 19951 37574
rect 25405 37634 25471 37637
rect 26200 37634 27000 37664
rect 25405 37632 27000 37634
rect 25405 37576 25410 37632
rect 25466 37576 27000 37632
rect 25405 37574 27000 37576
rect 25405 37571 25471 37574
rect 2946 37568 3262 37569
rect 2946 37504 2952 37568
rect 3016 37504 3032 37568
rect 3096 37504 3112 37568
rect 3176 37504 3192 37568
rect 3256 37504 3262 37568
rect 2946 37503 3262 37504
rect 12946 37568 13262 37569
rect 12946 37504 12952 37568
rect 13016 37504 13032 37568
rect 13096 37504 13112 37568
rect 13176 37504 13192 37568
rect 13256 37504 13262 37568
rect 12946 37503 13262 37504
rect 22946 37568 23262 37569
rect 22946 37504 22952 37568
rect 23016 37504 23032 37568
rect 23096 37504 23112 37568
rect 23176 37504 23192 37568
rect 23256 37504 23262 37568
rect 26200 37544 27000 37574
rect 22946 37503 23262 37504
rect 17769 37364 17835 37365
rect 17718 37300 17724 37364
rect 17788 37362 17835 37364
rect 17788 37360 17880 37362
rect 17830 37304 17880 37360
rect 17788 37302 17880 37304
rect 17788 37300 17835 37302
rect 17769 37299 17835 37300
rect 12065 37226 12131 37229
rect 19742 37226 19748 37228
rect 12065 37224 19748 37226
rect 12065 37168 12070 37224
rect 12126 37168 19748 37224
rect 12065 37166 19748 37168
rect 12065 37163 12131 37166
rect 19742 37164 19748 37166
rect 19812 37226 19818 37228
rect 23657 37226 23723 37229
rect 19812 37224 23723 37226
rect 19812 37168 23662 37224
rect 23718 37168 23723 37224
rect 19812 37166 23723 37168
rect 19812 37164 19818 37166
rect 23657 37163 23723 37166
rect 7946 37024 8262 37025
rect 7946 36960 7952 37024
rect 8016 36960 8032 37024
rect 8096 36960 8112 37024
rect 8176 36960 8192 37024
rect 8256 36960 8262 37024
rect 7946 36959 8262 36960
rect 17946 37024 18262 37025
rect 17946 36960 17952 37024
rect 18016 36960 18032 37024
rect 18096 36960 18112 37024
rect 18176 36960 18192 37024
rect 18256 36960 18262 37024
rect 17946 36959 18262 36960
rect 9857 36954 9923 36957
rect 17125 36954 17191 36957
rect 9857 36952 17191 36954
rect 9857 36896 9862 36952
rect 9918 36896 17130 36952
rect 17186 36896 17191 36952
rect 9857 36894 17191 36896
rect 9857 36891 9923 36894
rect 17125 36891 17191 36894
rect 24945 36954 25011 36957
rect 26200 36954 27000 36984
rect 24945 36952 27000 36954
rect 24945 36896 24950 36952
rect 25006 36896 27000 36952
rect 24945 36894 27000 36896
rect 24945 36891 25011 36894
rect 26200 36864 27000 36894
rect 14549 36818 14615 36821
rect 21541 36818 21607 36821
rect 23933 36818 23999 36821
rect 14549 36816 23999 36818
rect 14549 36760 14554 36816
rect 14610 36760 21546 36816
rect 21602 36760 23938 36816
rect 23994 36760 23999 36816
rect 14549 36758 23999 36760
rect 14549 36755 14615 36758
rect 21541 36755 21607 36758
rect 23933 36755 23999 36758
rect 12014 36620 12020 36684
rect 12084 36682 12090 36684
rect 19609 36682 19675 36685
rect 12084 36680 19675 36682
rect 12084 36624 19614 36680
rect 19670 36624 19675 36680
rect 12084 36622 19675 36624
rect 12084 36620 12090 36622
rect 19609 36619 19675 36622
rect 0 36546 800 36576
rect 1301 36546 1367 36549
rect 0 36544 1367 36546
rect 0 36488 1306 36544
rect 1362 36488 1367 36544
rect 0 36486 1367 36488
rect 0 36456 800 36486
rect 1301 36483 1367 36486
rect 2946 36480 3262 36481
rect 2946 36416 2952 36480
rect 3016 36416 3032 36480
rect 3096 36416 3112 36480
rect 3176 36416 3192 36480
rect 3256 36416 3262 36480
rect 2946 36415 3262 36416
rect 12946 36480 13262 36481
rect 12946 36416 12952 36480
rect 13016 36416 13032 36480
rect 13096 36416 13112 36480
rect 13176 36416 13192 36480
rect 13256 36416 13262 36480
rect 12946 36415 13262 36416
rect 22946 36480 23262 36481
rect 22946 36416 22952 36480
rect 23016 36416 23032 36480
rect 23096 36416 23112 36480
rect 23176 36416 23192 36480
rect 23256 36416 23262 36480
rect 22946 36415 23262 36416
rect 17585 36274 17651 36277
rect 21265 36274 21331 36277
rect 17585 36272 21331 36274
rect 17585 36216 17590 36272
rect 17646 36216 21270 36272
rect 21326 36216 21331 36272
rect 17585 36214 21331 36216
rect 17585 36211 17651 36214
rect 21265 36211 21331 36214
rect 25313 36274 25379 36277
rect 26200 36274 27000 36304
rect 25313 36272 27000 36274
rect 25313 36216 25318 36272
rect 25374 36216 27000 36272
rect 25313 36214 27000 36216
rect 25313 36211 25379 36214
rect 26200 36184 27000 36214
rect 7946 35936 8262 35937
rect 7946 35872 7952 35936
rect 8016 35872 8032 35936
rect 8096 35872 8112 35936
rect 8176 35872 8192 35936
rect 8256 35872 8262 35936
rect 7946 35871 8262 35872
rect 17946 35936 18262 35937
rect 17946 35872 17952 35936
rect 18016 35872 18032 35936
rect 18096 35872 18112 35936
rect 18176 35872 18192 35936
rect 18256 35872 18262 35936
rect 17946 35871 18262 35872
rect 8753 35866 8819 35869
rect 15377 35866 15443 35869
rect 8753 35864 15443 35866
rect 8753 35808 8758 35864
rect 8814 35808 15382 35864
rect 15438 35808 15443 35864
rect 8753 35806 15443 35808
rect 8753 35803 8819 35806
rect 15377 35803 15443 35806
rect 24761 35594 24827 35597
rect 26200 35594 27000 35624
rect 24761 35592 27000 35594
rect 24761 35536 24766 35592
rect 24822 35536 27000 35592
rect 24761 35534 27000 35536
rect 24761 35531 24827 35534
rect 26200 35504 27000 35534
rect 2946 35392 3262 35393
rect 2946 35328 2952 35392
rect 3016 35328 3032 35392
rect 3096 35328 3112 35392
rect 3176 35328 3192 35392
rect 3256 35328 3262 35392
rect 2946 35327 3262 35328
rect 12946 35392 13262 35393
rect 12946 35328 12952 35392
rect 13016 35328 13032 35392
rect 13096 35328 13112 35392
rect 13176 35328 13192 35392
rect 13256 35328 13262 35392
rect 12946 35327 13262 35328
rect 22946 35392 23262 35393
rect 22946 35328 22952 35392
rect 23016 35328 23032 35392
rect 23096 35328 23112 35392
rect 23176 35328 23192 35392
rect 23256 35328 23262 35392
rect 22946 35327 23262 35328
rect 13670 35260 13676 35324
rect 13740 35322 13746 35324
rect 13997 35322 14063 35325
rect 13740 35320 14063 35322
rect 13740 35264 14002 35320
rect 14058 35264 14063 35320
rect 13740 35262 14063 35264
rect 13740 35260 13746 35262
rect 12709 35186 12775 35189
rect 13678 35186 13738 35260
rect 13997 35259 14063 35262
rect 12709 35184 13738 35186
rect 12709 35128 12714 35184
rect 12770 35128 13738 35184
rect 12709 35126 13738 35128
rect 12709 35123 12775 35126
rect 22502 35124 22508 35188
rect 22572 35186 22578 35188
rect 22737 35186 22803 35189
rect 22572 35184 22803 35186
rect 22572 35128 22742 35184
rect 22798 35128 22803 35184
rect 22572 35126 22803 35128
rect 22572 35124 22578 35126
rect 22737 35123 22803 35126
rect 25313 34914 25379 34917
rect 26200 34914 27000 34944
rect 25313 34912 27000 34914
rect 25313 34856 25318 34912
rect 25374 34856 27000 34912
rect 25313 34854 27000 34856
rect 25313 34851 25379 34854
rect 7946 34848 8262 34849
rect 7946 34784 7952 34848
rect 8016 34784 8032 34848
rect 8096 34784 8112 34848
rect 8176 34784 8192 34848
rect 8256 34784 8262 34848
rect 7946 34783 8262 34784
rect 17946 34848 18262 34849
rect 17946 34784 17952 34848
rect 18016 34784 18032 34848
rect 18096 34784 18112 34848
rect 18176 34784 18192 34848
rect 18256 34784 18262 34848
rect 26200 34824 27000 34854
rect 17946 34783 18262 34784
rect 14457 34506 14523 34509
rect 15142 34506 15148 34508
rect 14457 34504 15148 34506
rect 14457 34448 14462 34504
rect 14518 34448 15148 34504
rect 14457 34446 15148 34448
rect 14457 34443 14523 34446
rect 15142 34444 15148 34446
rect 15212 34444 15218 34508
rect 2946 34304 3262 34305
rect 0 34234 800 34264
rect 2946 34240 2952 34304
rect 3016 34240 3032 34304
rect 3096 34240 3112 34304
rect 3176 34240 3192 34304
rect 3256 34240 3262 34304
rect 2946 34239 3262 34240
rect 12946 34304 13262 34305
rect 12946 34240 12952 34304
rect 13016 34240 13032 34304
rect 13096 34240 13112 34304
rect 13176 34240 13192 34304
rect 13256 34240 13262 34304
rect 12946 34239 13262 34240
rect 22946 34304 23262 34305
rect 22946 34240 22952 34304
rect 23016 34240 23032 34304
rect 23096 34240 23112 34304
rect 23176 34240 23192 34304
rect 23256 34240 23262 34304
rect 22946 34239 23262 34240
rect 1577 34234 1643 34237
rect 0 34232 1643 34234
rect 0 34176 1582 34232
rect 1638 34176 1643 34232
rect 0 34174 1643 34176
rect 0 34144 800 34174
rect 1577 34171 1643 34174
rect 25405 34234 25471 34237
rect 26200 34234 27000 34264
rect 25405 34232 27000 34234
rect 25405 34176 25410 34232
rect 25466 34176 27000 34232
rect 25405 34174 27000 34176
rect 25405 34171 25471 34174
rect 26200 34144 27000 34174
rect 7946 33760 8262 33761
rect 7946 33696 7952 33760
rect 8016 33696 8032 33760
rect 8096 33696 8112 33760
rect 8176 33696 8192 33760
rect 8256 33696 8262 33760
rect 7946 33695 8262 33696
rect 17946 33760 18262 33761
rect 17946 33696 17952 33760
rect 18016 33696 18032 33760
rect 18096 33696 18112 33760
rect 18176 33696 18192 33760
rect 18256 33696 18262 33760
rect 17946 33695 18262 33696
rect 12065 33692 12131 33693
rect 12014 33628 12020 33692
rect 12084 33690 12131 33692
rect 12084 33688 12176 33690
rect 12126 33632 12176 33688
rect 12084 33630 12176 33632
rect 12084 33628 12131 33630
rect 12065 33627 12131 33628
rect 13854 33492 13860 33556
rect 13924 33554 13930 33556
rect 18965 33554 19031 33557
rect 13924 33552 19031 33554
rect 13924 33496 18970 33552
rect 19026 33496 19031 33552
rect 13924 33494 19031 33496
rect 13924 33492 13930 33494
rect 18965 33491 19031 33494
rect 25313 33554 25379 33557
rect 26200 33554 27000 33584
rect 25313 33552 27000 33554
rect 25313 33496 25318 33552
rect 25374 33496 27000 33552
rect 25313 33494 27000 33496
rect 25313 33491 25379 33494
rect 26200 33464 27000 33494
rect 13997 33418 14063 33421
rect 17534 33418 17540 33420
rect 13997 33416 17540 33418
rect 13997 33360 14002 33416
rect 14058 33360 17540 33416
rect 13997 33358 17540 33360
rect 13997 33355 14063 33358
rect 17534 33356 17540 33358
rect 17604 33356 17610 33420
rect 2946 33216 3262 33217
rect 2946 33152 2952 33216
rect 3016 33152 3032 33216
rect 3096 33152 3112 33216
rect 3176 33152 3192 33216
rect 3256 33152 3262 33216
rect 2946 33151 3262 33152
rect 12946 33216 13262 33217
rect 12946 33152 12952 33216
rect 13016 33152 13032 33216
rect 13096 33152 13112 33216
rect 13176 33152 13192 33216
rect 13256 33152 13262 33216
rect 12946 33151 13262 33152
rect 22946 33216 23262 33217
rect 22946 33152 22952 33216
rect 23016 33152 23032 33216
rect 23096 33152 23112 33216
rect 23176 33152 23192 33216
rect 23256 33152 23262 33216
rect 22946 33151 23262 33152
rect 25313 32874 25379 32877
rect 26200 32874 27000 32904
rect 25313 32872 27000 32874
rect 25313 32816 25318 32872
rect 25374 32816 27000 32872
rect 25313 32814 27000 32816
rect 25313 32811 25379 32814
rect 26200 32784 27000 32814
rect 7946 32672 8262 32673
rect 7946 32608 7952 32672
rect 8016 32608 8032 32672
rect 8096 32608 8112 32672
rect 8176 32608 8192 32672
rect 8256 32608 8262 32672
rect 7946 32607 8262 32608
rect 17946 32672 18262 32673
rect 17946 32608 17952 32672
rect 18016 32608 18032 32672
rect 18096 32608 18112 32672
rect 18176 32608 18192 32672
rect 18256 32608 18262 32672
rect 17946 32607 18262 32608
rect 25313 32194 25379 32197
rect 26200 32194 27000 32224
rect 25313 32192 27000 32194
rect 25313 32136 25318 32192
rect 25374 32136 27000 32192
rect 25313 32134 27000 32136
rect 25313 32131 25379 32134
rect 2946 32128 3262 32129
rect 2946 32064 2952 32128
rect 3016 32064 3032 32128
rect 3096 32064 3112 32128
rect 3176 32064 3192 32128
rect 3256 32064 3262 32128
rect 2946 32063 3262 32064
rect 12946 32128 13262 32129
rect 12946 32064 12952 32128
rect 13016 32064 13032 32128
rect 13096 32064 13112 32128
rect 13176 32064 13192 32128
rect 13256 32064 13262 32128
rect 12946 32063 13262 32064
rect 22946 32128 23262 32129
rect 22946 32064 22952 32128
rect 23016 32064 23032 32128
rect 23096 32064 23112 32128
rect 23176 32064 23192 32128
rect 23256 32064 23262 32128
rect 26200 32104 27000 32134
rect 22946 32063 23262 32064
rect 0 31922 800 31952
rect 1301 31922 1367 31925
rect 0 31920 1367 31922
rect 0 31864 1306 31920
rect 1362 31864 1367 31920
rect 0 31862 1367 31864
rect 0 31832 800 31862
rect 1301 31859 1367 31862
rect 14406 31860 14412 31924
rect 14476 31922 14482 31924
rect 17033 31922 17099 31925
rect 14476 31920 17099 31922
rect 14476 31864 17038 31920
rect 17094 31864 17099 31920
rect 14476 31862 17099 31864
rect 14476 31860 14482 31862
rect 17033 31859 17099 31862
rect 7189 31786 7255 31789
rect 7373 31786 7439 31789
rect 7189 31784 7439 31786
rect 7189 31728 7194 31784
rect 7250 31728 7378 31784
rect 7434 31728 7439 31784
rect 7189 31726 7439 31728
rect 7189 31723 7255 31726
rect 7373 31723 7439 31726
rect 10225 31786 10291 31789
rect 10869 31786 10935 31789
rect 10225 31784 10935 31786
rect 10225 31728 10230 31784
rect 10286 31728 10874 31784
rect 10930 31728 10935 31784
rect 10225 31726 10935 31728
rect 10225 31723 10291 31726
rect 10869 31723 10935 31726
rect 21633 31786 21699 31789
rect 22318 31786 22324 31788
rect 21633 31784 22324 31786
rect 21633 31728 21638 31784
rect 21694 31728 22324 31784
rect 21633 31726 22324 31728
rect 21633 31723 21699 31726
rect 22318 31724 22324 31726
rect 22388 31724 22394 31788
rect 7946 31584 8262 31585
rect 7946 31520 7952 31584
rect 8016 31520 8032 31584
rect 8096 31520 8112 31584
rect 8176 31520 8192 31584
rect 8256 31520 8262 31584
rect 7946 31519 8262 31520
rect 17946 31584 18262 31585
rect 17946 31520 17952 31584
rect 18016 31520 18032 31584
rect 18096 31520 18112 31584
rect 18176 31520 18192 31584
rect 18256 31520 18262 31584
rect 17946 31519 18262 31520
rect 25313 31514 25379 31517
rect 26200 31514 27000 31544
rect 25313 31512 27000 31514
rect 25313 31456 25318 31512
rect 25374 31456 27000 31512
rect 25313 31454 27000 31456
rect 25313 31451 25379 31454
rect 26200 31424 27000 31454
rect 9857 31380 9923 31381
rect 9806 31378 9812 31380
rect 9766 31318 9812 31378
rect 9876 31376 9923 31380
rect 9918 31320 9923 31376
rect 9806 31316 9812 31318
rect 9876 31316 9923 31320
rect 9857 31315 9923 31316
rect 2946 31040 3262 31041
rect 2946 30976 2952 31040
rect 3016 30976 3032 31040
rect 3096 30976 3112 31040
rect 3176 30976 3192 31040
rect 3256 30976 3262 31040
rect 2946 30975 3262 30976
rect 12946 31040 13262 31041
rect 12946 30976 12952 31040
rect 13016 30976 13032 31040
rect 13096 30976 13112 31040
rect 13176 30976 13192 31040
rect 13256 30976 13262 31040
rect 12946 30975 13262 30976
rect 22946 31040 23262 31041
rect 22946 30976 22952 31040
rect 23016 30976 23032 31040
rect 23096 30976 23112 31040
rect 23176 30976 23192 31040
rect 23256 30976 23262 31040
rect 22946 30975 23262 30976
rect 18137 30834 18203 30837
rect 18454 30834 18460 30836
rect 18137 30832 18460 30834
rect 18137 30776 18142 30832
rect 18198 30776 18460 30832
rect 18137 30774 18460 30776
rect 18137 30771 18203 30774
rect 18454 30772 18460 30774
rect 18524 30772 18530 30836
rect 25405 30834 25471 30837
rect 26200 30834 27000 30864
rect 25405 30832 27000 30834
rect 25405 30776 25410 30832
rect 25466 30776 27000 30832
rect 25405 30774 27000 30776
rect 25405 30771 25471 30774
rect 26200 30744 27000 30774
rect 10593 30698 10659 30701
rect 13854 30698 13860 30700
rect 10593 30696 13860 30698
rect 10593 30640 10598 30696
rect 10654 30640 13860 30696
rect 10593 30638 13860 30640
rect 10593 30635 10659 30638
rect 13854 30636 13860 30638
rect 13924 30636 13930 30700
rect 18965 30698 19031 30701
rect 20478 30698 20484 30700
rect 18965 30696 20484 30698
rect 18965 30640 18970 30696
rect 19026 30640 20484 30696
rect 18965 30638 20484 30640
rect 18965 30635 19031 30638
rect 20478 30636 20484 30638
rect 20548 30636 20554 30700
rect 7946 30496 8262 30497
rect 7946 30432 7952 30496
rect 8016 30432 8032 30496
rect 8096 30432 8112 30496
rect 8176 30432 8192 30496
rect 8256 30432 8262 30496
rect 7946 30431 8262 30432
rect 17946 30496 18262 30497
rect 17946 30432 17952 30496
rect 18016 30432 18032 30496
rect 18096 30432 18112 30496
rect 18176 30432 18192 30496
rect 18256 30432 18262 30496
rect 17946 30431 18262 30432
rect 12985 30426 13051 30429
rect 17718 30426 17724 30428
rect 12985 30424 17724 30426
rect 12985 30368 12990 30424
rect 13046 30368 17724 30424
rect 12985 30366 17724 30368
rect 12985 30363 13051 30366
rect 17718 30364 17724 30366
rect 17788 30364 17794 30428
rect 14590 30228 14596 30292
rect 14660 30290 14666 30292
rect 19425 30290 19491 30293
rect 14660 30288 19491 30290
rect 14660 30232 19430 30288
rect 19486 30232 19491 30288
rect 14660 30230 19491 30232
rect 14660 30228 14666 30230
rect 19425 30227 19491 30230
rect 19558 30092 19564 30156
rect 19628 30154 19634 30156
rect 19977 30154 20043 30157
rect 19628 30152 20043 30154
rect 19628 30096 19982 30152
rect 20038 30096 20043 30152
rect 19628 30094 20043 30096
rect 19628 30092 19634 30094
rect 19977 30091 20043 30094
rect 25313 30154 25379 30157
rect 26200 30154 27000 30184
rect 25313 30152 27000 30154
rect 25313 30096 25318 30152
rect 25374 30096 27000 30152
rect 25313 30094 27000 30096
rect 25313 30091 25379 30094
rect 26200 30064 27000 30094
rect 16113 30018 16179 30021
rect 16246 30018 16252 30020
rect 16113 30016 16252 30018
rect 16113 29960 16118 30016
rect 16174 29960 16252 30016
rect 16113 29958 16252 29960
rect 16113 29955 16179 29958
rect 16246 29956 16252 29958
rect 16316 29956 16322 30020
rect 2946 29952 3262 29953
rect 2946 29888 2952 29952
rect 3016 29888 3032 29952
rect 3096 29888 3112 29952
rect 3176 29888 3192 29952
rect 3256 29888 3262 29952
rect 2946 29887 3262 29888
rect 12946 29952 13262 29953
rect 12946 29888 12952 29952
rect 13016 29888 13032 29952
rect 13096 29888 13112 29952
rect 13176 29888 13192 29952
rect 13256 29888 13262 29952
rect 12946 29887 13262 29888
rect 22946 29952 23262 29953
rect 22946 29888 22952 29952
rect 23016 29888 23032 29952
rect 23096 29888 23112 29952
rect 23176 29888 23192 29952
rect 23256 29888 23262 29952
rect 22946 29887 23262 29888
rect 17718 29684 17724 29748
rect 17788 29746 17794 29748
rect 18229 29746 18295 29749
rect 19374 29746 19380 29748
rect 17788 29744 19380 29746
rect 17788 29688 18234 29744
rect 18290 29688 19380 29744
rect 17788 29686 19380 29688
rect 17788 29684 17794 29686
rect 18229 29683 18295 29686
rect 19374 29684 19380 29686
rect 19444 29684 19450 29748
rect 19742 29684 19748 29748
rect 19812 29746 19818 29748
rect 19885 29746 19951 29749
rect 19812 29744 19951 29746
rect 19812 29688 19890 29744
rect 19946 29688 19951 29744
rect 19812 29686 19951 29688
rect 19812 29684 19818 29686
rect 19885 29683 19951 29686
rect 22277 29746 22343 29749
rect 22502 29746 22508 29748
rect 22277 29744 22508 29746
rect 22277 29688 22282 29744
rect 22338 29688 22508 29744
rect 22277 29686 22508 29688
rect 22277 29683 22343 29686
rect 22502 29684 22508 29686
rect 22572 29684 22578 29748
rect 0 29610 800 29640
rect 1301 29610 1367 29613
rect 0 29608 1367 29610
rect 0 29552 1306 29608
rect 1362 29552 1367 29608
rect 0 29550 1367 29552
rect 0 29520 800 29550
rect 1301 29547 1367 29550
rect 12341 29474 12407 29477
rect 12750 29474 12756 29476
rect 12341 29472 12756 29474
rect 12341 29416 12346 29472
rect 12402 29416 12756 29472
rect 12341 29414 12756 29416
rect 12341 29411 12407 29414
rect 12750 29412 12756 29414
rect 12820 29412 12826 29476
rect 21725 29474 21791 29477
rect 23422 29474 23428 29476
rect 21725 29472 23428 29474
rect 21725 29416 21730 29472
rect 21786 29416 23428 29472
rect 21725 29414 23428 29416
rect 21725 29411 21791 29414
rect 23422 29412 23428 29414
rect 23492 29412 23498 29476
rect 25405 29474 25471 29477
rect 26200 29474 27000 29504
rect 25405 29472 27000 29474
rect 25405 29416 25410 29472
rect 25466 29416 27000 29472
rect 25405 29414 27000 29416
rect 25405 29411 25471 29414
rect 7946 29408 8262 29409
rect 7946 29344 7952 29408
rect 8016 29344 8032 29408
rect 8096 29344 8112 29408
rect 8176 29344 8192 29408
rect 8256 29344 8262 29408
rect 7946 29343 8262 29344
rect 17946 29408 18262 29409
rect 17946 29344 17952 29408
rect 18016 29344 18032 29408
rect 18096 29344 18112 29408
rect 18176 29344 18192 29408
rect 18256 29344 18262 29408
rect 26200 29384 27000 29414
rect 17946 29343 18262 29344
rect 14590 29004 14596 29068
rect 14660 29066 14666 29068
rect 14733 29066 14799 29069
rect 16757 29068 16823 29069
rect 17493 29068 17559 29069
rect 16757 29066 16804 29068
rect 14660 29064 14799 29066
rect 14660 29008 14738 29064
rect 14794 29008 14799 29064
rect 14660 29006 14799 29008
rect 16712 29064 16804 29066
rect 16712 29008 16762 29064
rect 16712 29006 16804 29008
rect 14660 29004 14666 29006
rect 14733 29003 14799 29006
rect 16757 29004 16804 29006
rect 16868 29004 16874 29068
rect 17493 29066 17540 29068
rect 17448 29064 17540 29066
rect 17448 29008 17498 29064
rect 17448 29006 17540 29008
rect 17493 29004 17540 29006
rect 17604 29004 17610 29068
rect 16757 29003 16823 29004
rect 17493 29003 17559 29004
rect 2946 28864 3262 28865
rect 2946 28800 2952 28864
rect 3016 28800 3032 28864
rect 3096 28800 3112 28864
rect 3176 28800 3192 28864
rect 3256 28800 3262 28864
rect 2946 28799 3262 28800
rect 12946 28864 13262 28865
rect 12946 28800 12952 28864
rect 13016 28800 13032 28864
rect 13096 28800 13112 28864
rect 13176 28800 13192 28864
rect 13256 28800 13262 28864
rect 12946 28799 13262 28800
rect 22946 28864 23262 28865
rect 22946 28800 22952 28864
rect 23016 28800 23032 28864
rect 23096 28800 23112 28864
rect 23176 28800 23192 28864
rect 23256 28800 23262 28864
rect 22946 28799 23262 28800
rect 24117 28794 24183 28797
rect 26200 28794 27000 28824
rect 24117 28792 27000 28794
rect 24117 28736 24122 28792
rect 24178 28736 27000 28792
rect 24117 28734 27000 28736
rect 24117 28731 24183 28734
rect 26200 28704 27000 28734
rect 20897 28388 20963 28389
rect 20846 28324 20852 28388
rect 20916 28386 20963 28388
rect 20916 28384 21008 28386
rect 20958 28328 21008 28384
rect 20916 28326 21008 28328
rect 20916 28324 20963 28326
rect 20897 28323 20963 28324
rect 7946 28320 8262 28321
rect 7946 28256 7952 28320
rect 8016 28256 8032 28320
rect 8096 28256 8112 28320
rect 8176 28256 8192 28320
rect 8256 28256 8262 28320
rect 7946 28255 8262 28256
rect 17946 28320 18262 28321
rect 17946 28256 17952 28320
rect 18016 28256 18032 28320
rect 18096 28256 18112 28320
rect 18176 28256 18192 28320
rect 18256 28256 18262 28320
rect 17946 28255 18262 28256
rect 16246 28052 16252 28116
rect 16316 28114 16322 28116
rect 20437 28114 20503 28117
rect 16316 28112 20503 28114
rect 16316 28056 20442 28112
rect 20498 28056 20503 28112
rect 16316 28054 20503 28056
rect 16316 28052 16322 28054
rect 20437 28051 20503 28054
rect 24853 28114 24919 28117
rect 26200 28114 27000 28144
rect 24853 28112 27000 28114
rect 24853 28056 24858 28112
rect 24914 28056 27000 28112
rect 24853 28054 27000 28056
rect 24853 28051 24919 28054
rect 26200 28024 27000 28054
rect 2946 27776 3262 27777
rect 2946 27712 2952 27776
rect 3016 27712 3032 27776
rect 3096 27712 3112 27776
rect 3176 27712 3192 27776
rect 3256 27712 3262 27776
rect 2946 27711 3262 27712
rect 12946 27776 13262 27777
rect 12946 27712 12952 27776
rect 13016 27712 13032 27776
rect 13096 27712 13112 27776
rect 13176 27712 13192 27776
rect 13256 27712 13262 27776
rect 12946 27711 13262 27712
rect 22946 27776 23262 27777
rect 22946 27712 22952 27776
rect 23016 27712 23032 27776
rect 23096 27712 23112 27776
rect 23176 27712 23192 27776
rect 23256 27712 23262 27776
rect 22946 27711 23262 27712
rect 18454 27508 18460 27572
rect 18524 27570 18530 27572
rect 19241 27570 19307 27573
rect 21214 27570 21220 27572
rect 18524 27568 21220 27570
rect 18524 27512 19246 27568
rect 19302 27512 21220 27568
rect 18524 27510 21220 27512
rect 18524 27508 18530 27510
rect 19241 27507 19307 27510
rect 21214 27508 21220 27510
rect 21284 27508 21290 27572
rect 25405 27434 25471 27437
rect 26200 27434 27000 27464
rect 25405 27432 27000 27434
rect 25405 27376 25410 27432
rect 25466 27376 27000 27432
rect 25405 27374 27000 27376
rect 25405 27371 25471 27374
rect 26200 27344 27000 27374
rect 0 27298 800 27328
rect 1301 27298 1367 27301
rect 0 27296 1367 27298
rect 0 27240 1306 27296
rect 1362 27240 1367 27296
rect 0 27238 1367 27240
rect 0 27208 800 27238
rect 1301 27235 1367 27238
rect 7946 27232 8262 27233
rect 7946 27168 7952 27232
rect 8016 27168 8032 27232
rect 8096 27168 8112 27232
rect 8176 27168 8192 27232
rect 8256 27168 8262 27232
rect 7946 27167 8262 27168
rect 17946 27232 18262 27233
rect 17946 27168 17952 27232
rect 18016 27168 18032 27232
rect 18096 27168 18112 27232
rect 18176 27168 18192 27232
rect 18256 27168 18262 27232
rect 17946 27167 18262 27168
rect 15745 27164 15811 27165
rect 15694 27100 15700 27164
rect 15764 27162 15811 27164
rect 19241 27162 19307 27165
rect 21398 27162 21404 27164
rect 15764 27160 15856 27162
rect 15806 27104 15856 27160
rect 15764 27102 15856 27104
rect 19241 27160 21404 27162
rect 19241 27104 19246 27160
rect 19302 27104 21404 27160
rect 19241 27102 21404 27104
rect 15764 27100 15811 27102
rect 15745 27099 15811 27100
rect 19241 27099 19307 27102
rect 21398 27100 21404 27102
rect 21468 27100 21474 27164
rect 24669 26754 24735 26757
rect 26200 26754 27000 26784
rect 24669 26752 27000 26754
rect 24669 26696 24674 26752
rect 24730 26696 27000 26752
rect 24669 26694 27000 26696
rect 24669 26691 24735 26694
rect 2946 26688 3262 26689
rect 2946 26624 2952 26688
rect 3016 26624 3032 26688
rect 3096 26624 3112 26688
rect 3176 26624 3192 26688
rect 3256 26624 3262 26688
rect 2946 26623 3262 26624
rect 12946 26688 13262 26689
rect 12946 26624 12952 26688
rect 13016 26624 13032 26688
rect 13096 26624 13112 26688
rect 13176 26624 13192 26688
rect 13256 26624 13262 26688
rect 12946 26623 13262 26624
rect 22946 26688 23262 26689
rect 22946 26624 22952 26688
rect 23016 26624 23032 26688
rect 23096 26624 23112 26688
rect 23176 26624 23192 26688
rect 23256 26624 23262 26688
rect 26200 26664 27000 26694
rect 22946 26623 23262 26624
rect 23422 26148 23428 26212
rect 23492 26210 23498 26212
rect 23565 26210 23631 26213
rect 23492 26208 23631 26210
rect 23492 26152 23570 26208
rect 23626 26152 23631 26208
rect 23492 26150 23631 26152
rect 23492 26148 23498 26150
rect 23565 26147 23631 26150
rect 7946 26144 8262 26145
rect 7946 26080 7952 26144
rect 8016 26080 8032 26144
rect 8096 26080 8112 26144
rect 8176 26080 8192 26144
rect 8256 26080 8262 26144
rect 7946 26079 8262 26080
rect 17946 26144 18262 26145
rect 17946 26080 17952 26144
rect 18016 26080 18032 26144
rect 18096 26080 18112 26144
rect 18176 26080 18192 26144
rect 18256 26080 18262 26144
rect 17946 26079 18262 26080
rect 22277 26074 22343 26077
rect 26200 26074 27000 26104
rect 22277 26072 27000 26074
rect 22277 26016 22282 26072
rect 22338 26016 27000 26072
rect 22277 26014 27000 26016
rect 22277 26011 22343 26014
rect 26200 25984 27000 26014
rect 16113 25668 16179 25669
rect 16062 25604 16068 25668
rect 16132 25666 16179 25668
rect 16132 25664 16224 25666
rect 16174 25608 16224 25664
rect 16132 25606 16224 25608
rect 16132 25604 16179 25606
rect 16113 25603 16179 25604
rect 2946 25600 3262 25601
rect 2946 25536 2952 25600
rect 3016 25536 3032 25600
rect 3096 25536 3112 25600
rect 3176 25536 3192 25600
rect 3256 25536 3262 25600
rect 2946 25535 3262 25536
rect 12946 25600 13262 25601
rect 12946 25536 12952 25600
rect 13016 25536 13032 25600
rect 13096 25536 13112 25600
rect 13176 25536 13192 25600
rect 13256 25536 13262 25600
rect 12946 25535 13262 25536
rect 22946 25600 23262 25601
rect 22946 25536 22952 25600
rect 23016 25536 23032 25600
rect 23096 25536 23112 25600
rect 23176 25536 23192 25600
rect 23256 25536 23262 25600
rect 22946 25535 23262 25536
rect 25313 25394 25379 25397
rect 26200 25394 27000 25424
rect 25313 25392 27000 25394
rect 25313 25336 25318 25392
rect 25374 25336 27000 25392
rect 25313 25334 27000 25336
rect 25313 25331 25379 25334
rect 26200 25304 27000 25334
rect 7946 25056 8262 25057
rect 0 24986 800 25016
rect 7946 24992 7952 25056
rect 8016 24992 8032 25056
rect 8096 24992 8112 25056
rect 8176 24992 8192 25056
rect 8256 24992 8262 25056
rect 7946 24991 8262 24992
rect 17946 25056 18262 25057
rect 17946 24992 17952 25056
rect 18016 24992 18032 25056
rect 18096 24992 18112 25056
rect 18176 24992 18192 25056
rect 18256 24992 18262 25056
rect 17946 24991 18262 24992
rect 1301 24986 1367 24989
rect 0 24984 1367 24986
rect 0 24928 1306 24984
rect 1362 24928 1367 24984
rect 0 24926 1367 24928
rect 0 24896 800 24926
rect 1301 24923 1367 24926
rect 25129 24714 25195 24717
rect 26200 24714 27000 24744
rect 25129 24712 27000 24714
rect 25129 24656 25134 24712
rect 25190 24656 27000 24712
rect 25129 24654 27000 24656
rect 25129 24651 25195 24654
rect 26200 24624 27000 24654
rect 19333 24578 19399 24581
rect 20846 24578 20852 24580
rect 19333 24576 20852 24578
rect 19333 24520 19338 24576
rect 19394 24520 20852 24576
rect 19333 24518 20852 24520
rect 19333 24515 19399 24518
rect 20846 24516 20852 24518
rect 20916 24516 20922 24580
rect 2946 24512 3262 24513
rect 2946 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3262 24512
rect 2946 24447 3262 24448
rect 12946 24512 13262 24513
rect 12946 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13262 24512
rect 12946 24447 13262 24448
rect 22946 24512 23262 24513
rect 22946 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23262 24512
rect 22946 24447 23262 24448
rect 11605 24170 11671 24173
rect 12566 24170 12572 24172
rect 11605 24168 12572 24170
rect 11605 24112 11610 24168
rect 11666 24112 12572 24168
rect 11605 24110 12572 24112
rect 11605 24107 11671 24110
rect 12566 24108 12572 24110
rect 12636 24108 12642 24172
rect 24853 24034 24919 24037
rect 26200 24034 27000 24064
rect 24853 24032 27000 24034
rect 24853 23976 24858 24032
rect 24914 23976 27000 24032
rect 24853 23974 27000 23976
rect 24853 23971 24919 23974
rect 7946 23968 8262 23969
rect 7946 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8262 23968
rect 7946 23903 8262 23904
rect 17946 23968 18262 23969
rect 17946 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18262 23968
rect 26200 23944 27000 23974
rect 17946 23903 18262 23904
rect 13486 23428 13492 23492
rect 13556 23490 13562 23492
rect 14406 23490 14412 23492
rect 13556 23430 14412 23490
rect 13556 23428 13562 23430
rect 14406 23428 14412 23430
rect 14476 23428 14482 23492
rect 2946 23424 3262 23425
rect 2946 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3262 23424
rect 2946 23359 3262 23360
rect 12946 23424 13262 23425
rect 12946 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13262 23424
rect 12946 23359 13262 23360
rect 22946 23424 23262 23425
rect 22946 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23262 23424
rect 22946 23359 23262 23360
rect 13721 23354 13787 23357
rect 17718 23354 17724 23356
rect 13721 23352 17724 23354
rect 13721 23296 13726 23352
rect 13782 23296 17724 23352
rect 13721 23294 17724 23296
rect 13721 23291 13787 23294
rect 17718 23292 17724 23294
rect 17788 23292 17794 23356
rect 23381 23354 23447 23357
rect 26200 23354 27000 23384
rect 23381 23352 27000 23354
rect 23381 23296 23386 23352
rect 23442 23296 27000 23352
rect 23381 23294 27000 23296
rect 23381 23291 23447 23294
rect 26200 23264 27000 23294
rect 7946 22880 8262 22881
rect 7946 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8262 22880
rect 7946 22815 8262 22816
rect 17946 22880 18262 22881
rect 17946 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18262 22880
rect 17946 22815 18262 22816
rect 0 22674 800 22704
rect 933 22674 999 22677
rect 0 22672 999 22674
rect 0 22616 938 22672
rect 994 22616 999 22672
rect 0 22614 999 22616
rect 0 22584 800 22614
rect 933 22611 999 22614
rect 10174 22612 10180 22676
rect 10244 22674 10250 22676
rect 12525 22674 12591 22677
rect 12750 22674 12756 22676
rect 10244 22672 12756 22674
rect 10244 22616 12530 22672
rect 12586 22616 12756 22672
rect 10244 22614 12756 22616
rect 10244 22612 10250 22614
rect 12525 22611 12591 22614
rect 12750 22612 12756 22614
rect 12820 22612 12826 22676
rect 24853 22674 24919 22677
rect 26200 22674 27000 22704
rect 24853 22672 27000 22674
rect 24853 22616 24858 22672
rect 24914 22616 27000 22672
rect 24853 22614 27000 22616
rect 24853 22611 24919 22614
rect 26200 22584 27000 22614
rect 13169 22538 13235 22541
rect 13486 22538 13492 22540
rect 13169 22536 13492 22538
rect 13169 22480 13174 22536
rect 13230 22480 13492 22536
rect 13169 22478 13492 22480
rect 13169 22475 13235 22478
rect 13486 22476 13492 22478
rect 13556 22476 13562 22540
rect 2946 22336 3262 22337
rect 2946 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3262 22336
rect 2946 22271 3262 22272
rect 12946 22336 13262 22337
rect 12946 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13262 22336
rect 12946 22271 13262 22272
rect 22946 22336 23262 22337
rect 22946 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23262 22336
rect 22946 22271 23262 22272
rect 17718 22204 17724 22268
rect 17788 22266 17794 22268
rect 19057 22266 19123 22269
rect 17788 22264 19123 22266
rect 17788 22208 19062 22264
rect 19118 22208 19123 22264
rect 17788 22206 19123 22208
rect 17788 22204 17794 22206
rect 19057 22203 19123 22206
rect 24853 21994 24919 21997
rect 26200 21994 27000 22024
rect 24853 21992 27000 21994
rect 24853 21936 24858 21992
rect 24914 21936 27000 21992
rect 24853 21934 27000 21936
rect 24853 21931 24919 21934
rect 26200 21904 27000 21934
rect 13813 21860 13879 21861
rect 13813 21858 13860 21860
rect 13768 21856 13860 21858
rect 13924 21858 13930 21860
rect 14733 21858 14799 21861
rect 13924 21856 14799 21858
rect 13768 21800 13818 21856
rect 13924 21800 14738 21856
rect 14794 21800 14799 21856
rect 13768 21798 13860 21800
rect 13813 21796 13860 21798
rect 13924 21798 14799 21800
rect 13924 21796 13930 21798
rect 13813 21795 13879 21796
rect 14733 21795 14799 21798
rect 7946 21792 8262 21793
rect 7946 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8262 21792
rect 7946 21727 8262 21728
rect 17946 21792 18262 21793
rect 17946 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18262 21792
rect 17946 21727 18262 21728
rect 11053 21722 11119 21725
rect 15561 21722 15627 21725
rect 11053 21720 15627 21722
rect 11053 21664 11058 21720
rect 11114 21664 15566 21720
rect 15622 21664 15627 21720
rect 11053 21662 15627 21664
rect 11053 21659 11119 21662
rect 15561 21659 15627 21662
rect 11697 21586 11763 21589
rect 15469 21586 15535 21589
rect 11697 21584 15535 21586
rect 11697 21528 11702 21584
rect 11758 21528 15474 21584
rect 15530 21528 15535 21584
rect 11697 21526 15535 21528
rect 11697 21523 11763 21526
rect 15469 21523 15535 21526
rect 12893 21450 12959 21453
rect 14549 21450 14615 21453
rect 12893 21448 14615 21450
rect 12893 21392 12898 21448
rect 12954 21392 14554 21448
rect 14610 21392 14615 21448
rect 12893 21390 14615 21392
rect 12893 21387 12959 21390
rect 14549 21387 14615 21390
rect 24485 21314 24551 21317
rect 26200 21314 27000 21344
rect 24485 21312 27000 21314
rect 24485 21256 24490 21312
rect 24546 21256 27000 21312
rect 24485 21254 27000 21256
rect 24485 21251 24551 21254
rect 2946 21248 3262 21249
rect 2946 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3262 21248
rect 2946 21183 3262 21184
rect 12946 21248 13262 21249
rect 12946 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13262 21248
rect 12946 21183 13262 21184
rect 22946 21248 23262 21249
rect 22946 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23262 21248
rect 26200 21224 27000 21254
rect 22946 21183 23262 21184
rect 11697 21042 11763 21045
rect 13445 21042 13511 21045
rect 11697 21040 13511 21042
rect 11697 20984 11702 21040
rect 11758 20984 13450 21040
rect 13506 20984 13511 21040
rect 11697 20982 13511 20984
rect 11697 20979 11763 20982
rect 13445 20979 13511 20982
rect 7946 20704 8262 20705
rect 7946 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8262 20704
rect 7946 20639 8262 20640
rect 17946 20704 18262 20705
rect 17946 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18262 20704
rect 17946 20639 18262 20640
rect 16062 20572 16068 20636
rect 16132 20634 16138 20636
rect 16389 20634 16455 20637
rect 16132 20632 16455 20634
rect 16132 20576 16394 20632
rect 16450 20576 16455 20632
rect 16132 20574 16455 20576
rect 16132 20572 16138 20574
rect 16389 20571 16455 20574
rect 25129 20634 25195 20637
rect 26200 20634 27000 20664
rect 25129 20632 27000 20634
rect 25129 20576 25134 20632
rect 25190 20576 27000 20632
rect 25129 20574 27000 20576
rect 25129 20571 25195 20574
rect 26200 20544 27000 20574
rect 0 20362 800 20392
rect 1301 20362 1367 20365
rect 0 20360 1367 20362
rect 0 20304 1306 20360
rect 1362 20304 1367 20360
rect 0 20302 1367 20304
rect 0 20272 800 20302
rect 1301 20299 1367 20302
rect 14641 20226 14707 20229
rect 14958 20226 14964 20228
rect 14641 20224 14964 20226
rect 14641 20168 14646 20224
rect 14702 20168 14964 20224
rect 14641 20166 14964 20168
rect 14641 20163 14707 20166
rect 14958 20164 14964 20166
rect 15028 20164 15034 20228
rect 2946 20160 3262 20161
rect 2946 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3262 20160
rect 2946 20095 3262 20096
rect 12946 20160 13262 20161
rect 12946 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13262 20160
rect 12946 20095 13262 20096
rect 22946 20160 23262 20161
rect 22946 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23262 20160
rect 22946 20095 23262 20096
rect 17217 19954 17283 19957
rect 18638 19954 18644 19956
rect 17217 19952 18644 19954
rect 17217 19896 17222 19952
rect 17278 19896 18644 19952
rect 17217 19894 18644 19896
rect 17217 19891 17283 19894
rect 18638 19892 18644 19894
rect 18708 19892 18714 19956
rect 24853 19954 24919 19957
rect 26200 19954 27000 19984
rect 24853 19952 27000 19954
rect 24853 19896 24858 19952
rect 24914 19896 27000 19952
rect 24853 19894 27000 19896
rect 24853 19891 24919 19894
rect 26200 19864 27000 19894
rect 7946 19616 8262 19617
rect 7946 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8262 19616
rect 7946 19551 8262 19552
rect 17946 19616 18262 19617
rect 17946 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18262 19616
rect 17946 19551 18262 19552
rect 22093 19274 22159 19277
rect 26200 19274 27000 19304
rect 22093 19272 27000 19274
rect 22093 19216 22098 19272
rect 22154 19216 27000 19272
rect 22093 19214 27000 19216
rect 22093 19211 22159 19214
rect 26200 19184 27000 19214
rect 2946 19072 3262 19073
rect 2946 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3262 19072
rect 2946 19007 3262 19008
rect 12946 19072 13262 19073
rect 12946 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13262 19072
rect 12946 19007 13262 19008
rect 22946 19072 23262 19073
rect 22946 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23262 19072
rect 22946 19007 23262 19008
rect 17585 18868 17651 18869
rect 17534 18804 17540 18868
rect 17604 18866 17651 18868
rect 17604 18864 17696 18866
rect 17646 18808 17696 18864
rect 17604 18806 17696 18808
rect 17604 18804 17651 18806
rect 17585 18803 17651 18804
rect 23381 18594 23447 18597
rect 26200 18594 27000 18624
rect 23381 18592 27000 18594
rect 23381 18536 23386 18592
rect 23442 18536 27000 18592
rect 23381 18534 27000 18536
rect 23381 18531 23447 18534
rect 7946 18528 8262 18529
rect 7946 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8262 18528
rect 7946 18463 8262 18464
rect 17946 18528 18262 18529
rect 17946 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18262 18528
rect 26200 18504 27000 18534
rect 17946 18463 18262 18464
rect 18505 18324 18571 18325
rect 18454 18322 18460 18324
rect 18414 18262 18460 18322
rect 18524 18320 18571 18324
rect 18566 18264 18571 18320
rect 18454 18260 18460 18262
rect 18524 18260 18571 18264
rect 18505 18259 18571 18260
rect 0 18050 800 18080
rect 1301 18050 1367 18053
rect 0 18048 1367 18050
rect 0 17992 1306 18048
rect 1362 17992 1367 18048
rect 0 17990 1367 17992
rect 0 17960 800 17990
rect 1301 17987 1367 17990
rect 2946 17984 3262 17985
rect 2946 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3262 17984
rect 2946 17919 3262 17920
rect 12946 17984 13262 17985
rect 12946 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13262 17984
rect 12946 17919 13262 17920
rect 22946 17984 23262 17985
rect 22946 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23262 17984
rect 22946 17919 23262 17920
rect 12566 17852 12572 17916
rect 12636 17914 12642 17916
rect 12801 17914 12867 17917
rect 12636 17912 12867 17914
rect 12636 17856 12806 17912
rect 12862 17856 12867 17912
rect 12636 17854 12867 17856
rect 12636 17852 12642 17854
rect 12801 17851 12867 17854
rect 24761 17914 24827 17917
rect 26200 17914 27000 17944
rect 24761 17912 27000 17914
rect 24761 17856 24766 17912
rect 24822 17856 27000 17912
rect 24761 17854 27000 17856
rect 24761 17851 24827 17854
rect 26200 17824 27000 17854
rect 16205 17644 16271 17645
rect 16205 17642 16252 17644
rect 16160 17640 16252 17642
rect 16160 17584 16210 17640
rect 16160 17582 16252 17584
rect 16205 17580 16252 17582
rect 16316 17580 16322 17644
rect 17861 17642 17927 17645
rect 19558 17642 19564 17644
rect 17861 17640 19564 17642
rect 17861 17584 17866 17640
rect 17922 17584 19564 17640
rect 17861 17582 19564 17584
rect 16205 17579 16271 17580
rect 17861 17579 17927 17582
rect 19558 17580 19564 17582
rect 19628 17580 19634 17644
rect 7946 17440 8262 17441
rect 7946 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8262 17440
rect 7946 17375 8262 17376
rect 17946 17440 18262 17441
rect 17946 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18262 17440
rect 17946 17375 18262 17376
rect 24669 17234 24735 17237
rect 26200 17234 27000 17264
rect 24669 17232 27000 17234
rect 24669 17176 24674 17232
rect 24730 17176 27000 17232
rect 24669 17174 27000 17176
rect 24669 17171 24735 17174
rect 26200 17144 27000 17174
rect 2946 16896 3262 16897
rect 2946 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3262 16896
rect 2946 16831 3262 16832
rect 12946 16896 13262 16897
rect 12946 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13262 16896
rect 12946 16831 13262 16832
rect 22946 16896 23262 16897
rect 22946 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23262 16896
rect 22946 16831 23262 16832
rect 24853 16554 24919 16557
rect 26200 16554 27000 16584
rect 24853 16552 27000 16554
rect 24853 16496 24858 16552
rect 24914 16496 27000 16552
rect 24853 16494 27000 16496
rect 24853 16491 24919 16494
rect 26200 16464 27000 16494
rect 7946 16352 8262 16353
rect 7946 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8262 16352
rect 7946 16287 8262 16288
rect 17946 16352 18262 16353
rect 17946 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18262 16352
rect 17946 16287 18262 16288
rect 12801 16010 12867 16013
rect 13486 16010 13492 16012
rect 12801 16008 13492 16010
rect 12801 15952 12806 16008
rect 12862 15952 13492 16008
rect 12801 15950 13492 15952
rect 12801 15947 12867 15950
rect 13486 15948 13492 15950
rect 13556 15948 13562 16012
rect 24853 15874 24919 15877
rect 26200 15874 27000 15904
rect 24853 15872 27000 15874
rect 24853 15816 24858 15872
rect 24914 15816 27000 15872
rect 24853 15814 27000 15816
rect 24853 15811 24919 15814
rect 2946 15808 3262 15809
rect 0 15738 800 15768
rect 2946 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3262 15808
rect 2946 15743 3262 15744
rect 12946 15808 13262 15809
rect 12946 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13262 15808
rect 12946 15743 13262 15744
rect 22946 15808 23262 15809
rect 22946 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23262 15808
rect 26200 15784 27000 15814
rect 22946 15743 23262 15744
rect 1301 15738 1367 15741
rect 0 15736 1367 15738
rect 0 15680 1306 15736
rect 1362 15680 1367 15736
rect 0 15678 1367 15680
rect 0 15648 800 15678
rect 1301 15675 1367 15678
rect 19977 15602 20043 15605
rect 21633 15602 21699 15605
rect 19977 15600 21699 15602
rect 19977 15544 19982 15600
rect 20038 15544 21638 15600
rect 21694 15544 21699 15600
rect 19977 15542 21699 15544
rect 19977 15539 20043 15542
rect 21633 15539 21699 15542
rect 12065 15330 12131 15333
rect 13854 15330 13860 15332
rect 12065 15328 13860 15330
rect 12065 15272 12070 15328
rect 12126 15272 13860 15328
rect 12065 15270 13860 15272
rect 12065 15267 12131 15270
rect 13854 15268 13860 15270
rect 13924 15268 13930 15332
rect 15694 15268 15700 15332
rect 15764 15330 15770 15332
rect 16021 15330 16087 15333
rect 15764 15328 16087 15330
rect 15764 15272 16026 15328
rect 16082 15272 16087 15328
rect 15764 15270 16087 15272
rect 15764 15268 15770 15270
rect 16021 15267 16087 15270
rect 7946 15264 8262 15265
rect 7946 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8262 15264
rect 7946 15199 8262 15200
rect 17946 15264 18262 15265
rect 17946 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18262 15264
rect 17946 15199 18262 15200
rect 25129 15194 25195 15197
rect 26200 15194 27000 15224
rect 25129 15192 27000 15194
rect 25129 15136 25134 15192
rect 25190 15136 27000 15192
rect 25129 15134 27000 15136
rect 25129 15131 25195 15134
rect 26200 15104 27000 15134
rect 2946 14720 3262 14721
rect 2946 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3262 14720
rect 2946 14655 3262 14656
rect 12946 14720 13262 14721
rect 12946 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13262 14720
rect 12946 14655 13262 14656
rect 22946 14720 23262 14721
rect 22946 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23262 14720
rect 22946 14655 23262 14656
rect 24853 14514 24919 14517
rect 26200 14514 27000 14544
rect 24853 14512 27000 14514
rect 24853 14456 24858 14512
rect 24914 14456 27000 14512
rect 24853 14454 27000 14456
rect 24853 14451 24919 14454
rect 26200 14424 27000 14454
rect 7946 14176 8262 14177
rect 7946 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8262 14176
rect 7946 14111 8262 14112
rect 17946 14176 18262 14177
rect 17946 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18262 14176
rect 17946 14111 18262 14112
rect 24761 13834 24827 13837
rect 26200 13834 27000 13864
rect 24761 13832 27000 13834
rect 24761 13776 24766 13832
rect 24822 13776 27000 13832
rect 24761 13774 27000 13776
rect 24761 13771 24827 13774
rect 26200 13744 27000 13774
rect 2946 13632 3262 13633
rect 2946 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3262 13632
rect 2946 13567 3262 13568
rect 12946 13632 13262 13633
rect 12946 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13262 13632
rect 12946 13567 13262 13568
rect 22946 13632 23262 13633
rect 22946 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23262 13632
rect 22946 13567 23262 13568
rect 19333 13562 19399 13565
rect 19558 13562 19564 13564
rect 19333 13560 19564 13562
rect 19333 13504 19338 13560
rect 19394 13504 19564 13560
rect 19333 13502 19564 13504
rect 19333 13499 19399 13502
rect 19558 13500 19564 13502
rect 19628 13500 19634 13564
rect 0 13426 800 13456
rect 1761 13426 1827 13429
rect 0 13424 1827 13426
rect 0 13368 1766 13424
rect 1822 13368 1827 13424
rect 0 13366 1827 13368
rect 0 13336 800 13366
rect 1761 13363 1827 13366
rect 24669 13154 24735 13157
rect 26200 13154 27000 13184
rect 24669 13152 27000 13154
rect 24669 13096 24674 13152
rect 24730 13096 27000 13152
rect 24669 13094 27000 13096
rect 24669 13091 24735 13094
rect 7946 13088 8262 13089
rect 7946 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8262 13088
rect 7946 13023 8262 13024
rect 17946 13088 18262 13089
rect 17946 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18262 13088
rect 26200 13064 27000 13094
rect 17946 13023 18262 13024
rect 2946 12544 3262 12545
rect 2946 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3262 12544
rect 2946 12479 3262 12480
rect 12946 12544 13262 12545
rect 12946 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13262 12544
rect 12946 12479 13262 12480
rect 22946 12544 23262 12545
rect 22946 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23262 12544
rect 22946 12479 23262 12480
rect 24853 12474 24919 12477
rect 26200 12474 27000 12504
rect 24853 12472 27000 12474
rect 24853 12416 24858 12472
rect 24914 12416 27000 12472
rect 24853 12414 27000 12416
rect 24853 12411 24919 12414
rect 26200 12384 27000 12414
rect 7946 12000 8262 12001
rect 7946 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8262 12000
rect 7946 11935 8262 11936
rect 17946 12000 18262 12001
rect 17946 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18262 12000
rect 17946 11935 18262 11936
rect 24945 11794 25011 11797
rect 26200 11794 27000 11824
rect 24945 11792 27000 11794
rect 24945 11736 24950 11792
rect 25006 11736 27000 11792
rect 24945 11734 27000 11736
rect 24945 11731 25011 11734
rect 26200 11704 27000 11734
rect 2946 11456 3262 11457
rect 2946 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3262 11456
rect 2946 11391 3262 11392
rect 12946 11456 13262 11457
rect 12946 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13262 11456
rect 12946 11391 13262 11392
rect 22946 11456 23262 11457
rect 22946 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23262 11456
rect 22946 11391 23262 11392
rect 0 11114 800 11144
rect 3325 11114 3391 11117
rect 0 11112 3391 11114
rect 0 11056 3330 11112
rect 3386 11056 3391 11112
rect 0 11054 3391 11056
rect 0 11024 800 11054
rect 3325 11051 3391 11054
rect 24761 11114 24827 11117
rect 26200 11114 27000 11144
rect 24761 11112 27000 11114
rect 24761 11056 24766 11112
rect 24822 11056 27000 11112
rect 24761 11054 27000 11056
rect 24761 11051 24827 11054
rect 26200 11024 27000 11054
rect 7946 10912 8262 10913
rect 7946 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8262 10912
rect 7946 10847 8262 10848
rect 17946 10912 18262 10913
rect 17946 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18262 10912
rect 17946 10847 18262 10848
rect 24761 10434 24827 10437
rect 26200 10434 27000 10464
rect 24761 10432 27000 10434
rect 24761 10376 24766 10432
rect 24822 10376 27000 10432
rect 24761 10374 27000 10376
rect 24761 10371 24827 10374
rect 2946 10368 3262 10369
rect 2946 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3262 10368
rect 2946 10303 3262 10304
rect 12946 10368 13262 10369
rect 12946 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13262 10368
rect 12946 10303 13262 10304
rect 22946 10368 23262 10369
rect 22946 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23262 10368
rect 26200 10344 27000 10374
rect 22946 10303 23262 10304
rect 7946 9824 8262 9825
rect 7946 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8262 9824
rect 7946 9759 8262 9760
rect 17946 9824 18262 9825
rect 17946 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18262 9824
rect 17946 9759 18262 9760
rect 24853 9754 24919 9757
rect 26200 9754 27000 9784
rect 24853 9752 27000 9754
rect 24853 9696 24858 9752
rect 24914 9696 27000 9752
rect 24853 9694 27000 9696
rect 24853 9691 24919 9694
rect 26200 9664 27000 9694
rect 2946 9280 3262 9281
rect 2946 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3262 9280
rect 2946 9215 3262 9216
rect 12946 9280 13262 9281
rect 12946 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13262 9280
rect 12946 9215 13262 9216
rect 22946 9280 23262 9281
rect 22946 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23262 9280
rect 22946 9215 23262 9216
rect 25129 9074 25195 9077
rect 26200 9074 27000 9104
rect 25129 9072 27000 9074
rect 25129 9016 25134 9072
rect 25190 9016 27000 9072
rect 25129 9014 27000 9016
rect 25129 9011 25195 9014
rect 26200 8984 27000 9014
rect 0 8802 800 8832
rect 2865 8802 2931 8805
rect 0 8800 2931 8802
rect 0 8744 2870 8800
rect 2926 8744 2931 8800
rect 0 8742 2931 8744
rect 0 8712 800 8742
rect 2865 8739 2931 8742
rect 7946 8736 8262 8737
rect 7946 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8262 8736
rect 7946 8671 8262 8672
rect 17946 8736 18262 8737
rect 17946 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18262 8736
rect 17946 8671 18262 8672
rect 24761 8394 24827 8397
rect 26200 8394 27000 8424
rect 24761 8392 27000 8394
rect 24761 8336 24766 8392
rect 24822 8336 27000 8392
rect 24761 8334 27000 8336
rect 24761 8331 24827 8334
rect 26200 8304 27000 8334
rect 2946 8192 3262 8193
rect 2946 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3262 8192
rect 2946 8127 3262 8128
rect 12946 8192 13262 8193
rect 12946 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13262 8192
rect 12946 8127 13262 8128
rect 22946 8192 23262 8193
rect 22946 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23262 8192
rect 22946 8127 23262 8128
rect 24945 7714 25011 7717
rect 26200 7714 27000 7744
rect 24945 7712 27000 7714
rect 24945 7656 24950 7712
rect 25006 7656 27000 7712
rect 24945 7654 27000 7656
rect 24945 7651 25011 7654
rect 7946 7648 8262 7649
rect 7946 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8262 7648
rect 7946 7583 8262 7584
rect 17946 7648 18262 7649
rect 17946 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18262 7648
rect 26200 7624 27000 7654
rect 17946 7583 18262 7584
rect 2946 7104 3262 7105
rect 2946 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3262 7104
rect 2946 7039 3262 7040
rect 12946 7104 13262 7105
rect 12946 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13262 7104
rect 12946 7039 13262 7040
rect 22946 7104 23262 7105
rect 22946 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23262 7104
rect 22946 7039 23262 7040
rect 24761 7034 24827 7037
rect 26200 7034 27000 7064
rect 24761 7032 27000 7034
rect 24761 6976 24766 7032
rect 24822 6976 27000 7032
rect 24761 6974 27000 6976
rect 24761 6971 24827 6974
rect 26200 6944 27000 6974
rect 7946 6560 8262 6561
rect 0 6490 800 6520
rect 7946 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8262 6560
rect 7946 6495 8262 6496
rect 17946 6560 18262 6561
rect 17946 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18262 6560
rect 17946 6495 18262 6496
rect 3141 6490 3207 6493
rect 0 6488 3207 6490
rect 0 6432 3146 6488
rect 3202 6432 3207 6488
rect 0 6430 3207 6432
rect 0 6400 800 6430
rect 3141 6427 3207 6430
rect 24853 6354 24919 6357
rect 26200 6354 27000 6384
rect 24853 6352 27000 6354
rect 24853 6296 24858 6352
rect 24914 6296 27000 6352
rect 24853 6294 27000 6296
rect 24853 6291 24919 6294
rect 26200 6264 27000 6294
rect 2946 6016 3262 6017
rect 2946 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3262 6016
rect 2946 5951 3262 5952
rect 12946 6016 13262 6017
rect 12946 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13262 6016
rect 12946 5951 13262 5952
rect 22946 6016 23262 6017
rect 22946 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23262 6016
rect 22946 5951 23262 5952
rect 7833 5810 7899 5813
rect 14958 5810 14964 5812
rect 7833 5808 14964 5810
rect 7833 5752 7838 5808
rect 7894 5752 14964 5808
rect 7833 5750 14964 5752
rect 7833 5747 7899 5750
rect 14958 5748 14964 5750
rect 15028 5748 15034 5812
rect 7741 5674 7807 5677
rect 10174 5674 10180 5676
rect 7741 5672 10180 5674
rect 7741 5616 7746 5672
rect 7802 5616 10180 5672
rect 7741 5614 10180 5616
rect 7741 5611 7807 5614
rect 10174 5612 10180 5614
rect 10244 5612 10250 5676
rect 24761 5674 24827 5677
rect 26200 5674 27000 5704
rect 24761 5672 27000 5674
rect 24761 5616 24766 5672
rect 24822 5616 27000 5672
rect 24761 5614 27000 5616
rect 24761 5611 24827 5614
rect 26200 5584 27000 5614
rect 7946 5472 8262 5473
rect 7946 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8262 5472
rect 7946 5407 8262 5408
rect 17946 5472 18262 5473
rect 17946 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18262 5472
rect 17946 5407 18262 5408
rect 25313 4994 25379 4997
rect 26200 4994 27000 5024
rect 25313 4992 27000 4994
rect 25313 4936 25318 4992
rect 25374 4936 27000 4992
rect 25313 4934 27000 4936
rect 25313 4931 25379 4934
rect 2946 4928 3262 4929
rect 2946 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3262 4928
rect 2946 4863 3262 4864
rect 12946 4928 13262 4929
rect 12946 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13262 4928
rect 12946 4863 13262 4864
rect 22946 4928 23262 4929
rect 22946 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23262 4928
rect 26200 4904 27000 4934
rect 22946 4863 23262 4864
rect 7946 4384 8262 4385
rect 7946 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8262 4384
rect 7946 4319 8262 4320
rect 17946 4384 18262 4385
rect 17946 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18262 4384
rect 17946 4319 18262 4320
rect 23381 4314 23447 4317
rect 26200 4314 27000 4344
rect 23381 4312 27000 4314
rect 23381 4256 23386 4312
rect 23442 4256 27000 4312
rect 23381 4254 27000 4256
rect 23381 4251 23447 4254
rect 26200 4224 27000 4254
rect 0 4178 800 4208
rect 3233 4178 3299 4181
rect 0 4176 3299 4178
rect 0 4120 3238 4176
rect 3294 4120 3299 4176
rect 0 4118 3299 4120
rect 0 4088 800 4118
rect 3233 4115 3299 4118
rect 2946 3840 3262 3841
rect 2946 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3262 3840
rect 2946 3775 3262 3776
rect 12946 3840 13262 3841
rect 12946 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13262 3840
rect 12946 3775 13262 3776
rect 22946 3840 23262 3841
rect 22946 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23262 3840
rect 22946 3775 23262 3776
rect 16798 3436 16804 3500
rect 16868 3498 16874 3500
rect 23289 3498 23355 3501
rect 16868 3496 23355 3498
rect 16868 3440 23294 3496
rect 23350 3440 23355 3496
rect 16868 3438 23355 3440
rect 16868 3436 16874 3438
rect 23289 3435 23355 3438
rect 7946 3296 8262 3297
rect 7946 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8262 3296
rect 7946 3231 8262 3232
rect 17946 3296 18262 3297
rect 17946 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18262 3296
rect 17946 3231 18262 3232
rect 2946 2752 3262 2753
rect 2946 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3262 2752
rect 2946 2687 3262 2688
rect 12946 2752 13262 2753
rect 12946 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13262 2752
rect 12946 2687 13262 2688
rect 22946 2752 23262 2753
rect 22946 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23262 2752
rect 22946 2687 23262 2688
rect 15653 2684 15719 2685
rect 15653 2680 15700 2684
rect 15764 2682 15770 2684
rect 15653 2624 15658 2680
rect 15653 2620 15700 2624
rect 15764 2622 15810 2682
rect 15764 2620 15770 2622
rect 15653 2619 15719 2620
rect 7946 2208 8262 2209
rect 7946 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8262 2208
rect 7946 2143 8262 2144
rect 17946 2208 18262 2209
rect 17946 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18262 2208
rect 17946 2143 18262 2144
rect 0 1866 800 1896
rect 2773 1866 2839 1869
rect 0 1864 2839 1866
rect 0 1808 2778 1864
rect 2834 1808 2839 1864
rect 0 1806 2839 1808
rect 0 1776 800 1806
rect 2773 1803 2839 1806
<< via3 >>
rect 7952 54428 8016 54432
rect 7952 54372 7956 54428
rect 7956 54372 8012 54428
rect 8012 54372 8016 54428
rect 7952 54368 8016 54372
rect 8032 54428 8096 54432
rect 8032 54372 8036 54428
rect 8036 54372 8092 54428
rect 8092 54372 8096 54428
rect 8032 54368 8096 54372
rect 8112 54428 8176 54432
rect 8112 54372 8116 54428
rect 8116 54372 8172 54428
rect 8172 54372 8176 54428
rect 8112 54368 8176 54372
rect 8192 54428 8256 54432
rect 8192 54372 8196 54428
rect 8196 54372 8252 54428
rect 8252 54372 8256 54428
rect 8192 54368 8256 54372
rect 17952 54428 18016 54432
rect 17952 54372 17956 54428
rect 17956 54372 18012 54428
rect 18012 54372 18016 54428
rect 17952 54368 18016 54372
rect 18032 54428 18096 54432
rect 18032 54372 18036 54428
rect 18036 54372 18092 54428
rect 18092 54372 18096 54428
rect 18032 54368 18096 54372
rect 18112 54428 18176 54432
rect 18112 54372 18116 54428
rect 18116 54372 18172 54428
rect 18172 54372 18176 54428
rect 18112 54368 18176 54372
rect 18192 54428 18256 54432
rect 18192 54372 18196 54428
rect 18196 54372 18252 54428
rect 18252 54372 18256 54428
rect 18192 54368 18256 54372
rect 15884 53892 15948 53956
rect 2952 53884 3016 53888
rect 2952 53828 2956 53884
rect 2956 53828 3012 53884
rect 3012 53828 3016 53884
rect 2952 53824 3016 53828
rect 3032 53884 3096 53888
rect 3032 53828 3036 53884
rect 3036 53828 3092 53884
rect 3092 53828 3096 53884
rect 3032 53824 3096 53828
rect 3112 53884 3176 53888
rect 3112 53828 3116 53884
rect 3116 53828 3172 53884
rect 3172 53828 3176 53884
rect 3112 53824 3176 53828
rect 3192 53884 3256 53888
rect 3192 53828 3196 53884
rect 3196 53828 3252 53884
rect 3252 53828 3256 53884
rect 3192 53824 3256 53828
rect 12952 53884 13016 53888
rect 12952 53828 12956 53884
rect 12956 53828 13012 53884
rect 13012 53828 13016 53884
rect 12952 53824 13016 53828
rect 13032 53884 13096 53888
rect 13032 53828 13036 53884
rect 13036 53828 13092 53884
rect 13092 53828 13096 53884
rect 13032 53824 13096 53828
rect 13112 53884 13176 53888
rect 13112 53828 13116 53884
rect 13116 53828 13172 53884
rect 13172 53828 13176 53884
rect 13112 53824 13176 53828
rect 13192 53884 13256 53888
rect 13192 53828 13196 53884
rect 13196 53828 13252 53884
rect 13252 53828 13256 53884
rect 13192 53824 13256 53828
rect 22952 53884 23016 53888
rect 22952 53828 22956 53884
rect 22956 53828 23012 53884
rect 23012 53828 23016 53884
rect 22952 53824 23016 53828
rect 23032 53884 23096 53888
rect 23032 53828 23036 53884
rect 23036 53828 23092 53884
rect 23092 53828 23096 53884
rect 23032 53824 23096 53828
rect 23112 53884 23176 53888
rect 23112 53828 23116 53884
rect 23116 53828 23172 53884
rect 23172 53828 23176 53884
rect 23112 53824 23176 53828
rect 23192 53884 23256 53888
rect 23192 53828 23196 53884
rect 23196 53828 23252 53884
rect 23252 53828 23256 53884
rect 23192 53824 23256 53828
rect 7952 53340 8016 53344
rect 7952 53284 7956 53340
rect 7956 53284 8012 53340
rect 8012 53284 8016 53340
rect 7952 53280 8016 53284
rect 8032 53340 8096 53344
rect 8032 53284 8036 53340
rect 8036 53284 8092 53340
rect 8092 53284 8096 53340
rect 8032 53280 8096 53284
rect 8112 53340 8176 53344
rect 8112 53284 8116 53340
rect 8116 53284 8172 53340
rect 8172 53284 8176 53340
rect 8112 53280 8176 53284
rect 8192 53340 8256 53344
rect 8192 53284 8196 53340
rect 8196 53284 8252 53340
rect 8252 53284 8256 53340
rect 8192 53280 8256 53284
rect 17952 53340 18016 53344
rect 17952 53284 17956 53340
rect 17956 53284 18012 53340
rect 18012 53284 18016 53340
rect 17952 53280 18016 53284
rect 18032 53340 18096 53344
rect 18032 53284 18036 53340
rect 18036 53284 18092 53340
rect 18092 53284 18096 53340
rect 18032 53280 18096 53284
rect 18112 53340 18176 53344
rect 18112 53284 18116 53340
rect 18116 53284 18172 53340
rect 18172 53284 18176 53340
rect 18112 53280 18176 53284
rect 18192 53340 18256 53344
rect 18192 53284 18196 53340
rect 18196 53284 18252 53340
rect 18252 53284 18256 53340
rect 18192 53280 18256 53284
rect 2952 52796 3016 52800
rect 2952 52740 2956 52796
rect 2956 52740 3012 52796
rect 3012 52740 3016 52796
rect 2952 52736 3016 52740
rect 3032 52796 3096 52800
rect 3032 52740 3036 52796
rect 3036 52740 3092 52796
rect 3092 52740 3096 52796
rect 3032 52736 3096 52740
rect 3112 52796 3176 52800
rect 3112 52740 3116 52796
rect 3116 52740 3172 52796
rect 3172 52740 3176 52796
rect 3112 52736 3176 52740
rect 3192 52796 3256 52800
rect 3192 52740 3196 52796
rect 3196 52740 3252 52796
rect 3252 52740 3256 52796
rect 3192 52736 3256 52740
rect 12952 52796 13016 52800
rect 12952 52740 12956 52796
rect 12956 52740 13012 52796
rect 13012 52740 13016 52796
rect 12952 52736 13016 52740
rect 13032 52796 13096 52800
rect 13032 52740 13036 52796
rect 13036 52740 13092 52796
rect 13092 52740 13096 52796
rect 13032 52736 13096 52740
rect 13112 52796 13176 52800
rect 13112 52740 13116 52796
rect 13116 52740 13172 52796
rect 13172 52740 13176 52796
rect 13112 52736 13176 52740
rect 13192 52796 13256 52800
rect 13192 52740 13196 52796
rect 13196 52740 13252 52796
rect 13252 52740 13256 52796
rect 13192 52736 13256 52740
rect 22952 52796 23016 52800
rect 22952 52740 22956 52796
rect 22956 52740 23012 52796
rect 23012 52740 23016 52796
rect 22952 52736 23016 52740
rect 23032 52796 23096 52800
rect 23032 52740 23036 52796
rect 23036 52740 23092 52796
rect 23092 52740 23096 52796
rect 23032 52736 23096 52740
rect 23112 52796 23176 52800
rect 23112 52740 23116 52796
rect 23116 52740 23172 52796
rect 23172 52740 23176 52796
rect 23112 52736 23176 52740
rect 23192 52796 23256 52800
rect 23192 52740 23196 52796
rect 23196 52740 23252 52796
rect 23252 52740 23256 52796
rect 23192 52736 23256 52740
rect 14412 52592 14476 52596
rect 14412 52536 14426 52592
rect 14426 52536 14476 52592
rect 14412 52532 14476 52536
rect 15700 52532 15764 52596
rect 22324 52532 22388 52596
rect 7952 52252 8016 52256
rect 7952 52196 7956 52252
rect 7956 52196 8012 52252
rect 8012 52196 8016 52252
rect 7952 52192 8016 52196
rect 8032 52252 8096 52256
rect 8032 52196 8036 52252
rect 8036 52196 8092 52252
rect 8092 52196 8096 52252
rect 8032 52192 8096 52196
rect 8112 52252 8176 52256
rect 8112 52196 8116 52252
rect 8116 52196 8172 52252
rect 8172 52196 8176 52252
rect 8112 52192 8176 52196
rect 8192 52252 8256 52256
rect 8192 52196 8196 52252
rect 8196 52196 8252 52252
rect 8252 52196 8256 52252
rect 8192 52192 8256 52196
rect 17952 52252 18016 52256
rect 17952 52196 17956 52252
rect 17956 52196 18012 52252
rect 18012 52196 18016 52252
rect 17952 52192 18016 52196
rect 18032 52252 18096 52256
rect 18032 52196 18036 52252
rect 18036 52196 18092 52252
rect 18092 52196 18096 52252
rect 18032 52192 18096 52196
rect 18112 52252 18176 52256
rect 18112 52196 18116 52252
rect 18116 52196 18172 52252
rect 18172 52196 18176 52252
rect 18112 52192 18176 52196
rect 18192 52252 18256 52256
rect 18192 52196 18196 52252
rect 18196 52196 18252 52252
rect 18252 52196 18256 52252
rect 18192 52192 18256 52196
rect 2952 51708 3016 51712
rect 2952 51652 2956 51708
rect 2956 51652 3012 51708
rect 3012 51652 3016 51708
rect 2952 51648 3016 51652
rect 3032 51708 3096 51712
rect 3032 51652 3036 51708
rect 3036 51652 3092 51708
rect 3092 51652 3096 51708
rect 3032 51648 3096 51652
rect 3112 51708 3176 51712
rect 3112 51652 3116 51708
rect 3116 51652 3172 51708
rect 3172 51652 3176 51708
rect 3112 51648 3176 51652
rect 3192 51708 3256 51712
rect 3192 51652 3196 51708
rect 3196 51652 3252 51708
rect 3252 51652 3256 51708
rect 3192 51648 3256 51652
rect 12952 51708 13016 51712
rect 12952 51652 12956 51708
rect 12956 51652 13012 51708
rect 13012 51652 13016 51708
rect 12952 51648 13016 51652
rect 13032 51708 13096 51712
rect 13032 51652 13036 51708
rect 13036 51652 13092 51708
rect 13092 51652 13096 51708
rect 13032 51648 13096 51652
rect 13112 51708 13176 51712
rect 13112 51652 13116 51708
rect 13116 51652 13172 51708
rect 13172 51652 13176 51708
rect 13112 51648 13176 51652
rect 13192 51708 13256 51712
rect 13192 51652 13196 51708
rect 13196 51652 13252 51708
rect 13252 51652 13256 51708
rect 13192 51648 13256 51652
rect 22952 51708 23016 51712
rect 22952 51652 22956 51708
rect 22956 51652 23012 51708
rect 23012 51652 23016 51708
rect 22952 51648 23016 51652
rect 23032 51708 23096 51712
rect 23032 51652 23036 51708
rect 23036 51652 23092 51708
rect 23092 51652 23096 51708
rect 23032 51648 23096 51652
rect 23112 51708 23176 51712
rect 23112 51652 23116 51708
rect 23116 51652 23172 51708
rect 23172 51652 23176 51708
rect 23112 51648 23176 51652
rect 23192 51708 23256 51712
rect 23192 51652 23196 51708
rect 23196 51652 23252 51708
rect 23252 51652 23256 51708
rect 23192 51648 23256 51652
rect 7952 51164 8016 51168
rect 7952 51108 7956 51164
rect 7956 51108 8012 51164
rect 8012 51108 8016 51164
rect 7952 51104 8016 51108
rect 8032 51164 8096 51168
rect 8032 51108 8036 51164
rect 8036 51108 8092 51164
rect 8092 51108 8096 51164
rect 8032 51104 8096 51108
rect 8112 51164 8176 51168
rect 8112 51108 8116 51164
rect 8116 51108 8172 51164
rect 8172 51108 8176 51164
rect 8112 51104 8176 51108
rect 8192 51164 8256 51168
rect 8192 51108 8196 51164
rect 8196 51108 8252 51164
rect 8252 51108 8256 51164
rect 8192 51104 8256 51108
rect 17952 51164 18016 51168
rect 17952 51108 17956 51164
rect 17956 51108 18012 51164
rect 18012 51108 18016 51164
rect 17952 51104 18016 51108
rect 18032 51164 18096 51168
rect 18032 51108 18036 51164
rect 18036 51108 18092 51164
rect 18092 51108 18096 51164
rect 18032 51104 18096 51108
rect 18112 51164 18176 51168
rect 18112 51108 18116 51164
rect 18116 51108 18172 51164
rect 18172 51108 18176 51164
rect 18112 51104 18176 51108
rect 18192 51164 18256 51168
rect 18192 51108 18196 51164
rect 18196 51108 18252 51164
rect 18252 51108 18256 51164
rect 18192 51104 18256 51108
rect 2952 50620 3016 50624
rect 2952 50564 2956 50620
rect 2956 50564 3012 50620
rect 3012 50564 3016 50620
rect 2952 50560 3016 50564
rect 3032 50620 3096 50624
rect 3032 50564 3036 50620
rect 3036 50564 3092 50620
rect 3092 50564 3096 50620
rect 3032 50560 3096 50564
rect 3112 50620 3176 50624
rect 3112 50564 3116 50620
rect 3116 50564 3172 50620
rect 3172 50564 3176 50620
rect 3112 50560 3176 50564
rect 3192 50620 3256 50624
rect 3192 50564 3196 50620
rect 3196 50564 3252 50620
rect 3252 50564 3256 50620
rect 3192 50560 3256 50564
rect 12952 50620 13016 50624
rect 12952 50564 12956 50620
rect 12956 50564 13012 50620
rect 13012 50564 13016 50620
rect 12952 50560 13016 50564
rect 13032 50620 13096 50624
rect 13032 50564 13036 50620
rect 13036 50564 13092 50620
rect 13092 50564 13096 50620
rect 13032 50560 13096 50564
rect 13112 50620 13176 50624
rect 13112 50564 13116 50620
rect 13116 50564 13172 50620
rect 13172 50564 13176 50620
rect 13112 50560 13176 50564
rect 13192 50620 13256 50624
rect 13192 50564 13196 50620
rect 13196 50564 13252 50620
rect 13252 50564 13256 50620
rect 13192 50560 13256 50564
rect 22952 50620 23016 50624
rect 22952 50564 22956 50620
rect 22956 50564 23012 50620
rect 23012 50564 23016 50620
rect 22952 50560 23016 50564
rect 23032 50620 23096 50624
rect 23032 50564 23036 50620
rect 23036 50564 23092 50620
rect 23092 50564 23096 50620
rect 23032 50560 23096 50564
rect 23112 50620 23176 50624
rect 23112 50564 23116 50620
rect 23116 50564 23172 50620
rect 23172 50564 23176 50620
rect 23112 50560 23176 50564
rect 23192 50620 23256 50624
rect 23192 50564 23196 50620
rect 23196 50564 23252 50620
rect 23252 50564 23256 50620
rect 23192 50560 23256 50564
rect 7952 50076 8016 50080
rect 7952 50020 7956 50076
rect 7956 50020 8012 50076
rect 8012 50020 8016 50076
rect 7952 50016 8016 50020
rect 8032 50076 8096 50080
rect 8032 50020 8036 50076
rect 8036 50020 8092 50076
rect 8092 50020 8096 50076
rect 8032 50016 8096 50020
rect 8112 50076 8176 50080
rect 8112 50020 8116 50076
rect 8116 50020 8172 50076
rect 8172 50020 8176 50076
rect 8112 50016 8176 50020
rect 8192 50076 8256 50080
rect 8192 50020 8196 50076
rect 8196 50020 8252 50076
rect 8252 50020 8256 50076
rect 8192 50016 8256 50020
rect 17952 50076 18016 50080
rect 17952 50020 17956 50076
rect 17956 50020 18012 50076
rect 18012 50020 18016 50076
rect 17952 50016 18016 50020
rect 18032 50076 18096 50080
rect 18032 50020 18036 50076
rect 18036 50020 18092 50076
rect 18092 50020 18096 50076
rect 18032 50016 18096 50020
rect 18112 50076 18176 50080
rect 18112 50020 18116 50076
rect 18116 50020 18172 50076
rect 18172 50020 18176 50076
rect 18112 50016 18176 50020
rect 18192 50076 18256 50080
rect 18192 50020 18196 50076
rect 18196 50020 18252 50076
rect 18252 50020 18256 50076
rect 18192 50016 18256 50020
rect 2952 49532 3016 49536
rect 2952 49476 2956 49532
rect 2956 49476 3012 49532
rect 3012 49476 3016 49532
rect 2952 49472 3016 49476
rect 3032 49532 3096 49536
rect 3032 49476 3036 49532
rect 3036 49476 3092 49532
rect 3092 49476 3096 49532
rect 3032 49472 3096 49476
rect 3112 49532 3176 49536
rect 3112 49476 3116 49532
rect 3116 49476 3172 49532
rect 3172 49476 3176 49532
rect 3112 49472 3176 49476
rect 3192 49532 3256 49536
rect 3192 49476 3196 49532
rect 3196 49476 3252 49532
rect 3252 49476 3256 49532
rect 3192 49472 3256 49476
rect 12952 49532 13016 49536
rect 12952 49476 12956 49532
rect 12956 49476 13012 49532
rect 13012 49476 13016 49532
rect 12952 49472 13016 49476
rect 13032 49532 13096 49536
rect 13032 49476 13036 49532
rect 13036 49476 13092 49532
rect 13092 49476 13096 49532
rect 13032 49472 13096 49476
rect 13112 49532 13176 49536
rect 13112 49476 13116 49532
rect 13116 49476 13172 49532
rect 13172 49476 13176 49532
rect 13112 49472 13176 49476
rect 13192 49532 13256 49536
rect 13192 49476 13196 49532
rect 13196 49476 13252 49532
rect 13252 49476 13256 49532
rect 13192 49472 13256 49476
rect 22952 49532 23016 49536
rect 22952 49476 22956 49532
rect 22956 49476 23012 49532
rect 23012 49476 23016 49532
rect 22952 49472 23016 49476
rect 23032 49532 23096 49536
rect 23032 49476 23036 49532
rect 23036 49476 23092 49532
rect 23092 49476 23096 49532
rect 23032 49472 23096 49476
rect 23112 49532 23176 49536
rect 23112 49476 23116 49532
rect 23116 49476 23172 49532
rect 23172 49476 23176 49532
rect 23112 49472 23176 49476
rect 23192 49532 23256 49536
rect 23192 49476 23196 49532
rect 23196 49476 23252 49532
rect 23252 49476 23256 49532
rect 23192 49472 23256 49476
rect 7952 48988 8016 48992
rect 7952 48932 7956 48988
rect 7956 48932 8012 48988
rect 8012 48932 8016 48988
rect 7952 48928 8016 48932
rect 8032 48988 8096 48992
rect 8032 48932 8036 48988
rect 8036 48932 8092 48988
rect 8092 48932 8096 48988
rect 8032 48928 8096 48932
rect 8112 48988 8176 48992
rect 8112 48932 8116 48988
rect 8116 48932 8172 48988
rect 8172 48932 8176 48988
rect 8112 48928 8176 48932
rect 8192 48988 8256 48992
rect 8192 48932 8196 48988
rect 8196 48932 8252 48988
rect 8252 48932 8256 48988
rect 8192 48928 8256 48932
rect 17952 48988 18016 48992
rect 17952 48932 17956 48988
rect 17956 48932 18012 48988
rect 18012 48932 18016 48988
rect 17952 48928 18016 48932
rect 18032 48988 18096 48992
rect 18032 48932 18036 48988
rect 18036 48932 18092 48988
rect 18092 48932 18096 48988
rect 18032 48928 18096 48932
rect 18112 48988 18176 48992
rect 18112 48932 18116 48988
rect 18116 48932 18172 48988
rect 18172 48932 18176 48988
rect 18112 48928 18176 48932
rect 18192 48988 18256 48992
rect 18192 48932 18196 48988
rect 18196 48932 18252 48988
rect 18252 48932 18256 48988
rect 18192 48928 18256 48932
rect 2952 48444 3016 48448
rect 2952 48388 2956 48444
rect 2956 48388 3012 48444
rect 3012 48388 3016 48444
rect 2952 48384 3016 48388
rect 3032 48444 3096 48448
rect 3032 48388 3036 48444
rect 3036 48388 3092 48444
rect 3092 48388 3096 48444
rect 3032 48384 3096 48388
rect 3112 48444 3176 48448
rect 3112 48388 3116 48444
rect 3116 48388 3172 48444
rect 3172 48388 3176 48444
rect 3112 48384 3176 48388
rect 3192 48444 3256 48448
rect 3192 48388 3196 48444
rect 3196 48388 3252 48444
rect 3252 48388 3256 48444
rect 3192 48384 3256 48388
rect 12952 48444 13016 48448
rect 12952 48388 12956 48444
rect 12956 48388 13012 48444
rect 13012 48388 13016 48444
rect 12952 48384 13016 48388
rect 13032 48444 13096 48448
rect 13032 48388 13036 48444
rect 13036 48388 13092 48444
rect 13092 48388 13096 48444
rect 13032 48384 13096 48388
rect 13112 48444 13176 48448
rect 13112 48388 13116 48444
rect 13116 48388 13172 48444
rect 13172 48388 13176 48444
rect 13112 48384 13176 48388
rect 13192 48444 13256 48448
rect 13192 48388 13196 48444
rect 13196 48388 13252 48444
rect 13252 48388 13256 48444
rect 13192 48384 13256 48388
rect 22952 48444 23016 48448
rect 22952 48388 22956 48444
rect 22956 48388 23012 48444
rect 23012 48388 23016 48444
rect 22952 48384 23016 48388
rect 23032 48444 23096 48448
rect 23032 48388 23036 48444
rect 23036 48388 23092 48444
rect 23092 48388 23096 48444
rect 23032 48384 23096 48388
rect 23112 48444 23176 48448
rect 23112 48388 23116 48444
rect 23116 48388 23172 48444
rect 23172 48388 23176 48444
rect 23112 48384 23176 48388
rect 23192 48444 23256 48448
rect 23192 48388 23196 48444
rect 23196 48388 23252 48444
rect 23252 48388 23256 48444
rect 23192 48384 23256 48388
rect 7952 47900 8016 47904
rect 7952 47844 7956 47900
rect 7956 47844 8012 47900
rect 8012 47844 8016 47900
rect 7952 47840 8016 47844
rect 8032 47900 8096 47904
rect 8032 47844 8036 47900
rect 8036 47844 8092 47900
rect 8092 47844 8096 47900
rect 8032 47840 8096 47844
rect 8112 47900 8176 47904
rect 8112 47844 8116 47900
rect 8116 47844 8172 47900
rect 8172 47844 8176 47900
rect 8112 47840 8176 47844
rect 8192 47900 8256 47904
rect 8192 47844 8196 47900
rect 8196 47844 8252 47900
rect 8252 47844 8256 47900
rect 8192 47840 8256 47844
rect 17952 47900 18016 47904
rect 17952 47844 17956 47900
rect 17956 47844 18012 47900
rect 18012 47844 18016 47900
rect 17952 47840 18016 47844
rect 18032 47900 18096 47904
rect 18032 47844 18036 47900
rect 18036 47844 18092 47900
rect 18092 47844 18096 47900
rect 18032 47840 18096 47844
rect 18112 47900 18176 47904
rect 18112 47844 18116 47900
rect 18116 47844 18172 47900
rect 18172 47844 18176 47900
rect 18112 47840 18176 47844
rect 18192 47900 18256 47904
rect 18192 47844 18196 47900
rect 18196 47844 18252 47900
rect 18252 47844 18256 47900
rect 18192 47840 18256 47844
rect 2952 47356 3016 47360
rect 2952 47300 2956 47356
rect 2956 47300 3012 47356
rect 3012 47300 3016 47356
rect 2952 47296 3016 47300
rect 3032 47356 3096 47360
rect 3032 47300 3036 47356
rect 3036 47300 3092 47356
rect 3092 47300 3096 47356
rect 3032 47296 3096 47300
rect 3112 47356 3176 47360
rect 3112 47300 3116 47356
rect 3116 47300 3172 47356
rect 3172 47300 3176 47356
rect 3112 47296 3176 47300
rect 3192 47356 3256 47360
rect 3192 47300 3196 47356
rect 3196 47300 3252 47356
rect 3252 47300 3256 47356
rect 3192 47296 3256 47300
rect 12952 47356 13016 47360
rect 12952 47300 12956 47356
rect 12956 47300 13012 47356
rect 13012 47300 13016 47356
rect 12952 47296 13016 47300
rect 13032 47356 13096 47360
rect 13032 47300 13036 47356
rect 13036 47300 13092 47356
rect 13092 47300 13096 47356
rect 13032 47296 13096 47300
rect 13112 47356 13176 47360
rect 13112 47300 13116 47356
rect 13116 47300 13172 47356
rect 13172 47300 13176 47356
rect 13112 47296 13176 47300
rect 13192 47356 13256 47360
rect 13192 47300 13196 47356
rect 13196 47300 13252 47356
rect 13252 47300 13256 47356
rect 13192 47296 13256 47300
rect 22952 47356 23016 47360
rect 22952 47300 22956 47356
rect 22956 47300 23012 47356
rect 23012 47300 23016 47356
rect 22952 47296 23016 47300
rect 23032 47356 23096 47360
rect 23032 47300 23036 47356
rect 23036 47300 23092 47356
rect 23092 47300 23096 47356
rect 23032 47296 23096 47300
rect 23112 47356 23176 47360
rect 23112 47300 23116 47356
rect 23116 47300 23172 47356
rect 23172 47300 23176 47356
rect 23112 47296 23176 47300
rect 23192 47356 23256 47360
rect 23192 47300 23196 47356
rect 23196 47300 23252 47356
rect 23252 47300 23256 47356
rect 23192 47296 23256 47300
rect 7952 46812 8016 46816
rect 7952 46756 7956 46812
rect 7956 46756 8012 46812
rect 8012 46756 8016 46812
rect 7952 46752 8016 46756
rect 8032 46812 8096 46816
rect 8032 46756 8036 46812
rect 8036 46756 8092 46812
rect 8092 46756 8096 46812
rect 8032 46752 8096 46756
rect 8112 46812 8176 46816
rect 8112 46756 8116 46812
rect 8116 46756 8172 46812
rect 8172 46756 8176 46812
rect 8112 46752 8176 46756
rect 8192 46812 8256 46816
rect 8192 46756 8196 46812
rect 8196 46756 8252 46812
rect 8252 46756 8256 46812
rect 8192 46752 8256 46756
rect 17952 46812 18016 46816
rect 17952 46756 17956 46812
rect 17956 46756 18012 46812
rect 18012 46756 18016 46812
rect 17952 46752 18016 46756
rect 18032 46812 18096 46816
rect 18032 46756 18036 46812
rect 18036 46756 18092 46812
rect 18092 46756 18096 46812
rect 18032 46752 18096 46756
rect 18112 46812 18176 46816
rect 18112 46756 18116 46812
rect 18116 46756 18172 46812
rect 18172 46756 18176 46812
rect 18112 46752 18176 46756
rect 18192 46812 18256 46816
rect 18192 46756 18196 46812
rect 18196 46756 18252 46812
rect 18252 46756 18256 46812
rect 18192 46752 18256 46756
rect 2952 46268 3016 46272
rect 2952 46212 2956 46268
rect 2956 46212 3012 46268
rect 3012 46212 3016 46268
rect 2952 46208 3016 46212
rect 3032 46268 3096 46272
rect 3032 46212 3036 46268
rect 3036 46212 3092 46268
rect 3092 46212 3096 46268
rect 3032 46208 3096 46212
rect 3112 46268 3176 46272
rect 3112 46212 3116 46268
rect 3116 46212 3172 46268
rect 3172 46212 3176 46268
rect 3112 46208 3176 46212
rect 3192 46268 3256 46272
rect 3192 46212 3196 46268
rect 3196 46212 3252 46268
rect 3252 46212 3256 46268
rect 3192 46208 3256 46212
rect 12952 46268 13016 46272
rect 12952 46212 12956 46268
rect 12956 46212 13012 46268
rect 13012 46212 13016 46268
rect 12952 46208 13016 46212
rect 13032 46268 13096 46272
rect 13032 46212 13036 46268
rect 13036 46212 13092 46268
rect 13092 46212 13096 46268
rect 13032 46208 13096 46212
rect 13112 46268 13176 46272
rect 13112 46212 13116 46268
rect 13116 46212 13172 46268
rect 13172 46212 13176 46268
rect 13112 46208 13176 46212
rect 13192 46268 13256 46272
rect 13192 46212 13196 46268
rect 13196 46212 13252 46268
rect 13252 46212 13256 46268
rect 13192 46208 13256 46212
rect 22952 46268 23016 46272
rect 22952 46212 22956 46268
rect 22956 46212 23012 46268
rect 23012 46212 23016 46268
rect 22952 46208 23016 46212
rect 23032 46268 23096 46272
rect 23032 46212 23036 46268
rect 23036 46212 23092 46268
rect 23092 46212 23096 46268
rect 23032 46208 23096 46212
rect 23112 46268 23176 46272
rect 23112 46212 23116 46268
rect 23116 46212 23172 46268
rect 23172 46212 23176 46268
rect 23112 46208 23176 46212
rect 23192 46268 23256 46272
rect 23192 46212 23196 46268
rect 23196 46212 23252 46268
rect 23252 46212 23256 46268
rect 23192 46208 23256 46212
rect 20484 45792 20548 45796
rect 20484 45736 20534 45792
rect 20534 45736 20548 45792
rect 20484 45732 20548 45736
rect 7952 45724 8016 45728
rect 7952 45668 7956 45724
rect 7956 45668 8012 45724
rect 8012 45668 8016 45724
rect 7952 45664 8016 45668
rect 8032 45724 8096 45728
rect 8032 45668 8036 45724
rect 8036 45668 8092 45724
rect 8092 45668 8096 45724
rect 8032 45664 8096 45668
rect 8112 45724 8176 45728
rect 8112 45668 8116 45724
rect 8116 45668 8172 45724
rect 8172 45668 8176 45724
rect 8112 45664 8176 45668
rect 8192 45724 8256 45728
rect 8192 45668 8196 45724
rect 8196 45668 8252 45724
rect 8252 45668 8256 45724
rect 8192 45664 8256 45668
rect 17952 45724 18016 45728
rect 17952 45668 17956 45724
rect 17956 45668 18012 45724
rect 18012 45668 18016 45724
rect 17952 45664 18016 45668
rect 18032 45724 18096 45728
rect 18032 45668 18036 45724
rect 18036 45668 18092 45724
rect 18092 45668 18096 45724
rect 18032 45664 18096 45668
rect 18112 45724 18176 45728
rect 18112 45668 18116 45724
rect 18116 45668 18172 45724
rect 18172 45668 18176 45724
rect 18112 45664 18176 45668
rect 18192 45724 18256 45728
rect 18192 45668 18196 45724
rect 18196 45668 18252 45724
rect 18252 45668 18256 45724
rect 18192 45664 18256 45668
rect 21404 45520 21468 45524
rect 21404 45464 21454 45520
rect 21454 45464 21468 45520
rect 21404 45460 21468 45464
rect 12020 45188 12084 45252
rect 2952 45180 3016 45184
rect 2952 45124 2956 45180
rect 2956 45124 3012 45180
rect 3012 45124 3016 45180
rect 2952 45120 3016 45124
rect 3032 45180 3096 45184
rect 3032 45124 3036 45180
rect 3036 45124 3092 45180
rect 3092 45124 3096 45180
rect 3032 45120 3096 45124
rect 3112 45180 3176 45184
rect 3112 45124 3116 45180
rect 3116 45124 3172 45180
rect 3172 45124 3176 45180
rect 3112 45120 3176 45124
rect 3192 45180 3256 45184
rect 3192 45124 3196 45180
rect 3196 45124 3252 45180
rect 3252 45124 3256 45180
rect 3192 45120 3256 45124
rect 12952 45180 13016 45184
rect 12952 45124 12956 45180
rect 12956 45124 13012 45180
rect 13012 45124 13016 45180
rect 12952 45120 13016 45124
rect 13032 45180 13096 45184
rect 13032 45124 13036 45180
rect 13036 45124 13092 45180
rect 13092 45124 13096 45180
rect 13032 45120 13096 45124
rect 13112 45180 13176 45184
rect 13112 45124 13116 45180
rect 13116 45124 13172 45180
rect 13172 45124 13176 45180
rect 13112 45120 13176 45124
rect 13192 45180 13256 45184
rect 13192 45124 13196 45180
rect 13196 45124 13252 45180
rect 13252 45124 13256 45180
rect 13192 45120 13256 45124
rect 22952 45180 23016 45184
rect 22952 45124 22956 45180
rect 22956 45124 23012 45180
rect 23012 45124 23016 45180
rect 22952 45120 23016 45124
rect 23032 45180 23096 45184
rect 23032 45124 23036 45180
rect 23036 45124 23092 45180
rect 23092 45124 23096 45180
rect 23032 45120 23096 45124
rect 23112 45180 23176 45184
rect 23112 45124 23116 45180
rect 23116 45124 23172 45180
rect 23172 45124 23176 45180
rect 23112 45120 23176 45124
rect 23192 45180 23256 45184
rect 23192 45124 23196 45180
rect 23196 45124 23252 45180
rect 23252 45124 23256 45180
rect 23192 45120 23256 45124
rect 9812 44644 9876 44708
rect 7952 44636 8016 44640
rect 7952 44580 7956 44636
rect 7956 44580 8012 44636
rect 8012 44580 8016 44636
rect 7952 44576 8016 44580
rect 8032 44636 8096 44640
rect 8032 44580 8036 44636
rect 8036 44580 8092 44636
rect 8092 44580 8096 44636
rect 8032 44576 8096 44580
rect 8112 44636 8176 44640
rect 8112 44580 8116 44636
rect 8116 44580 8172 44636
rect 8172 44580 8176 44636
rect 8112 44576 8176 44580
rect 8192 44636 8256 44640
rect 8192 44580 8196 44636
rect 8196 44580 8252 44636
rect 8252 44580 8256 44636
rect 8192 44576 8256 44580
rect 17952 44636 18016 44640
rect 17952 44580 17956 44636
rect 17956 44580 18012 44636
rect 18012 44580 18016 44636
rect 17952 44576 18016 44580
rect 18032 44636 18096 44640
rect 18032 44580 18036 44636
rect 18036 44580 18092 44636
rect 18092 44580 18096 44636
rect 18032 44576 18096 44580
rect 18112 44636 18176 44640
rect 18112 44580 18116 44636
rect 18116 44580 18172 44636
rect 18172 44580 18176 44636
rect 18112 44576 18176 44580
rect 18192 44636 18256 44640
rect 18192 44580 18196 44636
rect 18196 44580 18252 44636
rect 18252 44580 18256 44636
rect 18192 44576 18256 44580
rect 19380 44236 19444 44300
rect 21036 44236 21100 44300
rect 2952 44092 3016 44096
rect 2952 44036 2956 44092
rect 2956 44036 3012 44092
rect 3012 44036 3016 44092
rect 2952 44032 3016 44036
rect 3032 44092 3096 44096
rect 3032 44036 3036 44092
rect 3036 44036 3092 44092
rect 3092 44036 3096 44092
rect 3032 44032 3096 44036
rect 3112 44092 3176 44096
rect 3112 44036 3116 44092
rect 3116 44036 3172 44092
rect 3172 44036 3176 44092
rect 3112 44032 3176 44036
rect 3192 44092 3256 44096
rect 3192 44036 3196 44092
rect 3196 44036 3252 44092
rect 3252 44036 3256 44092
rect 3192 44032 3256 44036
rect 12952 44092 13016 44096
rect 12952 44036 12956 44092
rect 12956 44036 13012 44092
rect 13012 44036 13016 44092
rect 12952 44032 13016 44036
rect 13032 44092 13096 44096
rect 13032 44036 13036 44092
rect 13036 44036 13092 44092
rect 13092 44036 13096 44092
rect 13032 44032 13096 44036
rect 13112 44092 13176 44096
rect 13112 44036 13116 44092
rect 13116 44036 13172 44092
rect 13172 44036 13176 44092
rect 13112 44032 13176 44036
rect 13192 44092 13256 44096
rect 13192 44036 13196 44092
rect 13196 44036 13252 44092
rect 13252 44036 13256 44092
rect 13192 44032 13256 44036
rect 22952 44092 23016 44096
rect 22952 44036 22956 44092
rect 22956 44036 23012 44092
rect 23012 44036 23016 44092
rect 22952 44032 23016 44036
rect 23032 44092 23096 44096
rect 23032 44036 23036 44092
rect 23036 44036 23092 44092
rect 23092 44036 23096 44092
rect 23032 44032 23096 44036
rect 23112 44092 23176 44096
rect 23112 44036 23116 44092
rect 23116 44036 23172 44092
rect 23172 44036 23176 44092
rect 23112 44032 23176 44036
rect 23192 44092 23256 44096
rect 23192 44036 23196 44092
rect 23196 44036 23252 44092
rect 23252 44036 23256 44092
rect 23192 44032 23256 44036
rect 7952 43548 8016 43552
rect 7952 43492 7956 43548
rect 7956 43492 8012 43548
rect 8012 43492 8016 43548
rect 7952 43488 8016 43492
rect 8032 43548 8096 43552
rect 8032 43492 8036 43548
rect 8036 43492 8092 43548
rect 8092 43492 8096 43548
rect 8032 43488 8096 43492
rect 8112 43548 8176 43552
rect 8112 43492 8116 43548
rect 8116 43492 8172 43548
rect 8172 43492 8176 43548
rect 8112 43488 8176 43492
rect 8192 43548 8256 43552
rect 8192 43492 8196 43548
rect 8196 43492 8252 43548
rect 8252 43492 8256 43548
rect 8192 43488 8256 43492
rect 17952 43548 18016 43552
rect 17952 43492 17956 43548
rect 17956 43492 18012 43548
rect 18012 43492 18016 43548
rect 17952 43488 18016 43492
rect 18032 43548 18096 43552
rect 18032 43492 18036 43548
rect 18036 43492 18092 43548
rect 18092 43492 18096 43548
rect 18032 43488 18096 43492
rect 18112 43548 18176 43552
rect 18112 43492 18116 43548
rect 18116 43492 18172 43548
rect 18172 43492 18176 43548
rect 18112 43488 18176 43492
rect 18192 43548 18256 43552
rect 18192 43492 18196 43548
rect 18196 43492 18252 43548
rect 18252 43492 18256 43548
rect 18192 43488 18256 43492
rect 2952 43004 3016 43008
rect 2952 42948 2956 43004
rect 2956 42948 3012 43004
rect 3012 42948 3016 43004
rect 2952 42944 3016 42948
rect 3032 43004 3096 43008
rect 3032 42948 3036 43004
rect 3036 42948 3092 43004
rect 3092 42948 3096 43004
rect 3032 42944 3096 42948
rect 3112 43004 3176 43008
rect 3112 42948 3116 43004
rect 3116 42948 3172 43004
rect 3172 42948 3176 43004
rect 3112 42944 3176 42948
rect 3192 43004 3256 43008
rect 3192 42948 3196 43004
rect 3196 42948 3252 43004
rect 3252 42948 3256 43004
rect 3192 42944 3256 42948
rect 12952 43004 13016 43008
rect 12952 42948 12956 43004
rect 12956 42948 13012 43004
rect 13012 42948 13016 43004
rect 12952 42944 13016 42948
rect 13032 43004 13096 43008
rect 13032 42948 13036 43004
rect 13036 42948 13092 43004
rect 13092 42948 13096 43004
rect 13032 42944 13096 42948
rect 13112 43004 13176 43008
rect 13112 42948 13116 43004
rect 13116 42948 13172 43004
rect 13172 42948 13176 43004
rect 13112 42944 13176 42948
rect 13192 43004 13256 43008
rect 13192 42948 13196 43004
rect 13196 42948 13252 43004
rect 13252 42948 13256 43004
rect 13192 42944 13256 42948
rect 22952 43004 23016 43008
rect 22952 42948 22956 43004
rect 22956 42948 23012 43004
rect 23012 42948 23016 43004
rect 22952 42944 23016 42948
rect 23032 43004 23096 43008
rect 23032 42948 23036 43004
rect 23036 42948 23092 43004
rect 23092 42948 23096 43004
rect 23032 42944 23096 42948
rect 23112 43004 23176 43008
rect 23112 42948 23116 43004
rect 23116 42948 23172 43004
rect 23172 42948 23176 43004
rect 23112 42944 23176 42948
rect 23192 43004 23256 43008
rect 23192 42948 23196 43004
rect 23196 42948 23252 43004
rect 23252 42948 23256 43004
rect 23192 42944 23256 42948
rect 7952 42460 8016 42464
rect 7952 42404 7956 42460
rect 7956 42404 8012 42460
rect 8012 42404 8016 42460
rect 7952 42400 8016 42404
rect 8032 42460 8096 42464
rect 8032 42404 8036 42460
rect 8036 42404 8092 42460
rect 8092 42404 8096 42460
rect 8032 42400 8096 42404
rect 8112 42460 8176 42464
rect 8112 42404 8116 42460
rect 8116 42404 8172 42460
rect 8172 42404 8176 42460
rect 8112 42400 8176 42404
rect 8192 42460 8256 42464
rect 8192 42404 8196 42460
rect 8196 42404 8252 42460
rect 8252 42404 8256 42460
rect 8192 42400 8256 42404
rect 17952 42460 18016 42464
rect 17952 42404 17956 42460
rect 17956 42404 18012 42460
rect 18012 42404 18016 42460
rect 17952 42400 18016 42404
rect 18032 42460 18096 42464
rect 18032 42404 18036 42460
rect 18036 42404 18092 42460
rect 18092 42404 18096 42460
rect 18032 42400 18096 42404
rect 18112 42460 18176 42464
rect 18112 42404 18116 42460
rect 18116 42404 18172 42460
rect 18172 42404 18176 42460
rect 18112 42400 18176 42404
rect 18192 42460 18256 42464
rect 18192 42404 18196 42460
rect 18196 42404 18252 42460
rect 18252 42404 18256 42460
rect 18192 42400 18256 42404
rect 2952 41916 3016 41920
rect 2952 41860 2956 41916
rect 2956 41860 3012 41916
rect 3012 41860 3016 41916
rect 2952 41856 3016 41860
rect 3032 41916 3096 41920
rect 3032 41860 3036 41916
rect 3036 41860 3092 41916
rect 3092 41860 3096 41916
rect 3032 41856 3096 41860
rect 3112 41916 3176 41920
rect 3112 41860 3116 41916
rect 3116 41860 3172 41916
rect 3172 41860 3176 41916
rect 3112 41856 3176 41860
rect 3192 41916 3256 41920
rect 3192 41860 3196 41916
rect 3196 41860 3252 41916
rect 3252 41860 3256 41916
rect 3192 41856 3256 41860
rect 12952 41916 13016 41920
rect 12952 41860 12956 41916
rect 12956 41860 13012 41916
rect 13012 41860 13016 41916
rect 12952 41856 13016 41860
rect 13032 41916 13096 41920
rect 13032 41860 13036 41916
rect 13036 41860 13092 41916
rect 13092 41860 13096 41916
rect 13032 41856 13096 41860
rect 13112 41916 13176 41920
rect 13112 41860 13116 41916
rect 13116 41860 13172 41916
rect 13172 41860 13176 41916
rect 13112 41856 13176 41860
rect 13192 41916 13256 41920
rect 13192 41860 13196 41916
rect 13196 41860 13252 41916
rect 13252 41860 13256 41916
rect 13192 41856 13256 41860
rect 22952 41916 23016 41920
rect 22952 41860 22956 41916
rect 22956 41860 23012 41916
rect 23012 41860 23016 41916
rect 22952 41856 23016 41860
rect 23032 41916 23096 41920
rect 23032 41860 23036 41916
rect 23036 41860 23092 41916
rect 23092 41860 23096 41916
rect 23032 41856 23096 41860
rect 23112 41916 23176 41920
rect 23112 41860 23116 41916
rect 23116 41860 23172 41916
rect 23172 41860 23176 41916
rect 23112 41856 23176 41860
rect 23192 41916 23256 41920
rect 23192 41860 23196 41916
rect 23196 41860 23252 41916
rect 23252 41860 23256 41916
rect 23192 41856 23256 41860
rect 21220 41440 21284 41444
rect 21220 41384 21234 41440
rect 21234 41384 21284 41440
rect 21220 41380 21284 41384
rect 7952 41372 8016 41376
rect 7952 41316 7956 41372
rect 7956 41316 8012 41372
rect 8012 41316 8016 41372
rect 7952 41312 8016 41316
rect 8032 41372 8096 41376
rect 8032 41316 8036 41372
rect 8036 41316 8092 41372
rect 8092 41316 8096 41372
rect 8032 41312 8096 41316
rect 8112 41372 8176 41376
rect 8112 41316 8116 41372
rect 8116 41316 8172 41372
rect 8172 41316 8176 41372
rect 8112 41312 8176 41316
rect 8192 41372 8256 41376
rect 8192 41316 8196 41372
rect 8196 41316 8252 41372
rect 8252 41316 8256 41372
rect 8192 41312 8256 41316
rect 17952 41372 18016 41376
rect 17952 41316 17956 41372
rect 17956 41316 18012 41372
rect 18012 41316 18016 41372
rect 17952 41312 18016 41316
rect 18032 41372 18096 41376
rect 18032 41316 18036 41372
rect 18036 41316 18092 41372
rect 18092 41316 18096 41372
rect 18032 41312 18096 41316
rect 18112 41372 18176 41376
rect 18112 41316 18116 41372
rect 18116 41316 18172 41372
rect 18172 41316 18176 41372
rect 18112 41312 18176 41316
rect 18192 41372 18256 41376
rect 18192 41316 18196 41372
rect 18196 41316 18252 41372
rect 18252 41316 18256 41372
rect 18192 41312 18256 41316
rect 13676 41244 13740 41308
rect 2952 40828 3016 40832
rect 2952 40772 2956 40828
rect 2956 40772 3012 40828
rect 3012 40772 3016 40828
rect 2952 40768 3016 40772
rect 3032 40828 3096 40832
rect 3032 40772 3036 40828
rect 3036 40772 3092 40828
rect 3092 40772 3096 40828
rect 3032 40768 3096 40772
rect 3112 40828 3176 40832
rect 3112 40772 3116 40828
rect 3116 40772 3172 40828
rect 3172 40772 3176 40828
rect 3112 40768 3176 40772
rect 3192 40828 3256 40832
rect 3192 40772 3196 40828
rect 3196 40772 3252 40828
rect 3252 40772 3256 40828
rect 3192 40768 3256 40772
rect 12952 40828 13016 40832
rect 12952 40772 12956 40828
rect 12956 40772 13012 40828
rect 13012 40772 13016 40828
rect 12952 40768 13016 40772
rect 13032 40828 13096 40832
rect 13032 40772 13036 40828
rect 13036 40772 13092 40828
rect 13092 40772 13096 40828
rect 13032 40768 13096 40772
rect 13112 40828 13176 40832
rect 13112 40772 13116 40828
rect 13116 40772 13172 40828
rect 13172 40772 13176 40828
rect 13112 40768 13176 40772
rect 13192 40828 13256 40832
rect 13192 40772 13196 40828
rect 13196 40772 13252 40828
rect 13252 40772 13256 40828
rect 13192 40768 13256 40772
rect 22952 40828 23016 40832
rect 22952 40772 22956 40828
rect 22956 40772 23012 40828
rect 23012 40772 23016 40828
rect 22952 40768 23016 40772
rect 23032 40828 23096 40832
rect 23032 40772 23036 40828
rect 23036 40772 23092 40828
rect 23092 40772 23096 40828
rect 23032 40768 23096 40772
rect 23112 40828 23176 40832
rect 23112 40772 23116 40828
rect 23116 40772 23172 40828
rect 23172 40772 23176 40828
rect 23112 40768 23176 40772
rect 23192 40828 23256 40832
rect 23192 40772 23196 40828
rect 23196 40772 23252 40828
rect 23252 40772 23256 40828
rect 23192 40768 23256 40772
rect 14596 40700 14660 40764
rect 7952 40284 8016 40288
rect 7952 40228 7956 40284
rect 7956 40228 8012 40284
rect 8012 40228 8016 40284
rect 7952 40224 8016 40228
rect 8032 40284 8096 40288
rect 8032 40228 8036 40284
rect 8036 40228 8092 40284
rect 8092 40228 8096 40284
rect 8032 40224 8096 40228
rect 8112 40284 8176 40288
rect 8112 40228 8116 40284
rect 8116 40228 8172 40284
rect 8172 40228 8176 40284
rect 8112 40224 8176 40228
rect 8192 40284 8256 40288
rect 8192 40228 8196 40284
rect 8196 40228 8252 40284
rect 8252 40228 8256 40284
rect 8192 40224 8256 40228
rect 17952 40284 18016 40288
rect 17952 40228 17956 40284
rect 17956 40228 18012 40284
rect 18012 40228 18016 40284
rect 17952 40224 18016 40228
rect 18032 40284 18096 40288
rect 18032 40228 18036 40284
rect 18036 40228 18092 40284
rect 18092 40228 18096 40284
rect 18032 40224 18096 40228
rect 18112 40284 18176 40288
rect 18112 40228 18116 40284
rect 18116 40228 18172 40284
rect 18172 40228 18176 40284
rect 18112 40224 18176 40228
rect 18192 40284 18256 40288
rect 18192 40228 18196 40284
rect 18196 40228 18252 40284
rect 18252 40228 18256 40284
rect 18192 40224 18256 40228
rect 2952 39740 3016 39744
rect 2952 39684 2956 39740
rect 2956 39684 3012 39740
rect 3012 39684 3016 39740
rect 2952 39680 3016 39684
rect 3032 39740 3096 39744
rect 3032 39684 3036 39740
rect 3036 39684 3092 39740
rect 3092 39684 3096 39740
rect 3032 39680 3096 39684
rect 3112 39740 3176 39744
rect 3112 39684 3116 39740
rect 3116 39684 3172 39740
rect 3172 39684 3176 39740
rect 3112 39680 3176 39684
rect 3192 39740 3256 39744
rect 3192 39684 3196 39740
rect 3196 39684 3252 39740
rect 3252 39684 3256 39740
rect 3192 39680 3256 39684
rect 12952 39740 13016 39744
rect 12952 39684 12956 39740
rect 12956 39684 13012 39740
rect 13012 39684 13016 39740
rect 12952 39680 13016 39684
rect 13032 39740 13096 39744
rect 13032 39684 13036 39740
rect 13036 39684 13092 39740
rect 13092 39684 13096 39740
rect 13032 39680 13096 39684
rect 13112 39740 13176 39744
rect 13112 39684 13116 39740
rect 13116 39684 13172 39740
rect 13172 39684 13176 39740
rect 13112 39680 13176 39684
rect 13192 39740 13256 39744
rect 13192 39684 13196 39740
rect 13196 39684 13252 39740
rect 13252 39684 13256 39740
rect 13192 39680 13256 39684
rect 22952 39740 23016 39744
rect 22952 39684 22956 39740
rect 22956 39684 23012 39740
rect 23012 39684 23016 39740
rect 22952 39680 23016 39684
rect 23032 39740 23096 39744
rect 23032 39684 23036 39740
rect 23036 39684 23092 39740
rect 23092 39684 23096 39740
rect 23032 39680 23096 39684
rect 23112 39740 23176 39744
rect 23112 39684 23116 39740
rect 23116 39684 23172 39740
rect 23172 39684 23176 39740
rect 23112 39680 23176 39684
rect 23192 39740 23256 39744
rect 23192 39684 23196 39740
rect 23196 39684 23252 39740
rect 23252 39684 23256 39740
rect 23192 39680 23256 39684
rect 7952 39196 8016 39200
rect 7952 39140 7956 39196
rect 7956 39140 8012 39196
rect 8012 39140 8016 39196
rect 7952 39136 8016 39140
rect 8032 39196 8096 39200
rect 8032 39140 8036 39196
rect 8036 39140 8092 39196
rect 8092 39140 8096 39196
rect 8032 39136 8096 39140
rect 8112 39196 8176 39200
rect 8112 39140 8116 39196
rect 8116 39140 8172 39196
rect 8172 39140 8176 39196
rect 8112 39136 8176 39140
rect 8192 39196 8256 39200
rect 8192 39140 8196 39196
rect 8196 39140 8252 39196
rect 8252 39140 8256 39196
rect 8192 39136 8256 39140
rect 17952 39196 18016 39200
rect 17952 39140 17956 39196
rect 17956 39140 18012 39196
rect 18012 39140 18016 39196
rect 17952 39136 18016 39140
rect 18032 39196 18096 39200
rect 18032 39140 18036 39196
rect 18036 39140 18092 39196
rect 18092 39140 18096 39196
rect 18032 39136 18096 39140
rect 18112 39196 18176 39200
rect 18112 39140 18116 39196
rect 18116 39140 18172 39196
rect 18172 39140 18176 39196
rect 18112 39136 18176 39140
rect 18192 39196 18256 39200
rect 18192 39140 18196 39196
rect 18196 39140 18252 39196
rect 18252 39140 18256 39196
rect 18192 39136 18256 39140
rect 17540 38932 17604 38996
rect 15148 38660 15212 38724
rect 18460 38720 18524 38724
rect 18460 38664 18474 38720
rect 18474 38664 18524 38720
rect 18460 38660 18524 38664
rect 2952 38652 3016 38656
rect 2952 38596 2956 38652
rect 2956 38596 3012 38652
rect 3012 38596 3016 38652
rect 2952 38592 3016 38596
rect 3032 38652 3096 38656
rect 3032 38596 3036 38652
rect 3036 38596 3092 38652
rect 3092 38596 3096 38652
rect 3032 38592 3096 38596
rect 3112 38652 3176 38656
rect 3112 38596 3116 38652
rect 3116 38596 3172 38652
rect 3172 38596 3176 38652
rect 3112 38592 3176 38596
rect 3192 38652 3256 38656
rect 3192 38596 3196 38652
rect 3196 38596 3252 38652
rect 3252 38596 3256 38652
rect 3192 38592 3256 38596
rect 12952 38652 13016 38656
rect 12952 38596 12956 38652
rect 12956 38596 13012 38652
rect 13012 38596 13016 38652
rect 12952 38592 13016 38596
rect 13032 38652 13096 38656
rect 13032 38596 13036 38652
rect 13036 38596 13092 38652
rect 13092 38596 13096 38652
rect 13032 38592 13096 38596
rect 13112 38652 13176 38656
rect 13112 38596 13116 38652
rect 13116 38596 13172 38652
rect 13172 38596 13176 38652
rect 13112 38592 13176 38596
rect 13192 38652 13256 38656
rect 13192 38596 13196 38652
rect 13196 38596 13252 38652
rect 13252 38596 13256 38652
rect 13192 38592 13256 38596
rect 22952 38652 23016 38656
rect 22952 38596 22956 38652
rect 22956 38596 23012 38652
rect 23012 38596 23016 38652
rect 22952 38592 23016 38596
rect 23032 38652 23096 38656
rect 23032 38596 23036 38652
rect 23036 38596 23092 38652
rect 23092 38596 23096 38652
rect 23032 38592 23096 38596
rect 23112 38652 23176 38656
rect 23112 38596 23116 38652
rect 23116 38596 23172 38652
rect 23172 38596 23176 38652
rect 23112 38592 23176 38596
rect 23192 38652 23256 38656
rect 23192 38596 23196 38652
rect 23196 38596 23252 38652
rect 23252 38596 23256 38652
rect 23192 38592 23256 38596
rect 7952 38108 8016 38112
rect 7952 38052 7956 38108
rect 7956 38052 8012 38108
rect 8012 38052 8016 38108
rect 7952 38048 8016 38052
rect 8032 38108 8096 38112
rect 8032 38052 8036 38108
rect 8036 38052 8092 38108
rect 8092 38052 8096 38108
rect 8032 38048 8096 38052
rect 8112 38108 8176 38112
rect 8112 38052 8116 38108
rect 8116 38052 8172 38108
rect 8172 38052 8176 38108
rect 8112 38048 8176 38052
rect 8192 38108 8256 38112
rect 8192 38052 8196 38108
rect 8196 38052 8252 38108
rect 8252 38052 8256 38108
rect 8192 38048 8256 38052
rect 17952 38108 18016 38112
rect 17952 38052 17956 38108
rect 17956 38052 18012 38108
rect 18012 38052 18016 38108
rect 17952 38048 18016 38052
rect 18032 38108 18096 38112
rect 18032 38052 18036 38108
rect 18036 38052 18092 38108
rect 18092 38052 18096 38108
rect 18032 38048 18096 38052
rect 18112 38108 18176 38112
rect 18112 38052 18116 38108
rect 18116 38052 18172 38108
rect 18172 38052 18176 38108
rect 18112 38048 18176 38052
rect 18192 38108 18256 38112
rect 18192 38052 18196 38108
rect 18196 38052 18252 38108
rect 18252 38052 18256 38108
rect 18192 38048 18256 38052
rect 18644 37572 18708 37636
rect 2952 37564 3016 37568
rect 2952 37508 2956 37564
rect 2956 37508 3012 37564
rect 3012 37508 3016 37564
rect 2952 37504 3016 37508
rect 3032 37564 3096 37568
rect 3032 37508 3036 37564
rect 3036 37508 3092 37564
rect 3092 37508 3096 37564
rect 3032 37504 3096 37508
rect 3112 37564 3176 37568
rect 3112 37508 3116 37564
rect 3116 37508 3172 37564
rect 3172 37508 3176 37564
rect 3112 37504 3176 37508
rect 3192 37564 3256 37568
rect 3192 37508 3196 37564
rect 3196 37508 3252 37564
rect 3252 37508 3256 37564
rect 3192 37504 3256 37508
rect 12952 37564 13016 37568
rect 12952 37508 12956 37564
rect 12956 37508 13012 37564
rect 13012 37508 13016 37564
rect 12952 37504 13016 37508
rect 13032 37564 13096 37568
rect 13032 37508 13036 37564
rect 13036 37508 13092 37564
rect 13092 37508 13096 37564
rect 13032 37504 13096 37508
rect 13112 37564 13176 37568
rect 13112 37508 13116 37564
rect 13116 37508 13172 37564
rect 13172 37508 13176 37564
rect 13112 37504 13176 37508
rect 13192 37564 13256 37568
rect 13192 37508 13196 37564
rect 13196 37508 13252 37564
rect 13252 37508 13256 37564
rect 13192 37504 13256 37508
rect 22952 37564 23016 37568
rect 22952 37508 22956 37564
rect 22956 37508 23012 37564
rect 23012 37508 23016 37564
rect 22952 37504 23016 37508
rect 23032 37564 23096 37568
rect 23032 37508 23036 37564
rect 23036 37508 23092 37564
rect 23092 37508 23096 37564
rect 23032 37504 23096 37508
rect 23112 37564 23176 37568
rect 23112 37508 23116 37564
rect 23116 37508 23172 37564
rect 23172 37508 23176 37564
rect 23112 37504 23176 37508
rect 23192 37564 23256 37568
rect 23192 37508 23196 37564
rect 23196 37508 23252 37564
rect 23252 37508 23256 37564
rect 23192 37504 23256 37508
rect 17724 37360 17788 37364
rect 17724 37304 17774 37360
rect 17774 37304 17788 37360
rect 17724 37300 17788 37304
rect 19748 37164 19812 37228
rect 7952 37020 8016 37024
rect 7952 36964 7956 37020
rect 7956 36964 8012 37020
rect 8012 36964 8016 37020
rect 7952 36960 8016 36964
rect 8032 37020 8096 37024
rect 8032 36964 8036 37020
rect 8036 36964 8092 37020
rect 8092 36964 8096 37020
rect 8032 36960 8096 36964
rect 8112 37020 8176 37024
rect 8112 36964 8116 37020
rect 8116 36964 8172 37020
rect 8172 36964 8176 37020
rect 8112 36960 8176 36964
rect 8192 37020 8256 37024
rect 8192 36964 8196 37020
rect 8196 36964 8252 37020
rect 8252 36964 8256 37020
rect 8192 36960 8256 36964
rect 17952 37020 18016 37024
rect 17952 36964 17956 37020
rect 17956 36964 18012 37020
rect 18012 36964 18016 37020
rect 17952 36960 18016 36964
rect 18032 37020 18096 37024
rect 18032 36964 18036 37020
rect 18036 36964 18092 37020
rect 18092 36964 18096 37020
rect 18032 36960 18096 36964
rect 18112 37020 18176 37024
rect 18112 36964 18116 37020
rect 18116 36964 18172 37020
rect 18172 36964 18176 37020
rect 18112 36960 18176 36964
rect 18192 37020 18256 37024
rect 18192 36964 18196 37020
rect 18196 36964 18252 37020
rect 18252 36964 18256 37020
rect 18192 36960 18256 36964
rect 12020 36620 12084 36684
rect 2952 36476 3016 36480
rect 2952 36420 2956 36476
rect 2956 36420 3012 36476
rect 3012 36420 3016 36476
rect 2952 36416 3016 36420
rect 3032 36476 3096 36480
rect 3032 36420 3036 36476
rect 3036 36420 3092 36476
rect 3092 36420 3096 36476
rect 3032 36416 3096 36420
rect 3112 36476 3176 36480
rect 3112 36420 3116 36476
rect 3116 36420 3172 36476
rect 3172 36420 3176 36476
rect 3112 36416 3176 36420
rect 3192 36476 3256 36480
rect 3192 36420 3196 36476
rect 3196 36420 3252 36476
rect 3252 36420 3256 36476
rect 3192 36416 3256 36420
rect 12952 36476 13016 36480
rect 12952 36420 12956 36476
rect 12956 36420 13012 36476
rect 13012 36420 13016 36476
rect 12952 36416 13016 36420
rect 13032 36476 13096 36480
rect 13032 36420 13036 36476
rect 13036 36420 13092 36476
rect 13092 36420 13096 36476
rect 13032 36416 13096 36420
rect 13112 36476 13176 36480
rect 13112 36420 13116 36476
rect 13116 36420 13172 36476
rect 13172 36420 13176 36476
rect 13112 36416 13176 36420
rect 13192 36476 13256 36480
rect 13192 36420 13196 36476
rect 13196 36420 13252 36476
rect 13252 36420 13256 36476
rect 13192 36416 13256 36420
rect 22952 36476 23016 36480
rect 22952 36420 22956 36476
rect 22956 36420 23012 36476
rect 23012 36420 23016 36476
rect 22952 36416 23016 36420
rect 23032 36476 23096 36480
rect 23032 36420 23036 36476
rect 23036 36420 23092 36476
rect 23092 36420 23096 36476
rect 23032 36416 23096 36420
rect 23112 36476 23176 36480
rect 23112 36420 23116 36476
rect 23116 36420 23172 36476
rect 23172 36420 23176 36476
rect 23112 36416 23176 36420
rect 23192 36476 23256 36480
rect 23192 36420 23196 36476
rect 23196 36420 23252 36476
rect 23252 36420 23256 36476
rect 23192 36416 23256 36420
rect 7952 35932 8016 35936
rect 7952 35876 7956 35932
rect 7956 35876 8012 35932
rect 8012 35876 8016 35932
rect 7952 35872 8016 35876
rect 8032 35932 8096 35936
rect 8032 35876 8036 35932
rect 8036 35876 8092 35932
rect 8092 35876 8096 35932
rect 8032 35872 8096 35876
rect 8112 35932 8176 35936
rect 8112 35876 8116 35932
rect 8116 35876 8172 35932
rect 8172 35876 8176 35932
rect 8112 35872 8176 35876
rect 8192 35932 8256 35936
rect 8192 35876 8196 35932
rect 8196 35876 8252 35932
rect 8252 35876 8256 35932
rect 8192 35872 8256 35876
rect 17952 35932 18016 35936
rect 17952 35876 17956 35932
rect 17956 35876 18012 35932
rect 18012 35876 18016 35932
rect 17952 35872 18016 35876
rect 18032 35932 18096 35936
rect 18032 35876 18036 35932
rect 18036 35876 18092 35932
rect 18092 35876 18096 35932
rect 18032 35872 18096 35876
rect 18112 35932 18176 35936
rect 18112 35876 18116 35932
rect 18116 35876 18172 35932
rect 18172 35876 18176 35932
rect 18112 35872 18176 35876
rect 18192 35932 18256 35936
rect 18192 35876 18196 35932
rect 18196 35876 18252 35932
rect 18252 35876 18256 35932
rect 18192 35872 18256 35876
rect 2952 35388 3016 35392
rect 2952 35332 2956 35388
rect 2956 35332 3012 35388
rect 3012 35332 3016 35388
rect 2952 35328 3016 35332
rect 3032 35388 3096 35392
rect 3032 35332 3036 35388
rect 3036 35332 3092 35388
rect 3092 35332 3096 35388
rect 3032 35328 3096 35332
rect 3112 35388 3176 35392
rect 3112 35332 3116 35388
rect 3116 35332 3172 35388
rect 3172 35332 3176 35388
rect 3112 35328 3176 35332
rect 3192 35388 3256 35392
rect 3192 35332 3196 35388
rect 3196 35332 3252 35388
rect 3252 35332 3256 35388
rect 3192 35328 3256 35332
rect 12952 35388 13016 35392
rect 12952 35332 12956 35388
rect 12956 35332 13012 35388
rect 13012 35332 13016 35388
rect 12952 35328 13016 35332
rect 13032 35388 13096 35392
rect 13032 35332 13036 35388
rect 13036 35332 13092 35388
rect 13092 35332 13096 35388
rect 13032 35328 13096 35332
rect 13112 35388 13176 35392
rect 13112 35332 13116 35388
rect 13116 35332 13172 35388
rect 13172 35332 13176 35388
rect 13112 35328 13176 35332
rect 13192 35388 13256 35392
rect 13192 35332 13196 35388
rect 13196 35332 13252 35388
rect 13252 35332 13256 35388
rect 13192 35328 13256 35332
rect 22952 35388 23016 35392
rect 22952 35332 22956 35388
rect 22956 35332 23012 35388
rect 23012 35332 23016 35388
rect 22952 35328 23016 35332
rect 23032 35388 23096 35392
rect 23032 35332 23036 35388
rect 23036 35332 23092 35388
rect 23092 35332 23096 35388
rect 23032 35328 23096 35332
rect 23112 35388 23176 35392
rect 23112 35332 23116 35388
rect 23116 35332 23172 35388
rect 23172 35332 23176 35388
rect 23112 35328 23176 35332
rect 23192 35388 23256 35392
rect 23192 35332 23196 35388
rect 23196 35332 23252 35388
rect 23252 35332 23256 35388
rect 23192 35328 23256 35332
rect 13676 35260 13740 35324
rect 22508 35124 22572 35188
rect 7952 34844 8016 34848
rect 7952 34788 7956 34844
rect 7956 34788 8012 34844
rect 8012 34788 8016 34844
rect 7952 34784 8016 34788
rect 8032 34844 8096 34848
rect 8032 34788 8036 34844
rect 8036 34788 8092 34844
rect 8092 34788 8096 34844
rect 8032 34784 8096 34788
rect 8112 34844 8176 34848
rect 8112 34788 8116 34844
rect 8116 34788 8172 34844
rect 8172 34788 8176 34844
rect 8112 34784 8176 34788
rect 8192 34844 8256 34848
rect 8192 34788 8196 34844
rect 8196 34788 8252 34844
rect 8252 34788 8256 34844
rect 8192 34784 8256 34788
rect 17952 34844 18016 34848
rect 17952 34788 17956 34844
rect 17956 34788 18012 34844
rect 18012 34788 18016 34844
rect 17952 34784 18016 34788
rect 18032 34844 18096 34848
rect 18032 34788 18036 34844
rect 18036 34788 18092 34844
rect 18092 34788 18096 34844
rect 18032 34784 18096 34788
rect 18112 34844 18176 34848
rect 18112 34788 18116 34844
rect 18116 34788 18172 34844
rect 18172 34788 18176 34844
rect 18112 34784 18176 34788
rect 18192 34844 18256 34848
rect 18192 34788 18196 34844
rect 18196 34788 18252 34844
rect 18252 34788 18256 34844
rect 18192 34784 18256 34788
rect 15148 34444 15212 34508
rect 2952 34300 3016 34304
rect 2952 34244 2956 34300
rect 2956 34244 3012 34300
rect 3012 34244 3016 34300
rect 2952 34240 3016 34244
rect 3032 34300 3096 34304
rect 3032 34244 3036 34300
rect 3036 34244 3092 34300
rect 3092 34244 3096 34300
rect 3032 34240 3096 34244
rect 3112 34300 3176 34304
rect 3112 34244 3116 34300
rect 3116 34244 3172 34300
rect 3172 34244 3176 34300
rect 3112 34240 3176 34244
rect 3192 34300 3256 34304
rect 3192 34244 3196 34300
rect 3196 34244 3252 34300
rect 3252 34244 3256 34300
rect 3192 34240 3256 34244
rect 12952 34300 13016 34304
rect 12952 34244 12956 34300
rect 12956 34244 13012 34300
rect 13012 34244 13016 34300
rect 12952 34240 13016 34244
rect 13032 34300 13096 34304
rect 13032 34244 13036 34300
rect 13036 34244 13092 34300
rect 13092 34244 13096 34300
rect 13032 34240 13096 34244
rect 13112 34300 13176 34304
rect 13112 34244 13116 34300
rect 13116 34244 13172 34300
rect 13172 34244 13176 34300
rect 13112 34240 13176 34244
rect 13192 34300 13256 34304
rect 13192 34244 13196 34300
rect 13196 34244 13252 34300
rect 13252 34244 13256 34300
rect 13192 34240 13256 34244
rect 22952 34300 23016 34304
rect 22952 34244 22956 34300
rect 22956 34244 23012 34300
rect 23012 34244 23016 34300
rect 22952 34240 23016 34244
rect 23032 34300 23096 34304
rect 23032 34244 23036 34300
rect 23036 34244 23092 34300
rect 23092 34244 23096 34300
rect 23032 34240 23096 34244
rect 23112 34300 23176 34304
rect 23112 34244 23116 34300
rect 23116 34244 23172 34300
rect 23172 34244 23176 34300
rect 23112 34240 23176 34244
rect 23192 34300 23256 34304
rect 23192 34244 23196 34300
rect 23196 34244 23252 34300
rect 23252 34244 23256 34300
rect 23192 34240 23256 34244
rect 7952 33756 8016 33760
rect 7952 33700 7956 33756
rect 7956 33700 8012 33756
rect 8012 33700 8016 33756
rect 7952 33696 8016 33700
rect 8032 33756 8096 33760
rect 8032 33700 8036 33756
rect 8036 33700 8092 33756
rect 8092 33700 8096 33756
rect 8032 33696 8096 33700
rect 8112 33756 8176 33760
rect 8112 33700 8116 33756
rect 8116 33700 8172 33756
rect 8172 33700 8176 33756
rect 8112 33696 8176 33700
rect 8192 33756 8256 33760
rect 8192 33700 8196 33756
rect 8196 33700 8252 33756
rect 8252 33700 8256 33756
rect 8192 33696 8256 33700
rect 17952 33756 18016 33760
rect 17952 33700 17956 33756
rect 17956 33700 18012 33756
rect 18012 33700 18016 33756
rect 17952 33696 18016 33700
rect 18032 33756 18096 33760
rect 18032 33700 18036 33756
rect 18036 33700 18092 33756
rect 18092 33700 18096 33756
rect 18032 33696 18096 33700
rect 18112 33756 18176 33760
rect 18112 33700 18116 33756
rect 18116 33700 18172 33756
rect 18172 33700 18176 33756
rect 18112 33696 18176 33700
rect 18192 33756 18256 33760
rect 18192 33700 18196 33756
rect 18196 33700 18252 33756
rect 18252 33700 18256 33756
rect 18192 33696 18256 33700
rect 12020 33688 12084 33692
rect 12020 33632 12070 33688
rect 12070 33632 12084 33688
rect 12020 33628 12084 33632
rect 13860 33492 13924 33556
rect 17540 33356 17604 33420
rect 2952 33212 3016 33216
rect 2952 33156 2956 33212
rect 2956 33156 3012 33212
rect 3012 33156 3016 33212
rect 2952 33152 3016 33156
rect 3032 33212 3096 33216
rect 3032 33156 3036 33212
rect 3036 33156 3092 33212
rect 3092 33156 3096 33212
rect 3032 33152 3096 33156
rect 3112 33212 3176 33216
rect 3112 33156 3116 33212
rect 3116 33156 3172 33212
rect 3172 33156 3176 33212
rect 3112 33152 3176 33156
rect 3192 33212 3256 33216
rect 3192 33156 3196 33212
rect 3196 33156 3252 33212
rect 3252 33156 3256 33212
rect 3192 33152 3256 33156
rect 12952 33212 13016 33216
rect 12952 33156 12956 33212
rect 12956 33156 13012 33212
rect 13012 33156 13016 33212
rect 12952 33152 13016 33156
rect 13032 33212 13096 33216
rect 13032 33156 13036 33212
rect 13036 33156 13092 33212
rect 13092 33156 13096 33212
rect 13032 33152 13096 33156
rect 13112 33212 13176 33216
rect 13112 33156 13116 33212
rect 13116 33156 13172 33212
rect 13172 33156 13176 33212
rect 13112 33152 13176 33156
rect 13192 33212 13256 33216
rect 13192 33156 13196 33212
rect 13196 33156 13252 33212
rect 13252 33156 13256 33212
rect 13192 33152 13256 33156
rect 22952 33212 23016 33216
rect 22952 33156 22956 33212
rect 22956 33156 23012 33212
rect 23012 33156 23016 33212
rect 22952 33152 23016 33156
rect 23032 33212 23096 33216
rect 23032 33156 23036 33212
rect 23036 33156 23092 33212
rect 23092 33156 23096 33212
rect 23032 33152 23096 33156
rect 23112 33212 23176 33216
rect 23112 33156 23116 33212
rect 23116 33156 23172 33212
rect 23172 33156 23176 33212
rect 23112 33152 23176 33156
rect 23192 33212 23256 33216
rect 23192 33156 23196 33212
rect 23196 33156 23252 33212
rect 23252 33156 23256 33212
rect 23192 33152 23256 33156
rect 7952 32668 8016 32672
rect 7952 32612 7956 32668
rect 7956 32612 8012 32668
rect 8012 32612 8016 32668
rect 7952 32608 8016 32612
rect 8032 32668 8096 32672
rect 8032 32612 8036 32668
rect 8036 32612 8092 32668
rect 8092 32612 8096 32668
rect 8032 32608 8096 32612
rect 8112 32668 8176 32672
rect 8112 32612 8116 32668
rect 8116 32612 8172 32668
rect 8172 32612 8176 32668
rect 8112 32608 8176 32612
rect 8192 32668 8256 32672
rect 8192 32612 8196 32668
rect 8196 32612 8252 32668
rect 8252 32612 8256 32668
rect 8192 32608 8256 32612
rect 17952 32668 18016 32672
rect 17952 32612 17956 32668
rect 17956 32612 18012 32668
rect 18012 32612 18016 32668
rect 17952 32608 18016 32612
rect 18032 32668 18096 32672
rect 18032 32612 18036 32668
rect 18036 32612 18092 32668
rect 18092 32612 18096 32668
rect 18032 32608 18096 32612
rect 18112 32668 18176 32672
rect 18112 32612 18116 32668
rect 18116 32612 18172 32668
rect 18172 32612 18176 32668
rect 18112 32608 18176 32612
rect 18192 32668 18256 32672
rect 18192 32612 18196 32668
rect 18196 32612 18252 32668
rect 18252 32612 18256 32668
rect 18192 32608 18256 32612
rect 2952 32124 3016 32128
rect 2952 32068 2956 32124
rect 2956 32068 3012 32124
rect 3012 32068 3016 32124
rect 2952 32064 3016 32068
rect 3032 32124 3096 32128
rect 3032 32068 3036 32124
rect 3036 32068 3092 32124
rect 3092 32068 3096 32124
rect 3032 32064 3096 32068
rect 3112 32124 3176 32128
rect 3112 32068 3116 32124
rect 3116 32068 3172 32124
rect 3172 32068 3176 32124
rect 3112 32064 3176 32068
rect 3192 32124 3256 32128
rect 3192 32068 3196 32124
rect 3196 32068 3252 32124
rect 3252 32068 3256 32124
rect 3192 32064 3256 32068
rect 12952 32124 13016 32128
rect 12952 32068 12956 32124
rect 12956 32068 13012 32124
rect 13012 32068 13016 32124
rect 12952 32064 13016 32068
rect 13032 32124 13096 32128
rect 13032 32068 13036 32124
rect 13036 32068 13092 32124
rect 13092 32068 13096 32124
rect 13032 32064 13096 32068
rect 13112 32124 13176 32128
rect 13112 32068 13116 32124
rect 13116 32068 13172 32124
rect 13172 32068 13176 32124
rect 13112 32064 13176 32068
rect 13192 32124 13256 32128
rect 13192 32068 13196 32124
rect 13196 32068 13252 32124
rect 13252 32068 13256 32124
rect 13192 32064 13256 32068
rect 22952 32124 23016 32128
rect 22952 32068 22956 32124
rect 22956 32068 23012 32124
rect 23012 32068 23016 32124
rect 22952 32064 23016 32068
rect 23032 32124 23096 32128
rect 23032 32068 23036 32124
rect 23036 32068 23092 32124
rect 23092 32068 23096 32124
rect 23032 32064 23096 32068
rect 23112 32124 23176 32128
rect 23112 32068 23116 32124
rect 23116 32068 23172 32124
rect 23172 32068 23176 32124
rect 23112 32064 23176 32068
rect 23192 32124 23256 32128
rect 23192 32068 23196 32124
rect 23196 32068 23252 32124
rect 23252 32068 23256 32124
rect 23192 32064 23256 32068
rect 14412 31860 14476 31924
rect 22324 31724 22388 31788
rect 7952 31580 8016 31584
rect 7952 31524 7956 31580
rect 7956 31524 8012 31580
rect 8012 31524 8016 31580
rect 7952 31520 8016 31524
rect 8032 31580 8096 31584
rect 8032 31524 8036 31580
rect 8036 31524 8092 31580
rect 8092 31524 8096 31580
rect 8032 31520 8096 31524
rect 8112 31580 8176 31584
rect 8112 31524 8116 31580
rect 8116 31524 8172 31580
rect 8172 31524 8176 31580
rect 8112 31520 8176 31524
rect 8192 31580 8256 31584
rect 8192 31524 8196 31580
rect 8196 31524 8252 31580
rect 8252 31524 8256 31580
rect 8192 31520 8256 31524
rect 17952 31580 18016 31584
rect 17952 31524 17956 31580
rect 17956 31524 18012 31580
rect 18012 31524 18016 31580
rect 17952 31520 18016 31524
rect 18032 31580 18096 31584
rect 18032 31524 18036 31580
rect 18036 31524 18092 31580
rect 18092 31524 18096 31580
rect 18032 31520 18096 31524
rect 18112 31580 18176 31584
rect 18112 31524 18116 31580
rect 18116 31524 18172 31580
rect 18172 31524 18176 31580
rect 18112 31520 18176 31524
rect 18192 31580 18256 31584
rect 18192 31524 18196 31580
rect 18196 31524 18252 31580
rect 18252 31524 18256 31580
rect 18192 31520 18256 31524
rect 9812 31376 9876 31380
rect 9812 31320 9862 31376
rect 9862 31320 9876 31376
rect 9812 31316 9876 31320
rect 2952 31036 3016 31040
rect 2952 30980 2956 31036
rect 2956 30980 3012 31036
rect 3012 30980 3016 31036
rect 2952 30976 3016 30980
rect 3032 31036 3096 31040
rect 3032 30980 3036 31036
rect 3036 30980 3092 31036
rect 3092 30980 3096 31036
rect 3032 30976 3096 30980
rect 3112 31036 3176 31040
rect 3112 30980 3116 31036
rect 3116 30980 3172 31036
rect 3172 30980 3176 31036
rect 3112 30976 3176 30980
rect 3192 31036 3256 31040
rect 3192 30980 3196 31036
rect 3196 30980 3252 31036
rect 3252 30980 3256 31036
rect 3192 30976 3256 30980
rect 12952 31036 13016 31040
rect 12952 30980 12956 31036
rect 12956 30980 13012 31036
rect 13012 30980 13016 31036
rect 12952 30976 13016 30980
rect 13032 31036 13096 31040
rect 13032 30980 13036 31036
rect 13036 30980 13092 31036
rect 13092 30980 13096 31036
rect 13032 30976 13096 30980
rect 13112 31036 13176 31040
rect 13112 30980 13116 31036
rect 13116 30980 13172 31036
rect 13172 30980 13176 31036
rect 13112 30976 13176 30980
rect 13192 31036 13256 31040
rect 13192 30980 13196 31036
rect 13196 30980 13252 31036
rect 13252 30980 13256 31036
rect 13192 30976 13256 30980
rect 22952 31036 23016 31040
rect 22952 30980 22956 31036
rect 22956 30980 23012 31036
rect 23012 30980 23016 31036
rect 22952 30976 23016 30980
rect 23032 31036 23096 31040
rect 23032 30980 23036 31036
rect 23036 30980 23092 31036
rect 23092 30980 23096 31036
rect 23032 30976 23096 30980
rect 23112 31036 23176 31040
rect 23112 30980 23116 31036
rect 23116 30980 23172 31036
rect 23172 30980 23176 31036
rect 23112 30976 23176 30980
rect 23192 31036 23256 31040
rect 23192 30980 23196 31036
rect 23196 30980 23252 31036
rect 23252 30980 23256 31036
rect 23192 30976 23256 30980
rect 18460 30772 18524 30836
rect 13860 30636 13924 30700
rect 20484 30636 20548 30700
rect 7952 30492 8016 30496
rect 7952 30436 7956 30492
rect 7956 30436 8012 30492
rect 8012 30436 8016 30492
rect 7952 30432 8016 30436
rect 8032 30492 8096 30496
rect 8032 30436 8036 30492
rect 8036 30436 8092 30492
rect 8092 30436 8096 30492
rect 8032 30432 8096 30436
rect 8112 30492 8176 30496
rect 8112 30436 8116 30492
rect 8116 30436 8172 30492
rect 8172 30436 8176 30492
rect 8112 30432 8176 30436
rect 8192 30492 8256 30496
rect 8192 30436 8196 30492
rect 8196 30436 8252 30492
rect 8252 30436 8256 30492
rect 8192 30432 8256 30436
rect 17952 30492 18016 30496
rect 17952 30436 17956 30492
rect 17956 30436 18012 30492
rect 18012 30436 18016 30492
rect 17952 30432 18016 30436
rect 18032 30492 18096 30496
rect 18032 30436 18036 30492
rect 18036 30436 18092 30492
rect 18092 30436 18096 30492
rect 18032 30432 18096 30436
rect 18112 30492 18176 30496
rect 18112 30436 18116 30492
rect 18116 30436 18172 30492
rect 18172 30436 18176 30492
rect 18112 30432 18176 30436
rect 18192 30492 18256 30496
rect 18192 30436 18196 30492
rect 18196 30436 18252 30492
rect 18252 30436 18256 30492
rect 18192 30432 18256 30436
rect 17724 30364 17788 30428
rect 14596 30228 14660 30292
rect 19564 30092 19628 30156
rect 16252 29956 16316 30020
rect 2952 29948 3016 29952
rect 2952 29892 2956 29948
rect 2956 29892 3012 29948
rect 3012 29892 3016 29948
rect 2952 29888 3016 29892
rect 3032 29948 3096 29952
rect 3032 29892 3036 29948
rect 3036 29892 3092 29948
rect 3092 29892 3096 29948
rect 3032 29888 3096 29892
rect 3112 29948 3176 29952
rect 3112 29892 3116 29948
rect 3116 29892 3172 29948
rect 3172 29892 3176 29948
rect 3112 29888 3176 29892
rect 3192 29948 3256 29952
rect 3192 29892 3196 29948
rect 3196 29892 3252 29948
rect 3252 29892 3256 29948
rect 3192 29888 3256 29892
rect 12952 29948 13016 29952
rect 12952 29892 12956 29948
rect 12956 29892 13012 29948
rect 13012 29892 13016 29948
rect 12952 29888 13016 29892
rect 13032 29948 13096 29952
rect 13032 29892 13036 29948
rect 13036 29892 13092 29948
rect 13092 29892 13096 29948
rect 13032 29888 13096 29892
rect 13112 29948 13176 29952
rect 13112 29892 13116 29948
rect 13116 29892 13172 29948
rect 13172 29892 13176 29948
rect 13112 29888 13176 29892
rect 13192 29948 13256 29952
rect 13192 29892 13196 29948
rect 13196 29892 13252 29948
rect 13252 29892 13256 29948
rect 13192 29888 13256 29892
rect 22952 29948 23016 29952
rect 22952 29892 22956 29948
rect 22956 29892 23012 29948
rect 23012 29892 23016 29948
rect 22952 29888 23016 29892
rect 23032 29948 23096 29952
rect 23032 29892 23036 29948
rect 23036 29892 23092 29948
rect 23092 29892 23096 29948
rect 23032 29888 23096 29892
rect 23112 29948 23176 29952
rect 23112 29892 23116 29948
rect 23116 29892 23172 29948
rect 23172 29892 23176 29948
rect 23112 29888 23176 29892
rect 23192 29948 23256 29952
rect 23192 29892 23196 29948
rect 23196 29892 23252 29948
rect 23252 29892 23256 29948
rect 23192 29888 23256 29892
rect 17724 29684 17788 29748
rect 19380 29684 19444 29748
rect 19748 29684 19812 29748
rect 22508 29684 22572 29748
rect 12756 29412 12820 29476
rect 23428 29412 23492 29476
rect 7952 29404 8016 29408
rect 7952 29348 7956 29404
rect 7956 29348 8012 29404
rect 8012 29348 8016 29404
rect 7952 29344 8016 29348
rect 8032 29404 8096 29408
rect 8032 29348 8036 29404
rect 8036 29348 8092 29404
rect 8092 29348 8096 29404
rect 8032 29344 8096 29348
rect 8112 29404 8176 29408
rect 8112 29348 8116 29404
rect 8116 29348 8172 29404
rect 8172 29348 8176 29404
rect 8112 29344 8176 29348
rect 8192 29404 8256 29408
rect 8192 29348 8196 29404
rect 8196 29348 8252 29404
rect 8252 29348 8256 29404
rect 8192 29344 8256 29348
rect 17952 29404 18016 29408
rect 17952 29348 17956 29404
rect 17956 29348 18012 29404
rect 18012 29348 18016 29404
rect 17952 29344 18016 29348
rect 18032 29404 18096 29408
rect 18032 29348 18036 29404
rect 18036 29348 18092 29404
rect 18092 29348 18096 29404
rect 18032 29344 18096 29348
rect 18112 29404 18176 29408
rect 18112 29348 18116 29404
rect 18116 29348 18172 29404
rect 18172 29348 18176 29404
rect 18112 29344 18176 29348
rect 18192 29404 18256 29408
rect 18192 29348 18196 29404
rect 18196 29348 18252 29404
rect 18252 29348 18256 29404
rect 18192 29344 18256 29348
rect 14596 29004 14660 29068
rect 16804 29064 16868 29068
rect 16804 29008 16818 29064
rect 16818 29008 16868 29064
rect 16804 29004 16868 29008
rect 17540 29064 17604 29068
rect 17540 29008 17554 29064
rect 17554 29008 17604 29064
rect 17540 29004 17604 29008
rect 2952 28860 3016 28864
rect 2952 28804 2956 28860
rect 2956 28804 3012 28860
rect 3012 28804 3016 28860
rect 2952 28800 3016 28804
rect 3032 28860 3096 28864
rect 3032 28804 3036 28860
rect 3036 28804 3092 28860
rect 3092 28804 3096 28860
rect 3032 28800 3096 28804
rect 3112 28860 3176 28864
rect 3112 28804 3116 28860
rect 3116 28804 3172 28860
rect 3172 28804 3176 28860
rect 3112 28800 3176 28804
rect 3192 28860 3256 28864
rect 3192 28804 3196 28860
rect 3196 28804 3252 28860
rect 3252 28804 3256 28860
rect 3192 28800 3256 28804
rect 12952 28860 13016 28864
rect 12952 28804 12956 28860
rect 12956 28804 13012 28860
rect 13012 28804 13016 28860
rect 12952 28800 13016 28804
rect 13032 28860 13096 28864
rect 13032 28804 13036 28860
rect 13036 28804 13092 28860
rect 13092 28804 13096 28860
rect 13032 28800 13096 28804
rect 13112 28860 13176 28864
rect 13112 28804 13116 28860
rect 13116 28804 13172 28860
rect 13172 28804 13176 28860
rect 13112 28800 13176 28804
rect 13192 28860 13256 28864
rect 13192 28804 13196 28860
rect 13196 28804 13252 28860
rect 13252 28804 13256 28860
rect 13192 28800 13256 28804
rect 22952 28860 23016 28864
rect 22952 28804 22956 28860
rect 22956 28804 23012 28860
rect 23012 28804 23016 28860
rect 22952 28800 23016 28804
rect 23032 28860 23096 28864
rect 23032 28804 23036 28860
rect 23036 28804 23092 28860
rect 23092 28804 23096 28860
rect 23032 28800 23096 28804
rect 23112 28860 23176 28864
rect 23112 28804 23116 28860
rect 23116 28804 23172 28860
rect 23172 28804 23176 28860
rect 23112 28800 23176 28804
rect 23192 28860 23256 28864
rect 23192 28804 23196 28860
rect 23196 28804 23252 28860
rect 23252 28804 23256 28860
rect 23192 28800 23256 28804
rect 20852 28384 20916 28388
rect 20852 28328 20902 28384
rect 20902 28328 20916 28384
rect 20852 28324 20916 28328
rect 7952 28316 8016 28320
rect 7952 28260 7956 28316
rect 7956 28260 8012 28316
rect 8012 28260 8016 28316
rect 7952 28256 8016 28260
rect 8032 28316 8096 28320
rect 8032 28260 8036 28316
rect 8036 28260 8092 28316
rect 8092 28260 8096 28316
rect 8032 28256 8096 28260
rect 8112 28316 8176 28320
rect 8112 28260 8116 28316
rect 8116 28260 8172 28316
rect 8172 28260 8176 28316
rect 8112 28256 8176 28260
rect 8192 28316 8256 28320
rect 8192 28260 8196 28316
rect 8196 28260 8252 28316
rect 8252 28260 8256 28316
rect 8192 28256 8256 28260
rect 17952 28316 18016 28320
rect 17952 28260 17956 28316
rect 17956 28260 18012 28316
rect 18012 28260 18016 28316
rect 17952 28256 18016 28260
rect 18032 28316 18096 28320
rect 18032 28260 18036 28316
rect 18036 28260 18092 28316
rect 18092 28260 18096 28316
rect 18032 28256 18096 28260
rect 18112 28316 18176 28320
rect 18112 28260 18116 28316
rect 18116 28260 18172 28316
rect 18172 28260 18176 28316
rect 18112 28256 18176 28260
rect 18192 28316 18256 28320
rect 18192 28260 18196 28316
rect 18196 28260 18252 28316
rect 18252 28260 18256 28316
rect 18192 28256 18256 28260
rect 16252 28052 16316 28116
rect 2952 27772 3016 27776
rect 2952 27716 2956 27772
rect 2956 27716 3012 27772
rect 3012 27716 3016 27772
rect 2952 27712 3016 27716
rect 3032 27772 3096 27776
rect 3032 27716 3036 27772
rect 3036 27716 3092 27772
rect 3092 27716 3096 27772
rect 3032 27712 3096 27716
rect 3112 27772 3176 27776
rect 3112 27716 3116 27772
rect 3116 27716 3172 27772
rect 3172 27716 3176 27772
rect 3112 27712 3176 27716
rect 3192 27772 3256 27776
rect 3192 27716 3196 27772
rect 3196 27716 3252 27772
rect 3252 27716 3256 27772
rect 3192 27712 3256 27716
rect 12952 27772 13016 27776
rect 12952 27716 12956 27772
rect 12956 27716 13012 27772
rect 13012 27716 13016 27772
rect 12952 27712 13016 27716
rect 13032 27772 13096 27776
rect 13032 27716 13036 27772
rect 13036 27716 13092 27772
rect 13092 27716 13096 27772
rect 13032 27712 13096 27716
rect 13112 27772 13176 27776
rect 13112 27716 13116 27772
rect 13116 27716 13172 27772
rect 13172 27716 13176 27772
rect 13112 27712 13176 27716
rect 13192 27772 13256 27776
rect 13192 27716 13196 27772
rect 13196 27716 13252 27772
rect 13252 27716 13256 27772
rect 13192 27712 13256 27716
rect 22952 27772 23016 27776
rect 22952 27716 22956 27772
rect 22956 27716 23012 27772
rect 23012 27716 23016 27772
rect 22952 27712 23016 27716
rect 23032 27772 23096 27776
rect 23032 27716 23036 27772
rect 23036 27716 23092 27772
rect 23092 27716 23096 27772
rect 23032 27712 23096 27716
rect 23112 27772 23176 27776
rect 23112 27716 23116 27772
rect 23116 27716 23172 27772
rect 23172 27716 23176 27772
rect 23112 27712 23176 27716
rect 23192 27772 23256 27776
rect 23192 27716 23196 27772
rect 23196 27716 23252 27772
rect 23252 27716 23256 27772
rect 23192 27712 23256 27716
rect 18460 27508 18524 27572
rect 21220 27508 21284 27572
rect 7952 27228 8016 27232
rect 7952 27172 7956 27228
rect 7956 27172 8012 27228
rect 8012 27172 8016 27228
rect 7952 27168 8016 27172
rect 8032 27228 8096 27232
rect 8032 27172 8036 27228
rect 8036 27172 8092 27228
rect 8092 27172 8096 27228
rect 8032 27168 8096 27172
rect 8112 27228 8176 27232
rect 8112 27172 8116 27228
rect 8116 27172 8172 27228
rect 8172 27172 8176 27228
rect 8112 27168 8176 27172
rect 8192 27228 8256 27232
rect 8192 27172 8196 27228
rect 8196 27172 8252 27228
rect 8252 27172 8256 27228
rect 8192 27168 8256 27172
rect 17952 27228 18016 27232
rect 17952 27172 17956 27228
rect 17956 27172 18012 27228
rect 18012 27172 18016 27228
rect 17952 27168 18016 27172
rect 18032 27228 18096 27232
rect 18032 27172 18036 27228
rect 18036 27172 18092 27228
rect 18092 27172 18096 27228
rect 18032 27168 18096 27172
rect 18112 27228 18176 27232
rect 18112 27172 18116 27228
rect 18116 27172 18172 27228
rect 18172 27172 18176 27228
rect 18112 27168 18176 27172
rect 18192 27228 18256 27232
rect 18192 27172 18196 27228
rect 18196 27172 18252 27228
rect 18252 27172 18256 27228
rect 18192 27168 18256 27172
rect 15700 27160 15764 27164
rect 15700 27104 15750 27160
rect 15750 27104 15764 27160
rect 15700 27100 15764 27104
rect 21404 27100 21468 27164
rect 2952 26684 3016 26688
rect 2952 26628 2956 26684
rect 2956 26628 3012 26684
rect 3012 26628 3016 26684
rect 2952 26624 3016 26628
rect 3032 26684 3096 26688
rect 3032 26628 3036 26684
rect 3036 26628 3092 26684
rect 3092 26628 3096 26684
rect 3032 26624 3096 26628
rect 3112 26684 3176 26688
rect 3112 26628 3116 26684
rect 3116 26628 3172 26684
rect 3172 26628 3176 26684
rect 3112 26624 3176 26628
rect 3192 26684 3256 26688
rect 3192 26628 3196 26684
rect 3196 26628 3252 26684
rect 3252 26628 3256 26684
rect 3192 26624 3256 26628
rect 12952 26684 13016 26688
rect 12952 26628 12956 26684
rect 12956 26628 13012 26684
rect 13012 26628 13016 26684
rect 12952 26624 13016 26628
rect 13032 26684 13096 26688
rect 13032 26628 13036 26684
rect 13036 26628 13092 26684
rect 13092 26628 13096 26684
rect 13032 26624 13096 26628
rect 13112 26684 13176 26688
rect 13112 26628 13116 26684
rect 13116 26628 13172 26684
rect 13172 26628 13176 26684
rect 13112 26624 13176 26628
rect 13192 26684 13256 26688
rect 13192 26628 13196 26684
rect 13196 26628 13252 26684
rect 13252 26628 13256 26684
rect 13192 26624 13256 26628
rect 22952 26684 23016 26688
rect 22952 26628 22956 26684
rect 22956 26628 23012 26684
rect 23012 26628 23016 26684
rect 22952 26624 23016 26628
rect 23032 26684 23096 26688
rect 23032 26628 23036 26684
rect 23036 26628 23092 26684
rect 23092 26628 23096 26684
rect 23032 26624 23096 26628
rect 23112 26684 23176 26688
rect 23112 26628 23116 26684
rect 23116 26628 23172 26684
rect 23172 26628 23176 26684
rect 23112 26624 23176 26628
rect 23192 26684 23256 26688
rect 23192 26628 23196 26684
rect 23196 26628 23252 26684
rect 23252 26628 23256 26684
rect 23192 26624 23256 26628
rect 23428 26148 23492 26212
rect 7952 26140 8016 26144
rect 7952 26084 7956 26140
rect 7956 26084 8012 26140
rect 8012 26084 8016 26140
rect 7952 26080 8016 26084
rect 8032 26140 8096 26144
rect 8032 26084 8036 26140
rect 8036 26084 8092 26140
rect 8092 26084 8096 26140
rect 8032 26080 8096 26084
rect 8112 26140 8176 26144
rect 8112 26084 8116 26140
rect 8116 26084 8172 26140
rect 8172 26084 8176 26140
rect 8112 26080 8176 26084
rect 8192 26140 8256 26144
rect 8192 26084 8196 26140
rect 8196 26084 8252 26140
rect 8252 26084 8256 26140
rect 8192 26080 8256 26084
rect 17952 26140 18016 26144
rect 17952 26084 17956 26140
rect 17956 26084 18012 26140
rect 18012 26084 18016 26140
rect 17952 26080 18016 26084
rect 18032 26140 18096 26144
rect 18032 26084 18036 26140
rect 18036 26084 18092 26140
rect 18092 26084 18096 26140
rect 18032 26080 18096 26084
rect 18112 26140 18176 26144
rect 18112 26084 18116 26140
rect 18116 26084 18172 26140
rect 18172 26084 18176 26140
rect 18112 26080 18176 26084
rect 18192 26140 18256 26144
rect 18192 26084 18196 26140
rect 18196 26084 18252 26140
rect 18252 26084 18256 26140
rect 18192 26080 18256 26084
rect 16068 25664 16132 25668
rect 16068 25608 16118 25664
rect 16118 25608 16132 25664
rect 16068 25604 16132 25608
rect 2952 25596 3016 25600
rect 2952 25540 2956 25596
rect 2956 25540 3012 25596
rect 3012 25540 3016 25596
rect 2952 25536 3016 25540
rect 3032 25596 3096 25600
rect 3032 25540 3036 25596
rect 3036 25540 3092 25596
rect 3092 25540 3096 25596
rect 3032 25536 3096 25540
rect 3112 25596 3176 25600
rect 3112 25540 3116 25596
rect 3116 25540 3172 25596
rect 3172 25540 3176 25596
rect 3112 25536 3176 25540
rect 3192 25596 3256 25600
rect 3192 25540 3196 25596
rect 3196 25540 3252 25596
rect 3252 25540 3256 25596
rect 3192 25536 3256 25540
rect 12952 25596 13016 25600
rect 12952 25540 12956 25596
rect 12956 25540 13012 25596
rect 13012 25540 13016 25596
rect 12952 25536 13016 25540
rect 13032 25596 13096 25600
rect 13032 25540 13036 25596
rect 13036 25540 13092 25596
rect 13092 25540 13096 25596
rect 13032 25536 13096 25540
rect 13112 25596 13176 25600
rect 13112 25540 13116 25596
rect 13116 25540 13172 25596
rect 13172 25540 13176 25596
rect 13112 25536 13176 25540
rect 13192 25596 13256 25600
rect 13192 25540 13196 25596
rect 13196 25540 13252 25596
rect 13252 25540 13256 25596
rect 13192 25536 13256 25540
rect 22952 25596 23016 25600
rect 22952 25540 22956 25596
rect 22956 25540 23012 25596
rect 23012 25540 23016 25596
rect 22952 25536 23016 25540
rect 23032 25596 23096 25600
rect 23032 25540 23036 25596
rect 23036 25540 23092 25596
rect 23092 25540 23096 25596
rect 23032 25536 23096 25540
rect 23112 25596 23176 25600
rect 23112 25540 23116 25596
rect 23116 25540 23172 25596
rect 23172 25540 23176 25596
rect 23112 25536 23176 25540
rect 23192 25596 23256 25600
rect 23192 25540 23196 25596
rect 23196 25540 23252 25596
rect 23252 25540 23256 25596
rect 23192 25536 23256 25540
rect 7952 25052 8016 25056
rect 7952 24996 7956 25052
rect 7956 24996 8012 25052
rect 8012 24996 8016 25052
rect 7952 24992 8016 24996
rect 8032 25052 8096 25056
rect 8032 24996 8036 25052
rect 8036 24996 8092 25052
rect 8092 24996 8096 25052
rect 8032 24992 8096 24996
rect 8112 25052 8176 25056
rect 8112 24996 8116 25052
rect 8116 24996 8172 25052
rect 8172 24996 8176 25052
rect 8112 24992 8176 24996
rect 8192 25052 8256 25056
rect 8192 24996 8196 25052
rect 8196 24996 8252 25052
rect 8252 24996 8256 25052
rect 8192 24992 8256 24996
rect 17952 25052 18016 25056
rect 17952 24996 17956 25052
rect 17956 24996 18012 25052
rect 18012 24996 18016 25052
rect 17952 24992 18016 24996
rect 18032 25052 18096 25056
rect 18032 24996 18036 25052
rect 18036 24996 18092 25052
rect 18092 24996 18096 25052
rect 18032 24992 18096 24996
rect 18112 25052 18176 25056
rect 18112 24996 18116 25052
rect 18116 24996 18172 25052
rect 18172 24996 18176 25052
rect 18112 24992 18176 24996
rect 18192 25052 18256 25056
rect 18192 24996 18196 25052
rect 18196 24996 18252 25052
rect 18252 24996 18256 25052
rect 18192 24992 18256 24996
rect 20852 24516 20916 24580
rect 2952 24508 3016 24512
rect 2952 24452 2956 24508
rect 2956 24452 3012 24508
rect 3012 24452 3016 24508
rect 2952 24448 3016 24452
rect 3032 24508 3096 24512
rect 3032 24452 3036 24508
rect 3036 24452 3092 24508
rect 3092 24452 3096 24508
rect 3032 24448 3096 24452
rect 3112 24508 3176 24512
rect 3112 24452 3116 24508
rect 3116 24452 3172 24508
rect 3172 24452 3176 24508
rect 3112 24448 3176 24452
rect 3192 24508 3256 24512
rect 3192 24452 3196 24508
rect 3196 24452 3252 24508
rect 3252 24452 3256 24508
rect 3192 24448 3256 24452
rect 12952 24508 13016 24512
rect 12952 24452 12956 24508
rect 12956 24452 13012 24508
rect 13012 24452 13016 24508
rect 12952 24448 13016 24452
rect 13032 24508 13096 24512
rect 13032 24452 13036 24508
rect 13036 24452 13092 24508
rect 13092 24452 13096 24508
rect 13032 24448 13096 24452
rect 13112 24508 13176 24512
rect 13112 24452 13116 24508
rect 13116 24452 13172 24508
rect 13172 24452 13176 24508
rect 13112 24448 13176 24452
rect 13192 24508 13256 24512
rect 13192 24452 13196 24508
rect 13196 24452 13252 24508
rect 13252 24452 13256 24508
rect 13192 24448 13256 24452
rect 22952 24508 23016 24512
rect 22952 24452 22956 24508
rect 22956 24452 23012 24508
rect 23012 24452 23016 24508
rect 22952 24448 23016 24452
rect 23032 24508 23096 24512
rect 23032 24452 23036 24508
rect 23036 24452 23092 24508
rect 23092 24452 23096 24508
rect 23032 24448 23096 24452
rect 23112 24508 23176 24512
rect 23112 24452 23116 24508
rect 23116 24452 23172 24508
rect 23172 24452 23176 24508
rect 23112 24448 23176 24452
rect 23192 24508 23256 24512
rect 23192 24452 23196 24508
rect 23196 24452 23252 24508
rect 23252 24452 23256 24508
rect 23192 24448 23256 24452
rect 12572 24108 12636 24172
rect 7952 23964 8016 23968
rect 7952 23908 7956 23964
rect 7956 23908 8012 23964
rect 8012 23908 8016 23964
rect 7952 23904 8016 23908
rect 8032 23964 8096 23968
rect 8032 23908 8036 23964
rect 8036 23908 8092 23964
rect 8092 23908 8096 23964
rect 8032 23904 8096 23908
rect 8112 23964 8176 23968
rect 8112 23908 8116 23964
rect 8116 23908 8172 23964
rect 8172 23908 8176 23964
rect 8112 23904 8176 23908
rect 8192 23964 8256 23968
rect 8192 23908 8196 23964
rect 8196 23908 8252 23964
rect 8252 23908 8256 23964
rect 8192 23904 8256 23908
rect 17952 23964 18016 23968
rect 17952 23908 17956 23964
rect 17956 23908 18012 23964
rect 18012 23908 18016 23964
rect 17952 23904 18016 23908
rect 18032 23964 18096 23968
rect 18032 23908 18036 23964
rect 18036 23908 18092 23964
rect 18092 23908 18096 23964
rect 18032 23904 18096 23908
rect 18112 23964 18176 23968
rect 18112 23908 18116 23964
rect 18116 23908 18172 23964
rect 18172 23908 18176 23964
rect 18112 23904 18176 23908
rect 18192 23964 18256 23968
rect 18192 23908 18196 23964
rect 18196 23908 18252 23964
rect 18252 23908 18256 23964
rect 18192 23904 18256 23908
rect 13492 23428 13556 23492
rect 14412 23428 14476 23492
rect 2952 23420 3016 23424
rect 2952 23364 2956 23420
rect 2956 23364 3012 23420
rect 3012 23364 3016 23420
rect 2952 23360 3016 23364
rect 3032 23420 3096 23424
rect 3032 23364 3036 23420
rect 3036 23364 3092 23420
rect 3092 23364 3096 23420
rect 3032 23360 3096 23364
rect 3112 23420 3176 23424
rect 3112 23364 3116 23420
rect 3116 23364 3172 23420
rect 3172 23364 3176 23420
rect 3112 23360 3176 23364
rect 3192 23420 3256 23424
rect 3192 23364 3196 23420
rect 3196 23364 3252 23420
rect 3252 23364 3256 23420
rect 3192 23360 3256 23364
rect 12952 23420 13016 23424
rect 12952 23364 12956 23420
rect 12956 23364 13012 23420
rect 13012 23364 13016 23420
rect 12952 23360 13016 23364
rect 13032 23420 13096 23424
rect 13032 23364 13036 23420
rect 13036 23364 13092 23420
rect 13092 23364 13096 23420
rect 13032 23360 13096 23364
rect 13112 23420 13176 23424
rect 13112 23364 13116 23420
rect 13116 23364 13172 23420
rect 13172 23364 13176 23420
rect 13112 23360 13176 23364
rect 13192 23420 13256 23424
rect 13192 23364 13196 23420
rect 13196 23364 13252 23420
rect 13252 23364 13256 23420
rect 13192 23360 13256 23364
rect 22952 23420 23016 23424
rect 22952 23364 22956 23420
rect 22956 23364 23012 23420
rect 23012 23364 23016 23420
rect 22952 23360 23016 23364
rect 23032 23420 23096 23424
rect 23032 23364 23036 23420
rect 23036 23364 23092 23420
rect 23092 23364 23096 23420
rect 23032 23360 23096 23364
rect 23112 23420 23176 23424
rect 23112 23364 23116 23420
rect 23116 23364 23172 23420
rect 23172 23364 23176 23420
rect 23112 23360 23176 23364
rect 23192 23420 23256 23424
rect 23192 23364 23196 23420
rect 23196 23364 23252 23420
rect 23252 23364 23256 23420
rect 23192 23360 23256 23364
rect 17724 23292 17788 23356
rect 7952 22876 8016 22880
rect 7952 22820 7956 22876
rect 7956 22820 8012 22876
rect 8012 22820 8016 22876
rect 7952 22816 8016 22820
rect 8032 22876 8096 22880
rect 8032 22820 8036 22876
rect 8036 22820 8092 22876
rect 8092 22820 8096 22876
rect 8032 22816 8096 22820
rect 8112 22876 8176 22880
rect 8112 22820 8116 22876
rect 8116 22820 8172 22876
rect 8172 22820 8176 22876
rect 8112 22816 8176 22820
rect 8192 22876 8256 22880
rect 8192 22820 8196 22876
rect 8196 22820 8252 22876
rect 8252 22820 8256 22876
rect 8192 22816 8256 22820
rect 17952 22876 18016 22880
rect 17952 22820 17956 22876
rect 17956 22820 18012 22876
rect 18012 22820 18016 22876
rect 17952 22816 18016 22820
rect 18032 22876 18096 22880
rect 18032 22820 18036 22876
rect 18036 22820 18092 22876
rect 18092 22820 18096 22876
rect 18032 22816 18096 22820
rect 18112 22876 18176 22880
rect 18112 22820 18116 22876
rect 18116 22820 18172 22876
rect 18172 22820 18176 22876
rect 18112 22816 18176 22820
rect 18192 22876 18256 22880
rect 18192 22820 18196 22876
rect 18196 22820 18252 22876
rect 18252 22820 18256 22876
rect 18192 22816 18256 22820
rect 10180 22612 10244 22676
rect 12756 22612 12820 22676
rect 13492 22476 13556 22540
rect 2952 22332 3016 22336
rect 2952 22276 2956 22332
rect 2956 22276 3012 22332
rect 3012 22276 3016 22332
rect 2952 22272 3016 22276
rect 3032 22332 3096 22336
rect 3032 22276 3036 22332
rect 3036 22276 3092 22332
rect 3092 22276 3096 22332
rect 3032 22272 3096 22276
rect 3112 22332 3176 22336
rect 3112 22276 3116 22332
rect 3116 22276 3172 22332
rect 3172 22276 3176 22332
rect 3112 22272 3176 22276
rect 3192 22332 3256 22336
rect 3192 22276 3196 22332
rect 3196 22276 3252 22332
rect 3252 22276 3256 22332
rect 3192 22272 3256 22276
rect 12952 22332 13016 22336
rect 12952 22276 12956 22332
rect 12956 22276 13012 22332
rect 13012 22276 13016 22332
rect 12952 22272 13016 22276
rect 13032 22332 13096 22336
rect 13032 22276 13036 22332
rect 13036 22276 13092 22332
rect 13092 22276 13096 22332
rect 13032 22272 13096 22276
rect 13112 22332 13176 22336
rect 13112 22276 13116 22332
rect 13116 22276 13172 22332
rect 13172 22276 13176 22332
rect 13112 22272 13176 22276
rect 13192 22332 13256 22336
rect 13192 22276 13196 22332
rect 13196 22276 13252 22332
rect 13252 22276 13256 22332
rect 13192 22272 13256 22276
rect 22952 22332 23016 22336
rect 22952 22276 22956 22332
rect 22956 22276 23012 22332
rect 23012 22276 23016 22332
rect 22952 22272 23016 22276
rect 23032 22332 23096 22336
rect 23032 22276 23036 22332
rect 23036 22276 23092 22332
rect 23092 22276 23096 22332
rect 23032 22272 23096 22276
rect 23112 22332 23176 22336
rect 23112 22276 23116 22332
rect 23116 22276 23172 22332
rect 23172 22276 23176 22332
rect 23112 22272 23176 22276
rect 23192 22332 23256 22336
rect 23192 22276 23196 22332
rect 23196 22276 23252 22332
rect 23252 22276 23256 22332
rect 23192 22272 23256 22276
rect 17724 22204 17788 22268
rect 13860 21856 13924 21860
rect 13860 21800 13874 21856
rect 13874 21800 13924 21856
rect 13860 21796 13924 21800
rect 7952 21788 8016 21792
rect 7952 21732 7956 21788
rect 7956 21732 8012 21788
rect 8012 21732 8016 21788
rect 7952 21728 8016 21732
rect 8032 21788 8096 21792
rect 8032 21732 8036 21788
rect 8036 21732 8092 21788
rect 8092 21732 8096 21788
rect 8032 21728 8096 21732
rect 8112 21788 8176 21792
rect 8112 21732 8116 21788
rect 8116 21732 8172 21788
rect 8172 21732 8176 21788
rect 8112 21728 8176 21732
rect 8192 21788 8256 21792
rect 8192 21732 8196 21788
rect 8196 21732 8252 21788
rect 8252 21732 8256 21788
rect 8192 21728 8256 21732
rect 17952 21788 18016 21792
rect 17952 21732 17956 21788
rect 17956 21732 18012 21788
rect 18012 21732 18016 21788
rect 17952 21728 18016 21732
rect 18032 21788 18096 21792
rect 18032 21732 18036 21788
rect 18036 21732 18092 21788
rect 18092 21732 18096 21788
rect 18032 21728 18096 21732
rect 18112 21788 18176 21792
rect 18112 21732 18116 21788
rect 18116 21732 18172 21788
rect 18172 21732 18176 21788
rect 18112 21728 18176 21732
rect 18192 21788 18256 21792
rect 18192 21732 18196 21788
rect 18196 21732 18252 21788
rect 18252 21732 18256 21788
rect 18192 21728 18256 21732
rect 2952 21244 3016 21248
rect 2952 21188 2956 21244
rect 2956 21188 3012 21244
rect 3012 21188 3016 21244
rect 2952 21184 3016 21188
rect 3032 21244 3096 21248
rect 3032 21188 3036 21244
rect 3036 21188 3092 21244
rect 3092 21188 3096 21244
rect 3032 21184 3096 21188
rect 3112 21244 3176 21248
rect 3112 21188 3116 21244
rect 3116 21188 3172 21244
rect 3172 21188 3176 21244
rect 3112 21184 3176 21188
rect 3192 21244 3256 21248
rect 3192 21188 3196 21244
rect 3196 21188 3252 21244
rect 3252 21188 3256 21244
rect 3192 21184 3256 21188
rect 12952 21244 13016 21248
rect 12952 21188 12956 21244
rect 12956 21188 13012 21244
rect 13012 21188 13016 21244
rect 12952 21184 13016 21188
rect 13032 21244 13096 21248
rect 13032 21188 13036 21244
rect 13036 21188 13092 21244
rect 13092 21188 13096 21244
rect 13032 21184 13096 21188
rect 13112 21244 13176 21248
rect 13112 21188 13116 21244
rect 13116 21188 13172 21244
rect 13172 21188 13176 21244
rect 13112 21184 13176 21188
rect 13192 21244 13256 21248
rect 13192 21188 13196 21244
rect 13196 21188 13252 21244
rect 13252 21188 13256 21244
rect 13192 21184 13256 21188
rect 22952 21244 23016 21248
rect 22952 21188 22956 21244
rect 22956 21188 23012 21244
rect 23012 21188 23016 21244
rect 22952 21184 23016 21188
rect 23032 21244 23096 21248
rect 23032 21188 23036 21244
rect 23036 21188 23092 21244
rect 23092 21188 23096 21244
rect 23032 21184 23096 21188
rect 23112 21244 23176 21248
rect 23112 21188 23116 21244
rect 23116 21188 23172 21244
rect 23172 21188 23176 21244
rect 23112 21184 23176 21188
rect 23192 21244 23256 21248
rect 23192 21188 23196 21244
rect 23196 21188 23252 21244
rect 23252 21188 23256 21244
rect 23192 21184 23256 21188
rect 7952 20700 8016 20704
rect 7952 20644 7956 20700
rect 7956 20644 8012 20700
rect 8012 20644 8016 20700
rect 7952 20640 8016 20644
rect 8032 20700 8096 20704
rect 8032 20644 8036 20700
rect 8036 20644 8092 20700
rect 8092 20644 8096 20700
rect 8032 20640 8096 20644
rect 8112 20700 8176 20704
rect 8112 20644 8116 20700
rect 8116 20644 8172 20700
rect 8172 20644 8176 20700
rect 8112 20640 8176 20644
rect 8192 20700 8256 20704
rect 8192 20644 8196 20700
rect 8196 20644 8252 20700
rect 8252 20644 8256 20700
rect 8192 20640 8256 20644
rect 17952 20700 18016 20704
rect 17952 20644 17956 20700
rect 17956 20644 18012 20700
rect 18012 20644 18016 20700
rect 17952 20640 18016 20644
rect 18032 20700 18096 20704
rect 18032 20644 18036 20700
rect 18036 20644 18092 20700
rect 18092 20644 18096 20700
rect 18032 20640 18096 20644
rect 18112 20700 18176 20704
rect 18112 20644 18116 20700
rect 18116 20644 18172 20700
rect 18172 20644 18176 20700
rect 18112 20640 18176 20644
rect 18192 20700 18256 20704
rect 18192 20644 18196 20700
rect 18196 20644 18252 20700
rect 18252 20644 18256 20700
rect 18192 20640 18256 20644
rect 16068 20572 16132 20636
rect 14964 20164 15028 20228
rect 2952 20156 3016 20160
rect 2952 20100 2956 20156
rect 2956 20100 3012 20156
rect 3012 20100 3016 20156
rect 2952 20096 3016 20100
rect 3032 20156 3096 20160
rect 3032 20100 3036 20156
rect 3036 20100 3092 20156
rect 3092 20100 3096 20156
rect 3032 20096 3096 20100
rect 3112 20156 3176 20160
rect 3112 20100 3116 20156
rect 3116 20100 3172 20156
rect 3172 20100 3176 20156
rect 3112 20096 3176 20100
rect 3192 20156 3256 20160
rect 3192 20100 3196 20156
rect 3196 20100 3252 20156
rect 3252 20100 3256 20156
rect 3192 20096 3256 20100
rect 12952 20156 13016 20160
rect 12952 20100 12956 20156
rect 12956 20100 13012 20156
rect 13012 20100 13016 20156
rect 12952 20096 13016 20100
rect 13032 20156 13096 20160
rect 13032 20100 13036 20156
rect 13036 20100 13092 20156
rect 13092 20100 13096 20156
rect 13032 20096 13096 20100
rect 13112 20156 13176 20160
rect 13112 20100 13116 20156
rect 13116 20100 13172 20156
rect 13172 20100 13176 20156
rect 13112 20096 13176 20100
rect 13192 20156 13256 20160
rect 13192 20100 13196 20156
rect 13196 20100 13252 20156
rect 13252 20100 13256 20156
rect 13192 20096 13256 20100
rect 22952 20156 23016 20160
rect 22952 20100 22956 20156
rect 22956 20100 23012 20156
rect 23012 20100 23016 20156
rect 22952 20096 23016 20100
rect 23032 20156 23096 20160
rect 23032 20100 23036 20156
rect 23036 20100 23092 20156
rect 23092 20100 23096 20156
rect 23032 20096 23096 20100
rect 23112 20156 23176 20160
rect 23112 20100 23116 20156
rect 23116 20100 23172 20156
rect 23172 20100 23176 20156
rect 23112 20096 23176 20100
rect 23192 20156 23256 20160
rect 23192 20100 23196 20156
rect 23196 20100 23252 20156
rect 23252 20100 23256 20156
rect 23192 20096 23256 20100
rect 18644 19892 18708 19956
rect 7952 19612 8016 19616
rect 7952 19556 7956 19612
rect 7956 19556 8012 19612
rect 8012 19556 8016 19612
rect 7952 19552 8016 19556
rect 8032 19612 8096 19616
rect 8032 19556 8036 19612
rect 8036 19556 8092 19612
rect 8092 19556 8096 19612
rect 8032 19552 8096 19556
rect 8112 19612 8176 19616
rect 8112 19556 8116 19612
rect 8116 19556 8172 19612
rect 8172 19556 8176 19612
rect 8112 19552 8176 19556
rect 8192 19612 8256 19616
rect 8192 19556 8196 19612
rect 8196 19556 8252 19612
rect 8252 19556 8256 19612
rect 8192 19552 8256 19556
rect 17952 19612 18016 19616
rect 17952 19556 17956 19612
rect 17956 19556 18012 19612
rect 18012 19556 18016 19612
rect 17952 19552 18016 19556
rect 18032 19612 18096 19616
rect 18032 19556 18036 19612
rect 18036 19556 18092 19612
rect 18092 19556 18096 19612
rect 18032 19552 18096 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 2952 19068 3016 19072
rect 2952 19012 2956 19068
rect 2956 19012 3012 19068
rect 3012 19012 3016 19068
rect 2952 19008 3016 19012
rect 3032 19068 3096 19072
rect 3032 19012 3036 19068
rect 3036 19012 3092 19068
rect 3092 19012 3096 19068
rect 3032 19008 3096 19012
rect 3112 19068 3176 19072
rect 3112 19012 3116 19068
rect 3116 19012 3172 19068
rect 3172 19012 3176 19068
rect 3112 19008 3176 19012
rect 3192 19068 3256 19072
rect 3192 19012 3196 19068
rect 3196 19012 3252 19068
rect 3252 19012 3256 19068
rect 3192 19008 3256 19012
rect 12952 19068 13016 19072
rect 12952 19012 12956 19068
rect 12956 19012 13012 19068
rect 13012 19012 13016 19068
rect 12952 19008 13016 19012
rect 13032 19068 13096 19072
rect 13032 19012 13036 19068
rect 13036 19012 13092 19068
rect 13092 19012 13096 19068
rect 13032 19008 13096 19012
rect 13112 19068 13176 19072
rect 13112 19012 13116 19068
rect 13116 19012 13172 19068
rect 13172 19012 13176 19068
rect 13112 19008 13176 19012
rect 13192 19068 13256 19072
rect 13192 19012 13196 19068
rect 13196 19012 13252 19068
rect 13252 19012 13256 19068
rect 13192 19008 13256 19012
rect 22952 19068 23016 19072
rect 22952 19012 22956 19068
rect 22956 19012 23012 19068
rect 23012 19012 23016 19068
rect 22952 19008 23016 19012
rect 23032 19068 23096 19072
rect 23032 19012 23036 19068
rect 23036 19012 23092 19068
rect 23092 19012 23096 19068
rect 23032 19008 23096 19012
rect 23112 19068 23176 19072
rect 23112 19012 23116 19068
rect 23116 19012 23172 19068
rect 23172 19012 23176 19068
rect 23112 19008 23176 19012
rect 23192 19068 23256 19072
rect 23192 19012 23196 19068
rect 23196 19012 23252 19068
rect 23252 19012 23256 19068
rect 23192 19008 23256 19012
rect 17540 18864 17604 18868
rect 17540 18808 17590 18864
rect 17590 18808 17604 18864
rect 17540 18804 17604 18808
rect 7952 18524 8016 18528
rect 7952 18468 7956 18524
rect 7956 18468 8012 18524
rect 8012 18468 8016 18524
rect 7952 18464 8016 18468
rect 8032 18524 8096 18528
rect 8032 18468 8036 18524
rect 8036 18468 8092 18524
rect 8092 18468 8096 18524
rect 8032 18464 8096 18468
rect 8112 18524 8176 18528
rect 8112 18468 8116 18524
rect 8116 18468 8172 18524
rect 8172 18468 8176 18524
rect 8112 18464 8176 18468
rect 8192 18524 8256 18528
rect 8192 18468 8196 18524
rect 8196 18468 8252 18524
rect 8252 18468 8256 18524
rect 8192 18464 8256 18468
rect 17952 18524 18016 18528
rect 17952 18468 17956 18524
rect 17956 18468 18012 18524
rect 18012 18468 18016 18524
rect 17952 18464 18016 18468
rect 18032 18524 18096 18528
rect 18032 18468 18036 18524
rect 18036 18468 18092 18524
rect 18092 18468 18096 18524
rect 18032 18464 18096 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 18460 18320 18524 18324
rect 18460 18264 18510 18320
rect 18510 18264 18524 18320
rect 18460 18260 18524 18264
rect 2952 17980 3016 17984
rect 2952 17924 2956 17980
rect 2956 17924 3012 17980
rect 3012 17924 3016 17980
rect 2952 17920 3016 17924
rect 3032 17980 3096 17984
rect 3032 17924 3036 17980
rect 3036 17924 3092 17980
rect 3092 17924 3096 17980
rect 3032 17920 3096 17924
rect 3112 17980 3176 17984
rect 3112 17924 3116 17980
rect 3116 17924 3172 17980
rect 3172 17924 3176 17980
rect 3112 17920 3176 17924
rect 3192 17980 3256 17984
rect 3192 17924 3196 17980
rect 3196 17924 3252 17980
rect 3252 17924 3256 17980
rect 3192 17920 3256 17924
rect 12952 17980 13016 17984
rect 12952 17924 12956 17980
rect 12956 17924 13012 17980
rect 13012 17924 13016 17980
rect 12952 17920 13016 17924
rect 13032 17980 13096 17984
rect 13032 17924 13036 17980
rect 13036 17924 13092 17980
rect 13092 17924 13096 17980
rect 13032 17920 13096 17924
rect 13112 17980 13176 17984
rect 13112 17924 13116 17980
rect 13116 17924 13172 17980
rect 13172 17924 13176 17980
rect 13112 17920 13176 17924
rect 13192 17980 13256 17984
rect 13192 17924 13196 17980
rect 13196 17924 13252 17980
rect 13252 17924 13256 17980
rect 13192 17920 13256 17924
rect 22952 17980 23016 17984
rect 22952 17924 22956 17980
rect 22956 17924 23012 17980
rect 23012 17924 23016 17980
rect 22952 17920 23016 17924
rect 23032 17980 23096 17984
rect 23032 17924 23036 17980
rect 23036 17924 23092 17980
rect 23092 17924 23096 17980
rect 23032 17920 23096 17924
rect 23112 17980 23176 17984
rect 23112 17924 23116 17980
rect 23116 17924 23172 17980
rect 23172 17924 23176 17980
rect 23112 17920 23176 17924
rect 23192 17980 23256 17984
rect 23192 17924 23196 17980
rect 23196 17924 23252 17980
rect 23252 17924 23256 17980
rect 23192 17920 23256 17924
rect 12572 17852 12636 17916
rect 16252 17640 16316 17644
rect 16252 17584 16266 17640
rect 16266 17584 16316 17640
rect 16252 17580 16316 17584
rect 19564 17580 19628 17644
rect 7952 17436 8016 17440
rect 7952 17380 7956 17436
rect 7956 17380 8012 17436
rect 8012 17380 8016 17436
rect 7952 17376 8016 17380
rect 8032 17436 8096 17440
rect 8032 17380 8036 17436
rect 8036 17380 8092 17436
rect 8092 17380 8096 17436
rect 8032 17376 8096 17380
rect 8112 17436 8176 17440
rect 8112 17380 8116 17436
rect 8116 17380 8172 17436
rect 8172 17380 8176 17436
rect 8112 17376 8176 17380
rect 8192 17436 8256 17440
rect 8192 17380 8196 17436
rect 8196 17380 8252 17436
rect 8252 17380 8256 17436
rect 8192 17376 8256 17380
rect 17952 17436 18016 17440
rect 17952 17380 17956 17436
rect 17956 17380 18012 17436
rect 18012 17380 18016 17436
rect 17952 17376 18016 17380
rect 18032 17436 18096 17440
rect 18032 17380 18036 17436
rect 18036 17380 18092 17436
rect 18092 17380 18096 17436
rect 18032 17376 18096 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 2952 16892 3016 16896
rect 2952 16836 2956 16892
rect 2956 16836 3012 16892
rect 3012 16836 3016 16892
rect 2952 16832 3016 16836
rect 3032 16892 3096 16896
rect 3032 16836 3036 16892
rect 3036 16836 3092 16892
rect 3092 16836 3096 16892
rect 3032 16832 3096 16836
rect 3112 16892 3176 16896
rect 3112 16836 3116 16892
rect 3116 16836 3172 16892
rect 3172 16836 3176 16892
rect 3112 16832 3176 16836
rect 3192 16892 3256 16896
rect 3192 16836 3196 16892
rect 3196 16836 3252 16892
rect 3252 16836 3256 16892
rect 3192 16832 3256 16836
rect 12952 16892 13016 16896
rect 12952 16836 12956 16892
rect 12956 16836 13012 16892
rect 13012 16836 13016 16892
rect 12952 16832 13016 16836
rect 13032 16892 13096 16896
rect 13032 16836 13036 16892
rect 13036 16836 13092 16892
rect 13092 16836 13096 16892
rect 13032 16832 13096 16836
rect 13112 16892 13176 16896
rect 13112 16836 13116 16892
rect 13116 16836 13172 16892
rect 13172 16836 13176 16892
rect 13112 16832 13176 16836
rect 13192 16892 13256 16896
rect 13192 16836 13196 16892
rect 13196 16836 13252 16892
rect 13252 16836 13256 16892
rect 13192 16832 13256 16836
rect 22952 16892 23016 16896
rect 22952 16836 22956 16892
rect 22956 16836 23012 16892
rect 23012 16836 23016 16892
rect 22952 16832 23016 16836
rect 23032 16892 23096 16896
rect 23032 16836 23036 16892
rect 23036 16836 23092 16892
rect 23092 16836 23096 16892
rect 23032 16832 23096 16836
rect 23112 16892 23176 16896
rect 23112 16836 23116 16892
rect 23116 16836 23172 16892
rect 23172 16836 23176 16892
rect 23112 16832 23176 16836
rect 23192 16892 23256 16896
rect 23192 16836 23196 16892
rect 23196 16836 23252 16892
rect 23252 16836 23256 16892
rect 23192 16832 23256 16836
rect 7952 16348 8016 16352
rect 7952 16292 7956 16348
rect 7956 16292 8012 16348
rect 8012 16292 8016 16348
rect 7952 16288 8016 16292
rect 8032 16348 8096 16352
rect 8032 16292 8036 16348
rect 8036 16292 8092 16348
rect 8092 16292 8096 16348
rect 8032 16288 8096 16292
rect 8112 16348 8176 16352
rect 8112 16292 8116 16348
rect 8116 16292 8172 16348
rect 8172 16292 8176 16348
rect 8112 16288 8176 16292
rect 8192 16348 8256 16352
rect 8192 16292 8196 16348
rect 8196 16292 8252 16348
rect 8252 16292 8256 16348
rect 8192 16288 8256 16292
rect 17952 16348 18016 16352
rect 17952 16292 17956 16348
rect 17956 16292 18012 16348
rect 18012 16292 18016 16348
rect 17952 16288 18016 16292
rect 18032 16348 18096 16352
rect 18032 16292 18036 16348
rect 18036 16292 18092 16348
rect 18092 16292 18096 16348
rect 18032 16288 18096 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 13492 15948 13556 16012
rect 2952 15804 3016 15808
rect 2952 15748 2956 15804
rect 2956 15748 3012 15804
rect 3012 15748 3016 15804
rect 2952 15744 3016 15748
rect 3032 15804 3096 15808
rect 3032 15748 3036 15804
rect 3036 15748 3092 15804
rect 3092 15748 3096 15804
rect 3032 15744 3096 15748
rect 3112 15804 3176 15808
rect 3112 15748 3116 15804
rect 3116 15748 3172 15804
rect 3172 15748 3176 15804
rect 3112 15744 3176 15748
rect 3192 15804 3256 15808
rect 3192 15748 3196 15804
rect 3196 15748 3252 15804
rect 3252 15748 3256 15804
rect 3192 15744 3256 15748
rect 12952 15804 13016 15808
rect 12952 15748 12956 15804
rect 12956 15748 13012 15804
rect 13012 15748 13016 15804
rect 12952 15744 13016 15748
rect 13032 15804 13096 15808
rect 13032 15748 13036 15804
rect 13036 15748 13092 15804
rect 13092 15748 13096 15804
rect 13032 15744 13096 15748
rect 13112 15804 13176 15808
rect 13112 15748 13116 15804
rect 13116 15748 13172 15804
rect 13172 15748 13176 15804
rect 13112 15744 13176 15748
rect 13192 15804 13256 15808
rect 13192 15748 13196 15804
rect 13196 15748 13252 15804
rect 13252 15748 13256 15804
rect 13192 15744 13256 15748
rect 22952 15804 23016 15808
rect 22952 15748 22956 15804
rect 22956 15748 23012 15804
rect 23012 15748 23016 15804
rect 22952 15744 23016 15748
rect 23032 15804 23096 15808
rect 23032 15748 23036 15804
rect 23036 15748 23092 15804
rect 23092 15748 23096 15804
rect 23032 15744 23096 15748
rect 23112 15804 23176 15808
rect 23112 15748 23116 15804
rect 23116 15748 23172 15804
rect 23172 15748 23176 15804
rect 23112 15744 23176 15748
rect 23192 15804 23256 15808
rect 23192 15748 23196 15804
rect 23196 15748 23252 15804
rect 23252 15748 23256 15804
rect 23192 15744 23256 15748
rect 13860 15268 13924 15332
rect 15700 15268 15764 15332
rect 7952 15260 8016 15264
rect 7952 15204 7956 15260
rect 7956 15204 8012 15260
rect 8012 15204 8016 15260
rect 7952 15200 8016 15204
rect 8032 15260 8096 15264
rect 8032 15204 8036 15260
rect 8036 15204 8092 15260
rect 8092 15204 8096 15260
rect 8032 15200 8096 15204
rect 8112 15260 8176 15264
rect 8112 15204 8116 15260
rect 8116 15204 8172 15260
rect 8172 15204 8176 15260
rect 8112 15200 8176 15204
rect 8192 15260 8256 15264
rect 8192 15204 8196 15260
rect 8196 15204 8252 15260
rect 8252 15204 8256 15260
rect 8192 15200 8256 15204
rect 17952 15260 18016 15264
rect 17952 15204 17956 15260
rect 17956 15204 18012 15260
rect 18012 15204 18016 15260
rect 17952 15200 18016 15204
rect 18032 15260 18096 15264
rect 18032 15204 18036 15260
rect 18036 15204 18092 15260
rect 18092 15204 18096 15260
rect 18032 15200 18096 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 2952 14716 3016 14720
rect 2952 14660 2956 14716
rect 2956 14660 3012 14716
rect 3012 14660 3016 14716
rect 2952 14656 3016 14660
rect 3032 14716 3096 14720
rect 3032 14660 3036 14716
rect 3036 14660 3092 14716
rect 3092 14660 3096 14716
rect 3032 14656 3096 14660
rect 3112 14716 3176 14720
rect 3112 14660 3116 14716
rect 3116 14660 3172 14716
rect 3172 14660 3176 14716
rect 3112 14656 3176 14660
rect 3192 14716 3256 14720
rect 3192 14660 3196 14716
rect 3196 14660 3252 14716
rect 3252 14660 3256 14716
rect 3192 14656 3256 14660
rect 12952 14716 13016 14720
rect 12952 14660 12956 14716
rect 12956 14660 13012 14716
rect 13012 14660 13016 14716
rect 12952 14656 13016 14660
rect 13032 14716 13096 14720
rect 13032 14660 13036 14716
rect 13036 14660 13092 14716
rect 13092 14660 13096 14716
rect 13032 14656 13096 14660
rect 13112 14716 13176 14720
rect 13112 14660 13116 14716
rect 13116 14660 13172 14716
rect 13172 14660 13176 14716
rect 13112 14656 13176 14660
rect 13192 14716 13256 14720
rect 13192 14660 13196 14716
rect 13196 14660 13252 14716
rect 13252 14660 13256 14716
rect 13192 14656 13256 14660
rect 22952 14716 23016 14720
rect 22952 14660 22956 14716
rect 22956 14660 23012 14716
rect 23012 14660 23016 14716
rect 22952 14656 23016 14660
rect 23032 14716 23096 14720
rect 23032 14660 23036 14716
rect 23036 14660 23092 14716
rect 23092 14660 23096 14716
rect 23032 14656 23096 14660
rect 23112 14716 23176 14720
rect 23112 14660 23116 14716
rect 23116 14660 23172 14716
rect 23172 14660 23176 14716
rect 23112 14656 23176 14660
rect 23192 14716 23256 14720
rect 23192 14660 23196 14716
rect 23196 14660 23252 14716
rect 23252 14660 23256 14716
rect 23192 14656 23256 14660
rect 7952 14172 8016 14176
rect 7952 14116 7956 14172
rect 7956 14116 8012 14172
rect 8012 14116 8016 14172
rect 7952 14112 8016 14116
rect 8032 14172 8096 14176
rect 8032 14116 8036 14172
rect 8036 14116 8092 14172
rect 8092 14116 8096 14172
rect 8032 14112 8096 14116
rect 8112 14172 8176 14176
rect 8112 14116 8116 14172
rect 8116 14116 8172 14172
rect 8172 14116 8176 14172
rect 8112 14112 8176 14116
rect 8192 14172 8256 14176
rect 8192 14116 8196 14172
rect 8196 14116 8252 14172
rect 8252 14116 8256 14172
rect 8192 14112 8256 14116
rect 17952 14172 18016 14176
rect 17952 14116 17956 14172
rect 17956 14116 18012 14172
rect 18012 14116 18016 14172
rect 17952 14112 18016 14116
rect 18032 14172 18096 14176
rect 18032 14116 18036 14172
rect 18036 14116 18092 14172
rect 18092 14116 18096 14172
rect 18032 14112 18096 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 2952 13628 3016 13632
rect 2952 13572 2956 13628
rect 2956 13572 3012 13628
rect 3012 13572 3016 13628
rect 2952 13568 3016 13572
rect 3032 13628 3096 13632
rect 3032 13572 3036 13628
rect 3036 13572 3092 13628
rect 3092 13572 3096 13628
rect 3032 13568 3096 13572
rect 3112 13628 3176 13632
rect 3112 13572 3116 13628
rect 3116 13572 3172 13628
rect 3172 13572 3176 13628
rect 3112 13568 3176 13572
rect 3192 13628 3256 13632
rect 3192 13572 3196 13628
rect 3196 13572 3252 13628
rect 3252 13572 3256 13628
rect 3192 13568 3256 13572
rect 12952 13628 13016 13632
rect 12952 13572 12956 13628
rect 12956 13572 13012 13628
rect 13012 13572 13016 13628
rect 12952 13568 13016 13572
rect 13032 13628 13096 13632
rect 13032 13572 13036 13628
rect 13036 13572 13092 13628
rect 13092 13572 13096 13628
rect 13032 13568 13096 13572
rect 13112 13628 13176 13632
rect 13112 13572 13116 13628
rect 13116 13572 13172 13628
rect 13172 13572 13176 13628
rect 13112 13568 13176 13572
rect 13192 13628 13256 13632
rect 13192 13572 13196 13628
rect 13196 13572 13252 13628
rect 13252 13572 13256 13628
rect 13192 13568 13256 13572
rect 22952 13628 23016 13632
rect 22952 13572 22956 13628
rect 22956 13572 23012 13628
rect 23012 13572 23016 13628
rect 22952 13568 23016 13572
rect 23032 13628 23096 13632
rect 23032 13572 23036 13628
rect 23036 13572 23092 13628
rect 23092 13572 23096 13628
rect 23032 13568 23096 13572
rect 23112 13628 23176 13632
rect 23112 13572 23116 13628
rect 23116 13572 23172 13628
rect 23172 13572 23176 13628
rect 23112 13568 23176 13572
rect 23192 13628 23256 13632
rect 23192 13572 23196 13628
rect 23196 13572 23252 13628
rect 23252 13572 23256 13628
rect 23192 13568 23256 13572
rect 19564 13500 19628 13564
rect 7952 13084 8016 13088
rect 7952 13028 7956 13084
rect 7956 13028 8012 13084
rect 8012 13028 8016 13084
rect 7952 13024 8016 13028
rect 8032 13084 8096 13088
rect 8032 13028 8036 13084
rect 8036 13028 8092 13084
rect 8092 13028 8096 13084
rect 8032 13024 8096 13028
rect 8112 13084 8176 13088
rect 8112 13028 8116 13084
rect 8116 13028 8172 13084
rect 8172 13028 8176 13084
rect 8112 13024 8176 13028
rect 8192 13084 8256 13088
rect 8192 13028 8196 13084
rect 8196 13028 8252 13084
rect 8252 13028 8256 13084
rect 8192 13024 8256 13028
rect 17952 13084 18016 13088
rect 17952 13028 17956 13084
rect 17956 13028 18012 13084
rect 18012 13028 18016 13084
rect 17952 13024 18016 13028
rect 18032 13084 18096 13088
rect 18032 13028 18036 13084
rect 18036 13028 18092 13084
rect 18092 13028 18096 13084
rect 18032 13024 18096 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 2952 12540 3016 12544
rect 2952 12484 2956 12540
rect 2956 12484 3012 12540
rect 3012 12484 3016 12540
rect 2952 12480 3016 12484
rect 3032 12540 3096 12544
rect 3032 12484 3036 12540
rect 3036 12484 3092 12540
rect 3092 12484 3096 12540
rect 3032 12480 3096 12484
rect 3112 12540 3176 12544
rect 3112 12484 3116 12540
rect 3116 12484 3172 12540
rect 3172 12484 3176 12540
rect 3112 12480 3176 12484
rect 3192 12540 3256 12544
rect 3192 12484 3196 12540
rect 3196 12484 3252 12540
rect 3252 12484 3256 12540
rect 3192 12480 3256 12484
rect 12952 12540 13016 12544
rect 12952 12484 12956 12540
rect 12956 12484 13012 12540
rect 13012 12484 13016 12540
rect 12952 12480 13016 12484
rect 13032 12540 13096 12544
rect 13032 12484 13036 12540
rect 13036 12484 13092 12540
rect 13092 12484 13096 12540
rect 13032 12480 13096 12484
rect 13112 12540 13176 12544
rect 13112 12484 13116 12540
rect 13116 12484 13172 12540
rect 13172 12484 13176 12540
rect 13112 12480 13176 12484
rect 13192 12540 13256 12544
rect 13192 12484 13196 12540
rect 13196 12484 13252 12540
rect 13252 12484 13256 12540
rect 13192 12480 13256 12484
rect 22952 12540 23016 12544
rect 22952 12484 22956 12540
rect 22956 12484 23012 12540
rect 23012 12484 23016 12540
rect 22952 12480 23016 12484
rect 23032 12540 23096 12544
rect 23032 12484 23036 12540
rect 23036 12484 23092 12540
rect 23092 12484 23096 12540
rect 23032 12480 23096 12484
rect 23112 12540 23176 12544
rect 23112 12484 23116 12540
rect 23116 12484 23172 12540
rect 23172 12484 23176 12540
rect 23112 12480 23176 12484
rect 23192 12540 23256 12544
rect 23192 12484 23196 12540
rect 23196 12484 23252 12540
rect 23252 12484 23256 12540
rect 23192 12480 23256 12484
rect 7952 11996 8016 12000
rect 7952 11940 7956 11996
rect 7956 11940 8012 11996
rect 8012 11940 8016 11996
rect 7952 11936 8016 11940
rect 8032 11996 8096 12000
rect 8032 11940 8036 11996
rect 8036 11940 8092 11996
rect 8092 11940 8096 11996
rect 8032 11936 8096 11940
rect 8112 11996 8176 12000
rect 8112 11940 8116 11996
rect 8116 11940 8172 11996
rect 8172 11940 8176 11996
rect 8112 11936 8176 11940
rect 8192 11996 8256 12000
rect 8192 11940 8196 11996
rect 8196 11940 8252 11996
rect 8252 11940 8256 11996
rect 8192 11936 8256 11940
rect 17952 11996 18016 12000
rect 17952 11940 17956 11996
rect 17956 11940 18012 11996
rect 18012 11940 18016 11996
rect 17952 11936 18016 11940
rect 18032 11996 18096 12000
rect 18032 11940 18036 11996
rect 18036 11940 18092 11996
rect 18092 11940 18096 11996
rect 18032 11936 18096 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 2952 11452 3016 11456
rect 2952 11396 2956 11452
rect 2956 11396 3012 11452
rect 3012 11396 3016 11452
rect 2952 11392 3016 11396
rect 3032 11452 3096 11456
rect 3032 11396 3036 11452
rect 3036 11396 3092 11452
rect 3092 11396 3096 11452
rect 3032 11392 3096 11396
rect 3112 11452 3176 11456
rect 3112 11396 3116 11452
rect 3116 11396 3172 11452
rect 3172 11396 3176 11452
rect 3112 11392 3176 11396
rect 3192 11452 3256 11456
rect 3192 11396 3196 11452
rect 3196 11396 3252 11452
rect 3252 11396 3256 11452
rect 3192 11392 3256 11396
rect 12952 11452 13016 11456
rect 12952 11396 12956 11452
rect 12956 11396 13012 11452
rect 13012 11396 13016 11452
rect 12952 11392 13016 11396
rect 13032 11452 13096 11456
rect 13032 11396 13036 11452
rect 13036 11396 13092 11452
rect 13092 11396 13096 11452
rect 13032 11392 13096 11396
rect 13112 11452 13176 11456
rect 13112 11396 13116 11452
rect 13116 11396 13172 11452
rect 13172 11396 13176 11452
rect 13112 11392 13176 11396
rect 13192 11452 13256 11456
rect 13192 11396 13196 11452
rect 13196 11396 13252 11452
rect 13252 11396 13256 11452
rect 13192 11392 13256 11396
rect 22952 11452 23016 11456
rect 22952 11396 22956 11452
rect 22956 11396 23012 11452
rect 23012 11396 23016 11452
rect 22952 11392 23016 11396
rect 23032 11452 23096 11456
rect 23032 11396 23036 11452
rect 23036 11396 23092 11452
rect 23092 11396 23096 11452
rect 23032 11392 23096 11396
rect 23112 11452 23176 11456
rect 23112 11396 23116 11452
rect 23116 11396 23172 11452
rect 23172 11396 23176 11452
rect 23112 11392 23176 11396
rect 23192 11452 23256 11456
rect 23192 11396 23196 11452
rect 23196 11396 23252 11452
rect 23252 11396 23256 11452
rect 23192 11392 23256 11396
rect 7952 10908 8016 10912
rect 7952 10852 7956 10908
rect 7956 10852 8012 10908
rect 8012 10852 8016 10908
rect 7952 10848 8016 10852
rect 8032 10908 8096 10912
rect 8032 10852 8036 10908
rect 8036 10852 8092 10908
rect 8092 10852 8096 10908
rect 8032 10848 8096 10852
rect 8112 10908 8176 10912
rect 8112 10852 8116 10908
rect 8116 10852 8172 10908
rect 8172 10852 8176 10908
rect 8112 10848 8176 10852
rect 8192 10908 8256 10912
rect 8192 10852 8196 10908
rect 8196 10852 8252 10908
rect 8252 10852 8256 10908
rect 8192 10848 8256 10852
rect 17952 10908 18016 10912
rect 17952 10852 17956 10908
rect 17956 10852 18012 10908
rect 18012 10852 18016 10908
rect 17952 10848 18016 10852
rect 18032 10908 18096 10912
rect 18032 10852 18036 10908
rect 18036 10852 18092 10908
rect 18092 10852 18096 10908
rect 18032 10848 18096 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 2952 10364 3016 10368
rect 2952 10308 2956 10364
rect 2956 10308 3012 10364
rect 3012 10308 3016 10364
rect 2952 10304 3016 10308
rect 3032 10364 3096 10368
rect 3032 10308 3036 10364
rect 3036 10308 3092 10364
rect 3092 10308 3096 10364
rect 3032 10304 3096 10308
rect 3112 10364 3176 10368
rect 3112 10308 3116 10364
rect 3116 10308 3172 10364
rect 3172 10308 3176 10364
rect 3112 10304 3176 10308
rect 3192 10364 3256 10368
rect 3192 10308 3196 10364
rect 3196 10308 3252 10364
rect 3252 10308 3256 10364
rect 3192 10304 3256 10308
rect 12952 10364 13016 10368
rect 12952 10308 12956 10364
rect 12956 10308 13012 10364
rect 13012 10308 13016 10364
rect 12952 10304 13016 10308
rect 13032 10364 13096 10368
rect 13032 10308 13036 10364
rect 13036 10308 13092 10364
rect 13092 10308 13096 10364
rect 13032 10304 13096 10308
rect 13112 10364 13176 10368
rect 13112 10308 13116 10364
rect 13116 10308 13172 10364
rect 13172 10308 13176 10364
rect 13112 10304 13176 10308
rect 13192 10364 13256 10368
rect 13192 10308 13196 10364
rect 13196 10308 13252 10364
rect 13252 10308 13256 10364
rect 13192 10304 13256 10308
rect 22952 10364 23016 10368
rect 22952 10308 22956 10364
rect 22956 10308 23012 10364
rect 23012 10308 23016 10364
rect 22952 10304 23016 10308
rect 23032 10364 23096 10368
rect 23032 10308 23036 10364
rect 23036 10308 23092 10364
rect 23092 10308 23096 10364
rect 23032 10304 23096 10308
rect 23112 10364 23176 10368
rect 23112 10308 23116 10364
rect 23116 10308 23172 10364
rect 23172 10308 23176 10364
rect 23112 10304 23176 10308
rect 23192 10364 23256 10368
rect 23192 10308 23196 10364
rect 23196 10308 23252 10364
rect 23252 10308 23256 10364
rect 23192 10304 23256 10308
rect 7952 9820 8016 9824
rect 7952 9764 7956 9820
rect 7956 9764 8012 9820
rect 8012 9764 8016 9820
rect 7952 9760 8016 9764
rect 8032 9820 8096 9824
rect 8032 9764 8036 9820
rect 8036 9764 8092 9820
rect 8092 9764 8096 9820
rect 8032 9760 8096 9764
rect 8112 9820 8176 9824
rect 8112 9764 8116 9820
rect 8116 9764 8172 9820
rect 8172 9764 8176 9820
rect 8112 9760 8176 9764
rect 8192 9820 8256 9824
rect 8192 9764 8196 9820
rect 8196 9764 8252 9820
rect 8252 9764 8256 9820
rect 8192 9760 8256 9764
rect 17952 9820 18016 9824
rect 17952 9764 17956 9820
rect 17956 9764 18012 9820
rect 18012 9764 18016 9820
rect 17952 9760 18016 9764
rect 18032 9820 18096 9824
rect 18032 9764 18036 9820
rect 18036 9764 18092 9820
rect 18092 9764 18096 9820
rect 18032 9760 18096 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 2952 9276 3016 9280
rect 2952 9220 2956 9276
rect 2956 9220 3012 9276
rect 3012 9220 3016 9276
rect 2952 9216 3016 9220
rect 3032 9276 3096 9280
rect 3032 9220 3036 9276
rect 3036 9220 3092 9276
rect 3092 9220 3096 9276
rect 3032 9216 3096 9220
rect 3112 9276 3176 9280
rect 3112 9220 3116 9276
rect 3116 9220 3172 9276
rect 3172 9220 3176 9276
rect 3112 9216 3176 9220
rect 3192 9276 3256 9280
rect 3192 9220 3196 9276
rect 3196 9220 3252 9276
rect 3252 9220 3256 9276
rect 3192 9216 3256 9220
rect 12952 9276 13016 9280
rect 12952 9220 12956 9276
rect 12956 9220 13012 9276
rect 13012 9220 13016 9276
rect 12952 9216 13016 9220
rect 13032 9276 13096 9280
rect 13032 9220 13036 9276
rect 13036 9220 13092 9276
rect 13092 9220 13096 9276
rect 13032 9216 13096 9220
rect 13112 9276 13176 9280
rect 13112 9220 13116 9276
rect 13116 9220 13172 9276
rect 13172 9220 13176 9276
rect 13112 9216 13176 9220
rect 13192 9276 13256 9280
rect 13192 9220 13196 9276
rect 13196 9220 13252 9276
rect 13252 9220 13256 9276
rect 13192 9216 13256 9220
rect 22952 9276 23016 9280
rect 22952 9220 22956 9276
rect 22956 9220 23012 9276
rect 23012 9220 23016 9276
rect 22952 9216 23016 9220
rect 23032 9276 23096 9280
rect 23032 9220 23036 9276
rect 23036 9220 23092 9276
rect 23092 9220 23096 9276
rect 23032 9216 23096 9220
rect 23112 9276 23176 9280
rect 23112 9220 23116 9276
rect 23116 9220 23172 9276
rect 23172 9220 23176 9276
rect 23112 9216 23176 9220
rect 23192 9276 23256 9280
rect 23192 9220 23196 9276
rect 23196 9220 23252 9276
rect 23252 9220 23256 9276
rect 23192 9216 23256 9220
rect 7952 8732 8016 8736
rect 7952 8676 7956 8732
rect 7956 8676 8012 8732
rect 8012 8676 8016 8732
rect 7952 8672 8016 8676
rect 8032 8732 8096 8736
rect 8032 8676 8036 8732
rect 8036 8676 8092 8732
rect 8092 8676 8096 8732
rect 8032 8672 8096 8676
rect 8112 8732 8176 8736
rect 8112 8676 8116 8732
rect 8116 8676 8172 8732
rect 8172 8676 8176 8732
rect 8112 8672 8176 8676
rect 8192 8732 8256 8736
rect 8192 8676 8196 8732
rect 8196 8676 8252 8732
rect 8252 8676 8256 8732
rect 8192 8672 8256 8676
rect 17952 8732 18016 8736
rect 17952 8676 17956 8732
rect 17956 8676 18012 8732
rect 18012 8676 18016 8732
rect 17952 8672 18016 8676
rect 18032 8732 18096 8736
rect 18032 8676 18036 8732
rect 18036 8676 18092 8732
rect 18092 8676 18096 8732
rect 18032 8672 18096 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 2952 8188 3016 8192
rect 2952 8132 2956 8188
rect 2956 8132 3012 8188
rect 3012 8132 3016 8188
rect 2952 8128 3016 8132
rect 3032 8188 3096 8192
rect 3032 8132 3036 8188
rect 3036 8132 3092 8188
rect 3092 8132 3096 8188
rect 3032 8128 3096 8132
rect 3112 8188 3176 8192
rect 3112 8132 3116 8188
rect 3116 8132 3172 8188
rect 3172 8132 3176 8188
rect 3112 8128 3176 8132
rect 3192 8188 3256 8192
rect 3192 8132 3196 8188
rect 3196 8132 3252 8188
rect 3252 8132 3256 8188
rect 3192 8128 3256 8132
rect 12952 8188 13016 8192
rect 12952 8132 12956 8188
rect 12956 8132 13012 8188
rect 13012 8132 13016 8188
rect 12952 8128 13016 8132
rect 13032 8188 13096 8192
rect 13032 8132 13036 8188
rect 13036 8132 13092 8188
rect 13092 8132 13096 8188
rect 13032 8128 13096 8132
rect 13112 8188 13176 8192
rect 13112 8132 13116 8188
rect 13116 8132 13172 8188
rect 13172 8132 13176 8188
rect 13112 8128 13176 8132
rect 13192 8188 13256 8192
rect 13192 8132 13196 8188
rect 13196 8132 13252 8188
rect 13252 8132 13256 8188
rect 13192 8128 13256 8132
rect 22952 8188 23016 8192
rect 22952 8132 22956 8188
rect 22956 8132 23012 8188
rect 23012 8132 23016 8188
rect 22952 8128 23016 8132
rect 23032 8188 23096 8192
rect 23032 8132 23036 8188
rect 23036 8132 23092 8188
rect 23092 8132 23096 8188
rect 23032 8128 23096 8132
rect 23112 8188 23176 8192
rect 23112 8132 23116 8188
rect 23116 8132 23172 8188
rect 23172 8132 23176 8188
rect 23112 8128 23176 8132
rect 23192 8188 23256 8192
rect 23192 8132 23196 8188
rect 23196 8132 23252 8188
rect 23252 8132 23256 8188
rect 23192 8128 23256 8132
rect 7952 7644 8016 7648
rect 7952 7588 7956 7644
rect 7956 7588 8012 7644
rect 8012 7588 8016 7644
rect 7952 7584 8016 7588
rect 8032 7644 8096 7648
rect 8032 7588 8036 7644
rect 8036 7588 8092 7644
rect 8092 7588 8096 7644
rect 8032 7584 8096 7588
rect 8112 7644 8176 7648
rect 8112 7588 8116 7644
rect 8116 7588 8172 7644
rect 8172 7588 8176 7644
rect 8112 7584 8176 7588
rect 8192 7644 8256 7648
rect 8192 7588 8196 7644
rect 8196 7588 8252 7644
rect 8252 7588 8256 7644
rect 8192 7584 8256 7588
rect 17952 7644 18016 7648
rect 17952 7588 17956 7644
rect 17956 7588 18012 7644
rect 18012 7588 18016 7644
rect 17952 7584 18016 7588
rect 18032 7644 18096 7648
rect 18032 7588 18036 7644
rect 18036 7588 18092 7644
rect 18092 7588 18096 7644
rect 18032 7584 18096 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 2952 7100 3016 7104
rect 2952 7044 2956 7100
rect 2956 7044 3012 7100
rect 3012 7044 3016 7100
rect 2952 7040 3016 7044
rect 3032 7100 3096 7104
rect 3032 7044 3036 7100
rect 3036 7044 3092 7100
rect 3092 7044 3096 7100
rect 3032 7040 3096 7044
rect 3112 7100 3176 7104
rect 3112 7044 3116 7100
rect 3116 7044 3172 7100
rect 3172 7044 3176 7100
rect 3112 7040 3176 7044
rect 3192 7100 3256 7104
rect 3192 7044 3196 7100
rect 3196 7044 3252 7100
rect 3252 7044 3256 7100
rect 3192 7040 3256 7044
rect 12952 7100 13016 7104
rect 12952 7044 12956 7100
rect 12956 7044 13012 7100
rect 13012 7044 13016 7100
rect 12952 7040 13016 7044
rect 13032 7100 13096 7104
rect 13032 7044 13036 7100
rect 13036 7044 13092 7100
rect 13092 7044 13096 7100
rect 13032 7040 13096 7044
rect 13112 7100 13176 7104
rect 13112 7044 13116 7100
rect 13116 7044 13172 7100
rect 13172 7044 13176 7100
rect 13112 7040 13176 7044
rect 13192 7100 13256 7104
rect 13192 7044 13196 7100
rect 13196 7044 13252 7100
rect 13252 7044 13256 7100
rect 13192 7040 13256 7044
rect 22952 7100 23016 7104
rect 22952 7044 22956 7100
rect 22956 7044 23012 7100
rect 23012 7044 23016 7100
rect 22952 7040 23016 7044
rect 23032 7100 23096 7104
rect 23032 7044 23036 7100
rect 23036 7044 23092 7100
rect 23092 7044 23096 7100
rect 23032 7040 23096 7044
rect 23112 7100 23176 7104
rect 23112 7044 23116 7100
rect 23116 7044 23172 7100
rect 23172 7044 23176 7100
rect 23112 7040 23176 7044
rect 23192 7100 23256 7104
rect 23192 7044 23196 7100
rect 23196 7044 23252 7100
rect 23252 7044 23256 7100
rect 23192 7040 23256 7044
rect 7952 6556 8016 6560
rect 7952 6500 7956 6556
rect 7956 6500 8012 6556
rect 8012 6500 8016 6556
rect 7952 6496 8016 6500
rect 8032 6556 8096 6560
rect 8032 6500 8036 6556
rect 8036 6500 8092 6556
rect 8092 6500 8096 6556
rect 8032 6496 8096 6500
rect 8112 6556 8176 6560
rect 8112 6500 8116 6556
rect 8116 6500 8172 6556
rect 8172 6500 8176 6556
rect 8112 6496 8176 6500
rect 8192 6556 8256 6560
rect 8192 6500 8196 6556
rect 8196 6500 8252 6556
rect 8252 6500 8256 6556
rect 8192 6496 8256 6500
rect 17952 6556 18016 6560
rect 17952 6500 17956 6556
rect 17956 6500 18012 6556
rect 18012 6500 18016 6556
rect 17952 6496 18016 6500
rect 18032 6556 18096 6560
rect 18032 6500 18036 6556
rect 18036 6500 18092 6556
rect 18092 6500 18096 6556
rect 18032 6496 18096 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 2952 6012 3016 6016
rect 2952 5956 2956 6012
rect 2956 5956 3012 6012
rect 3012 5956 3016 6012
rect 2952 5952 3016 5956
rect 3032 6012 3096 6016
rect 3032 5956 3036 6012
rect 3036 5956 3092 6012
rect 3092 5956 3096 6012
rect 3032 5952 3096 5956
rect 3112 6012 3176 6016
rect 3112 5956 3116 6012
rect 3116 5956 3172 6012
rect 3172 5956 3176 6012
rect 3112 5952 3176 5956
rect 3192 6012 3256 6016
rect 3192 5956 3196 6012
rect 3196 5956 3252 6012
rect 3252 5956 3256 6012
rect 3192 5952 3256 5956
rect 12952 6012 13016 6016
rect 12952 5956 12956 6012
rect 12956 5956 13012 6012
rect 13012 5956 13016 6012
rect 12952 5952 13016 5956
rect 13032 6012 13096 6016
rect 13032 5956 13036 6012
rect 13036 5956 13092 6012
rect 13092 5956 13096 6012
rect 13032 5952 13096 5956
rect 13112 6012 13176 6016
rect 13112 5956 13116 6012
rect 13116 5956 13172 6012
rect 13172 5956 13176 6012
rect 13112 5952 13176 5956
rect 13192 6012 13256 6016
rect 13192 5956 13196 6012
rect 13196 5956 13252 6012
rect 13252 5956 13256 6012
rect 13192 5952 13256 5956
rect 22952 6012 23016 6016
rect 22952 5956 22956 6012
rect 22956 5956 23012 6012
rect 23012 5956 23016 6012
rect 22952 5952 23016 5956
rect 23032 6012 23096 6016
rect 23032 5956 23036 6012
rect 23036 5956 23092 6012
rect 23092 5956 23096 6012
rect 23032 5952 23096 5956
rect 23112 6012 23176 6016
rect 23112 5956 23116 6012
rect 23116 5956 23172 6012
rect 23172 5956 23176 6012
rect 23112 5952 23176 5956
rect 23192 6012 23256 6016
rect 23192 5956 23196 6012
rect 23196 5956 23252 6012
rect 23252 5956 23256 6012
rect 23192 5952 23256 5956
rect 14964 5748 15028 5812
rect 10180 5612 10244 5676
rect 7952 5468 8016 5472
rect 7952 5412 7956 5468
rect 7956 5412 8012 5468
rect 8012 5412 8016 5468
rect 7952 5408 8016 5412
rect 8032 5468 8096 5472
rect 8032 5412 8036 5468
rect 8036 5412 8092 5468
rect 8092 5412 8096 5468
rect 8032 5408 8096 5412
rect 8112 5468 8176 5472
rect 8112 5412 8116 5468
rect 8116 5412 8172 5468
rect 8172 5412 8176 5468
rect 8112 5408 8176 5412
rect 8192 5468 8256 5472
rect 8192 5412 8196 5468
rect 8196 5412 8252 5468
rect 8252 5412 8256 5468
rect 8192 5408 8256 5412
rect 17952 5468 18016 5472
rect 17952 5412 17956 5468
rect 17956 5412 18012 5468
rect 18012 5412 18016 5468
rect 17952 5408 18016 5412
rect 18032 5468 18096 5472
rect 18032 5412 18036 5468
rect 18036 5412 18092 5468
rect 18092 5412 18096 5468
rect 18032 5408 18096 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 2952 4924 3016 4928
rect 2952 4868 2956 4924
rect 2956 4868 3012 4924
rect 3012 4868 3016 4924
rect 2952 4864 3016 4868
rect 3032 4924 3096 4928
rect 3032 4868 3036 4924
rect 3036 4868 3092 4924
rect 3092 4868 3096 4924
rect 3032 4864 3096 4868
rect 3112 4924 3176 4928
rect 3112 4868 3116 4924
rect 3116 4868 3172 4924
rect 3172 4868 3176 4924
rect 3112 4864 3176 4868
rect 3192 4924 3256 4928
rect 3192 4868 3196 4924
rect 3196 4868 3252 4924
rect 3252 4868 3256 4924
rect 3192 4864 3256 4868
rect 12952 4924 13016 4928
rect 12952 4868 12956 4924
rect 12956 4868 13012 4924
rect 13012 4868 13016 4924
rect 12952 4864 13016 4868
rect 13032 4924 13096 4928
rect 13032 4868 13036 4924
rect 13036 4868 13092 4924
rect 13092 4868 13096 4924
rect 13032 4864 13096 4868
rect 13112 4924 13176 4928
rect 13112 4868 13116 4924
rect 13116 4868 13172 4924
rect 13172 4868 13176 4924
rect 13112 4864 13176 4868
rect 13192 4924 13256 4928
rect 13192 4868 13196 4924
rect 13196 4868 13252 4924
rect 13252 4868 13256 4924
rect 13192 4864 13256 4868
rect 22952 4924 23016 4928
rect 22952 4868 22956 4924
rect 22956 4868 23012 4924
rect 23012 4868 23016 4924
rect 22952 4864 23016 4868
rect 23032 4924 23096 4928
rect 23032 4868 23036 4924
rect 23036 4868 23092 4924
rect 23092 4868 23096 4924
rect 23032 4864 23096 4868
rect 23112 4924 23176 4928
rect 23112 4868 23116 4924
rect 23116 4868 23172 4924
rect 23172 4868 23176 4924
rect 23112 4864 23176 4868
rect 23192 4924 23256 4928
rect 23192 4868 23196 4924
rect 23196 4868 23252 4924
rect 23252 4868 23256 4924
rect 23192 4864 23256 4868
rect 7952 4380 8016 4384
rect 7952 4324 7956 4380
rect 7956 4324 8012 4380
rect 8012 4324 8016 4380
rect 7952 4320 8016 4324
rect 8032 4380 8096 4384
rect 8032 4324 8036 4380
rect 8036 4324 8092 4380
rect 8092 4324 8096 4380
rect 8032 4320 8096 4324
rect 8112 4380 8176 4384
rect 8112 4324 8116 4380
rect 8116 4324 8172 4380
rect 8172 4324 8176 4380
rect 8112 4320 8176 4324
rect 8192 4380 8256 4384
rect 8192 4324 8196 4380
rect 8196 4324 8252 4380
rect 8252 4324 8256 4380
rect 8192 4320 8256 4324
rect 17952 4380 18016 4384
rect 17952 4324 17956 4380
rect 17956 4324 18012 4380
rect 18012 4324 18016 4380
rect 17952 4320 18016 4324
rect 18032 4380 18096 4384
rect 18032 4324 18036 4380
rect 18036 4324 18092 4380
rect 18092 4324 18096 4380
rect 18032 4320 18096 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 2952 3836 3016 3840
rect 2952 3780 2956 3836
rect 2956 3780 3012 3836
rect 3012 3780 3016 3836
rect 2952 3776 3016 3780
rect 3032 3836 3096 3840
rect 3032 3780 3036 3836
rect 3036 3780 3092 3836
rect 3092 3780 3096 3836
rect 3032 3776 3096 3780
rect 3112 3836 3176 3840
rect 3112 3780 3116 3836
rect 3116 3780 3172 3836
rect 3172 3780 3176 3836
rect 3112 3776 3176 3780
rect 3192 3836 3256 3840
rect 3192 3780 3196 3836
rect 3196 3780 3252 3836
rect 3252 3780 3256 3836
rect 3192 3776 3256 3780
rect 12952 3836 13016 3840
rect 12952 3780 12956 3836
rect 12956 3780 13012 3836
rect 13012 3780 13016 3836
rect 12952 3776 13016 3780
rect 13032 3836 13096 3840
rect 13032 3780 13036 3836
rect 13036 3780 13092 3836
rect 13092 3780 13096 3836
rect 13032 3776 13096 3780
rect 13112 3836 13176 3840
rect 13112 3780 13116 3836
rect 13116 3780 13172 3836
rect 13172 3780 13176 3836
rect 13112 3776 13176 3780
rect 13192 3836 13256 3840
rect 13192 3780 13196 3836
rect 13196 3780 13252 3836
rect 13252 3780 13256 3836
rect 13192 3776 13256 3780
rect 22952 3836 23016 3840
rect 22952 3780 22956 3836
rect 22956 3780 23012 3836
rect 23012 3780 23016 3836
rect 22952 3776 23016 3780
rect 23032 3836 23096 3840
rect 23032 3780 23036 3836
rect 23036 3780 23092 3836
rect 23092 3780 23096 3836
rect 23032 3776 23096 3780
rect 23112 3836 23176 3840
rect 23112 3780 23116 3836
rect 23116 3780 23172 3836
rect 23172 3780 23176 3836
rect 23112 3776 23176 3780
rect 23192 3836 23256 3840
rect 23192 3780 23196 3836
rect 23196 3780 23252 3836
rect 23252 3780 23256 3836
rect 23192 3776 23256 3780
rect 16804 3436 16868 3500
rect 7952 3292 8016 3296
rect 7952 3236 7956 3292
rect 7956 3236 8012 3292
rect 8012 3236 8016 3292
rect 7952 3232 8016 3236
rect 8032 3292 8096 3296
rect 8032 3236 8036 3292
rect 8036 3236 8092 3292
rect 8092 3236 8096 3292
rect 8032 3232 8096 3236
rect 8112 3292 8176 3296
rect 8112 3236 8116 3292
rect 8116 3236 8172 3292
rect 8172 3236 8176 3292
rect 8112 3232 8176 3236
rect 8192 3292 8256 3296
rect 8192 3236 8196 3292
rect 8196 3236 8252 3292
rect 8252 3236 8256 3292
rect 8192 3232 8256 3236
rect 17952 3292 18016 3296
rect 17952 3236 17956 3292
rect 17956 3236 18012 3292
rect 18012 3236 18016 3292
rect 17952 3232 18016 3236
rect 18032 3292 18096 3296
rect 18032 3236 18036 3292
rect 18036 3236 18092 3292
rect 18092 3236 18096 3292
rect 18032 3232 18096 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 2952 2748 3016 2752
rect 2952 2692 2956 2748
rect 2956 2692 3012 2748
rect 3012 2692 3016 2748
rect 2952 2688 3016 2692
rect 3032 2748 3096 2752
rect 3032 2692 3036 2748
rect 3036 2692 3092 2748
rect 3092 2692 3096 2748
rect 3032 2688 3096 2692
rect 3112 2748 3176 2752
rect 3112 2692 3116 2748
rect 3116 2692 3172 2748
rect 3172 2692 3176 2748
rect 3112 2688 3176 2692
rect 3192 2748 3256 2752
rect 3192 2692 3196 2748
rect 3196 2692 3252 2748
rect 3252 2692 3256 2748
rect 3192 2688 3256 2692
rect 12952 2748 13016 2752
rect 12952 2692 12956 2748
rect 12956 2692 13012 2748
rect 13012 2692 13016 2748
rect 12952 2688 13016 2692
rect 13032 2748 13096 2752
rect 13032 2692 13036 2748
rect 13036 2692 13092 2748
rect 13092 2692 13096 2748
rect 13032 2688 13096 2692
rect 13112 2748 13176 2752
rect 13112 2692 13116 2748
rect 13116 2692 13172 2748
rect 13172 2692 13176 2748
rect 13112 2688 13176 2692
rect 13192 2748 13256 2752
rect 13192 2692 13196 2748
rect 13196 2692 13252 2748
rect 13252 2692 13256 2748
rect 13192 2688 13256 2692
rect 22952 2748 23016 2752
rect 22952 2692 22956 2748
rect 22956 2692 23012 2748
rect 23012 2692 23016 2748
rect 22952 2688 23016 2692
rect 23032 2748 23096 2752
rect 23032 2692 23036 2748
rect 23036 2692 23092 2748
rect 23092 2692 23096 2748
rect 23032 2688 23096 2692
rect 23112 2748 23176 2752
rect 23112 2692 23116 2748
rect 23116 2692 23172 2748
rect 23172 2692 23176 2748
rect 23112 2688 23176 2692
rect 23192 2748 23256 2752
rect 23192 2692 23196 2748
rect 23196 2692 23252 2748
rect 23252 2692 23256 2748
rect 23192 2688 23256 2692
rect 15700 2680 15764 2684
rect 15700 2624 15714 2680
rect 15714 2624 15764 2680
rect 15700 2620 15764 2624
rect 7952 2204 8016 2208
rect 7952 2148 7956 2204
rect 7956 2148 8012 2204
rect 8012 2148 8016 2204
rect 7952 2144 8016 2148
rect 8032 2204 8096 2208
rect 8032 2148 8036 2204
rect 8036 2148 8092 2204
rect 8092 2148 8096 2204
rect 8032 2144 8096 2148
rect 8112 2204 8176 2208
rect 8112 2148 8116 2204
rect 8116 2148 8172 2204
rect 8172 2148 8176 2204
rect 8112 2144 8176 2148
rect 8192 2204 8256 2208
rect 8192 2148 8196 2204
rect 8196 2148 8252 2204
rect 8252 2148 8256 2204
rect 8192 2144 8256 2148
rect 17952 2204 18016 2208
rect 17952 2148 17956 2204
rect 17956 2148 18012 2204
rect 18012 2148 18016 2204
rect 17952 2144 18016 2148
rect 18032 2204 18096 2208
rect 18032 2148 18036 2204
rect 18036 2148 18092 2204
rect 18092 2148 18096 2204
rect 18032 2144 18096 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
<< metal4 >>
rect 2944 53888 3264 54448
rect 2944 53824 2952 53888
rect 3016 53824 3032 53888
rect 3096 53824 3112 53888
rect 3176 53824 3192 53888
rect 3256 53824 3264 53888
rect 2944 52800 3264 53824
rect 2944 52736 2952 52800
rect 3016 52736 3032 52800
rect 3096 52736 3112 52800
rect 3176 52736 3192 52800
rect 3256 52736 3264 52800
rect 2944 51712 3264 52736
rect 2944 51648 2952 51712
rect 3016 51648 3032 51712
rect 3096 51648 3112 51712
rect 3176 51648 3192 51712
rect 3256 51648 3264 51712
rect 2944 50624 3264 51648
rect 2944 50560 2952 50624
rect 3016 50560 3032 50624
rect 3096 50560 3112 50624
rect 3176 50560 3192 50624
rect 3256 50560 3264 50624
rect 2944 49536 3264 50560
rect 2944 49472 2952 49536
rect 3016 49472 3032 49536
rect 3096 49472 3112 49536
rect 3176 49472 3192 49536
rect 3256 49472 3264 49536
rect 2944 48448 3264 49472
rect 2944 48384 2952 48448
rect 3016 48384 3032 48448
rect 3096 48384 3112 48448
rect 3176 48384 3192 48448
rect 3256 48384 3264 48448
rect 2944 47360 3264 48384
rect 2944 47296 2952 47360
rect 3016 47296 3032 47360
rect 3096 47296 3112 47360
rect 3176 47296 3192 47360
rect 3256 47296 3264 47360
rect 2944 46272 3264 47296
rect 2944 46208 2952 46272
rect 3016 46208 3032 46272
rect 3096 46208 3112 46272
rect 3176 46208 3192 46272
rect 3256 46208 3264 46272
rect 2944 45184 3264 46208
rect 2944 45120 2952 45184
rect 3016 45120 3032 45184
rect 3096 45120 3112 45184
rect 3176 45120 3192 45184
rect 3256 45120 3264 45184
rect 2944 44096 3264 45120
rect 2944 44032 2952 44096
rect 3016 44032 3032 44096
rect 3096 44032 3112 44096
rect 3176 44032 3192 44096
rect 3256 44032 3264 44096
rect 2944 43008 3264 44032
rect 2944 42944 2952 43008
rect 3016 42944 3032 43008
rect 3096 42944 3112 43008
rect 3176 42944 3192 43008
rect 3256 42944 3264 43008
rect 2944 41920 3264 42944
rect 2944 41856 2952 41920
rect 3016 41856 3032 41920
rect 3096 41856 3112 41920
rect 3176 41856 3192 41920
rect 3256 41856 3264 41920
rect 2944 40832 3264 41856
rect 2944 40768 2952 40832
rect 3016 40768 3032 40832
rect 3096 40768 3112 40832
rect 3176 40768 3192 40832
rect 3256 40768 3264 40832
rect 2944 39744 3264 40768
rect 2944 39680 2952 39744
rect 3016 39680 3032 39744
rect 3096 39680 3112 39744
rect 3176 39680 3192 39744
rect 3256 39680 3264 39744
rect 2944 38656 3264 39680
rect 2944 38592 2952 38656
rect 3016 38592 3032 38656
rect 3096 38592 3112 38656
rect 3176 38592 3192 38656
rect 3256 38592 3264 38656
rect 2944 37568 3264 38592
rect 2944 37504 2952 37568
rect 3016 37504 3032 37568
rect 3096 37504 3112 37568
rect 3176 37504 3192 37568
rect 3256 37504 3264 37568
rect 2944 36480 3264 37504
rect 2944 36416 2952 36480
rect 3016 36416 3032 36480
rect 3096 36416 3112 36480
rect 3176 36416 3192 36480
rect 3256 36416 3264 36480
rect 2944 35392 3264 36416
rect 2944 35328 2952 35392
rect 3016 35328 3032 35392
rect 3096 35328 3112 35392
rect 3176 35328 3192 35392
rect 3256 35328 3264 35392
rect 2944 34304 3264 35328
rect 2944 34240 2952 34304
rect 3016 34240 3032 34304
rect 3096 34240 3112 34304
rect 3176 34240 3192 34304
rect 3256 34240 3264 34304
rect 2944 33216 3264 34240
rect 2944 33152 2952 33216
rect 3016 33152 3032 33216
rect 3096 33152 3112 33216
rect 3176 33152 3192 33216
rect 3256 33152 3264 33216
rect 2944 32128 3264 33152
rect 2944 32064 2952 32128
rect 3016 32064 3032 32128
rect 3096 32064 3112 32128
rect 3176 32064 3192 32128
rect 3256 32064 3264 32128
rect 2944 31040 3264 32064
rect 2944 30976 2952 31040
rect 3016 30976 3032 31040
rect 3096 30976 3112 31040
rect 3176 30976 3192 31040
rect 3256 30976 3264 31040
rect 2944 29952 3264 30976
rect 2944 29888 2952 29952
rect 3016 29888 3032 29952
rect 3096 29888 3112 29952
rect 3176 29888 3192 29952
rect 3256 29888 3264 29952
rect 2944 28864 3264 29888
rect 2944 28800 2952 28864
rect 3016 28800 3032 28864
rect 3096 28800 3112 28864
rect 3176 28800 3192 28864
rect 3256 28800 3264 28864
rect 2944 27776 3264 28800
rect 2944 27712 2952 27776
rect 3016 27712 3032 27776
rect 3096 27712 3112 27776
rect 3176 27712 3192 27776
rect 3256 27712 3264 27776
rect 2944 26688 3264 27712
rect 2944 26624 2952 26688
rect 3016 26624 3032 26688
rect 3096 26624 3112 26688
rect 3176 26624 3192 26688
rect 3256 26624 3264 26688
rect 2944 25600 3264 26624
rect 2944 25536 2952 25600
rect 3016 25536 3032 25600
rect 3096 25536 3112 25600
rect 3176 25536 3192 25600
rect 3256 25536 3264 25600
rect 2944 24512 3264 25536
rect 2944 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3264 24512
rect 2944 23424 3264 24448
rect 2944 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3264 23424
rect 2944 22336 3264 23360
rect 2944 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3264 22336
rect 2944 21248 3264 22272
rect 2944 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3264 21248
rect 2944 20160 3264 21184
rect 2944 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3264 20160
rect 2944 19072 3264 20096
rect 2944 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3264 19072
rect 2944 17984 3264 19008
rect 2944 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3264 17984
rect 2944 16896 3264 17920
rect 2944 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3264 16896
rect 2944 15808 3264 16832
rect 2944 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3264 15808
rect 2944 14720 3264 15744
rect 2944 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3264 14720
rect 2944 13632 3264 14656
rect 2944 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3264 13632
rect 2944 12544 3264 13568
rect 2944 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3264 12544
rect 2944 11456 3264 12480
rect 2944 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3264 11456
rect 2944 10368 3264 11392
rect 2944 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3264 10368
rect 2944 9280 3264 10304
rect 2944 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3264 9280
rect 2944 8192 3264 9216
rect 2944 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3264 8192
rect 2944 7104 3264 8128
rect 2944 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3264 7104
rect 2944 6016 3264 7040
rect 2944 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3264 6016
rect 2944 4928 3264 5952
rect 2944 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3264 4928
rect 2944 3840 3264 4864
rect 2944 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3264 3840
rect 2944 2752 3264 3776
rect 2944 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3264 2752
rect 2944 2128 3264 2688
rect 7944 54432 8264 54448
rect 7944 54368 7952 54432
rect 8016 54368 8032 54432
rect 8096 54368 8112 54432
rect 8176 54368 8192 54432
rect 8256 54368 8264 54432
rect 7944 53344 8264 54368
rect 7944 53280 7952 53344
rect 8016 53280 8032 53344
rect 8096 53280 8112 53344
rect 8176 53280 8192 53344
rect 8256 53280 8264 53344
rect 7944 52256 8264 53280
rect 7944 52192 7952 52256
rect 8016 52192 8032 52256
rect 8096 52192 8112 52256
rect 8176 52192 8192 52256
rect 8256 52192 8264 52256
rect 7944 51168 8264 52192
rect 7944 51104 7952 51168
rect 8016 51104 8032 51168
rect 8096 51104 8112 51168
rect 8176 51104 8192 51168
rect 8256 51104 8264 51168
rect 7944 50080 8264 51104
rect 7944 50016 7952 50080
rect 8016 50016 8032 50080
rect 8096 50016 8112 50080
rect 8176 50016 8192 50080
rect 8256 50016 8264 50080
rect 7944 48992 8264 50016
rect 7944 48928 7952 48992
rect 8016 48928 8032 48992
rect 8096 48928 8112 48992
rect 8176 48928 8192 48992
rect 8256 48928 8264 48992
rect 7944 47904 8264 48928
rect 7944 47840 7952 47904
rect 8016 47840 8032 47904
rect 8096 47840 8112 47904
rect 8176 47840 8192 47904
rect 8256 47840 8264 47904
rect 7944 46816 8264 47840
rect 7944 46752 7952 46816
rect 8016 46752 8032 46816
rect 8096 46752 8112 46816
rect 8176 46752 8192 46816
rect 8256 46752 8264 46816
rect 7944 45728 8264 46752
rect 7944 45664 7952 45728
rect 8016 45664 8032 45728
rect 8096 45664 8112 45728
rect 8176 45664 8192 45728
rect 8256 45664 8264 45728
rect 7944 44640 8264 45664
rect 12944 53888 13264 54448
rect 17944 54432 18264 54448
rect 17944 54368 17952 54432
rect 18016 54368 18032 54432
rect 18096 54368 18112 54432
rect 18176 54368 18192 54432
rect 18256 54368 18264 54432
rect 15883 53956 15949 53957
rect 15883 53892 15884 53956
rect 15948 53892 15949 53956
rect 15883 53891 15949 53892
rect 12944 53824 12952 53888
rect 13016 53824 13032 53888
rect 13096 53824 13112 53888
rect 13176 53824 13192 53888
rect 13256 53824 13264 53888
rect 12944 52800 13264 53824
rect 12944 52736 12952 52800
rect 13016 52736 13032 52800
rect 13096 52736 13112 52800
rect 13176 52736 13192 52800
rect 13256 52736 13264 52800
rect 12944 51712 13264 52736
rect 14411 52596 14477 52597
rect 14411 52532 14412 52596
rect 14476 52532 14477 52596
rect 14411 52531 14477 52532
rect 15699 52596 15765 52597
rect 15699 52532 15700 52596
rect 15764 52532 15765 52596
rect 15699 52531 15765 52532
rect 12944 51648 12952 51712
rect 13016 51648 13032 51712
rect 13096 51648 13112 51712
rect 13176 51648 13192 51712
rect 13256 51648 13264 51712
rect 12944 50624 13264 51648
rect 12944 50560 12952 50624
rect 13016 50560 13032 50624
rect 13096 50560 13112 50624
rect 13176 50560 13192 50624
rect 13256 50560 13264 50624
rect 12944 49536 13264 50560
rect 12944 49472 12952 49536
rect 13016 49472 13032 49536
rect 13096 49472 13112 49536
rect 13176 49472 13192 49536
rect 13256 49472 13264 49536
rect 12944 48448 13264 49472
rect 12944 48384 12952 48448
rect 13016 48384 13032 48448
rect 13096 48384 13112 48448
rect 13176 48384 13192 48448
rect 13256 48384 13264 48448
rect 12944 47360 13264 48384
rect 12944 47296 12952 47360
rect 13016 47296 13032 47360
rect 13096 47296 13112 47360
rect 13176 47296 13192 47360
rect 13256 47296 13264 47360
rect 12944 46272 13264 47296
rect 12944 46208 12952 46272
rect 13016 46208 13032 46272
rect 13096 46208 13112 46272
rect 13176 46208 13192 46272
rect 13256 46208 13264 46272
rect 12019 45252 12085 45253
rect 12019 45188 12020 45252
rect 12084 45188 12085 45252
rect 12019 45187 12085 45188
rect 9811 44708 9877 44709
rect 9811 44644 9812 44708
rect 9876 44644 9877 44708
rect 9811 44643 9877 44644
rect 7944 44576 7952 44640
rect 8016 44576 8032 44640
rect 8096 44576 8112 44640
rect 8176 44576 8192 44640
rect 8256 44576 8264 44640
rect 7944 43552 8264 44576
rect 7944 43488 7952 43552
rect 8016 43488 8032 43552
rect 8096 43488 8112 43552
rect 8176 43488 8192 43552
rect 8256 43488 8264 43552
rect 7944 42464 8264 43488
rect 7944 42400 7952 42464
rect 8016 42400 8032 42464
rect 8096 42400 8112 42464
rect 8176 42400 8192 42464
rect 8256 42400 8264 42464
rect 7944 41376 8264 42400
rect 7944 41312 7952 41376
rect 8016 41312 8032 41376
rect 8096 41312 8112 41376
rect 8176 41312 8192 41376
rect 8256 41312 8264 41376
rect 7944 40288 8264 41312
rect 7944 40224 7952 40288
rect 8016 40224 8032 40288
rect 8096 40224 8112 40288
rect 8176 40224 8192 40288
rect 8256 40224 8264 40288
rect 7944 39200 8264 40224
rect 7944 39136 7952 39200
rect 8016 39136 8032 39200
rect 8096 39136 8112 39200
rect 8176 39136 8192 39200
rect 8256 39136 8264 39200
rect 7944 38112 8264 39136
rect 7944 38048 7952 38112
rect 8016 38048 8032 38112
rect 8096 38048 8112 38112
rect 8176 38048 8192 38112
rect 8256 38048 8264 38112
rect 7944 37024 8264 38048
rect 7944 36960 7952 37024
rect 8016 36960 8032 37024
rect 8096 36960 8112 37024
rect 8176 36960 8192 37024
rect 8256 36960 8264 37024
rect 7944 35936 8264 36960
rect 7944 35872 7952 35936
rect 8016 35872 8032 35936
rect 8096 35872 8112 35936
rect 8176 35872 8192 35936
rect 8256 35872 8264 35936
rect 7944 34848 8264 35872
rect 7944 34784 7952 34848
rect 8016 34784 8032 34848
rect 8096 34784 8112 34848
rect 8176 34784 8192 34848
rect 8256 34784 8264 34848
rect 7944 33760 8264 34784
rect 7944 33696 7952 33760
rect 8016 33696 8032 33760
rect 8096 33696 8112 33760
rect 8176 33696 8192 33760
rect 8256 33696 8264 33760
rect 7944 32672 8264 33696
rect 7944 32608 7952 32672
rect 8016 32608 8032 32672
rect 8096 32608 8112 32672
rect 8176 32608 8192 32672
rect 8256 32608 8264 32672
rect 7944 31584 8264 32608
rect 7944 31520 7952 31584
rect 8016 31520 8032 31584
rect 8096 31520 8112 31584
rect 8176 31520 8192 31584
rect 8256 31520 8264 31584
rect 7944 30496 8264 31520
rect 9814 31381 9874 44643
rect 12022 36685 12082 45187
rect 12944 45184 13264 46208
rect 12944 45120 12952 45184
rect 13016 45120 13032 45184
rect 13096 45120 13112 45184
rect 13176 45120 13192 45184
rect 13256 45120 13264 45184
rect 12944 44096 13264 45120
rect 12944 44032 12952 44096
rect 13016 44032 13032 44096
rect 13096 44032 13112 44096
rect 13176 44032 13192 44096
rect 13256 44032 13264 44096
rect 12944 43008 13264 44032
rect 12944 42944 12952 43008
rect 13016 42944 13032 43008
rect 13096 42944 13112 43008
rect 13176 42944 13192 43008
rect 13256 42944 13264 43008
rect 12944 41920 13264 42944
rect 12944 41856 12952 41920
rect 13016 41856 13032 41920
rect 13096 41856 13112 41920
rect 13176 41856 13192 41920
rect 13256 41856 13264 41920
rect 12944 40832 13264 41856
rect 13675 41308 13741 41309
rect 13675 41244 13676 41308
rect 13740 41244 13741 41308
rect 13675 41243 13741 41244
rect 12944 40768 12952 40832
rect 13016 40768 13032 40832
rect 13096 40768 13112 40832
rect 13176 40768 13192 40832
rect 13256 40768 13264 40832
rect 12944 39744 13264 40768
rect 12944 39680 12952 39744
rect 13016 39680 13032 39744
rect 13096 39680 13112 39744
rect 13176 39680 13192 39744
rect 13256 39680 13264 39744
rect 12944 38656 13264 39680
rect 12944 38592 12952 38656
rect 13016 38592 13032 38656
rect 13096 38592 13112 38656
rect 13176 38592 13192 38656
rect 13256 38592 13264 38656
rect 12944 37568 13264 38592
rect 12944 37504 12952 37568
rect 13016 37504 13032 37568
rect 13096 37504 13112 37568
rect 13176 37504 13192 37568
rect 13256 37504 13264 37568
rect 12019 36684 12085 36685
rect 12019 36620 12020 36684
rect 12084 36620 12085 36684
rect 12019 36619 12085 36620
rect 12022 33693 12082 36619
rect 12944 36480 13264 37504
rect 12944 36416 12952 36480
rect 13016 36416 13032 36480
rect 13096 36416 13112 36480
rect 13176 36416 13192 36480
rect 13256 36416 13264 36480
rect 12944 35392 13264 36416
rect 12944 35328 12952 35392
rect 13016 35328 13032 35392
rect 13096 35328 13112 35392
rect 13176 35328 13192 35392
rect 13256 35328 13264 35392
rect 12944 34304 13264 35328
rect 13678 35325 13738 41243
rect 13675 35324 13741 35325
rect 13675 35260 13676 35324
rect 13740 35260 13741 35324
rect 13675 35259 13741 35260
rect 12944 34240 12952 34304
rect 13016 34240 13032 34304
rect 13096 34240 13112 34304
rect 13176 34240 13192 34304
rect 13256 34240 13264 34304
rect 12019 33692 12085 33693
rect 12019 33628 12020 33692
rect 12084 33628 12085 33692
rect 12019 33627 12085 33628
rect 12944 33216 13264 34240
rect 13859 33556 13925 33557
rect 13859 33492 13860 33556
rect 13924 33492 13925 33556
rect 13859 33491 13925 33492
rect 12944 33152 12952 33216
rect 13016 33152 13032 33216
rect 13096 33152 13112 33216
rect 13176 33152 13192 33216
rect 13256 33152 13264 33216
rect 12944 32128 13264 33152
rect 12944 32064 12952 32128
rect 13016 32064 13032 32128
rect 13096 32064 13112 32128
rect 13176 32064 13192 32128
rect 13256 32064 13264 32128
rect 9811 31380 9877 31381
rect 9811 31316 9812 31380
rect 9876 31316 9877 31380
rect 9811 31315 9877 31316
rect 7944 30432 7952 30496
rect 8016 30432 8032 30496
rect 8096 30432 8112 30496
rect 8176 30432 8192 30496
rect 8256 30432 8264 30496
rect 7944 29408 8264 30432
rect 12944 31040 13264 32064
rect 12944 30976 12952 31040
rect 13016 30976 13032 31040
rect 13096 30976 13112 31040
rect 13176 30976 13192 31040
rect 13256 30976 13264 31040
rect 12944 29952 13264 30976
rect 13862 30701 13922 33491
rect 14414 31925 14474 52531
rect 14595 40764 14661 40765
rect 14595 40700 14596 40764
rect 14660 40700 14661 40764
rect 14595 40699 14661 40700
rect 14411 31924 14477 31925
rect 14411 31860 14412 31924
rect 14476 31860 14477 31924
rect 14411 31859 14477 31860
rect 13859 30700 13925 30701
rect 13859 30636 13860 30700
rect 13924 30636 13925 30700
rect 13859 30635 13925 30636
rect 12944 29888 12952 29952
rect 13016 29888 13032 29952
rect 13096 29888 13112 29952
rect 13176 29888 13192 29952
rect 13256 29888 13264 29952
rect 12755 29476 12821 29477
rect 12755 29412 12756 29476
rect 12820 29412 12821 29476
rect 12755 29411 12821 29412
rect 7944 29344 7952 29408
rect 8016 29344 8032 29408
rect 8096 29344 8112 29408
rect 8176 29344 8192 29408
rect 8256 29344 8264 29408
rect 7944 28320 8264 29344
rect 7944 28256 7952 28320
rect 8016 28256 8032 28320
rect 8096 28256 8112 28320
rect 8176 28256 8192 28320
rect 8256 28256 8264 28320
rect 7944 27232 8264 28256
rect 7944 27168 7952 27232
rect 8016 27168 8032 27232
rect 8096 27168 8112 27232
rect 8176 27168 8192 27232
rect 8256 27168 8264 27232
rect 7944 26144 8264 27168
rect 7944 26080 7952 26144
rect 8016 26080 8032 26144
rect 8096 26080 8112 26144
rect 8176 26080 8192 26144
rect 8256 26080 8264 26144
rect 7944 25056 8264 26080
rect 7944 24992 7952 25056
rect 8016 24992 8032 25056
rect 8096 24992 8112 25056
rect 8176 24992 8192 25056
rect 8256 24992 8264 25056
rect 7944 23968 8264 24992
rect 12571 24172 12637 24173
rect 12571 24108 12572 24172
rect 12636 24108 12637 24172
rect 12571 24107 12637 24108
rect 7944 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8264 23968
rect 7944 22880 8264 23904
rect 7944 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8264 22880
rect 7944 21792 8264 22816
rect 10179 22676 10245 22677
rect 10179 22612 10180 22676
rect 10244 22612 10245 22676
rect 10179 22611 10245 22612
rect 7944 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8264 21792
rect 7944 20704 8264 21728
rect 7944 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8264 20704
rect 7944 19616 8264 20640
rect 7944 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8264 19616
rect 7944 18528 8264 19552
rect 7944 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8264 18528
rect 7944 17440 8264 18464
rect 7944 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8264 17440
rect 7944 16352 8264 17376
rect 7944 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8264 16352
rect 7944 15264 8264 16288
rect 7944 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8264 15264
rect 7944 14176 8264 15200
rect 7944 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8264 14176
rect 7944 13088 8264 14112
rect 7944 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8264 13088
rect 7944 12000 8264 13024
rect 7944 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8264 12000
rect 7944 10912 8264 11936
rect 7944 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8264 10912
rect 7944 9824 8264 10848
rect 7944 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8264 9824
rect 7944 8736 8264 9760
rect 7944 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8264 8736
rect 7944 7648 8264 8672
rect 7944 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8264 7648
rect 7944 6560 8264 7584
rect 7944 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8264 6560
rect 7944 5472 8264 6496
rect 10182 5677 10242 22611
rect 12574 17917 12634 24107
rect 12758 22677 12818 29411
rect 12944 28864 13264 29888
rect 12944 28800 12952 28864
rect 13016 28800 13032 28864
rect 13096 28800 13112 28864
rect 13176 28800 13192 28864
rect 13256 28800 13264 28864
rect 12944 27776 13264 28800
rect 12944 27712 12952 27776
rect 13016 27712 13032 27776
rect 13096 27712 13112 27776
rect 13176 27712 13192 27776
rect 13256 27712 13264 27776
rect 12944 26688 13264 27712
rect 12944 26624 12952 26688
rect 13016 26624 13032 26688
rect 13096 26624 13112 26688
rect 13176 26624 13192 26688
rect 13256 26624 13264 26688
rect 12944 25600 13264 26624
rect 12944 25536 12952 25600
rect 13016 25536 13032 25600
rect 13096 25536 13112 25600
rect 13176 25536 13192 25600
rect 13256 25536 13264 25600
rect 12944 24512 13264 25536
rect 12944 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13264 24512
rect 12944 23424 13264 24448
rect 13491 23492 13557 23493
rect 13491 23428 13492 23492
rect 13556 23428 13557 23492
rect 13491 23427 13557 23428
rect 12944 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13264 23424
rect 12755 22676 12821 22677
rect 12755 22612 12756 22676
rect 12820 22612 12821 22676
rect 12755 22611 12821 22612
rect 12944 22336 13264 23360
rect 13494 22541 13554 23427
rect 13491 22540 13557 22541
rect 13491 22476 13492 22540
rect 13556 22476 13557 22540
rect 13491 22475 13557 22476
rect 12944 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13264 22336
rect 12944 21248 13264 22272
rect 12944 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13264 21248
rect 12944 20160 13264 21184
rect 12944 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13264 20160
rect 12944 19072 13264 20096
rect 12944 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13264 19072
rect 12944 17984 13264 19008
rect 12944 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13264 17984
rect 12571 17916 12637 17917
rect 12571 17852 12572 17916
rect 12636 17852 12637 17916
rect 12571 17851 12637 17852
rect 12944 16896 13264 17920
rect 12944 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13264 16896
rect 12944 15808 13264 16832
rect 13494 16013 13554 22475
rect 13862 21861 13922 30635
rect 14414 23493 14474 31859
rect 14598 30293 14658 40699
rect 15147 38724 15213 38725
rect 15147 38660 15148 38724
rect 15212 38660 15213 38724
rect 15147 38659 15213 38660
rect 15150 34509 15210 38659
rect 15147 34508 15213 34509
rect 15147 34444 15148 34508
rect 15212 34444 15213 34508
rect 15147 34443 15213 34444
rect 14595 30292 14661 30293
rect 14595 30228 14596 30292
rect 14660 30228 14661 30292
rect 14595 30227 14661 30228
rect 14598 29069 14658 30227
rect 14595 29068 14661 29069
rect 14595 29004 14596 29068
rect 14660 29004 14661 29068
rect 14595 29003 14661 29004
rect 15702 27165 15762 52531
rect 15886 31770 15946 53891
rect 17944 53344 18264 54368
rect 17944 53280 17952 53344
rect 18016 53280 18032 53344
rect 18096 53280 18112 53344
rect 18176 53280 18192 53344
rect 18256 53280 18264 53344
rect 17944 52256 18264 53280
rect 22944 53888 23264 54448
rect 22944 53824 22952 53888
rect 23016 53824 23032 53888
rect 23096 53824 23112 53888
rect 23176 53824 23192 53888
rect 23256 53824 23264 53888
rect 22944 52800 23264 53824
rect 22944 52736 22952 52800
rect 23016 52736 23032 52800
rect 23096 52736 23112 52800
rect 23176 52736 23192 52800
rect 23256 52736 23264 52800
rect 22323 52596 22389 52597
rect 22323 52532 22324 52596
rect 22388 52532 22389 52596
rect 22323 52531 22389 52532
rect 17944 52192 17952 52256
rect 18016 52192 18032 52256
rect 18096 52192 18112 52256
rect 18176 52192 18192 52256
rect 18256 52192 18264 52256
rect 17944 51168 18264 52192
rect 17944 51104 17952 51168
rect 18016 51104 18032 51168
rect 18096 51104 18112 51168
rect 18176 51104 18192 51168
rect 18256 51104 18264 51168
rect 17944 50080 18264 51104
rect 17944 50016 17952 50080
rect 18016 50016 18032 50080
rect 18096 50016 18112 50080
rect 18176 50016 18192 50080
rect 18256 50016 18264 50080
rect 17944 48992 18264 50016
rect 17944 48928 17952 48992
rect 18016 48928 18032 48992
rect 18096 48928 18112 48992
rect 18176 48928 18192 48992
rect 18256 48928 18264 48992
rect 17944 47904 18264 48928
rect 17944 47840 17952 47904
rect 18016 47840 18032 47904
rect 18096 47840 18112 47904
rect 18176 47840 18192 47904
rect 18256 47840 18264 47904
rect 17944 46816 18264 47840
rect 17944 46752 17952 46816
rect 18016 46752 18032 46816
rect 18096 46752 18112 46816
rect 18176 46752 18192 46816
rect 18256 46752 18264 46816
rect 17944 45728 18264 46752
rect 20483 45796 20549 45797
rect 20483 45732 20484 45796
rect 20548 45732 20549 45796
rect 20483 45731 20549 45732
rect 17944 45664 17952 45728
rect 18016 45664 18032 45728
rect 18096 45664 18112 45728
rect 18176 45664 18192 45728
rect 18256 45664 18264 45728
rect 17944 44640 18264 45664
rect 17944 44576 17952 44640
rect 18016 44576 18032 44640
rect 18096 44576 18112 44640
rect 18176 44576 18192 44640
rect 18256 44576 18264 44640
rect 17944 43552 18264 44576
rect 19379 44300 19445 44301
rect 19379 44236 19380 44300
rect 19444 44236 19445 44300
rect 19379 44235 19445 44236
rect 17944 43488 17952 43552
rect 18016 43488 18032 43552
rect 18096 43488 18112 43552
rect 18176 43488 18192 43552
rect 18256 43488 18264 43552
rect 17944 42464 18264 43488
rect 17944 42400 17952 42464
rect 18016 42400 18032 42464
rect 18096 42400 18112 42464
rect 18176 42400 18192 42464
rect 18256 42400 18264 42464
rect 17944 41376 18264 42400
rect 17944 41312 17952 41376
rect 18016 41312 18032 41376
rect 18096 41312 18112 41376
rect 18176 41312 18192 41376
rect 18256 41312 18264 41376
rect 17944 40288 18264 41312
rect 17944 40224 17952 40288
rect 18016 40224 18032 40288
rect 18096 40224 18112 40288
rect 18176 40224 18192 40288
rect 18256 40224 18264 40288
rect 17944 39200 18264 40224
rect 17944 39136 17952 39200
rect 18016 39136 18032 39200
rect 18096 39136 18112 39200
rect 18176 39136 18192 39200
rect 18256 39136 18264 39200
rect 17539 38996 17605 38997
rect 17539 38932 17540 38996
rect 17604 38932 17605 38996
rect 17539 38931 17605 38932
rect 17542 33421 17602 38931
rect 17944 38112 18264 39136
rect 18459 38724 18525 38725
rect 18459 38660 18460 38724
rect 18524 38660 18525 38724
rect 18459 38659 18525 38660
rect 17944 38048 17952 38112
rect 18016 38048 18032 38112
rect 18096 38048 18112 38112
rect 18176 38048 18192 38112
rect 18256 38048 18264 38112
rect 17723 37364 17789 37365
rect 17723 37300 17724 37364
rect 17788 37300 17789 37364
rect 17723 37299 17789 37300
rect 17539 33420 17605 33421
rect 17539 33356 17540 33420
rect 17604 33356 17605 33420
rect 17539 33355 17605 33356
rect 15886 31710 16314 31770
rect 16254 30021 16314 31710
rect 17726 30429 17786 37299
rect 17944 37024 18264 38048
rect 17944 36960 17952 37024
rect 18016 36960 18032 37024
rect 18096 36960 18112 37024
rect 18176 36960 18192 37024
rect 18256 36960 18264 37024
rect 17944 35936 18264 36960
rect 17944 35872 17952 35936
rect 18016 35872 18032 35936
rect 18096 35872 18112 35936
rect 18176 35872 18192 35936
rect 18256 35872 18264 35936
rect 17944 34848 18264 35872
rect 17944 34784 17952 34848
rect 18016 34784 18032 34848
rect 18096 34784 18112 34848
rect 18176 34784 18192 34848
rect 18256 34784 18264 34848
rect 17944 33760 18264 34784
rect 17944 33696 17952 33760
rect 18016 33696 18032 33760
rect 18096 33696 18112 33760
rect 18176 33696 18192 33760
rect 18256 33696 18264 33760
rect 17944 32672 18264 33696
rect 17944 32608 17952 32672
rect 18016 32608 18032 32672
rect 18096 32608 18112 32672
rect 18176 32608 18192 32672
rect 18256 32608 18264 32672
rect 17944 31584 18264 32608
rect 17944 31520 17952 31584
rect 18016 31520 18032 31584
rect 18096 31520 18112 31584
rect 18176 31520 18192 31584
rect 18256 31520 18264 31584
rect 17944 30496 18264 31520
rect 18462 30837 18522 38659
rect 18643 37636 18709 37637
rect 18643 37572 18644 37636
rect 18708 37572 18709 37636
rect 18643 37571 18709 37572
rect 18459 30836 18525 30837
rect 18459 30772 18460 30836
rect 18524 30772 18525 30836
rect 18459 30771 18525 30772
rect 17944 30432 17952 30496
rect 18016 30432 18032 30496
rect 18096 30432 18112 30496
rect 18176 30432 18192 30496
rect 18256 30432 18264 30496
rect 17723 30428 17789 30429
rect 17723 30364 17724 30428
rect 17788 30364 17789 30428
rect 17723 30363 17789 30364
rect 16251 30020 16317 30021
rect 16251 29956 16252 30020
rect 16316 29956 16317 30020
rect 16251 29955 16317 29956
rect 16254 28117 16314 29955
rect 17723 29748 17789 29749
rect 17723 29684 17724 29748
rect 17788 29684 17789 29748
rect 17723 29683 17789 29684
rect 16803 29068 16869 29069
rect 16803 29004 16804 29068
rect 16868 29004 16869 29068
rect 16803 29003 16869 29004
rect 17539 29068 17605 29069
rect 17539 29004 17540 29068
rect 17604 29004 17605 29068
rect 17539 29003 17605 29004
rect 16251 28116 16317 28117
rect 16251 28052 16252 28116
rect 16316 28052 16317 28116
rect 16251 28051 16317 28052
rect 15699 27164 15765 27165
rect 15699 27100 15700 27164
rect 15764 27100 15765 27164
rect 15699 27099 15765 27100
rect 16067 25668 16133 25669
rect 16067 25604 16068 25668
rect 16132 25604 16133 25668
rect 16067 25603 16133 25604
rect 14411 23492 14477 23493
rect 14411 23428 14412 23492
rect 14476 23428 14477 23492
rect 14411 23427 14477 23428
rect 13859 21860 13925 21861
rect 13859 21796 13860 21860
rect 13924 21796 13925 21860
rect 13859 21795 13925 21796
rect 13491 16012 13557 16013
rect 13491 15948 13492 16012
rect 13556 15948 13557 16012
rect 13491 15947 13557 15948
rect 12944 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13264 15808
rect 12944 14720 13264 15744
rect 13862 15333 13922 21795
rect 16070 20637 16130 25603
rect 16067 20636 16133 20637
rect 16067 20572 16068 20636
rect 16132 20572 16133 20636
rect 16067 20571 16133 20572
rect 14963 20228 15029 20229
rect 14963 20164 14964 20228
rect 15028 20164 15029 20228
rect 14963 20163 15029 20164
rect 13859 15332 13925 15333
rect 13859 15268 13860 15332
rect 13924 15268 13925 15332
rect 13859 15267 13925 15268
rect 12944 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13264 14720
rect 12944 13632 13264 14656
rect 12944 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13264 13632
rect 12944 12544 13264 13568
rect 12944 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13264 12544
rect 12944 11456 13264 12480
rect 12944 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13264 11456
rect 12944 10368 13264 11392
rect 12944 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13264 10368
rect 12944 9280 13264 10304
rect 12944 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13264 9280
rect 12944 8192 13264 9216
rect 12944 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13264 8192
rect 12944 7104 13264 8128
rect 12944 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13264 7104
rect 12944 6016 13264 7040
rect 12944 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13264 6016
rect 10179 5676 10245 5677
rect 10179 5612 10180 5676
rect 10244 5612 10245 5676
rect 10179 5611 10245 5612
rect 7944 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8264 5472
rect 7944 4384 8264 5408
rect 7944 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8264 4384
rect 7944 3296 8264 4320
rect 7944 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8264 3296
rect 7944 2208 8264 3232
rect 7944 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8264 2208
rect 7944 2128 8264 2144
rect 12944 4928 13264 5952
rect 14966 5813 15026 20163
rect 16254 17645 16314 28051
rect 16251 17644 16317 17645
rect 16251 17580 16252 17644
rect 16316 17580 16317 17644
rect 16251 17579 16317 17580
rect 15699 15332 15765 15333
rect 15699 15268 15700 15332
rect 15764 15268 15765 15332
rect 15699 15267 15765 15268
rect 14963 5812 15029 5813
rect 14963 5748 14964 5812
rect 15028 5748 15029 5812
rect 14963 5747 15029 5748
rect 12944 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13264 4928
rect 12944 3840 13264 4864
rect 12944 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13264 3840
rect 12944 2752 13264 3776
rect 12944 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13264 2752
rect 12944 2128 13264 2688
rect 15702 2685 15762 15267
rect 16806 3501 16866 29003
rect 17542 18869 17602 29003
rect 17726 23357 17786 29683
rect 17944 29408 18264 30432
rect 17944 29344 17952 29408
rect 18016 29344 18032 29408
rect 18096 29344 18112 29408
rect 18176 29344 18192 29408
rect 18256 29344 18264 29408
rect 17944 28320 18264 29344
rect 17944 28256 17952 28320
rect 18016 28256 18032 28320
rect 18096 28256 18112 28320
rect 18176 28256 18192 28320
rect 18256 28256 18264 28320
rect 17944 27232 18264 28256
rect 18459 27572 18525 27573
rect 18459 27508 18460 27572
rect 18524 27508 18525 27572
rect 18459 27507 18525 27508
rect 17944 27168 17952 27232
rect 18016 27168 18032 27232
rect 18096 27168 18112 27232
rect 18176 27168 18192 27232
rect 18256 27168 18264 27232
rect 17944 26144 18264 27168
rect 17944 26080 17952 26144
rect 18016 26080 18032 26144
rect 18096 26080 18112 26144
rect 18176 26080 18192 26144
rect 18256 26080 18264 26144
rect 17944 25056 18264 26080
rect 17944 24992 17952 25056
rect 18016 24992 18032 25056
rect 18096 24992 18112 25056
rect 18176 24992 18192 25056
rect 18256 24992 18264 25056
rect 17944 23968 18264 24992
rect 17944 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18264 23968
rect 17723 23356 17789 23357
rect 17723 23292 17724 23356
rect 17788 23292 17789 23356
rect 17723 23291 17789 23292
rect 17726 22269 17786 23291
rect 17944 22880 18264 23904
rect 17944 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18264 22880
rect 17723 22268 17789 22269
rect 17723 22204 17724 22268
rect 17788 22204 17789 22268
rect 17723 22203 17789 22204
rect 17944 21792 18264 22816
rect 17944 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18264 21792
rect 17944 20704 18264 21728
rect 17944 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18264 20704
rect 17944 19616 18264 20640
rect 17944 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18264 19616
rect 17539 18868 17605 18869
rect 17539 18804 17540 18868
rect 17604 18804 17605 18868
rect 17539 18803 17605 18804
rect 17944 18528 18264 19552
rect 17944 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18264 18528
rect 17944 17440 18264 18464
rect 18462 18325 18522 27507
rect 18646 19957 18706 37571
rect 19382 29749 19442 44235
rect 19747 37228 19813 37229
rect 19747 37164 19748 37228
rect 19812 37164 19813 37228
rect 19747 37163 19813 37164
rect 19563 30156 19629 30157
rect 19563 30092 19564 30156
rect 19628 30092 19629 30156
rect 19563 30091 19629 30092
rect 19379 29748 19445 29749
rect 19379 29684 19380 29748
rect 19444 29684 19445 29748
rect 19379 29683 19445 29684
rect 18643 19956 18709 19957
rect 18643 19892 18644 19956
rect 18708 19892 18709 19956
rect 18643 19891 18709 19892
rect 18459 18324 18525 18325
rect 18459 18260 18460 18324
rect 18524 18260 18525 18324
rect 18459 18259 18525 18260
rect 19566 17645 19626 30091
rect 19750 29749 19810 37163
rect 20486 30701 20546 45731
rect 21403 45524 21469 45525
rect 21403 45460 21404 45524
rect 21468 45460 21469 45524
rect 21403 45459 21469 45460
rect 21035 44300 21101 44301
rect 21035 44236 21036 44300
rect 21100 44236 21101 44300
rect 21035 44235 21101 44236
rect 21038 31770 21098 44235
rect 21219 41444 21285 41445
rect 21219 41380 21220 41444
rect 21284 41380 21285 41444
rect 21219 41379 21285 41380
rect 20854 31710 21098 31770
rect 20483 30700 20549 30701
rect 20483 30636 20484 30700
rect 20548 30636 20549 30700
rect 20483 30635 20549 30636
rect 19747 29748 19813 29749
rect 19747 29684 19748 29748
rect 19812 29684 19813 29748
rect 19747 29683 19813 29684
rect 20854 28389 20914 31710
rect 20851 28388 20917 28389
rect 20851 28324 20852 28388
rect 20916 28324 20917 28388
rect 20851 28323 20917 28324
rect 20854 24581 20914 28323
rect 21222 27573 21282 41379
rect 21219 27572 21285 27573
rect 21219 27508 21220 27572
rect 21284 27508 21285 27572
rect 21219 27507 21285 27508
rect 21406 27165 21466 45459
rect 22326 31789 22386 52531
rect 22944 51712 23264 52736
rect 22944 51648 22952 51712
rect 23016 51648 23032 51712
rect 23096 51648 23112 51712
rect 23176 51648 23192 51712
rect 23256 51648 23264 51712
rect 22944 50624 23264 51648
rect 22944 50560 22952 50624
rect 23016 50560 23032 50624
rect 23096 50560 23112 50624
rect 23176 50560 23192 50624
rect 23256 50560 23264 50624
rect 22944 49536 23264 50560
rect 22944 49472 22952 49536
rect 23016 49472 23032 49536
rect 23096 49472 23112 49536
rect 23176 49472 23192 49536
rect 23256 49472 23264 49536
rect 22944 48448 23264 49472
rect 22944 48384 22952 48448
rect 23016 48384 23032 48448
rect 23096 48384 23112 48448
rect 23176 48384 23192 48448
rect 23256 48384 23264 48448
rect 22944 47360 23264 48384
rect 22944 47296 22952 47360
rect 23016 47296 23032 47360
rect 23096 47296 23112 47360
rect 23176 47296 23192 47360
rect 23256 47296 23264 47360
rect 22944 46272 23264 47296
rect 22944 46208 22952 46272
rect 23016 46208 23032 46272
rect 23096 46208 23112 46272
rect 23176 46208 23192 46272
rect 23256 46208 23264 46272
rect 22944 45184 23264 46208
rect 22944 45120 22952 45184
rect 23016 45120 23032 45184
rect 23096 45120 23112 45184
rect 23176 45120 23192 45184
rect 23256 45120 23264 45184
rect 22944 44096 23264 45120
rect 22944 44032 22952 44096
rect 23016 44032 23032 44096
rect 23096 44032 23112 44096
rect 23176 44032 23192 44096
rect 23256 44032 23264 44096
rect 22944 43008 23264 44032
rect 22944 42944 22952 43008
rect 23016 42944 23032 43008
rect 23096 42944 23112 43008
rect 23176 42944 23192 43008
rect 23256 42944 23264 43008
rect 22944 41920 23264 42944
rect 22944 41856 22952 41920
rect 23016 41856 23032 41920
rect 23096 41856 23112 41920
rect 23176 41856 23192 41920
rect 23256 41856 23264 41920
rect 22944 40832 23264 41856
rect 22944 40768 22952 40832
rect 23016 40768 23032 40832
rect 23096 40768 23112 40832
rect 23176 40768 23192 40832
rect 23256 40768 23264 40832
rect 22944 39744 23264 40768
rect 22944 39680 22952 39744
rect 23016 39680 23032 39744
rect 23096 39680 23112 39744
rect 23176 39680 23192 39744
rect 23256 39680 23264 39744
rect 22944 38656 23264 39680
rect 22944 38592 22952 38656
rect 23016 38592 23032 38656
rect 23096 38592 23112 38656
rect 23176 38592 23192 38656
rect 23256 38592 23264 38656
rect 22944 37568 23264 38592
rect 22944 37504 22952 37568
rect 23016 37504 23032 37568
rect 23096 37504 23112 37568
rect 23176 37504 23192 37568
rect 23256 37504 23264 37568
rect 22944 36480 23264 37504
rect 22944 36416 22952 36480
rect 23016 36416 23032 36480
rect 23096 36416 23112 36480
rect 23176 36416 23192 36480
rect 23256 36416 23264 36480
rect 22944 35392 23264 36416
rect 22944 35328 22952 35392
rect 23016 35328 23032 35392
rect 23096 35328 23112 35392
rect 23176 35328 23192 35392
rect 23256 35328 23264 35392
rect 22507 35188 22573 35189
rect 22507 35124 22508 35188
rect 22572 35124 22573 35188
rect 22507 35123 22573 35124
rect 22323 31788 22389 31789
rect 22323 31724 22324 31788
rect 22388 31724 22389 31788
rect 22323 31723 22389 31724
rect 22510 29749 22570 35123
rect 22944 34304 23264 35328
rect 22944 34240 22952 34304
rect 23016 34240 23032 34304
rect 23096 34240 23112 34304
rect 23176 34240 23192 34304
rect 23256 34240 23264 34304
rect 22944 33216 23264 34240
rect 22944 33152 22952 33216
rect 23016 33152 23032 33216
rect 23096 33152 23112 33216
rect 23176 33152 23192 33216
rect 23256 33152 23264 33216
rect 22944 32128 23264 33152
rect 22944 32064 22952 32128
rect 23016 32064 23032 32128
rect 23096 32064 23112 32128
rect 23176 32064 23192 32128
rect 23256 32064 23264 32128
rect 22944 31040 23264 32064
rect 22944 30976 22952 31040
rect 23016 30976 23032 31040
rect 23096 30976 23112 31040
rect 23176 30976 23192 31040
rect 23256 30976 23264 31040
rect 22944 29952 23264 30976
rect 22944 29888 22952 29952
rect 23016 29888 23032 29952
rect 23096 29888 23112 29952
rect 23176 29888 23192 29952
rect 23256 29888 23264 29952
rect 22507 29748 22573 29749
rect 22507 29684 22508 29748
rect 22572 29684 22573 29748
rect 22507 29683 22573 29684
rect 22944 28864 23264 29888
rect 23427 29476 23493 29477
rect 23427 29412 23428 29476
rect 23492 29412 23493 29476
rect 23427 29411 23493 29412
rect 22944 28800 22952 28864
rect 23016 28800 23032 28864
rect 23096 28800 23112 28864
rect 23176 28800 23192 28864
rect 23256 28800 23264 28864
rect 22944 27776 23264 28800
rect 22944 27712 22952 27776
rect 23016 27712 23032 27776
rect 23096 27712 23112 27776
rect 23176 27712 23192 27776
rect 23256 27712 23264 27776
rect 21403 27164 21469 27165
rect 21403 27100 21404 27164
rect 21468 27100 21469 27164
rect 21403 27099 21469 27100
rect 22944 26688 23264 27712
rect 22944 26624 22952 26688
rect 23016 26624 23032 26688
rect 23096 26624 23112 26688
rect 23176 26624 23192 26688
rect 23256 26624 23264 26688
rect 22944 25600 23264 26624
rect 23430 26213 23490 29411
rect 23427 26212 23493 26213
rect 23427 26148 23428 26212
rect 23492 26148 23493 26212
rect 23427 26147 23493 26148
rect 22944 25536 22952 25600
rect 23016 25536 23032 25600
rect 23096 25536 23112 25600
rect 23176 25536 23192 25600
rect 23256 25536 23264 25600
rect 20851 24580 20917 24581
rect 20851 24516 20852 24580
rect 20916 24516 20917 24580
rect 20851 24515 20917 24516
rect 22944 24512 23264 25536
rect 22944 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23264 24512
rect 22944 23424 23264 24448
rect 22944 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23264 23424
rect 22944 22336 23264 23360
rect 22944 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23264 22336
rect 22944 21248 23264 22272
rect 22944 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23264 21248
rect 22944 20160 23264 21184
rect 22944 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23264 20160
rect 22944 19072 23264 20096
rect 22944 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23264 19072
rect 22944 17984 23264 19008
rect 22944 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23264 17984
rect 19563 17644 19629 17645
rect 19563 17580 19564 17644
rect 19628 17580 19629 17644
rect 19563 17579 19629 17580
rect 17944 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18264 17440
rect 17944 16352 18264 17376
rect 17944 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18264 16352
rect 17944 15264 18264 16288
rect 17944 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18264 15264
rect 17944 14176 18264 15200
rect 17944 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18264 14176
rect 17944 13088 18264 14112
rect 19566 13565 19626 17579
rect 22944 16896 23264 17920
rect 22944 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23264 16896
rect 22944 15808 23264 16832
rect 22944 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23264 15808
rect 22944 14720 23264 15744
rect 22944 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23264 14720
rect 22944 13632 23264 14656
rect 22944 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23264 13632
rect 19563 13564 19629 13565
rect 19563 13500 19564 13564
rect 19628 13500 19629 13564
rect 19563 13499 19629 13500
rect 17944 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18264 13088
rect 17944 12000 18264 13024
rect 17944 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18264 12000
rect 17944 10912 18264 11936
rect 17944 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18264 10912
rect 17944 9824 18264 10848
rect 17944 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18264 9824
rect 17944 8736 18264 9760
rect 17944 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18264 8736
rect 17944 7648 18264 8672
rect 17944 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18264 7648
rect 17944 6560 18264 7584
rect 17944 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18264 6560
rect 17944 5472 18264 6496
rect 17944 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18264 5472
rect 17944 4384 18264 5408
rect 17944 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18264 4384
rect 16803 3500 16869 3501
rect 16803 3436 16804 3500
rect 16868 3436 16869 3500
rect 16803 3435 16869 3436
rect 17944 3296 18264 4320
rect 17944 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18264 3296
rect 15699 2684 15765 2685
rect 15699 2620 15700 2684
rect 15764 2620 15765 2684
rect 15699 2619 15765 2620
rect 17944 2208 18264 3232
rect 17944 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18264 2208
rect 17944 2128 18264 2144
rect 22944 12544 23264 13568
rect 22944 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23264 12544
rect 22944 11456 23264 12480
rect 22944 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23264 11456
rect 22944 10368 23264 11392
rect 22944 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23264 10368
rect 22944 9280 23264 10304
rect 22944 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23264 9280
rect 22944 8192 23264 9216
rect 22944 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23264 8192
rect 22944 7104 23264 8128
rect 22944 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23264 7104
rect 22944 6016 23264 7040
rect 22944 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23264 6016
rect 22944 4928 23264 5952
rect 22944 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23264 4928
rect 22944 3840 23264 4864
rect 22944 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23264 3840
rect 22944 2752 23264 3776
rect 22944 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23264 2752
rect 22944 2128 23264 2688
use sky130_fd_sc_hd__clkbuf_1  _109_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24656 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _110_
timestamp 1676037725
transform 1 0 24564 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _111_
timestamp 1676037725
transform -1 0 23368 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _112_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 24932 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _113_
timestamp 1676037725
transform 1 0 24564 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _114_
timestamp 1676037725
transform -1 0 24104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _115_
timestamp 1676037725
transform 1 0 24564 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _116_
timestamp 1676037725
transform 1 0 15916 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _117_
timestamp 1676037725
transform -1 0 23460 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _118_
timestamp 1676037725
transform -1 0 22724 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _119_
timestamp 1676037725
transform -1 0 21068 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _120_
timestamp 1676037725
transform 1 0 20424 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _121_
timestamp 1676037725
transform 1 0 21160 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _122_
timestamp 1676037725
transform 1 0 21620 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _123_
timestamp 1676037725
transform 1 0 21160 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _124_
timestamp 1676037725
transform 1 0 21896 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _125_
timestamp 1676037725
transform -1 0 24932 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _126_
timestamp 1676037725
transform 1 0 22816 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _127_
timestamp 1676037725
transform 1 0 22172 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _128_
timestamp 1676037725
transform -1 0 24932 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _129_
timestamp 1676037725
transform -1 0 23736 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _130_
timestamp 1676037725
transform -1 0 24472 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _131_
timestamp 1676037725
transform -1 0 25208 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _132_
timestamp 1676037725
transform 1 0 24564 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _133_
timestamp 1676037725
transform -1 0 24932 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _134_
timestamp 1676037725
transform -1 0 24932 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _135_
timestamp 1676037725
transform -1 0 24932 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _136_
timestamp 1676037725
transform -1 0 24932 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _137_
timestamp 1676037725
transform 1 0 24564 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _138_
timestamp 1676037725
transform -1 0 12696 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _139_
timestamp 1676037725
transform -1 0 14628 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _140_
timestamp 1676037725
transform 1 0 12696 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _141_
timestamp 1676037725
transform 1 0 11500 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _142_
timestamp 1676037725
transform 1 0 13432 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _143_
timestamp 1676037725
transform 1 0 13432 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _144_
timestamp 1676037725
transform -1 0 16376 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _145_
timestamp 1676037725
transform -1 0 17204 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _146_
timestamp 1676037725
transform 1 0 15456 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _147_
timestamp 1676037725
transform 1 0 14812 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _148_
timestamp 1676037725
transform 1 0 15180 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _149_
timestamp 1676037725
transform 1 0 14260 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _150_
timestamp 1676037725
transform 1 0 17112 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _151_
timestamp 1676037725
transform 1 0 17204 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _152_
timestamp 1676037725
transform 1 0 16008 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _153_
timestamp 1676037725
transform 1 0 16008 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _154_
timestamp 1676037725
transform 1 0 17388 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _155_
timestamp 1676037725
transform 1 0 17940 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _156_
timestamp 1676037725
transform 1 0 18216 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _157_
timestamp 1676037725
transform 1 0 20240 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _158_
timestamp 1676037725
transform 1 0 19412 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _159_
timestamp 1676037725
transform 1 0 19596 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _160_
timestamp 1676037725
transform 1 0 19780 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _161_
timestamp 1676037725
transform 1 0 18400 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _162_
timestamp 1676037725
transform 1 0 18124 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _163_
timestamp 1676037725
transform 1 0 20240 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _164_
timestamp 1676037725
transform 1 0 18584 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _165_
timestamp 1676037725
transform -1 0 20240 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _166_
timestamp 1676037725
transform 1 0 19320 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _167_
timestamp 1676037725
transform -1 0 19688 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _168_
timestamp 1676037725
transform 1 0 2668 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _169_
timestamp 1676037725
transform -1 0 4048 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _170_
timestamp 1676037725
transform -1 0 4232 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _171_
timestamp 1676037725
transform -1 0 7084 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _172_
timestamp 1676037725
transform -1 0 4508 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _173_
timestamp 1676037725
transform -1 0 4692 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _174_
timestamp 1676037725
transform -1 0 5612 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _175_
timestamp 1676037725
transform 1 0 6624 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _176_
timestamp 1676037725
transform -1 0 6624 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _177_
timestamp 1676037725
transform -1 0 6716 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _178_
timestamp 1676037725
transform -1 0 7452 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _179_
timestamp 1676037725
transform 1 0 5888 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _180_
timestamp 1676037725
transform -1 0 7728 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _181_
timestamp 1676037725
transform -1 0 7912 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _182_
timestamp 1676037725
transform -1 0 8648 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _183_
timestamp 1676037725
transform -1 0 6808 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _184_
timestamp 1676037725
transform -1 0 8832 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _185_
timestamp 1676037725
transform -1 0 8648 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _186_
timestamp 1676037725
transform -1 0 10028 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _187_
timestamp 1676037725
transform 1 0 7820 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _188_
timestamp 1676037725
transform -1 0 10764 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _189_
timestamp 1676037725
transform 1 0 9936 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _190_
timestamp 1676037725
transform -1 0 12052 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _191_
timestamp 1676037725
transform 1 0 9292 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _192_
timestamp 1676037725
transform 1 0 9108 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _193_
timestamp 1676037725
transform -1 0 13248 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _194_
timestamp 1676037725
transform 1 0 9660 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _195_
timestamp 1676037725
transform -1 0 10764 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _196_
timestamp 1676037725
transform -1 0 11960 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _197_
timestamp 1676037725
transform -1 0 12052 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _198_
timestamp 1676037725
transform -1 0 2760 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _199_
timestamp 1676037725
transform 1 0 2024 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _200_
timestamp 1676037725
transform 1 0 2024 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _201_
timestamp 1676037725
transform 1 0 2024 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _202_
timestamp 1676037725
transform 1 0 2668 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _203_
timestamp 1676037725
transform 1 0 1932 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _204_
timestamp 1676037725
transform 1 0 2024 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _205_
timestamp 1676037725
transform 1 0 2024 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _206_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23184 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _207_
timestamp 1676037725
transform 1 0 2024 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _208_
timestamp 1676037725
transform 1 0 24564 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _209_
timestamp 1676037725
transform 1 0 24564 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _210_
timestamp 1676037725
transform -1 0 24012 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _211_
timestamp 1676037725
transform 1 0 24656 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _212_
timestamp 1676037725
transform 1 0 24564 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _213_
timestamp 1676037725
transform 1 0 23828 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _214_
timestamp 1676037725
transform 1 0 24564 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _215_
timestamp 1676037725
transform -1 0 24104 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _216_
timestamp 1676037725
transform -1 0 24196 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _217_
timestamp 1676037725
transform -1 0 23552 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _218_
timestamp 1676037725
transform -1 0 24932 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__138__A pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12696 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__139__A
timestamp 1676037725
transform 1 0 14812 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__140__A
timestamp 1676037725
transform 1 0 13064 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__142__A
timestamp 1676037725
transform -1 0 13984 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__143__A
timestamp 1676037725
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__144__A
timestamp 1676037725
transform 1 0 16192 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__146__A
timestamp 1676037725
transform 1 0 16652 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__147__A
timestamp 1676037725
transform 1 0 15364 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__148__A
timestamp 1676037725
transform -1 0 16100 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__150__A
timestamp 1676037725
transform -1 0 16928 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__151__A
timestamp 1676037725
transform -1 0 17020 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__152__A
timestamp 1676037725
transform -1 0 16836 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__154__A
timestamp 1676037725
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__155__A
timestamp 1676037725
transform 1 0 18676 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__156__A
timestamp 1676037725
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__158__A
timestamp 1676037725
transform 1 0 19964 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__159__A
timestamp 1676037725
transform 1 0 20148 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__160__A
timestamp 1676037725
transform -1 0 20516 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__163__A
timestamp 1676037725
transform -1 0 20976 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__168__A
timestamp 1676037725
transform -1 0 3404 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__169__A
timestamp 1676037725
transform 1 0 4232 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__170__A
timestamp 1676037725
transform 1 0 4416 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__172__A
timestamp 1676037725
transform -1 0 4876 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__173__A
timestamp 1676037725
transform -1 0 5060 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__174__A
timestamp 1676037725
transform -1 0 5980 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__176__A
timestamp 1676037725
transform -1 0 6072 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__177__A
timestamp 1676037725
transform -1 0 7084 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__178__A
timestamp 1676037725
transform 1 0 6716 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__180__A
timestamp 1676037725
transform -1 0 8096 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__181__A
timestamp 1676037725
transform 1 0 7176 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__182__A
timestamp 1676037725
transform -1 0 9108 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__184__A
timestamp 1676037725
transform -1 0 8464 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__185__A
timestamp 1676037725
transform -1 0 8280 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__186__A
timestamp 1676037725
transform -1 0 9476 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__188__A
timestamp 1676037725
transform -1 0 11132 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__189__A
timestamp 1676037725
transform -1 0 9752 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__190__A
timestamp 1676037725
transform 1 0 12236 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__193__A
timestamp 1676037725
transform 1 0 13432 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__206__A
timestamp 1676037725
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__207__A
timestamp 1676037725
transform 1 0 2484 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__208__A
timestamp 1676037725
transform 1 0 25024 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__209__A
timestamp 1676037725
transform 1 0 25208 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__210__A
timestamp 1676037725
transform 1 0 25024 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__211__A
timestamp 1676037725
transform -1 0 25484 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__212__A
timestamp 1676037725
transform 1 0 25024 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__213__A
timestamp 1676037725
transform -1 0 23644 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__214__A
timestamp 1676037725
transform -1 0 25300 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__215__A
timestamp 1676037725
transform 1 0 25116 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__216__A
timestamp 1676037725
transform -1 0 24564 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__217__A
timestamp 1676037725
transform -1 0 23736 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__218__A
timestamp 1676037725
transform 1 0 25116 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 11500 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 6808 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1676037725
transform 1 0 6992 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 9476 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 14076 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 10856 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1676037725
transform 1 0 8464 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 11132 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 12328 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 8188 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1676037725
transform 1 0 6808 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 7912 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 10488 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 7544 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1676037725
transform 1 0 6348 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 12880 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 13524 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_3__A0
timestamp 1676037725
transform 1 0 13616 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 12420 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_4__A1
timestamp 1676037725
transform 1 0 10304 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_2__A0
timestamp 1676037725
transform 1 0 6992 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_3__A1
timestamp 1676037725
transform 1 0 10672 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 15272 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_3__A0
timestamp 1676037725
transform 1 0 15272 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_4__A0
timestamp 1676037725
transform 1 0 12788 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_4__A1
timestamp 1676037725
transform 1 0 11684 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_3__A1
timestamp 1676037725
transform 1 0 12328 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 15272 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 14904 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 15088 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 12328 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_4__A0
timestamp 1676037725
transform 1 0 10948 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_4__A1
timestamp 1676037725
transform 1 0 9568 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_2__A0
timestamp 1676037725
transform 1 0 7452 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 12052 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 14076 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 12696 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_3__A0
timestamp 1676037725
transform 1 0 13156 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 11132 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_4__A0
timestamp 1676037725
transform 1 0 11316 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_2__A0
timestamp 1676037725
transform 1 0 7268 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3__A1
timestamp 1676037725
transform 1 0 9016 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1676037725
transform 1 0 3496 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 5060 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1676037725
transform 1 0 2484 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 4416 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1676037725
transform 1 0 4232 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 5888 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1676037725
transform -1 0 10028 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 12328 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1676037725
transform 1 0 16652 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_0_0_prog_clk_A
timestamp 1676037725
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_1_0_prog_clk_A
timestamp 1676037725
transform 1 0 11500 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_2_0_prog_clk_A
timestamp 1676037725
transform 1 0 8280 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_3_0_prog_clk_A
timestamp 1676037725
transform 1 0 11500 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_4_0_prog_clk_A
timestamp 1676037725
transform 1 0 17572 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_5_0_prog_clk_A
timestamp 1676037725
transform 1 0 19964 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_6_0_prog_clk_A
timestamp 1676037725
transform 1 0 17756 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_7_0_prog_clk_A
timestamp 1676037725
transform -1 0 21988 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_8_0_prog_clk_A
timestamp 1676037725
transform 1 0 8648 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_9_0_prog_clk_A
timestamp 1676037725
transform 1 0 12420 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_10_0_prog_clk_A
timestamp 1676037725
transform 1 0 10120 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_11_0_prog_clk_A
timestamp 1676037725
transform 1 0 12512 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_12_0_prog_clk_A
timestamp 1676037725
transform 1 0 19228 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_13_0_prog_clk_A
timestamp 1676037725
transform 1 0 21068 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_14_0_prog_clk_A
timestamp 1676037725
transform 1 0 17572 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_15_0_prog_clk_A
timestamp 1676037725
transform 1 0 20148 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1676037725
transform -1 0 2208 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1676037725
transform -1 0 2300 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1676037725
transform -1 0 25576 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1676037725
transform -1 0 24932 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1676037725
transform -1 0 24932 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1676037725
transform -1 0 25392 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1676037725
transform -1 0 24932 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1676037725
transform -1 0 24932 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1676037725
transform -1 0 24748 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1676037725
transform -1 0 25392 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1676037725
transform -1 0 24564 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1676037725
transform -1 0 24932 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1676037725
transform -1 0 24932 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1676037725
transform -1 0 21068 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1676037725
transform -1 0 25576 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1676037725
transform -1 0 24288 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1676037725
transform -1 0 23644 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1676037725
transform -1 0 24564 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1676037725
transform 1 0 25392 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1676037725
transform -1 0 24932 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1676037725
transform 1 0 25392 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1676037725
transform 1 0 25392 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1676037725
transform 1 0 25024 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1676037725
transform 1 0 23736 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1676037725
transform -1 0 24564 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1676037725
transform 1 0 25300 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1676037725
transform -1 0 24748 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1676037725
transform -1 0 23736 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1676037725
transform -1 0 25576 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1676037725
transform -1 0 25576 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1676037725
transform -1 0 24932 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1676037725
transform -1 0 25576 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1676037725
transform -1 0 1564 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1676037725
transform -1 0 4692 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1676037725
transform -1 0 5520 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1676037725
transform -1 0 5612 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1676037725
transform -1 0 6532 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1676037725
transform -1 0 7084 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1676037725
transform -1 0 6532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1676037725
transform -1 0 6900 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1676037725
transform -1 0 7268 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1676037725
transform -1 0 6808 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1676037725
transform -1 0 8372 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1676037725
transform -1 0 1564 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1676037725
transform -1 0 9108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1676037725
transform 1 0 8372 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1676037725
transform -1 0 10028 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1676037725
transform -1 0 9844 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1676037725
transform -1 0 10028 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1676037725
transform -1 0 11408 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1676037725
transform -1 0 12052 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1676037725
transform -1 0 9292 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1676037725
transform -1 0 14260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1676037725
transform -1 0 12788 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1676037725
transform -1 0 1748 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1676037725
transform -1 0 1656 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1676037725
transform -1 0 4232 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1676037725
transform -1 0 3036 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1676037725
transform -1 0 3312 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1676037725
transform -1 0 4048 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1676037725
transform -1 0 3956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1676037725
transform -1 0 4508 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 1676037725
transform -1 0 12420 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 1676037725
transform -1 0 16836 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 1676037725
transform -1 0 16468 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 1676037725
transform -1 0 17204 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 1676037725
transform -1 0 19044 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input68_A
timestamp 1676037725
transform -1 0 18308 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 1676037725
transform -1 0 17940 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input70_A
timestamp 1676037725
transform -1 0 18676 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input71_A
timestamp 1676037725
transform -1 0 19412 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input72_A
timestamp 1676037725
transform -1 0 20148 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input73_A
timestamp 1676037725
transform -1 0 21620 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input74_A
timestamp 1676037725
transform -1 0 14996 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input75_A
timestamp 1676037725
transform -1 0 20424 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input76_A
timestamp 1676037725
transform -1 0 20884 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input77_A
timestamp 1676037725
transform -1 0 20332 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input78_A
timestamp 1676037725
transform -1 0 21252 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input79_A
timestamp 1676037725
transform -1 0 21988 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input80_A
timestamp 1676037725
transform -1 0 21528 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input81_A
timestamp 1676037725
transform -1 0 21712 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input82_A
timestamp 1676037725
transform -1 0 23368 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input83_A
timestamp 1676037725
transform -1 0 25208 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input84_A
timestamp 1676037725
transform -1 0 25208 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input85_A
timestamp 1676037725
transform -1 0 13892 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input86_A
timestamp 1676037725
transform -1 0 14260 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input87_A
timestamp 1676037725
transform -1 0 13984 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input88_A
timestamp 1676037725
transform -1 0 14996 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input89_A
timestamp 1676037725
transform -1 0 14444 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input90_A
timestamp 1676037725
transform -1 0 15364 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input91_A
timestamp 1676037725
transform -1 0 16100 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input92_A
timestamp 1676037725
transform -1 0 15548 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input93_A
timestamp 1676037725
transform -1 0 2208 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input94_A
timestamp 1676037725
transform -1 0 2208 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input95_A
timestamp 1676037725
transform -1 0 2208 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input96_A
timestamp 1676037725
transform -1 0 2208 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input97_A
timestamp 1676037725
transform -1 0 2300 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input98_A
timestamp 1676037725
transform -1 0 25576 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input99_A
timestamp 1676037725
transform -1 0 2208 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input100_A
timestamp 1676037725
transform -1 0 23368 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input101_A
timestamp 1676037725
transform -1 0 25300 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input102_A
timestamp 1676037725
transform -1 0 24288 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input103_A
timestamp 1676037725
transform -1 0 23552 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input104_A
timestamp 1676037725
transform 1 0 25392 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input105_A
timestamp 1676037725
transform -1 0 24840 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input106_A
timestamp 1676037725
transform -1 0 24840 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input107_A
timestamp 1676037725
transform -1 0 24840 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input108_A
timestamp 1676037725
transform -1 0 24840 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input109_A
timestamp 1676037725
transform -1 0 24840 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input110_A
timestamp 1676037725
transform -1 0 25576 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input111_A
timestamp 1676037725
transform -1 0 25576 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input112_A
timestamp 1676037725
transform -1 0 24840 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input113_A
timestamp 1676037725
transform -1 0 24840 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input114_A
timestamp 1676037725
transform 1 0 24380 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input115_A
timestamp 1676037725
transform -1 0 1564 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input116_A
timestamp 1676037725
transform -1 0 2300 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input117_A
timestamp 1676037725
transform -1 0 1564 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input118_A
timestamp 1676037725
transform -1 0 3956 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 18768 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 16008 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 16284 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 17480 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 20700 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 23368 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 24748 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 25300 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 24932 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 22172 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 21988 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 21344 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 16560 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 16652 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 18860 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21436 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 23000 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 25116 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 24196 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 25208 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 25116 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 19780 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 16560 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 17204 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 16284 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 16100 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 18860 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 22816 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 22264 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 18676 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 10672 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 20700 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 24104 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 25208 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 25392 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 25208 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 24104 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 25300 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 23828 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 23460 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 24656 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 25392 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 24564 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 24380 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 24288 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 24012 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 24012 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21712 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 20424 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 21436 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21252 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 19872 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 19688 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 18860 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 17848 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 17848 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 16928 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 16284 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 15732 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 15364 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 16284 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 15640 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 15364 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 14076 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 13892 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 13524 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 12512 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 13248 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 13800 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 13708 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 11224 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 10212 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 8280 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 8556 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 8280 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 8280 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 8372 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 9936 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 11500 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 10856 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 9660 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 11316 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 13248 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 14444 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 16192 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 18492 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 17756 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 19320 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21528 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 22172 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 24012 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 24656 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 23092 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 21528 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 20056 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 18952 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 18860 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 6716 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1676037725
transform 1 0 9016 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 11224 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 12696 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 14076 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 14076 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 12696 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 12788 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 11500 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 9384 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 11500 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 8096 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 6900 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 8924 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 7268 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 6348 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 8648 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 11132 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 10120 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 11224 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 9660 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 6992 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 7544 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 6900 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 5520 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 6348 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 8372 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 8556 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 9844 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 13248 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 17204 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 20884 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 18860 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 16376 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_1.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 16652 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_1.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 11316 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_1.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 11500 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_3.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 17020 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_3.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 18584 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_3.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 16376 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 20424 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_5.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 21436 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_5.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 20516 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_7.mux_l1_in_0__A0
timestamp 1676037725
transform -1 0 18584 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_7.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 18952 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_7.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 17388 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_7.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_11.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 16284 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_11.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 18676 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_11.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 16100 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_11.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 12604 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_13.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 16744 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_13.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 18124 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_13.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 17020 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_21.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 19320 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_21.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 19504 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_21.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 19412 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_29.mux_l1_in_0__A0
timestamp 1676037725
transform -1 0 17572 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_29.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 17664 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_29.mux_l1_in_2__A0
timestamp 1676037725
transform -1 0 18860 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_37.mux_l1_in_0__A1
timestamp 1676037725
transform -1 0 19228 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_37.mux_l2_in_1__A1
timestamp 1676037725
transform -1 0 12512 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_45.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 19872 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_53.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 16008 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_0.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 22448 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_0.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 21528 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_0.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 23736 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_0.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 23552 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_0.mux_l2_in_1__A1
timestamp 1676037725
transform -1 0 23000 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_2.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 22632 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_2.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 23000 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_2.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 22632 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_2.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 19596 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_2.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 20976 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_4.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 21436 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_4.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 22908 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_4.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 21528 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_4.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 18952 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_6.mux_l1_in_0__A0
timestamp 1676037725
transform -1 0 21712 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_6.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 22632 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_6.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 22448 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_6.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 18952 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_6.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 20332 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_8.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 20516 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_8.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 20148 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_8.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 20792 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_8.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 17756 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_8.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 19044 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_10.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 19320 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_10.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 21068 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_10.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 20332 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_10.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 15548 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_12.mux_l1_in_0__A0
timestamp 1676037725
transform -1 0 20424 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_12.mux_l2_in_0__A0
timestamp 1676037725
transform 1 0 20424 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_12.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 16284 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_14.mux_l1_in_0__A0
timestamp 1676037725
transform -1 0 19228 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_14.mux_l2_in_0__A0
timestamp 1676037725
transform 1 0 18492 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_14.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 15088 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_16.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 18032 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_16.mux_l2_in_0__A0
timestamp 1676037725
transform 1 0 17848 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_16.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 13340 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_18.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 18308 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_18.mux_l2_in_0__A0
timestamp 1676037725
transform 1 0 17848 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_18.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 12696 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_20.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 15180 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_20.mux_l2_in_0__A0
timestamp 1676037725
transform 1 0 16652 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_20.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 12696 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_22.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 14260 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_22.mux_l2_in_0__A0
timestamp 1676037725
transform 1 0 14260 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_22.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 10212 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_24.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 15824 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_24.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 15640 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_24.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 11776 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_26.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 16652 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_26.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 15824 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_26.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 9108 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_28.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 12788 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_28.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 12972 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_28.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 7084 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_30.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 13156 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_30.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 13340 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_30.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 7176 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_32.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 13616 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_32.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 13432 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_32.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 7452 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_34.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 15272 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_34.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 13892 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_34.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 9200 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_36.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 12604 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_36.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 12236 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_36.mux_l2_in_0__A0
timestamp 1676037725
transform 1 0 7176 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_38.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 13064 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_40.mux_l1_in_0__A1
timestamp 1676037725
transform -1 0 15916 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_44.mux_l1_in_0__A1
timestamp 1676037725
transform -1 0 16836 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_46.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 16744 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_46.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 18124 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_48.mux_l1_in_0__A0
timestamp 1676037725
transform -1 0 19136 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_48.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 21712 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_50.mux_l1_in_0__A0
timestamp 1676037725
transform -1 0 25208 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_50.mux_l1_in_0__A1
timestamp 1676037725
transform -1 0 25576 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_52.mux_l1_in_0__A0
timestamp 1676037725
transform -1 0 20148 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_52.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 21068 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_54.mux_l1_in_0__A1
timestamp 1676037725
transform -1 0 19228 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_56.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 18032 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_0.mux_l1_in_0__S
timestamp 1676037725
transform 1 0 9016 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_0.mux_l1_in_1__S
timestamp 1676037725
transform 1 0 17020 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_0.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 14168 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_0.mux_l1_in_2__S
timestamp 1676037725
transform 1 0 15272 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_0.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 9200 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_0.mux_l1_in_3__S
timestamp 1676037725
transform 1 0 10764 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_2.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 14812 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_2.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 11224 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_2.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 11500 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_4.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 14076 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_4.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 9568 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_4.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 9752 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_6.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 8648 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_6.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 12788 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_6.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 6716 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_10.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 7360 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_10.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 12236 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_10.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 6624 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_12.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 8464 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_12.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 8648 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_20.mux_l1_in_0__A1
timestamp 1676037725
transform -1 0 13892 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_20.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 8464 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_20.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 8648 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_28.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 12328 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_28.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 11960 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_28.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 4140 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_36.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 7452 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_44.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 11132 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_52.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 14444 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3864 0 -1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 11224 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 7268 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 4968 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 7176 0 -1 19584
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 11868 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform -1 0 10672 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform -1 0 8648 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 8832 0 -1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 12328 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform -1 0 8004 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform -1 0 6624 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 5612 0 1 16320
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 8556 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform -1 0 7360 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform -1 0 6072 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12696 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_1_
timestamp 1676037725
transform 1 0 13248 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_2_
timestamp 1676037725
transform 1 0 13616 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_3_
timestamp 1676037725
transform 1 0 12604 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_4_
timestamp 1676037725
transform 1 0 10672 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_0_
timestamp 1676037725
transform 1 0 10120 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_1_
timestamp 1676037725
transform 1 0 11684 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_2_
timestamp 1676037725
transform -1 0 8188 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_3__271 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10764 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_3_
timestamp 1676037725
transform 1 0 9568 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l3_in_0_
timestamp 1676037725
transform 1 0 9108 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l3_in_1_
timestamp 1676037725
transform 1 0 7360 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l4_in_0_
timestamp 1676037725
transform 1 0 6532 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 4140 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14904 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_1_
timestamp 1676037725
transform 1 0 14812 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_2_
timestamp 1676037725
transform 1 0 14260 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_3_
timestamp 1676037725
transform 1 0 14260 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_4_
timestamp 1676037725
transform 1 0 11868 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_0_
timestamp 1676037725
transform 1 0 13064 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_1_
timestamp 1676037725
transform 1 0 12512 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_2_
timestamp 1676037725
transform 1 0 9200 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_3__272
timestamp 1676037725
transform -1 0 11224 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_3_
timestamp 1676037725
transform 1 0 11316 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l3_in_0_
timestamp 1676037725
transform 1 0 10396 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l3_in_1_
timestamp 1676037725
transform 1 0 9108 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l4_in_0_
timestamp 1676037725
transform 1 0 7544 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 4876 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15456 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_1_
timestamp 1676037725
transform 1 0 14260 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_2_
timestamp 1676037725
transform 1 0 13892 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_3_
timestamp 1676037725
transform 1 0 12696 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_4_
timestamp 1676037725
transform 1 0 9936 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11776 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_1_
timestamp 1676037725
transform 1 0 11684 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_2_
timestamp 1676037725
transform 1 0 7820 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_3__273
timestamp 1676037725
transform 1 0 9200 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_3_
timestamp 1676037725
transform 1 0 8740 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l3_in_0_
timestamp 1676037725
transform 1 0 8740 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l3_in_1_
timestamp 1676037725
transform 1 0 6992 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l4_in_0_
timestamp 1676037725
transform 1 0 5244 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 3956 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_0_
timestamp 1676037725
transform 1 0 12788 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_1_
timestamp 1676037725
transform 1 0 12420 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_2_
timestamp 1676037725
transform 1 0 13064 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_3_
timestamp 1676037725
transform 1 0 11500 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_4_
timestamp 1676037725
transform 1 0 10304 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_0_
timestamp 1676037725
transform 1 0 10396 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_1_
timestamp 1676037725
transform 1 0 10304 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_2_
timestamp 1676037725
transform 1 0 7636 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3__274
timestamp 1676037725
transform 1 0 9108 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3_
timestamp 1676037725
transform 1 0 8464 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l3_in_0_
timestamp 1676037725
transform 1 0 7728 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l3_in_1_
timestamp 1676037725
transform 1 0 6164 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l4_in_0_
timestamp 1676037725
transform 1 0 5152 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 3680 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3956 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3312 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 4508 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 3312 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 4876 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1676037725
transform 1 0 3956 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1676037725
transform 1 0 3680 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1676037725
transform -1 0 3404 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1676037725
transform -1 0 3312 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 3864 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1676037725
transform 1 0 3956 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1676037725
transform 1 0 3956 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1676037725
transform -1 0 4968 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1676037725
transform -1 0 3220 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 3864 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1676037725
transform 1 0 3956 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1676037725
transform 1 0 3864 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1676037725
transform -1 0 9660 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1676037725
transform -1 0 3496 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_2  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 10212 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 16376 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7912 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_prog_clk
timestamp 1676037725
transform -1 0 11316 0 1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_prog_clk
timestamp 1676037725
transform -1 0 8280 0 -1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_prog_clk
timestamp 1676037725
transform 1 0 10488 0 1 21760
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_prog_clk
timestamp 1676037725
transform -1 0 18952 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_prog_clk
timestamp 1676037725
transform 1 0 20332 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_prog_clk
timestamp 1676037725
transform 1 0 17940 0 1 21760
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_prog_clk
timestamp 1676037725
transform 1 0 20608 0 1 21760
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_prog_clk
timestamp 1676037725
transform -1 0 10120 0 1 35904
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_prog_clk
timestamp 1676037725
transform -1 0 12236 0 1 35904
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_prog_clk
timestamp 1676037725
transform -1 0 9936 0 -1 40256
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_prog_clk
timestamp 1676037725
transform 1 0 11316 0 1 40256
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_prog_clk
timestamp 1676037725
transform -1 0 20424 0 1 36992
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_prog_clk
timestamp 1676037725
transform 1 0 21436 0 1 38080
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_prog_clk
timestamp 1676037725
transform 1 0 17940 0 1 41344
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_prog_clk
timestamp 1676037725
transform -1 0 21528 0 -1 42432
box -38 -48 1050 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1656 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26
timestamp 1676037725
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31
timestamp 1676037725
transform 1 0 3956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5060 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48
timestamp 1676037725
transform 1 0 5520 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1676037725
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59
timestamp 1676037725
transform 1 0 6532 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62
timestamp 1676037725
transform 1 0 6808 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_68
timestamp 1676037725
transform 1 0 7360 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1676037725
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_89
timestamp 1676037725
transform 1 0 9292 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93
timestamp 1676037725
transform 1 0 9660 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1676037725
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1676037725
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_118
timestamp 1676037725
transform 1 0 11960 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1676037725
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_143
timestamp 1676037725
transform 1 0 14260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_161 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15916 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1676037725
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1676037725
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_187 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18308 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 1676037725
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1676037725
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_215
timestamp 1676037725
transform 1 0 20884 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp 1676037725
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1676037725
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_243
timestamp 1676037725
transform 1 0 23460 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251
timestamp 1676037725
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1676037725
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_259
timestamp 1676037725
transform 1 0 24932 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_263
timestamp 1676037725
transform 1 0 25300 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_7
timestamp 1676037725
transform 1 0 1748 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_13
timestamp 1676037725
transform 1 0 2300 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_17
timestamp 1676037725
transform 1 0 2668 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_22
timestamp 1676037725
transform 1 0 3128 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_30
timestamp 1676037725
transform 1 0 3864 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_38
timestamp 1676037725
transform 1 0 4600 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_46
timestamp 1676037725
transform 1 0 5336 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1676037725
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59
timestamp 1676037725
transform 1 0 6532 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_63
timestamp 1676037725
transform 1 0 6900 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_75
timestamp 1676037725
transform 1 0 8004 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_79
timestamp 1676037725
transform 1 0 8372 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_91
timestamp 1676037725
transform 1 0 9476 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_97
timestamp 1676037725
transform 1 0 10028 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1676037725
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_113
timestamp 1676037725
transform 1 0 11500 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_125
timestamp 1676037725
transform 1 0 12604 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_145
timestamp 1676037725
transform 1 0 14444 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_165
timestamp 1676037725
transform 1 0 16284 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1676037725
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_187
timestamp 1676037725
transform 1 0 18308 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_207 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20148 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_219
timestamp 1676037725
transform 1 0 21252 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1676037725
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1676037725
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_237
timestamp 1676037725
transform 1 0 22908 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_243
timestamp 1676037725
transform 1 0 23460 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_264
timestamp 1676037725
transform 1 0 25392 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_9
timestamp 1676037725
transform 1 0 1932 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_16
timestamp 1676037725
transform 1 0 2576 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_20
timestamp 1676037725
transform 1 0 2944 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_25
timestamp 1676037725
transform 1 0 3404 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_34
timestamp 1676037725
transform 1 0 4232 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_39
timestamp 1676037725
transform 1 0 4692 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_45
timestamp 1676037725
transform 1 0 5244 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_52
timestamp 1676037725
transform 1 0 5888 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_56
timestamp 1676037725
transform 1 0 6256 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_61
timestamp 1676037725
transform 1 0 6716 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_67
timestamp 1676037725
transform 1 0 7268 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_73
timestamp 1676037725
transform 1 0 7820 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_81
timestamp 1676037725
transform 1 0 8556 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_85
timestamp 1676037725
transform 1 0 8924 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_93
timestamp 1676037725
transform 1 0 9660 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_107
timestamp 1676037725
transform 1 0 10948 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_115
timestamp 1676037725
transform 1 0 11684 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_119
timestamp 1676037725
transform 1 0 12052 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1676037725
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_141
timestamp 1676037725
transform 1 0 14076 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_159
timestamp 1676037725
transform 1 0 15732 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_179
timestamp 1676037725
transform 1 0 17572 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_191
timestamp 1676037725
transform 1 0 18676 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1676037725
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1676037725
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_215
timestamp 1676037725
transform 1 0 20884 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_235
timestamp 1676037725
transform 1 0 22724 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_239
timestamp 1676037725
transform 1 0 23092 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_250
timestamp 1676037725
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_255
timestamp 1676037725
transform 1 0 24564 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_258
timestamp 1676037725
transform 1 0 24840 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_264
timestamp 1676037725
transform 1 0 25392 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_8
timestamp 1676037725
transform 1 0 1840 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_13
timestamp 1676037725
transform 1 0 2300 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_21
timestamp 1676037725
transform 1 0 3036 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_24
timestamp 1676037725
transform 1 0 3312 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_36
timestamp 1676037725
transform 1 0 4416 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_44
timestamp 1676037725
transform 1 0 5152 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_49
timestamp 1676037725
transform 1 0 5612 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1676037725
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_69
timestamp 1676037725
transform 1 0 7452 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_77
timestamp 1676037725
transform 1 0 8188 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_81
timestamp 1676037725
transform 1 0 8556 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_93
timestamp 1676037725
transform 1 0 9660 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_97
timestamp 1676037725
transform 1 0 10028 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_109
timestamp 1676037725
transform 1 0 11132 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1676037725
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_127
timestamp 1676037725
transform 1 0 12788 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_145
timestamp 1676037725
transform 1 0 14444 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_157
timestamp 1676037725
transform 1 0 15548 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_165
timestamp 1676037725
transform 1 0 16284 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_169
timestamp 1676037725
transform 1 0 16652 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_187
timestamp 1676037725
transform 1 0 18308 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_207
timestamp 1676037725
transform 1 0 20148 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_219
timestamp 1676037725
transform 1 0 21252 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1676037725
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_225
timestamp 1676037725
transform 1 0 21804 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_243
timestamp 1676037725
transform 1 0 23460 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_263
timestamp 1676037725
transform 1 0 25300 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5
timestamp 1676037725
transform 1 0 1564 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_17
timestamp 1676037725
transform 1 0 2668 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_25
timestamp 1676037725
transform 1 0 3404 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1676037725
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1676037725
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1676037725
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1676037725
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1676037725
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1676037725
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1676037725
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1676037725
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1676037725
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1676037725
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1676037725
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1676037725
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1676037725
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_193
timestamp 1676037725
transform 1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_197
timestamp 1676037725
transform 1 0 19228 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_215
timestamp 1676037725
transform 1 0 20884 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_235
timestamp 1676037725
transform 1 0 22724 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_247
timestamp 1676037725
transform 1 0 23828 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1676037725
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_253
timestamp 1676037725
transform 1 0 24380 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_264
timestamp 1676037725
transform 1 0 25392 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1676037725
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1676037725
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1676037725
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1676037725
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1676037725
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1676037725
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1676037725
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1676037725
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1676037725
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1676037725
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1676037725
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1676037725
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1676037725
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1676037725
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_165
timestamp 1676037725
transform 1 0 16284 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1676037725
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_197
timestamp 1676037725
transform 1 0 19228 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1676037725
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1676037725
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_225
timestamp 1676037725
transform 1 0 21804 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_243
timestamp 1676037725
transform 1 0 23460 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_247
timestamp 1676037725
transform 1 0 23828 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_264
timestamp 1676037725
transform 1 0 25392 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1676037725
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1676037725
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1676037725
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1676037725
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1676037725
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1676037725
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1676037725
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1676037725
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1676037725
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1676037725
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1676037725
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1676037725
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1676037725
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1676037725
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1676037725
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1676037725
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1676037725
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1676037725
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_197
timestamp 1676037725
transform 1 0 19228 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_208
timestamp 1676037725
transform 1 0 20240 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_212
timestamp 1676037725
transform 1 0 20608 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_229
timestamp 1676037725
transform 1 0 22172 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_249
timestamp 1676037725
transform 1 0 24012 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1676037725
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_265
timestamp 1676037725
transform 1 0 25484 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1676037725
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1676037725
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1676037725
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1676037725
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1676037725
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1676037725
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1676037725
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1676037725
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1676037725
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1676037725
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1676037725
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1676037725
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1676037725
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1676037725
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1676037725
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1676037725
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1676037725
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1676037725
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_193
timestamp 1676037725
transform 1 0 18860 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_197
timestamp 1676037725
transform 1 0 19228 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_202
timestamp 1676037725
transform 1 0 19688 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_222
timestamp 1676037725
transform 1 0 21528 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_225
timestamp 1676037725
transform 1 0 21804 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_244
timestamp 1676037725
transform 1 0 23552 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_264
timestamp 1676037725
transform 1 0 25392 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1676037725
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1676037725
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1676037725
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1676037725
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1676037725
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1676037725
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1676037725
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1676037725
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1676037725
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1676037725
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1676037725
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1676037725
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1676037725
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1676037725
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1676037725
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_177
timestamp 1676037725
transform 1 0 17388 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1676037725
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1676037725
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_197
timestamp 1676037725
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_202
timestamp 1676037725
transform 1 0 19688 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_230
timestamp 1676037725
transform 1 0 22264 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp 1676037725
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_253
timestamp 1676037725
transform 1 0 24380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_258
timestamp 1676037725
transform 1 0 24840 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1676037725
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1676037725
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1676037725
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1676037725
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1676037725
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1676037725
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1676037725
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1676037725
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1676037725
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1676037725
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1676037725
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1676037725
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1676037725
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1676037725
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1676037725
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1676037725
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1676037725
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1676037725
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1676037725
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_205
timestamp 1676037725
transform 1 0 19964 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_222
timestamp 1676037725
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_225
timestamp 1676037725
transform 1 0 21804 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_244
timestamp 1676037725
transform 1 0 23552 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_264
timestamp 1676037725
transform 1 0 25392 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1676037725
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1676037725
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1676037725
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1676037725
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1676037725
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1676037725
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1676037725
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1676037725
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1676037725
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1676037725
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1676037725
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1676037725
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1676037725
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1676037725
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1676037725
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1676037725
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1676037725
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_189
timestamp 1676037725
transform 1 0 18492 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_194
timestamp 1676037725
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_197
timestamp 1676037725
transform 1 0 19228 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_205
timestamp 1676037725
transform 1 0 19964 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_212
timestamp 1676037725
transform 1 0 20608 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_224
timestamp 1676037725
transform 1 0 21712 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_232
timestamp 1676037725
transform 1 0 22448 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_250
timestamp 1676037725
transform 1 0 24104 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_253
timestamp 1676037725
transform 1 0 24380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_259
timestamp 1676037725
transform 1 0 24932 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_265
timestamp 1676037725
transform 1 0 25484 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1676037725
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1676037725
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_27
timestamp 1676037725
transform 1 0 3588 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_53
timestamp 1676037725
transform 1 0 5980 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_59
timestamp 1676037725
transform 1 0 6532 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_71
timestamp 1676037725
transform 1 0 7636 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_83
timestamp 1676037725
transform 1 0 8740 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_95
timestamp 1676037725
transform 1 0 9844 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_107
timestamp 1676037725
transform 1 0 10948 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1676037725
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1676037725
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1676037725
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1676037725
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1676037725
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1676037725
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1676037725
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1676037725
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1676037725
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1676037725
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1676037725
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1676037725
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1676037725
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_225
timestamp 1676037725
transform 1 0 21804 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_244
timestamp 1676037725
transform 1 0 23552 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_264
timestamp 1676037725
transform 1 0 25392 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1676037725
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1676037725
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1676037725
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1676037725
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1676037725
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1676037725
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1676037725
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1676037725
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1676037725
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1676037725
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1676037725
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1676037725
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1676037725
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1676037725
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1676037725
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1676037725
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_153
timestamp 1676037725
transform 1 0 15180 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_161
timestamp 1676037725
transform 1 0 15916 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_166
timestamp 1676037725
transform 1 0 16376 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_178
timestamp 1676037725
transform 1 0 17480 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_186
timestamp 1676037725
transform 1 0 18216 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_192
timestamp 1676037725
transform 1 0 18768 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1676037725
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1676037725
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1676037725
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_233
timestamp 1676037725
transform 1 0 22540 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_242
timestamp 1676037725
transform 1 0 23368 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_250
timestamp 1676037725
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_253
timestamp 1676037725
transform 1 0 24380 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_259
timestamp 1676037725
transform 1 0 24932 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_265
timestamp 1676037725
transform 1 0 25484 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1676037725
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1676037725
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1676037725
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1676037725
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1676037725
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_57
timestamp 1676037725
transform 1 0 6348 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_68
timestamp 1676037725
transform 1 0 7360 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_80
timestamp 1676037725
transform 1 0 8464 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_92
timestamp 1676037725
transform 1 0 9568 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_104
timestamp 1676037725
transform 1 0 10672 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1676037725
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1676037725
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_137
timestamp 1676037725
transform 1 0 13708 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_147
timestamp 1676037725
transform 1 0 14628 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_159
timestamp 1676037725
transform 1 0 15732 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1676037725
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1676037725
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1676037725
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1676037725
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1676037725
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1676037725
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1676037725
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_225
timestamp 1676037725
transform 1 0 21804 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_230
timestamp 1676037725
transform 1 0 22264 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_242
timestamp 1676037725
transform 1 0 23368 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_264
timestamp 1676037725
transform 1 0 25392 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1676037725
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1676037725
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1676037725
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1676037725
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1676037725
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1676037725
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1676037725
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1676037725
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1676037725
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1676037725
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1676037725
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_109
timestamp 1676037725
transform 1 0 11132 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_117
timestamp 1676037725
transform 1 0 11868 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_129
timestamp 1676037725
transform 1 0 12972 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_137
timestamp 1676037725
transform 1 0 13708 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1676037725
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1676037725
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_165
timestamp 1676037725
transform 1 0 16284 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_175
timestamp 1676037725
transform 1 0 17204 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_187
timestamp 1676037725
transform 1 0 18308 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1676037725
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1676037725
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1676037725
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_221
timestamp 1676037725
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_233
timestamp 1676037725
transform 1 0 22540 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_250
timestamp 1676037725
transform 1 0 24104 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1676037725
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_258
timestamp 1676037725
transform 1 0 24840 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1676037725
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1676037725
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1676037725
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1676037725
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1676037725
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1676037725
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1676037725
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1676037725
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1676037725
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1676037725
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1676037725
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1676037725
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1676037725
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1676037725
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_137
timestamp 1676037725
transform 1 0 13708 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_15_147
timestamp 1676037725
transform 1 0 14628 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_153
timestamp 1676037725
transform 1 0 15180 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_156
timestamp 1676037725
transform 1 0 15456 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1676037725
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_181
timestamp 1676037725
transform 1 0 17756 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_204
timestamp 1676037725
transform 1 0 19872 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_208
timestamp 1676037725
transform 1 0 20240 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_216
timestamp 1676037725
transform 1 0 20976 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_220
timestamp 1676037725
transform 1 0 21344 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1676037725
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_237
timestamp 1676037725
transform 1 0 22908 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_245
timestamp 1676037725
transform 1 0 23644 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_264
timestamp 1676037725
transform 1 0 25392 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1676037725
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1676037725
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1676037725
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1676037725
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1676037725
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1676037725
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1676037725
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1676037725
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1676037725
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1676037725
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1676037725
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_109
timestamp 1676037725
transform 1 0 11132 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_130
timestamp 1676037725
transform 1 0 13064 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_134
timestamp 1676037725
transform 1 0 13432 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1676037725
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_152
timestamp 1676037725
transform 1 0 15088 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1676037725
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_177
timestamp 1676037725
transform 1 0 17388 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_16_188
timestamp 1676037725
transform 1 0 18400 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_197
timestamp 1676037725
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_208
timestamp 1676037725
transform 1 0 20240 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_215
timestamp 1676037725
transform 1 0 20884 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_227
timestamp 1676037725
transform 1 0 21988 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_16_238
timestamp 1676037725
transform 1 0 23000 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_246
timestamp 1676037725
transform 1 0 23736 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_250
timestamp 1676037725
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_253
timestamp 1676037725
transform 1 0 24380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_259
timestamp 1676037725
transform 1 0 24932 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_265
timestamp 1676037725
transform 1 0 25484 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1676037725
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1676037725
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1676037725
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1676037725
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1676037725
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1676037725
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1676037725
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1676037725
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1676037725
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1676037725
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1676037725
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1676037725
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1676037725
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_145
timestamp 1676037725
transform 1 0 14444 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_149
timestamp 1676037725
transform 1 0 14812 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_159
timestamp 1676037725
transform 1 0 15732 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1676037725
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1676037725
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1676037725
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_193
timestamp 1676037725
transform 1 0 18860 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_196
timestamp 1676037725
transform 1 0 19136 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_200
timestamp 1676037725
transform 1 0 19504 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_204
timestamp 1676037725
transform 1 0 19872 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_212
timestamp 1676037725
transform 1 0 20608 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_216
timestamp 1676037725
transform 1 0 20976 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_17_225
timestamp 1676037725
transform 1 0 21804 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_231
timestamp 1676037725
transform 1 0 22356 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_235
timestamp 1676037725
transform 1 0 22724 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_239
timestamp 1676037725
transform 1 0 23092 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_243
timestamp 1676037725
transform 1 0 23460 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_247
timestamp 1676037725
transform 1 0 23828 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_264
timestamp 1676037725
transform 1 0 25392 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1676037725
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1676037725
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1676037725
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1676037725
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1676037725
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1676037725
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1676037725
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1676037725
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1676037725
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_85
timestamp 1676037725
transform 1 0 8924 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_109
timestamp 1676037725
transform 1 0 11132 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_113
timestamp 1676037725
transform 1 0 11500 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_125
timestamp 1676037725
transform 1 0 12604 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_130
timestamp 1676037725
transform 1 0 13064 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1676037725
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1676037725
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_152
timestamp 1676037725
transform 1 0 15088 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_160
timestamp 1676037725
transform 1 0 15824 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_167
timestamp 1676037725
transform 1 0 16468 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_171
timestamp 1676037725
transform 1 0 16836 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1676037725
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_197
timestamp 1676037725
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_203
timestamp 1676037725
transform 1 0 19780 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_207
timestamp 1676037725
transform 1 0 20148 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_213
timestamp 1676037725
transform 1 0 20700 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_217
timestamp 1676037725
transform 1 0 21068 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_221
timestamp 1676037725
transform 1 0 21436 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_224
timestamp 1676037725
transform 1 0 21712 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_232
timestamp 1676037725
transform 1 0 22448 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_250
timestamp 1676037725
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1676037725
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_258
timestamp 1676037725
transform 1 0 24840 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1676037725
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1676037725
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1676037725
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1676037725
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1676037725
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1676037725
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1676037725
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1676037725
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_81
timestamp 1676037725
transform 1 0 8556 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1676037725
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1676037725
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1676037725
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_113
timestamp 1676037725
transform 1 0 11500 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_125
timestamp 1676037725
transform 1 0 12604 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_129
timestamp 1676037725
transform 1 0 12972 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_132
timestamp 1676037725
transform 1 0 13248 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_138
timestamp 1676037725
transform 1 0 13800 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_162
timestamp 1676037725
transform 1 0 16008 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1676037725
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1676037725
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_180
timestamp 1676037725
transform 1 0 17664 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_193
timestamp 1676037725
transform 1 0 18860 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_197
timestamp 1676037725
transform 1 0 19228 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_201
timestamp 1676037725
transform 1 0 19596 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1676037725
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_225
timestamp 1676037725
transform 1 0 21804 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_244
timestamp 1676037725
transform 1 0 23552 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_264
timestamp 1676037725
transform 1 0 25392 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1676037725
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1676037725
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1676037725
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1676037725
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1676037725
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_53
timestamp 1676037725
transform 1 0 5980 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_61
timestamp 1676037725
transform 1 0 6716 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 1676037725
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_87
timestamp 1676037725
transform 1 0 9108 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_99
timestamp 1676037725
transform 1 0 10212 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_111
timestamp 1676037725
transform 1 0 11316 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_128
timestamp 1676037725
transform 1 0 12880 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_132
timestamp 1676037725
transform 1 0 13248 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_20_143
timestamp 1676037725
transform 1 0 14260 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_153
timestamp 1676037725
transform 1 0 15180 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_157
timestamp 1676037725
transform 1 0 15548 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_172
timestamp 1676037725
transform 1 0 16928 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_176
timestamp 1676037725
transform 1 0 17296 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_181
timestamp 1676037725
transform 1 0 17756 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1676037725
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_199
timestamp 1676037725
transform 1 0 19412 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_205
timestamp 1676037725
transform 1 0 19964 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_209
timestamp 1676037725
transform 1 0 20332 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_213
timestamp 1676037725
transform 1 0 20700 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_234
timestamp 1676037725
transform 1 0 22632 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_241
timestamp 1676037725
transform 1 0 23276 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_248
timestamp 1676037725
transform 1 0 23920 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1676037725
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_265
timestamp 1676037725
transform 1 0 25484 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1676037725
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_21
timestamp 1676037725
transform 1 0 3036 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_33
timestamp 1676037725
transform 1 0 4140 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_45
timestamp 1676037725
transform 1 0 5244 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_53
timestamp 1676037725
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1676037725
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_69
timestamp 1676037725
transform 1 0 7452 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_77
timestamp 1676037725
transform 1 0 8188 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_82
timestamp 1676037725
transform 1 0 8648 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_107
timestamp 1676037725
transform 1 0 10948 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1676037725
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_113
timestamp 1676037725
transform 1 0 11500 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_121
timestamp 1676037725
transform 1 0 12236 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_124
timestamp 1676037725
transform 1 0 12512 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_135
timestamp 1676037725
transform 1 0 13524 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_148
timestamp 1676037725
transform 1 0 14720 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_152
timestamp 1676037725
transform 1 0 15088 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_157
timestamp 1676037725
transform 1 0 15548 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_163
timestamp 1676037725
transform 1 0 16100 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1676037725
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1676037725
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_191
timestamp 1676037725
transform 1 0 18676 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_198
timestamp 1676037725
transform 1 0 19320 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_202
timestamp 1676037725
transform 1 0 19688 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_207
timestamp 1676037725
transform 1 0 20148 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_211
timestamp 1676037725
transform 1 0 20516 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1676037725
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_225
timestamp 1676037725
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_230
timestamp 1676037725
transform 1 0 22264 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_237
timestamp 1676037725
transform 1 0 22908 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_241
timestamp 1676037725
transform 1 0 23276 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_247
timestamp 1676037725
transform 1 0 23828 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_264
timestamp 1676037725
transform 1 0 25392 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1676037725
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1676037725
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1676037725
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1676037725
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1676037725
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_53
timestamp 1676037725
transform 1 0 5980 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_61
timestamp 1676037725
transform 1 0 6716 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1676037725
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_85
timestamp 1676037725
transform 1 0 8924 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_97
timestamp 1676037725
transform 1 0 10028 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_122
timestamp 1676037725
transform 1 0 12328 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_126
timestamp 1676037725
transform 1 0 12696 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_136
timestamp 1676037725
transform 1 0 13616 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_141
timestamp 1676037725
transform 1 0 14076 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_149
timestamp 1676037725
transform 1 0 14812 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_171
timestamp 1676037725
transform 1 0 16836 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_175
timestamp 1676037725
transform 1 0 17204 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_179
timestamp 1676037725
transform 1 0 17572 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_187
timestamp 1676037725
transform 1 0 18308 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1676037725
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1676037725
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1676037725
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_221
timestamp 1676037725
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_233
timestamp 1676037725
transform 1 0 22540 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_242
timestamp 1676037725
transform 1 0 23368 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_250
timestamp 1676037725
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1676037725
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_265
timestamp 1676037725
transform 1 0 25484 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1676037725
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1676037725
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1676037725
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1676037725
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1676037725
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1676037725
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1676037725
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1676037725
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_81
timestamp 1676037725
transform 1 0 8556 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_104
timestamp 1676037725
transform 1 0 10672 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_108
timestamp 1676037725
transform 1 0 11040 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_113
timestamp 1676037725
transform 1 0 11500 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_121
timestamp 1676037725
transform 1 0 12236 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_126
timestamp 1676037725
transform 1 0 12696 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_139
timestamp 1676037725
transform 1 0 13892 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_151
timestamp 1676037725
transform 1 0 14996 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_159
timestamp 1676037725
transform 1 0 15732 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1676037725
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_171
timestamp 1676037725
transform 1 0 16836 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_182
timestamp 1676037725
transform 1 0 17848 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_186
timestamp 1676037725
transform 1 0 18216 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_192
timestamp 1676037725
transform 1 0 18768 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_205
timestamp 1676037725
transform 1 0 19964 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_212
timestamp 1676037725
transform 1 0 20608 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_218
timestamp 1676037725
transform 1 0 21160 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_222
timestamp 1676037725
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_225
timestamp 1676037725
transform 1 0 21804 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_244
timestamp 1676037725
transform 1 0 23552 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_264
timestamp 1676037725
transform 1 0 25392 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1676037725
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1676037725
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1676037725
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1676037725
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1676037725
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_53
timestamp 1676037725
transform 1 0 5980 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_75
timestamp 1676037725
transform 1 0 8004 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_79
timestamp 1676037725
transform 1 0 8372 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1676037725
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1676037725
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_97
timestamp 1676037725
transform 1 0 10028 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_120
timestamp 1676037725
transform 1 0 12144 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_124
timestamp 1676037725
transform 1 0 12512 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_128
timestamp 1676037725
transform 1 0 12880 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1676037725
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_147
timestamp 1676037725
transform 1 0 14628 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_151
timestamp 1676037725
transform 1 0 14996 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_159
timestamp 1676037725
transform 1 0 15732 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_181
timestamp 1676037725
transform 1 0 17756 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_194
timestamp 1676037725
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_197
timestamp 1676037725
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_208
timestamp 1676037725
transform 1 0 20240 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_215
timestamp 1676037725
transform 1 0 20884 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_219
timestamp 1676037725
transform 1 0 21252 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_230
timestamp 1676037725
transform 1 0 22264 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_250
timestamp 1676037725
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1676037725
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_265
timestamp 1676037725
transform 1 0 25484 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1676037725
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_21
timestamp 1676037725
transform 1 0 3036 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_33
timestamp 1676037725
transform 1 0 4140 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_45
timestamp 1676037725
transform 1 0 5244 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_53
timestamp 1676037725
transform 1 0 5980 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1676037725
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_69
timestamp 1676037725
transform 1 0 7452 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_79
timestamp 1676037725
transform 1 0 8372 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_92
timestamp 1676037725
transform 1 0 9568 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_100
timestamp 1676037725
transform 1 0 10304 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1676037725
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1676037725
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1676037725
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1676037725
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_158
timestamp 1676037725
transform 1 0 15640 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1676037725
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_171
timestamp 1676037725
transform 1 0 16836 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_179
timestamp 1676037725
transform 1 0 17572 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_183
timestamp 1676037725
transform 1 0 17940 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_195
timestamp 1676037725
transform 1 0 19044 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_199
timestamp 1676037725
transform 1 0 19412 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_203
timestamp 1676037725
transform 1 0 19780 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_207
timestamp 1676037725
transform 1 0 20148 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_214
timestamp 1676037725
transform 1 0 20792 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_222
timestamp 1676037725
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_225
timestamp 1676037725
transform 1 0 21804 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_244
timestamp 1676037725
transform 1 0 23552 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_264
timestamp 1676037725
transform 1 0 25392 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_3
timestamp 1676037725
transform 1 0 1380 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_11
timestamp 1676037725
transform 1 0 2116 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_18
timestamp 1676037725
transform 1 0 2760 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_26
timestamp 1676037725
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1676037725
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_41
timestamp 1676037725
transform 1 0 4876 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_72
timestamp 1676037725
transform 1 0 7728 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_76
timestamp 1676037725
transform 1 0 8096 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_85
timestamp 1676037725
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_96
timestamp 1676037725
transform 1 0 9936 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_109
timestamp 1676037725
transform 1 0 11132 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_113
timestamp 1676037725
transform 1 0 11500 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1676037725
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_143
timestamp 1676037725
transform 1 0 14260 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_155
timestamp 1676037725
transform 1 0 15364 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_162
timestamp 1676037725
transform 1 0 16008 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_166
timestamp 1676037725
transform 1 0 16376 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_178
timestamp 1676037725
transform 1 0 17480 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_190
timestamp 1676037725
transform 1 0 18584 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_26_197
timestamp 1676037725
transform 1 0 19228 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_203
timestamp 1676037725
transform 1 0 19780 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_213
timestamp 1676037725
transform 1 0 20700 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_221
timestamp 1676037725
transform 1 0 21436 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_243
timestamp 1676037725
transform 1 0 23460 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_250
timestamp 1676037725
transform 1 0 24104 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_255
timestamp 1676037725
transform 1 0 24564 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_263
timestamp 1676037725
transform 1 0 25300 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1676037725
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1676037725
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1676037725
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_39
timestamp 1676037725
transform 1 0 4692 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1676037725
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_57
timestamp 1676037725
transform 1 0 6348 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_63
timestamp 1676037725
transform 1 0 6900 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_73
timestamp 1676037725
transform 1 0 7820 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_81
timestamp 1676037725
transform 1 0 8556 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_92
timestamp 1676037725
transform 1 0 9568 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_107
timestamp 1676037725
transform 1 0 10948 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1676037725
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 1676037725
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_124
timestamp 1676037725
transform 1 0 12512 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_130
timestamp 1676037725
transform 1 0 13064 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_141
timestamp 1676037725
transform 1 0 14076 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_27_151
timestamp 1676037725
transform 1 0 14996 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1676037725
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_171
timestamp 1676037725
transform 1 0 16836 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_175
timestamp 1676037725
transform 1 0 17204 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_196
timestamp 1676037725
transform 1 0 19136 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_200
timestamp 1676037725
transform 1 0 19504 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_222
timestamp 1676037725
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_225
timestamp 1676037725
transform 1 0 21804 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_247
timestamp 1676037725
transform 1 0 23828 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_251
timestamp 1676037725
transform 1 0 24196 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_263
timestamp 1676037725
transform 1 0 25300 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1676037725
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1676037725
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1676037725
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_29
timestamp 1676037725
transform 1 0 3772 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_37
timestamp 1676037725
transform 1 0 4508 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_60
timestamp 1676037725
transform 1 0 6624 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_64
timestamp 1676037725
transform 1 0 6992 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_68
timestamp 1676037725
transform 1 0 7360 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_79
timestamp 1676037725
transform 1 0 8372 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_85
timestamp 1676037725
transform 1 0 8924 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_93
timestamp 1676037725
transform 1 0 9660 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_97
timestamp 1676037725
transform 1 0 10028 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_111
timestamp 1676037725
transform 1 0 11316 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_115
timestamp 1676037725
transform 1 0 11684 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_123
timestamp 1676037725
transform 1 0 12420 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_133
timestamp 1676037725
transform 1 0 13340 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_137
timestamp 1676037725
transform 1 0 13708 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_141
timestamp 1676037725
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_152
timestamp 1676037725
transform 1 0 15088 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_156
timestamp 1676037725
transform 1 0 15456 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_160
timestamp 1676037725
transform 1 0 15824 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_182
timestamp 1676037725
transform 1 0 17848 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_190
timestamp 1676037725
transform 1 0 18584 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1676037725
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_219
timestamp 1676037725
transform 1 0 21252 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_227
timestamp 1676037725
transform 1 0 21988 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_231
timestamp 1676037725
transform 1 0 22356 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_250
timestamp 1676037725
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1676037725
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_265
timestamp 1676037725
transform 1 0 25484 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1676037725
transform 1 0 1380 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_21
timestamp 1676037725
transform 1 0 3036 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_33
timestamp 1676037725
transform 1 0 4140 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_45
timestamp 1676037725
transform 1 0 5244 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_53
timestamp 1676037725
transform 1 0 5980 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1676037725
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_69
timestamp 1676037725
transform 1 0 7452 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_73
timestamp 1676037725
transform 1 0 7820 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_85
timestamp 1676037725
transform 1 0 8924 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_110
timestamp 1676037725
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_115
timestamp 1676037725
transform 1 0 11684 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_121
timestamp 1676037725
transform 1 0 12236 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_132
timestamp 1676037725
transform 1 0 13248 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_145
timestamp 1676037725
transform 1 0 14444 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_157
timestamp 1676037725
transform 1 0 15548 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_165
timestamp 1676037725
transform 1 0 16284 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_169
timestamp 1676037725
transform 1 0 16652 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_176
timestamp 1676037725
transform 1 0 17296 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_181
timestamp 1676037725
transform 1 0 17756 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_194
timestamp 1676037725
transform 1 0 18952 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_202
timestamp 1676037725
transform 1 0 19688 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_207
timestamp 1676037725
transform 1 0 20148 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_220
timestamp 1676037725
transform 1 0 21344 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_225
timestamp 1676037725
transform 1 0 21804 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_233
timestamp 1676037725
transform 1 0 22540 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_254
timestamp 1676037725
transform 1 0 24472 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_258
timestamp 1676037725
transform 1 0 24840 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_30_3
timestamp 1676037725
transform 1 0 1380 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_9
timestamp 1676037725
transform 1 0 1932 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_13
timestamp 1676037725
transform 1 0 2300 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_25
timestamp 1676037725
transform 1 0 3404 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_29
timestamp 1676037725
transform 1 0 3772 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_34
timestamp 1676037725
transform 1 0 4232 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_46
timestamp 1676037725
transform 1 0 5336 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_58
timestamp 1676037725
transform 1 0 6440 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_82
timestamp 1676037725
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_85
timestamp 1676037725
transform 1 0 8924 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_91
timestamp 1676037725
transform 1 0 9476 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_95
timestamp 1676037725
transform 1 0 9844 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_99
timestamp 1676037725
transform 1 0 10212 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_102
timestamp 1676037725
transform 1 0 10488 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_113
timestamp 1676037725
transform 1 0 11500 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_121
timestamp 1676037725
transform 1 0 12236 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_124
timestamp 1676037725
transform 1 0 12512 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_135
timestamp 1676037725
transform 1 0 13524 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1676037725
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1676037725
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1676037725
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_165
timestamp 1676037725
transform 1 0 16284 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_169
timestamp 1676037725
transform 1 0 16652 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_172
timestamp 1676037725
transform 1 0 16928 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_183
timestamp 1676037725
transform 1 0 17940 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_187
timestamp 1676037725
transform 1 0 18308 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_193
timestamp 1676037725
transform 1 0 18860 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_197
timestamp 1676037725
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_208
timestamp 1676037725
transform 1 0 20240 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_212
timestamp 1676037725
transform 1 0 20608 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_222
timestamp 1676037725
transform 1 0 21528 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_226
timestamp 1676037725
transform 1 0 21896 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_248
timestamp 1676037725
transform 1 0 23920 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1676037725
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_259
timestamp 1676037725
transform 1 0 24932 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_265
timestamp 1676037725
transform 1 0 25484 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1676037725
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1676037725
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1676037725
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_39
timestamp 1676037725
transform 1 0 4692 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_44
timestamp 1676037725
transform 1 0 5152 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_57
timestamp 1676037725
transform 1 0 6348 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_61
timestamp 1676037725
transform 1 0 6716 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_64
timestamp 1676037725
transform 1 0 6992 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_89
timestamp 1676037725
transform 1 0 9292 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_93
timestamp 1676037725
transform 1 0 9660 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_110
timestamp 1676037725
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1676037725
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_125
timestamp 1676037725
transform 1 0 12604 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_128
timestamp 1676037725
transform 1 0 12880 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_139
timestamp 1676037725
transform 1 0 13892 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_143
timestamp 1676037725
transform 1 0 14260 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_155
timestamp 1676037725
transform 1 0 15364 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1676037725
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_169
timestamp 1676037725
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_173
timestamp 1676037725
transform 1 0 17020 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_179
timestamp 1676037725
transform 1 0 17572 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_186
timestamp 1676037725
transform 1 0 18216 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_193
timestamp 1676037725
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_205
timestamp 1676037725
transform 1 0 19964 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp 1676037725
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_225
timestamp 1676037725
transform 1 0 21804 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_244
timestamp 1676037725
transform 1 0 23552 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_264
timestamp 1676037725
transform 1 0 25392 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_3
timestamp 1676037725
transform 1 0 1380 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_9
timestamp 1676037725
transform 1 0 1932 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_13
timestamp 1676037725
transform 1 0 2300 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_25
timestamp 1676037725
transform 1 0 3404 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1676037725
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_41
timestamp 1676037725
transform 1 0 4876 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_32_67
timestamp 1676037725
transform 1 0 7268 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_71
timestamp 1676037725
transform 1 0 7636 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_82
timestamp 1676037725
transform 1 0 8648 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_85
timestamp 1676037725
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_96
timestamp 1676037725
transform 1 0 9936 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_32_104
timestamp 1676037725
transform 1 0 10672 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_110
timestamp 1676037725
transform 1 0 11224 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_120
timestamp 1676037725
transform 1 0 12144 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_124
timestamp 1676037725
transform 1 0 12512 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_136
timestamp 1676037725
transform 1 0 13616 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1676037725
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_153
timestamp 1676037725
transform 1 0 15180 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_32_164
timestamp 1676037725
transform 1 0 16192 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_32_172
timestamp 1676037725
transform 1 0 16928 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_178
timestamp 1676037725
transform 1 0 17480 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_191
timestamp 1676037725
transform 1 0 18676 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1676037725
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_197
timestamp 1676037725
transform 1 0 19228 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_202
timestamp 1676037725
transform 1 0 19688 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_214
timestamp 1676037725
transform 1 0 20792 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_222
timestamp 1676037725
transform 1 0 21528 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_230
timestamp 1676037725
transform 1 0 22264 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_250
timestamp 1676037725
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1676037725
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_265
timestamp 1676037725
transform 1 0 25484 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1676037725
transform 1 0 1380 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_21
timestamp 1676037725
transform 1 0 3036 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_29
timestamp 1676037725
transform 1 0 3772 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_50
timestamp 1676037725
transform 1 0 5704 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 1676037725
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_57
timestamp 1676037725
transform 1 0 6348 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_63
timestamp 1676037725
transform 1 0 6900 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_66
timestamp 1676037725
transform 1 0 7176 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_77
timestamp 1676037725
transform 1 0 8188 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_102
timestamp 1676037725
transform 1 0 10488 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_106
timestamp 1676037725
transform 1 0 10856 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1676037725
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_113
timestamp 1676037725
transform 1 0 11500 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_124
timestamp 1676037725
transform 1 0 12512 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_136
timestamp 1676037725
transform 1 0 13616 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_153
timestamp 1676037725
transform 1 0 15180 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_160
timestamp 1676037725
transform 1 0 15824 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_169
timestamp 1676037725
transform 1 0 16652 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_180
timestamp 1676037725
transform 1 0 17664 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_188
timestamp 1676037725
transform 1 0 18400 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_211
timestamp 1676037725
transform 1 0 20516 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_215
timestamp 1676037725
transform 1 0 20884 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1676037725
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_225
timestamp 1676037725
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_236
timestamp 1676037725
transform 1 0 22816 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_240
timestamp 1676037725
transform 1 0 23184 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_261
timestamp 1676037725
transform 1 0 25116 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_265
timestamp 1676037725
transform 1 0 25484 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1676037725
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_15
timestamp 1676037725
transform 1 0 2484 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_26
timestamp 1676037725
transform 1 0 3496 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_29
timestamp 1676037725
transform 1 0 3772 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_33
timestamp 1676037725
transform 1 0 4140 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_36
timestamp 1676037725
transform 1 0 4416 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_34_62
timestamp 1676037725
transform 1 0 6808 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_66
timestamp 1676037725
transform 1 0 7176 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_69
timestamp 1676037725
transform 1 0 7452 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_80
timestamp 1676037725
transform 1 0 8464 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1676037725
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_97
timestamp 1676037725
transform 1 0 10028 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_109
timestamp 1676037725
transform 1 0 11132 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_115
timestamp 1676037725
transform 1 0 11684 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_126
timestamp 1676037725
transform 1 0 12696 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_134
timestamp 1676037725
transform 1 0 13432 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_138
timestamp 1676037725
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_141
timestamp 1676037725
transform 1 0 14076 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_163
timestamp 1676037725
transform 1 0 16100 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_167
timestamp 1676037725
transform 1 0 16468 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_172
timestamp 1676037725
transform 1 0 16928 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_184
timestamp 1676037725
transform 1 0 18032 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_194
timestamp 1676037725
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_197
timestamp 1676037725
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_202
timestamp 1676037725
transform 1 0 19688 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_210
timestamp 1676037725
transform 1 0 20424 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_232
timestamp 1676037725
transform 1 0 22448 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_240
timestamp 1676037725
transform 1 0 23184 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_244
timestamp 1676037725
transform 1 0 23552 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1676037725
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_265
timestamp 1676037725
transform 1 0 25484 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1676037725
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_23
timestamp 1676037725
transform 1 0 3220 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_27
timestamp 1676037725
transform 1 0 3588 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_31
timestamp 1676037725
transform 1 0 3956 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_35
timestamp 1676037725
transform 1 0 4324 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_42
timestamp 1676037725
transform 1 0 4968 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_54
timestamp 1676037725
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_57
timestamp 1676037725
transform 1 0 6348 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_68
timestamp 1676037725
transform 1 0 7360 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_81
timestamp 1676037725
transform 1 0 8556 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_89
timestamp 1676037725
transform 1 0 9292 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_94
timestamp 1676037725
transform 1 0 9752 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_105
timestamp 1676037725
transform 1 0 10764 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_109
timestamp 1676037725
transform 1 0 11132 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_35_117
timestamp 1676037725
transform 1 0 11868 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_125
timestamp 1676037725
transform 1 0 12604 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_135
timestamp 1676037725
transform 1 0 13524 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_148
timestamp 1676037725
transform 1 0 14720 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_154
timestamp 1676037725
transform 1 0 15272 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_159
timestamp 1676037725
transform 1 0 15732 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1676037725
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_169
timestamp 1676037725
transform 1 0 16652 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_177
timestamp 1676037725
transform 1 0 17388 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_180
timestamp 1676037725
transform 1 0 17664 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_183
timestamp 1676037725
transform 1 0 17940 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_194
timestamp 1676037725
transform 1 0 18952 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_200
timestamp 1676037725
transform 1 0 19504 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_221
timestamp 1676037725
transform 1 0 21436 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1676037725
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_230
timestamp 1676037725
transform 1 0 22264 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_257
timestamp 1676037725
transform 1 0 24748 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_261
timestamp 1676037725
transform 1 0 25116 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_265
timestamp 1676037725
transform 1 0 25484 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_3
timestamp 1676037725
transform 1 0 1380 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_9
timestamp 1676037725
transform 1 0 1932 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_13
timestamp 1676037725
transform 1 0 2300 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_20
timestamp 1676037725
transform 1 0 2944 0 1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1676037725
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1676037725
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_53
timestamp 1676037725
transform 1 0 5980 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_64
timestamp 1676037725
transform 1 0 6992 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1676037725
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1676037725
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1676037725
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_97
timestamp 1676037725
transform 1 0 10028 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_101
timestamp 1676037725
transform 1 0 10396 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_113
timestamp 1676037725
transform 1 0 11500 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_126
timestamp 1676037725
transform 1 0 12696 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_130
timestamp 1676037725
transform 1 0 13064 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_134
timestamp 1676037725
transform 1 0 13432 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_141
timestamp 1676037725
transform 1 0 14076 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_152
timestamp 1676037725
transform 1 0 15088 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_156
timestamp 1676037725
transform 1 0 15456 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_178
timestamp 1676037725
transform 1 0 17480 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_182
timestamp 1676037725
transform 1 0 17848 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_194
timestamp 1676037725
transform 1 0 18952 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_197
timestamp 1676037725
transform 1 0 19228 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_208
timestamp 1676037725
transform 1 0 20240 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_223
timestamp 1676037725
transform 1 0 21620 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_229
timestamp 1676037725
transform 1 0 22172 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_233
timestamp 1676037725
transform 1 0 22540 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_250
timestamp 1676037725
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_253
timestamp 1676037725
transform 1 0 24380 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_259
timestamp 1676037725
transform 1 0 24932 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_263
timestamp 1676037725
transform 1 0 25300 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_3
timestamp 1676037725
transform 1 0 1380 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_12
timestamp 1676037725
transform 1 0 2208 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_24
timestamp 1676037725
transform 1 0 3312 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_37_33
timestamp 1676037725
transform 1 0 4140 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_41
timestamp 1676037725
transform 1 0 4876 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_37_53
timestamp 1676037725
transform 1 0 5980 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_37_57
timestamp 1676037725
transform 1 0 6348 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_65
timestamp 1676037725
transform 1 0 7084 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_78
timestamp 1676037725
transform 1 0 8280 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_102
timestamp 1676037725
transform 1 0 10488 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_108
timestamp 1676037725
transform 1 0 11040 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_113
timestamp 1676037725
transform 1 0 11500 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_129
timestamp 1676037725
transform 1 0 12972 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_153
timestamp 1676037725
transform 1 0 15180 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_160
timestamp 1676037725
transform 1 0 15824 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_164
timestamp 1676037725
transform 1 0 16192 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_169
timestamp 1676037725
transform 1 0 16652 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_180
timestamp 1676037725
transform 1 0 17664 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_187
timestamp 1676037725
transform 1 0 18308 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_218
timestamp 1676037725
transform 1 0 21160 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_222
timestamp 1676037725
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_225
timestamp 1676037725
transform 1 0 21804 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_233
timestamp 1676037725
transform 1 0 22540 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_257
timestamp 1676037725
transform 1 0 24748 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_264
timestamp 1676037725
transform 1 0 25392 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_3
timestamp 1676037725
transform 1 0 1380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_21
timestamp 1676037725
transform 1 0 3036 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1676037725
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_29
timestamp 1676037725
transform 1 0 3772 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_36
timestamp 1676037725
transform 1 0 4416 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_68
timestamp 1676037725
transform 1 0 7360 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_72
timestamp 1676037725
transform 1 0 7728 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_80
timestamp 1676037725
transform 1 0 8464 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_85
timestamp 1676037725
transform 1 0 8924 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_90
timestamp 1676037725
transform 1 0 9384 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_101
timestamp 1676037725
transform 1 0 10396 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_108
timestamp 1676037725
transform 1 0 11040 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_121
timestamp 1676037725
transform 1 0 12236 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_134
timestamp 1676037725
transform 1 0 13432 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_138
timestamp 1676037725
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1676037725
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1676037725
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_165
timestamp 1676037725
transform 1 0 16284 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_173
timestamp 1676037725
transform 1 0 17020 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_194
timestamp 1676037725
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_199
timestamp 1676037725
transform 1 0 19412 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_227
timestamp 1676037725
transform 1 0 21988 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_231
timestamp 1676037725
transform 1 0 22356 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_250
timestamp 1676037725
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_253
timestamp 1676037725
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_264
timestamp 1676037725
transform 1 0 25392 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_3
timestamp 1676037725
transform 1 0 1380 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_9
timestamp 1676037725
transform 1 0 1932 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_30
timestamp 1676037725
transform 1 0 3864 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_54
timestamp 1676037725
transform 1 0 6072 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_59
timestamp 1676037725
transform 1 0 6532 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_71
timestamp 1676037725
transform 1 0 7636 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_79
timestamp 1676037725
transform 1 0 8372 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_89
timestamp 1676037725
transform 1 0 9292 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_102
timestamp 1676037725
transform 1 0 10488 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_39_109
timestamp 1676037725
transform 1 0 11132 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_39_115
timestamp 1676037725
transform 1 0 11684 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_121
timestamp 1676037725
transform 1 0 12236 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_131
timestamp 1676037725
transform 1 0 13156 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_138
timestamp 1676037725
transform 1 0 13800 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_150
timestamp 1676037725
transform 1 0 14904 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_156
timestamp 1676037725
transform 1 0 15456 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_166
timestamp 1676037725
transform 1 0 16376 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_169
timestamp 1676037725
transform 1 0 16652 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_177
timestamp 1676037725
transform 1 0 17388 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_181
timestamp 1676037725
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_193
timestamp 1676037725
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_205
timestamp 1676037725
transform 1 0 19964 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_39_213
timestamp 1676037725
transform 1 0 20700 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_221
timestamp 1676037725
transform 1 0 21436 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_39_225
timestamp 1676037725
transform 1 0 21804 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_244
timestamp 1676037725
transform 1 0 23552 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_264
timestamp 1676037725
transform 1 0 25392 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1676037725
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_17
timestamp 1676037725
transform 1 0 2668 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_25
timestamp 1676037725
transform 1 0 3404 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_29
timestamp 1676037725
transform 1 0 3772 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_34
timestamp 1676037725
transform 1 0 4232 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_38
timestamp 1676037725
transform 1 0 4600 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_50
timestamp 1676037725
transform 1 0 5704 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_62
timestamp 1676037725
transform 1 0 6808 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_68
timestamp 1676037725
transform 1 0 7360 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_71
timestamp 1676037725
transform 1 0 7636 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_82
timestamp 1676037725
transform 1 0 8648 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_85
timestamp 1676037725
transform 1 0 8924 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_107
timestamp 1676037725
transform 1 0 10948 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_111
timestamp 1676037725
transform 1 0 11316 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_122
timestamp 1676037725
transform 1 0 12328 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_127
timestamp 1676037725
transform 1 0 12788 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_138
timestamp 1676037725
transform 1 0 13800 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_141
timestamp 1676037725
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_152
timestamp 1676037725
transform 1 0 15088 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_165
timestamp 1676037725
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_179
timestamp 1676037725
transform 1 0 17572 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_190
timestamp 1676037725
transform 1 0 18584 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_40_197
timestamp 1676037725
transform 1 0 19228 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_209
timestamp 1676037725
transform 1 0 20332 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_222
timestamp 1676037725
transform 1 0 21528 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_250
timestamp 1676037725
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_253
timestamp 1676037725
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_259
timestamp 1676037725
transform 1 0 24932 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_265
timestamp 1676037725
transform 1 0 25484 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_3
timestamp 1676037725
transform 1 0 1380 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_9
timestamp 1676037725
transform 1 0 1932 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_13
timestamp 1676037725
transform 1 0 2300 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_41
timestamp 1676037725
transform 1 0 4876 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_45
timestamp 1676037725
transform 1 0 5244 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_53
timestamp 1676037725
transform 1 0 5980 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_41_57
timestamp 1676037725
transform 1 0 6348 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_65
timestamp 1676037725
transform 1 0 7084 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_70
timestamp 1676037725
transform 1 0 7544 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_94
timestamp 1676037725
transform 1 0 9752 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_98
timestamp 1676037725
transform 1 0 10120 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_110
timestamp 1676037725
transform 1 0 11224 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_113
timestamp 1676037725
transform 1 0 11500 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_118
timestamp 1676037725
transform 1 0 11960 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_129
timestamp 1676037725
transform 1 0 12972 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_133
timestamp 1676037725
transform 1 0 13340 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_145
timestamp 1676037725
transform 1 0 14444 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_166
timestamp 1676037725
transform 1 0 16376 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_171
timestamp 1676037725
transform 1 0 16836 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_192
timestamp 1676037725
transform 1 0 18768 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_196
timestamp 1676037725
transform 1 0 19136 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_206
timestamp 1676037725
transform 1 0 20056 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_218
timestamp 1676037725
transform 1 0 21160 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_41_225
timestamp 1676037725
transform 1 0 21804 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_236
timestamp 1676037725
transform 1 0 22816 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_260
timestamp 1676037725
transform 1 0 25024 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_264
timestamp 1676037725
transform 1 0 25392 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_3
timestamp 1676037725
transform 1 0 1380 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_21
timestamp 1676037725
transform 1 0 3036 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_25
timestamp 1676037725
transform 1 0 3404 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_29
timestamp 1676037725
transform 1 0 3772 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_37
timestamp 1676037725
transform 1 0 4508 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_49
timestamp 1676037725
transform 1 0 5612 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_77
timestamp 1676037725
transform 1 0 8188 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_81
timestamp 1676037725
transform 1 0 8556 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_85
timestamp 1676037725
transform 1 0 8924 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_90
timestamp 1676037725
transform 1 0 9384 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_102
timestamp 1676037725
transform 1 0 10488 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_114
timestamp 1676037725
transform 1 0 11592 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_122
timestamp 1676037725
transform 1 0 12328 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_128
timestamp 1676037725
transform 1 0 12880 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_141
timestamp 1676037725
transform 1 0 14076 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_149
timestamp 1676037725
transform 1 0 14812 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_161
timestamp 1676037725
transform 1 0 15916 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_174
timestamp 1676037725
transform 1 0 17112 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_182
timestamp 1676037725
transform 1 0 17848 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_186
timestamp 1676037725
transform 1 0 18216 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_192
timestamp 1676037725
transform 1 0 18768 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1676037725
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1676037725
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_209
timestamp 1676037725
transform 1 0 20332 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_230
timestamp 1676037725
transform 1 0 22264 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_243
timestamp 1676037725
transform 1 0 23460 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_250
timestamp 1676037725
transform 1 0 24104 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_253
timestamp 1676037725
transform 1 0 24380 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_258
timestamp 1676037725
transform 1 0 24840 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_262
timestamp 1676037725
transform 1 0 25208 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1676037725
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_15
timestamp 1676037725
transform 1 0 2484 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_24
timestamp 1676037725
transform 1 0 3312 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_31
timestamp 1676037725
transform 1 0 3956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_43
timestamp 1676037725
transform 1 0 5060 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1676037725
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_57
timestamp 1676037725
transform 1 0 6348 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_67
timestamp 1676037725
transform 1 0 7268 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_78
timestamp 1676037725
transform 1 0 8280 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_85
timestamp 1676037725
transform 1 0 8924 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_93
timestamp 1676037725
transform 1 0 9660 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1676037725
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1676037725
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_43_113
timestamp 1676037725
transform 1 0 11500 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_136
timestamp 1676037725
transform 1 0 13616 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_140
timestamp 1676037725
transform 1 0 13984 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_152
timestamp 1676037725
transform 1 0 15088 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_160
timestamp 1676037725
transform 1 0 15824 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_43_165
timestamp 1676037725
transform 1 0 16284 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_43_169
timestamp 1676037725
transform 1 0 16652 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_193
timestamp 1676037725
transform 1 0 18860 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_206
timestamp 1676037725
transform 1 0 20056 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_213
timestamp 1676037725
transform 1 0 20700 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_217
timestamp 1676037725
transform 1 0 21068 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_222
timestamp 1676037725
transform 1 0 21528 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_225
timestamp 1676037725
transform 1 0 21804 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_236
timestamp 1676037725
transform 1 0 22816 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_240
timestamp 1676037725
transform 1 0 23184 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_246
timestamp 1676037725
transform 1 0 23736 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_254
timestamp 1676037725
transform 1 0 24472 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_262
timestamp 1676037725
transform 1 0 25208 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1676037725
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1676037725
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1676037725
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_29
timestamp 1676037725
transform 1 0 3772 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_52
timestamp 1676037725
transform 1 0 5888 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_76
timestamp 1676037725
transform 1 0 8096 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_80
timestamp 1676037725
transform 1 0 8464 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_85
timestamp 1676037725
transform 1 0 8924 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_89
timestamp 1676037725
transform 1 0 9292 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_95
timestamp 1676037725
transform 1 0 9844 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_108
timestamp 1676037725
transform 1 0 11040 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_120
timestamp 1676037725
transform 1 0 12144 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_126
timestamp 1676037725
transform 1 0 12696 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_136
timestamp 1676037725
transform 1 0 13616 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_141
timestamp 1676037725
transform 1 0 14076 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_145
timestamp 1676037725
transform 1 0 14444 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_166
timestamp 1676037725
transform 1 0 16376 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_44_170
timestamp 1676037725
transform 1 0 16744 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_175
timestamp 1676037725
transform 1 0 17204 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_186
timestamp 1676037725
transform 1 0 18216 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_194
timestamp 1676037725
transform 1 0 18952 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_197
timestamp 1676037725
transform 1 0 19228 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_201
timestamp 1676037725
transform 1 0 19596 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_212
timestamp 1676037725
transform 1 0 20608 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_220
timestamp 1676037725
transform 1 0 21344 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_242
timestamp 1676037725
transform 1 0 23368 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_246
timestamp 1676037725
transform 1 0 23736 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_250
timestamp 1676037725
transform 1 0 24104 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_253
timestamp 1676037725
transform 1 0 24380 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_259
timestamp 1676037725
transform 1 0 24932 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_44_263
timestamp 1676037725
transform 1 0 25300 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_45_3
timestamp 1676037725
transform 1 0 1380 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_9
timestamp 1676037725
transform 1 0 1932 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_13
timestamp 1676037725
transform 1 0 2300 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_21
timestamp 1676037725
transform 1 0 3036 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1676037725
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1676037725
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1676037725
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1676037725
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_57
timestamp 1676037725
transform 1 0 6348 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_65
timestamp 1676037725
transform 1 0 7084 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_68
timestamp 1676037725
transform 1 0 7360 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_79
timestamp 1676037725
transform 1 0 8372 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_86
timestamp 1676037725
transform 1 0 9016 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_94
timestamp 1676037725
transform 1 0 9752 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_45_106
timestamp 1676037725
transform 1 0 10856 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_45_113
timestamp 1676037725
transform 1 0 11500 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_135
timestamp 1676037725
transform 1 0 13524 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_139
timestamp 1676037725
transform 1 0 13892 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_156
timestamp 1676037725
transform 1 0 15456 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_162
timestamp 1676037725
transform 1 0 16008 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_171
timestamp 1676037725
transform 1 0 16836 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_175
timestamp 1676037725
transform 1 0 17204 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_186
timestamp 1676037725
transform 1 0 18216 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_192
timestamp 1676037725
transform 1 0 18768 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_204
timestamp 1676037725
transform 1 0 19872 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_216
timestamp 1676037725
transform 1 0 20976 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_225
timestamp 1676037725
transform 1 0 21804 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_249
timestamp 1676037725
transform 1 0 24012 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_253
timestamp 1676037725
transform 1 0 24380 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_259
timestamp 1676037725
transform 1 0 24932 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_45_265
timestamp 1676037725
transform 1 0 25484 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_3
timestamp 1676037725
transform 1 0 1380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_21
timestamp 1676037725
transform 1 0 3036 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1676037725
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_29
timestamp 1676037725
transform 1 0 3772 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_52
timestamp 1676037725
transform 1 0 5888 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_76
timestamp 1676037725
transform 1 0 8096 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_80
timestamp 1676037725
transform 1 0 8464 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1676037725
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_97
timestamp 1676037725
transform 1 0 10028 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_103
timestamp 1676037725
transform 1 0 10580 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_107
timestamp 1676037725
transform 1 0 10948 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_119
timestamp 1676037725
transform 1 0 12052 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_124
timestamp 1676037725
transform 1 0 12512 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_135
timestamp 1676037725
transform 1 0 13524 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1676037725
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_141
timestamp 1676037725
transform 1 0 14076 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_152
timestamp 1676037725
transform 1 0 15088 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_156
timestamp 1676037725
transform 1 0 15456 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_166
timestamp 1676037725
transform 1 0 16376 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_179
timestamp 1676037725
transform 1 0 17572 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_192
timestamp 1676037725
transform 1 0 18768 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_197
timestamp 1676037725
transform 1 0 19228 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_219
timestamp 1676037725
transform 1 0 21252 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_223
timestamp 1676037725
transform 1 0 21620 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_229
timestamp 1676037725
transform 1 0 22172 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_250
timestamp 1676037725
transform 1 0 24104 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_253
timestamp 1676037725
transform 1 0 24380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_259
timestamp 1676037725
transform 1 0 24932 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_265
timestamp 1676037725
transform 1 0 25484 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1676037725
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1676037725
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1676037725
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1676037725
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1676037725
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1676037725
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_57
timestamp 1676037725
transform 1 0 6348 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_79
timestamp 1676037725
transform 1 0 8372 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_83
timestamp 1676037725
transform 1 0 8740 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_87
timestamp 1676037725
transform 1 0 9108 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_108
timestamp 1676037725
transform 1 0 11040 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_113
timestamp 1676037725
transform 1 0 11500 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_126
timestamp 1676037725
transform 1 0 12696 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_130
timestamp 1676037725
transform 1 0 13064 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_134
timestamp 1676037725
transform 1 0 13432 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_47_138
timestamp 1676037725
transform 1 0 13800 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_141
timestamp 1676037725
transform 1 0 14076 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_152
timestamp 1676037725
transform 1 0 15088 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_156
timestamp 1676037725
transform 1 0 15456 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_169
timestamp 1676037725
transform 1 0 16652 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_180
timestamp 1676037725
transform 1 0 17664 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_193
timestamp 1676037725
transform 1 0 18860 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_200
timestamp 1676037725
transform 1 0 19504 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_208
timestamp 1676037725
transform 1 0 20240 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_212
timestamp 1676037725
transform 1 0 20608 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_220
timestamp 1676037725
transform 1 0 21344 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1676037725
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_225
timestamp 1676037725
transform 1 0 21804 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_236
timestamp 1676037725
transform 1 0 22816 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_240
timestamp 1676037725
transform 1 0 23184 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_244
timestamp 1676037725
transform 1 0 23552 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_251
timestamp 1676037725
transform 1 0 24196 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_259
timestamp 1676037725
transform 1 0 24932 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_263
timestamp 1676037725
transform 1 0 25300 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1676037725
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1676037725
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1676037725
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_29
timestamp 1676037725
transform 1 0 3772 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_52
timestamp 1676037725
transform 1 0 5888 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_76
timestamp 1676037725
transform 1 0 8096 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_85
timestamp 1676037725
transform 1 0 8924 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_96
timestamp 1676037725
transform 1 0 9936 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_108
timestamp 1676037725
transform 1 0 11040 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_130
timestamp 1676037725
transform 1 0 13064 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_136
timestamp 1676037725
transform 1 0 13616 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_141
timestamp 1676037725
transform 1 0 14076 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_145
timestamp 1676037725
transform 1 0 14444 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_166
timestamp 1676037725
transform 1 0 16376 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_48_170
timestamp 1676037725
transform 1 0 16744 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_182
timestamp 1676037725
transform 1 0 17848 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_189
timestamp 1676037725
transform 1 0 18492 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_48_193
timestamp 1676037725
transform 1 0 18860 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_48_197
timestamp 1676037725
transform 1 0 19228 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_208
timestamp 1676037725
transform 1 0 20240 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_221
timestamp 1676037725
transform 1 0 21436 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_234
timestamp 1676037725
transform 1 0 22632 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_238
timestamp 1676037725
transform 1 0 23000 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_246
timestamp 1676037725
transform 1 0 23736 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_250
timestamp 1676037725
transform 1 0 24104 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_257
timestamp 1676037725
transform 1 0 24748 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_264
timestamp 1676037725
transform 1 0 25392 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1676037725
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1676037725
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1676037725
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1676037725
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1676037725
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1676037725
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1676037725
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_69
timestamp 1676037725
transform 1 0 7452 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_97
timestamp 1676037725
transform 1 0 10028 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_101
timestamp 1676037725
transform 1 0 10396 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_109
timestamp 1676037725
transform 1 0 11132 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_49_113
timestamp 1676037725
transform 1 0 11500 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_49_125
timestamp 1676037725
transform 1 0 12604 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_135
timestamp 1676037725
transform 1 0 13524 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_143
timestamp 1676037725
transform 1 0 14260 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_49_166
timestamp 1676037725
transform 1 0 16376 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_171
timestamp 1676037725
transform 1 0 16836 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_179
timestamp 1676037725
transform 1 0 17572 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_201
timestamp 1676037725
transform 1 0 19596 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_205
timestamp 1676037725
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1676037725
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1676037725
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_225
timestamp 1676037725
transform 1 0 21804 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_230
timestamp 1676037725
transform 1 0 22264 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_242
timestamp 1676037725
transform 1 0 23368 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_246
timestamp 1676037725
transform 1 0 23736 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_251
timestamp 1676037725
transform 1 0 24196 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_259
timestamp 1676037725
transform 1 0 24932 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_263
timestamp 1676037725
transform 1 0 25300 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_3
timestamp 1676037725
transform 1 0 1380 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_21
timestamp 1676037725
transform 1 0 3036 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1676037725
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_29
timestamp 1676037725
transform 1 0 3772 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_52
timestamp 1676037725
transform 1 0 5888 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_64
timestamp 1676037725
transform 1 0 6992 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_76
timestamp 1676037725
transform 1 0 8096 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_85
timestamp 1676037725
transform 1 0 8924 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_50_96
timestamp 1676037725
transform 1 0 9936 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_50_101
timestamp 1676037725
transform 1 0 10396 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_112
timestamp 1676037725
transform 1 0 11408 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_125
timestamp 1676037725
transform 1 0 12604 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_138
timestamp 1676037725
transform 1 0 13800 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1676037725
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1676037725
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_165
timestamp 1676037725
transform 1 0 16284 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_169
timestamp 1676037725
transform 1 0 16652 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_172
timestamp 1676037725
transform 1 0 16928 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_183
timestamp 1676037725
transform 1 0 17940 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_187
timestamp 1676037725
transform 1 0 18308 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1676037725
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_197
timestamp 1676037725
transform 1 0 19228 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_208
timestamp 1676037725
transform 1 0 20240 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_223
timestamp 1676037725
transform 1 0 21620 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_236
timestamp 1676037725
transform 1 0 22816 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_50_249
timestamp 1676037725
transform 1 0 24012 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_50_253
timestamp 1676037725
transform 1 0 24380 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_264
timestamp 1676037725
transform 1 0 25392 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1676037725
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1676037725
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1676037725
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1676037725
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1676037725
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1676037725
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1676037725
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_69
timestamp 1676037725
transform 1 0 7452 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_91
timestamp 1676037725
transform 1 0 9476 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_95
timestamp 1676037725
transform 1 0 9844 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_107
timestamp 1676037725
transform 1 0 10948 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1676037725
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_113
timestamp 1676037725
transform 1 0 11500 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_51_118
timestamp 1676037725
transform 1 0 11960 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_51_123
timestamp 1676037725
transform 1 0 12420 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_134
timestamp 1676037725
transform 1 0 13432 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_146
timestamp 1676037725
transform 1 0 14536 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_51_158
timestamp 1676037725
transform 1 0 15640 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_51_162
timestamp 1676037725
transform 1 0 16008 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1676037725
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_171
timestamp 1676037725
transform 1 0 16836 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_175
timestamp 1676037725
transform 1 0 17204 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_185
timestamp 1676037725
transform 1 0 18124 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_198
timestamp 1676037725
transform 1 0 19320 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_211
timestamp 1676037725
transform 1 0 20516 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1676037725
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_225
timestamp 1676037725
transform 1 0 21804 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_51_236
timestamp 1676037725
transform 1 0 22816 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_242
timestamp 1676037725
transform 1 0 23368 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_51_263
timestamp 1676037725
transform 1 0 25300 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1676037725
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1676037725
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1676037725
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1676037725
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1676037725
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_53
timestamp 1676037725
transform 1 0 5980 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_63
timestamp 1676037725
transform 1 0 6900 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_74
timestamp 1676037725
transform 1 0 7912 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_82
timestamp 1676037725
transform 1 0 8648 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1676037725
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_97
timestamp 1676037725
transform 1 0 10028 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_103
timestamp 1676037725
transform 1 0 10580 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_124
timestamp 1676037725
transform 1 0 12512 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_128
timestamp 1676037725
transform 1 0 12880 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_138
timestamp 1676037725
transform 1 0 13800 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_141
timestamp 1676037725
transform 1 0 14076 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_163
timestamp 1676037725
transform 1 0 16100 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_176
timestamp 1676037725
transform 1 0 17296 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_189
timestamp 1676037725
transform 1 0 18492 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_52_193
timestamp 1676037725
transform 1 0 18860 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_52_197
timestamp 1676037725
transform 1 0 19228 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_202
timestamp 1676037725
transform 1 0 19688 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_52_219
timestamp 1676037725
transform 1 0 21252 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_227
timestamp 1676037725
transform 1 0 21988 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_52_250
timestamp 1676037725
transform 1 0 24104 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_253
timestamp 1676037725
transform 1 0 24380 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_258
timestamp 1676037725
transform 1 0 24840 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1676037725
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1676037725
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_27
timestamp 1676037725
transform 1 0 3588 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_53_35
timestamp 1676037725
transform 1 0 4324 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_46
timestamp 1676037725
transform 1 0 5336 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_54
timestamp 1676037725
transform 1 0 6072 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_53_57
timestamp 1676037725
transform 1 0 6348 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_53_62
timestamp 1676037725
transform 1 0 6808 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_73
timestamp 1676037725
transform 1 0 7820 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_80
timestamp 1676037725
transform 1 0 8464 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_87
timestamp 1676037725
transform 1 0 9108 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_91
timestamp 1676037725
transform 1 0 9476 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_96
timestamp 1676037725
transform 1 0 9936 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_107
timestamp 1676037725
transform 1 0 10948 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1676037725
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_113
timestamp 1676037725
transform 1 0 11500 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_121
timestamp 1676037725
transform 1 0 12236 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_53_126
timestamp 1676037725
transform 1 0 12696 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_129
timestamp 1676037725
transform 1 0 12972 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_141
timestamp 1676037725
transform 1 0 14076 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_153
timestamp 1676037725
transform 1 0 15180 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_165
timestamp 1676037725
transform 1 0 16284 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_53_169
timestamp 1676037725
transform 1 0 16652 0 -1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_53_184
timestamp 1676037725
transform 1 0 18032 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_196
timestamp 1676037725
transform 1 0 19136 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_53_202
timestamp 1676037725
transform 1 0 19688 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_208
timestamp 1676037725
transform 1 0 20240 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_211
timestamp 1676037725
transform 1 0 20516 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_219
timestamp 1676037725
transform 1 0 21252 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_53_225
timestamp 1676037725
transform 1 0 21804 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_230
timestamp 1676037725
transform 1 0 22264 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_234
timestamp 1676037725
transform 1 0 22632 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_245
timestamp 1676037725
transform 1 0 23644 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_249
timestamp 1676037725
transform 1 0 24012 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_252
timestamp 1676037725
transform 1 0 24288 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_264
timestamp 1676037725
transform 1 0 25392 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1676037725
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1676037725
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1676037725
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1676037725
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_41
timestamp 1676037725
transform 1 0 4876 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_64
timestamp 1676037725
transform 1 0 6992 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_68
timestamp 1676037725
transform 1 0 7360 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_78
timestamp 1676037725
transform 1 0 8280 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_54_85
timestamp 1676037725
transform 1 0 8924 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_107
timestamp 1676037725
transform 1 0 10948 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_54_111
timestamp 1676037725
transform 1 0 11316 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_117
timestamp 1676037725
transform 1 0 11868 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_120
timestamp 1676037725
transform 1 0 12144 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_131
timestamp 1676037725
transform 1 0 13156 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1676037725
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1676037725
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_173
timestamp 1676037725
transform 1 0 17020 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_54_179
timestamp 1676037725
transform 1 0 17572 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_182
timestamp 1676037725
transform 1 0 17848 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_197
timestamp 1676037725
transform 1 0 19228 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_209
timestamp 1676037725
transform 1 0 20332 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_222
timestamp 1676037725
transform 1 0 21528 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_235
timestamp 1676037725
transform 1 0 22724 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_242
timestamp 1676037725
transform 1 0 23368 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_248
timestamp 1676037725
transform 1 0 23920 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_253
timestamp 1676037725
transform 1 0 24380 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_259
timestamp 1676037725
transform 1 0 24932 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_264
timestamp 1676037725
transform 1 0 25392 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_3
timestamp 1676037725
transform 1 0 1380 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_8
timestamp 1676037725
transform 1 0 1840 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_12
timestamp 1676037725
transform 1 0 2208 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_24
timestamp 1676037725
transform 1 0 3312 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_36
timestamp 1676037725
transform 1 0 4416 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_55_45
timestamp 1676037725
transform 1 0 5244 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_53
timestamp 1676037725
transform 1 0 5980 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_55_57
timestamp 1676037725
transform 1 0 6348 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_63
timestamp 1676037725
transform 1 0 6900 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_55_66
timestamp 1676037725
transform 1 0 7176 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_55_72
timestamp 1676037725
transform 1 0 7728 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_55_83
timestamp 1676037725
transform 1 0 8740 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_108
timestamp 1676037725
transform 1 0 11040 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1676037725
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_125
timestamp 1676037725
transform 1 0 12604 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_128
timestamp 1676037725
transform 1 0 12880 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_132
timestamp 1676037725
transform 1 0 13248 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_136
timestamp 1676037725
transform 1 0 13616 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_144
timestamp 1676037725
transform 1 0 14352 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_55_165
timestamp 1676037725
transform 1 0 16284 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_55_169
timestamp 1676037725
transform 1 0 16652 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_180
timestamp 1676037725
transform 1 0 17664 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_193
timestamp 1676037725
transform 1 0 18860 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_206
timestamp 1676037725
transform 1 0 20056 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_55_221
timestamp 1676037725
transform 1 0 21436 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_55_225
timestamp 1676037725
transform 1 0 21804 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_230
timestamp 1676037725
transform 1 0 22264 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_243
timestamp 1676037725
transform 1 0 23460 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_250
timestamp 1676037725
transform 1 0 24104 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_256
timestamp 1676037725
transform 1 0 24656 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_259
timestamp 1676037725
transform 1 0 24932 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_264
timestamp 1676037725
transform 1 0 25392 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1676037725
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1676037725
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1676037725
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1676037725
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_41
timestamp 1676037725
transform 1 0 4876 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_47
timestamp 1676037725
transform 1 0 5428 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_68
timestamp 1676037725
transform 1 0 7360 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_72
timestamp 1676037725
transform 1 0 7728 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_85
timestamp 1676037725
transform 1 0 8924 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_96
timestamp 1676037725
transform 1 0 9936 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_100
timestamp 1676037725
transform 1 0 10304 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_112
timestamp 1676037725
transform 1 0 11408 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_124
timestamp 1676037725
transform 1 0 12512 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_56_137
timestamp 1676037725
transform 1 0 13708 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_56_141
timestamp 1676037725
transform 1 0 14076 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_145
timestamp 1676037725
transform 1 0 14444 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_157
timestamp 1676037725
transform 1 0 15548 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_56_167
timestamp 1676037725
transform 1 0 16468 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_191
timestamp 1676037725
transform 1 0 18676 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1676037725
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_56_197
timestamp 1676037725
transform 1 0 19228 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_56_203
timestamp 1676037725
transform 1 0 19780 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_209
timestamp 1676037725
transform 1 0 20332 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_230
timestamp 1676037725
transform 1 0 22264 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_243
timestamp 1676037725
transform 1 0 23460 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1676037725
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_253
timestamp 1676037725
transform 1 0 24380 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_259
timestamp 1676037725
transform 1 0 24932 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_264
timestamp 1676037725
transform 1 0 25392 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1676037725
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1676037725
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1676037725
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1676037725
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1676037725
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1676037725
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1676037725
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_69
timestamp 1676037725
transform 1 0 7452 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_92
timestamp 1676037725
transform 1 0 9568 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_105
timestamp 1676037725
transform 1 0 10764 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_109
timestamp 1676037725
transform 1 0 11132 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_115
timestamp 1676037725
transform 1 0 11684 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_57_126
timestamp 1676037725
transform 1 0 12696 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_57_143
timestamp 1676037725
transform 1 0 14260 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_156
timestamp 1676037725
transform 1 0 15456 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1676037725
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_181
timestamp 1676037725
transform 1 0 17756 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_185
timestamp 1676037725
transform 1 0 18124 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_195
timestamp 1676037725
transform 1 0 19044 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_207
timestamp 1676037725
transform 1 0 20148 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_219
timestamp 1676037725
transform 1 0 21252 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1676037725
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_225
timestamp 1676037725
transform 1 0 21804 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_229
timestamp 1676037725
transform 1 0 22172 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_232
timestamp 1676037725
transform 1 0 22448 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_240
timestamp 1676037725
transform 1 0 23184 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_57_264
timestamp 1676037725
transform 1 0 25392 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1676037725
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1676037725
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1676037725
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1676037725
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_61
timestamp 1676037725
transform 1 0 6716 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1676037725
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_77
timestamp 1676037725
transform 1 0 8188 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_81
timestamp 1676037725
transform 1 0 8556 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_85
timestamp 1676037725
transform 1 0 8924 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_96
timestamp 1676037725
transform 1 0 9936 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_108
timestamp 1676037725
transform 1 0 11040 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_120
timestamp 1676037725
transform 1 0 12144 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_130
timestamp 1676037725
transform 1 0 13064 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_134
timestamp 1676037725
transform 1 0 13432 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_58_137
timestamp 1676037725
transform 1 0 13708 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1676037725
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1676037725
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_165
timestamp 1676037725
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_177
timestamp 1676037725
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_189
timestamp 1676037725
transform 1 0 18492 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_58_193
timestamp 1676037725
transform 1 0 18860 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_197
timestamp 1676037725
transform 1 0 19228 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_58_208
timestamp 1676037725
transform 1 0 20240 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_58_234
timestamp 1676037725
transform 1 0 22632 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_58_238
timestamp 1676037725
transform 1 0 23000 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_58_247
timestamp 1676037725
transform 1 0 23828 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1676037725
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_253
timestamp 1676037725
transform 1 0 24380 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_258
timestamp 1676037725
transform 1 0 24840 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_3
timestamp 1676037725
transform 1 0 1380 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_8
timestamp 1676037725
transform 1 0 1840 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_12
timestamp 1676037725
transform 1 0 2208 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_24
timestamp 1676037725
transform 1 0 3312 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_46
timestamp 1676037725
transform 1 0 5336 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_59_50
timestamp 1676037725
transform 1 0 5704 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_59_57
timestamp 1676037725
transform 1 0 6348 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_82
timestamp 1676037725
transform 1 0 8648 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_95
timestamp 1676037725
transform 1 0 9844 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_107
timestamp 1676037725
transform 1 0 10948 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1676037725
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_113
timestamp 1676037725
transform 1 0 11500 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_135
timestamp 1676037725
transform 1 0 13524 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_139
timestamp 1676037725
transform 1 0 13892 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_150
timestamp 1676037725
transform 1 0 14904 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_162
timestamp 1676037725
transform 1 0 16008 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_59_169
timestamp 1676037725
transform 1 0 16652 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_191
timestamp 1676037725
transform 1 0 18676 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_204
timestamp 1676037725
transform 1 0 19872 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_211
timestamp 1676037725
transform 1 0 20516 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1676037725
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_225
timestamp 1676037725
transform 1 0 21804 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_236
timestamp 1676037725
transform 1 0 22816 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_243
timestamp 1676037725
transform 1 0 23460 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_255
timestamp 1676037725
transform 1 0 24564 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_59_264
timestamp 1676037725
transform 1 0 25392 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1676037725
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1676037725
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1676037725
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1676037725
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_41
timestamp 1676037725
transform 1 0 4876 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_65
timestamp 1676037725
transform 1 0 7084 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_69
timestamp 1676037725
transform 1 0 7452 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_80
timestamp 1676037725
transform 1 0 8464 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_85
timestamp 1676037725
transform 1 0 8924 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_91
timestamp 1676037725
transform 1 0 9476 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_101
timestamp 1676037725
transform 1 0 10396 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_113
timestamp 1676037725
transform 1 0 11500 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_117
timestamp 1676037725
transform 1 0 11868 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_138
timestamp 1676037725
transform 1 0 13800 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_143
timestamp 1676037725
transform 1 0 14260 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_147
timestamp 1676037725
transform 1 0 14628 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_158
timestamp 1676037725
transform 1 0 15640 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_170
timestamp 1676037725
transform 1 0 16744 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_60_182
timestamp 1676037725
transform 1 0 17848 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_60_194
timestamp 1676037725
transform 1 0 18952 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_60_197
timestamp 1676037725
transform 1 0 19228 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_60_214
timestamp 1676037725
transform 1 0 20792 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_231
timestamp 1676037725
transform 1 0 22356 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_244
timestamp 1676037725
transform 1 0 23552 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_253
timestamp 1676037725
transform 1 0 24380 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_259
timestamp 1676037725
transform 1 0 24932 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_264
timestamp 1676037725
transform 1 0 25392 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1676037725
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1676037725
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_27
timestamp 1676037725
transform 1 0 3588 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_33
timestamp 1676037725
transform 1 0 4140 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_54
timestamp 1676037725
transform 1 0 6072 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_59
timestamp 1676037725
transform 1 0 6532 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_71
timestamp 1676037725
transform 1 0 7636 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_83
timestamp 1676037725
transform 1 0 8740 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_89
timestamp 1676037725
transform 1 0 9292 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_110
timestamp 1676037725
transform 1 0 11224 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_115
timestamp 1676037725
transform 1 0 11684 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_137
timestamp 1676037725
transform 1 0 13708 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_61_141
timestamp 1676037725
transform 1 0 14076 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_144
timestamp 1676037725
transform 1 0 14352 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_149
timestamp 1676037725
transform 1 0 14812 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_162
timestamp 1676037725
transform 1 0 16008 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_61_169
timestamp 1676037725
transform 1 0 16652 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_180
timestamp 1676037725
transform 1 0 17664 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_188
timestamp 1676037725
transform 1 0 18400 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_61_211
timestamp 1676037725
transform 1 0 20516 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_215
timestamp 1676037725
transform 1 0 20884 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1676037725
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_225
timestamp 1676037725
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_237
timestamp 1676037725
transform 1 0 22908 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_243
timestamp 1676037725
transform 1 0 23460 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_264
timestamp 1676037725
transform 1 0 25392 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1676037725
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1676037725
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1676037725
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1676037725
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1676037725
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_53
timestamp 1676037725
transform 1 0 5980 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_74
timestamp 1676037725
transform 1 0 7912 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_78
timestamp 1676037725
transform 1 0 8280 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_85
timestamp 1676037725
transform 1 0 8924 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_98
timestamp 1676037725
transform 1 0 10120 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_105
timestamp 1676037725
transform 1 0 10764 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_109
timestamp 1676037725
transform 1 0 11132 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_121
timestamp 1676037725
transform 1 0 12236 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_125
timestamp 1676037725
transform 1 0 12604 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_137
timestamp 1676037725
transform 1 0 13708 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_62_141
timestamp 1676037725
transform 1 0 14076 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_152
timestamp 1676037725
transform 1 0 15088 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_62_156
timestamp 1676037725
transform 1 0 15456 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_159
timestamp 1676037725
transform 1 0 15732 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_170
timestamp 1676037725
transform 1 0 16744 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_183
timestamp 1676037725
transform 1 0 17940 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1676037725
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_197
timestamp 1676037725
transform 1 0 19228 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_203
timestamp 1676037725
transform 1 0 19780 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_214
timestamp 1676037725
transform 1 0 20792 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_62_218
timestamp 1676037725
transform 1 0 21160 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_62_230
timestamp 1676037725
transform 1 0 22264 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_236
timestamp 1676037725
transform 1 0 22816 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_240
timestamp 1676037725
transform 1 0 23184 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_250
timestamp 1676037725
transform 1 0 24104 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_253
timestamp 1676037725
transform 1 0 24380 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_259
timestamp 1676037725
transform 1 0 24932 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_264
timestamp 1676037725
transform 1 0 25392 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_3
timestamp 1676037725
transform 1 0 1380 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_8
timestamp 1676037725
transform 1 0 1840 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_12
timestamp 1676037725
transform 1 0 2208 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_24
timestamp 1676037725
transform 1 0 3312 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_36
timestamp 1676037725
transform 1 0 4416 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_53
timestamp 1676037725
transform 1 0 5980 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1676037725
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_69
timestamp 1676037725
transform 1 0 7452 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_90
timestamp 1676037725
transform 1 0 9384 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_103
timestamp 1676037725
transform 1 0 10580 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_110
timestamp 1676037725
transform 1 0 11224 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_113
timestamp 1676037725
transform 1 0 11500 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_124
timestamp 1676037725
transform 1 0 12512 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_128
timestamp 1676037725
transform 1 0 12880 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_138
timestamp 1676037725
transform 1 0 13800 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_146
timestamp 1676037725
transform 1 0 14536 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_150
timestamp 1676037725
transform 1 0 14904 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_163
timestamp 1676037725
transform 1 0 16100 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1676037725
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_169
timestamp 1676037725
transform 1 0 16652 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_174
timestamp 1676037725
transform 1 0 17112 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_182
timestamp 1676037725
transform 1 0 17848 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_193
timestamp 1676037725
transform 1 0 18860 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_63_199
timestamp 1676037725
transform 1 0 19412 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_211
timestamp 1676037725
transform 1 0 20516 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1676037725
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_225
timestamp 1676037725
transform 1 0 21804 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_233
timestamp 1676037725
transform 1 0 22540 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_256
timestamp 1676037725
transform 1 0 24656 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_260
timestamp 1676037725
transform 1 0 25024 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_264
timestamp 1676037725
transform 1 0 25392 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_3
timestamp 1676037725
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1676037725
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1676037725
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1676037725
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_41
timestamp 1676037725
transform 1 0 4876 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_68
timestamp 1676037725
transform 1 0 7360 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_64_81
timestamp 1676037725
transform 1 0 8556 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_64_87
timestamp 1676037725
transform 1 0 9108 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_92
timestamp 1676037725
transform 1 0 9568 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_103
timestamp 1676037725
transform 1 0 10580 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_107
timestamp 1676037725
transform 1 0 10948 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_120
timestamp 1676037725
transform 1 0 12144 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_124
timestamp 1676037725
transform 1 0 12512 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_128
timestamp 1676037725
transform 1 0 12880 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_141
timestamp 1676037725
transform 1 0 14076 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_149
timestamp 1676037725
transform 1 0 14812 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_160
timestamp 1676037725
transform 1 0 15824 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_64_164
timestamp 1676037725
transform 1 0 16192 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_176
timestamp 1676037725
transform 1 0 17296 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_180
timestamp 1676037725
transform 1 0 17664 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_183
timestamp 1676037725
transform 1 0 17940 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_194
timestamp 1676037725
transform 1 0 18952 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_197
timestamp 1676037725
transform 1 0 19228 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_210
timestamp 1676037725
transform 1 0 20424 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_218
timestamp 1676037725
transform 1 0 21160 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_241
timestamp 1676037725
transform 1 0 23276 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_245
timestamp 1676037725
transform 1 0 23644 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_250
timestamp 1676037725
transform 1 0 24104 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_64_255
timestamp 1676037725
transform 1 0 24564 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_64_258
timestamp 1676037725
transform 1 0 24840 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_264
timestamp 1676037725
transform 1 0 25392 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_65_3
timestamp 1676037725
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_15
timestamp 1676037725
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_27
timestamp 1676037725
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_39
timestamp 1676037725
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1676037725
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1676037725
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_57
timestamp 1676037725
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_65_69
timestamp 1676037725
transform 1 0 7452 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_94
timestamp 1676037725
transform 1 0 9752 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_107
timestamp 1676037725
transform 1 0 10948 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1676037725
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_65_115
timestamp 1676037725
transform 1 0 11684 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_65_124
timestamp 1676037725
transform 1 0 12512 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_137
timestamp 1676037725
transform 1 0 13708 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_65_144
timestamp 1676037725
transform 1 0 14352 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_65_159
timestamp 1676037725
transform 1 0 15732 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_166
timestamp 1676037725
transform 1 0 16376 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_171
timestamp 1676037725
transform 1 0 16836 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_193
timestamp 1676037725
transform 1 0 18860 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_197
timestamp 1676037725
transform 1 0 19228 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_202
timestamp 1676037725
transform 1 0 19688 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_206
timestamp 1676037725
transform 1 0 20056 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_65_217
timestamp 1676037725
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1676037725
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_225
timestamp 1676037725
transform 1 0 21804 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_236
timestamp 1676037725
transform 1 0 22816 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_260
timestamp 1676037725
transform 1 0 25024 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_66_3
timestamp 1676037725
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_15
timestamp 1676037725
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1676037725
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1676037725
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_66_61
timestamp 1676037725
transform 1 0 6716 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_65
timestamp 1676037725
transform 1 0 7084 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_71
timestamp 1676037725
transform 1 0 7636 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_82
timestamp 1676037725
transform 1 0 8648 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_66_85
timestamp 1676037725
transform 1 0 8924 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_66_100
timestamp 1676037725
transform 1 0 10304 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_113
timestamp 1676037725
transform 1 0 11500 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_117
timestamp 1676037725
transform 1 0 11868 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_127
timestamp 1676037725
transform 1 0 12788 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1676037725
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_143
timestamp 1676037725
transform 1 0 14260 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_154
timestamp 1676037725
transform 1 0 15272 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_167
timestamp 1676037725
transform 1 0 16468 0 1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_66_180
timestamp 1676037725
transform 1 0 17664 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_192
timestamp 1676037725
transform 1 0 18768 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1676037725
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_197
timestamp 1676037725
transform 1 0 19228 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_66_208
timestamp 1676037725
transform 1 0 20240 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_216
timestamp 1676037725
transform 1 0 20976 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_219
timestamp 1676037725
transform 1 0 21252 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_232
timestamp 1676037725
transform 1 0 22448 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_236
timestamp 1676037725
transform 1 0 22816 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_247
timestamp 1676037725
transform 1 0 23828 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1676037725
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_259
timestamp 1676037725
transform 1 0 24932 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_264
timestamp 1676037725
transform 1 0 25392 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_3
timestamp 1676037725
transform 1 0 1380 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_8
timestamp 1676037725
transform 1 0 1840 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_67_12
timestamp 1676037725
transform 1 0 2208 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_24
timestamp 1676037725
transform 1 0 3312 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_32
timestamp 1676037725
transform 1 0 4048 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_54
timestamp 1676037725
transform 1 0 6072 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_67_59
timestamp 1676037725
transform 1 0 6532 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_71
timestamp 1676037725
transform 1 0 7636 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_79
timestamp 1676037725
transform 1 0 8372 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_67_84
timestamp 1676037725
transform 1 0 8832 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_92
timestamp 1676037725
transform 1 0 9568 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_103
timestamp 1676037725
transform 1 0 10580 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_110
timestamp 1676037725
transform 1 0 11224 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_67_113
timestamp 1676037725
transform 1 0 11500 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_67_125
timestamp 1676037725
transform 1 0 12604 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_129
timestamp 1676037725
transform 1 0 12972 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_135
timestamp 1676037725
transform 1 0 13524 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_67_146
timestamp 1676037725
transform 1 0 14536 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_67_154
timestamp 1676037725
transform 1 0 15272 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_67_165
timestamp 1676037725
transform 1 0 16284 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_67_169
timestamp 1676037725
transform 1 0 16652 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_177
timestamp 1676037725
transform 1 0 17388 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_67_200
timestamp 1676037725
transform 1 0 19504 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_213
timestamp 1676037725
transform 1 0 20700 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_67_219
timestamp 1676037725
transform 1 0 21252 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_67_225
timestamp 1676037725
transform 1 0 21804 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_236
timestamp 1676037725
transform 1 0 22816 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_240
timestamp 1676037725
transform 1 0 23184 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_67_263
timestamp 1676037725
transform 1 0 25300 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1676037725
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1676037725
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1676037725
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1676037725
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_41
timestamp 1676037725
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_53
timestamp 1676037725
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_65
timestamp 1676037725
transform 1 0 7084 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_68_80
timestamp 1676037725
transform 1 0 8464 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_85
timestamp 1676037725
transform 1 0 8924 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_96
timestamp 1676037725
transform 1 0 9936 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_121
timestamp 1676037725
transform 1 0 12236 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_68_134
timestamp 1676037725
transform 1 0 13432 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_68_141
timestamp 1676037725
transform 1 0 14076 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_68_152
timestamp 1676037725
transform 1 0 15088 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_158
timestamp 1676037725
transform 1 0 15640 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_168
timestamp 1676037725
transform 1 0 16560 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_176
timestamp 1676037725
transform 1 0 17296 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_186
timestamp 1676037725
transform 1 0 18216 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_194
timestamp 1676037725
transform 1 0 18952 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_68_197
timestamp 1676037725
transform 1 0 19228 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_68_209
timestamp 1676037725
transform 1 0 20332 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_222
timestamp 1676037725
transform 1 0 21528 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_235
timestamp 1676037725
transform 1 0 22724 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_239
timestamp 1676037725
transform 1 0 23092 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_245
timestamp 1676037725
transform 1 0 23644 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_250
timestamp 1676037725
transform 1 0 24104 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_253
timestamp 1676037725
transform 1 0 24380 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_264
timestamp 1676037725
transform 1 0 25392 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_69_3
timestamp 1676037725
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_15
timestamp 1676037725
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_27
timestamp 1676037725
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_39
timestamp 1676037725
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1676037725
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1676037725
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_57
timestamp 1676037725
transform 1 0 6348 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_69_65
timestamp 1676037725
transform 1 0 7084 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_69_70
timestamp 1676037725
transform 1 0 7544 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_81
timestamp 1676037725
transform 1 0 8556 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_69_96
timestamp 1676037725
transform 1 0 9936 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_69_100
timestamp 1676037725
transform 1 0 10304 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_113
timestamp 1676037725
transform 1 0 11500 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_119
timestamp 1676037725
transform 1 0 12052 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_140
timestamp 1676037725
transform 1 0 13984 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_69_147
timestamp 1676037725
transform 1 0 14628 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_151
timestamp 1676037725
transform 1 0 14996 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_69_162
timestamp 1676037725
transform 1 0 16008 0 -1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_69_169
timestamp 1676037725
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_181
timestamp 1676037725
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_193
timestamp 1676037725
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_69_205
timestamp 1676037725
transform 1 0 19964 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_211
timestamp 1676037725
transform 1 0 20516 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_222
timestamp 1676037725
transform 1 0 21528 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_225
timestamp 1676037725
transform 1 0 21804 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_236
timestamp 1676037725
transform 1 0 22816 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_250
timestamp 1676037725
transform 1 0 24104 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_69_264
timestamp 1676037725
transform 1 0 25392 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_70_3
timestamp 1676037725
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_70_15
timestamp 1676037725
transform 1 0 2484 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_21
timestamp 1676037725
transform 1 0 3036 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_70_25
timestamp 1676037725
transform 1 0 3404 0 1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1676037725
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1676037725
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_53
timestamp 1676037725
transform 1 0 5980 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_70_77
timestamp 1676037725
transform 1 0 8188 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_70_81
timestamp 1676037725
transform 1 0 8556 0 1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_70_85
timestamp 1676037725
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_97
timestamp 1676037725
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_70_109
timestamp 1676037725
transform 1 0 11132 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_122
timestamp 1676037725
transform 1 0 12328 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_126
timestamp 1676037725
transform 1 0 12696 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_70_137
timestamp 1676037725
transform 1 0 13708 0 1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_70_145
timestamp 1676037725
transform 1 0 14444 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_70_157
timestamp 1676037725
transform 1 0 15548 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_70_169
timestamp 1676037725
transform 1 0 16652 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_70_175
timestamp 1676037725
transform 1 0 17204 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_70_186
timestamp 1676037725
transform 1 0 18216 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_70_194
timestamp 1676037725
transform 1 0 18952 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_197
timestamp 1676037725
transform 1 0 19228 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_208
timestamp 1676037725
transform 1 0 20240 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_212
timestamp 1676037725
transform 1 0 20608 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_216
timestamp 1676037725
transform 1 0 20976 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_70_238
timestamp 1676037725
transform 1 0 23000 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_70_245
timestamp 1676037725
transform 1 0 23644 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_70_249
timestamp 1676037725
transform 1 0 24012 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_70_255
timestamp 1676037725
transform 1 0 24564 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_259
timestamp 1676037725
transform 1 0 24932 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_264
timestamp 1676037725
transform 1 0 25392 0 1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_71_3
timestamp 1676037725
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_15
timestamp 1676037725
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_71_27
timestamp 1676037725
transform 1 0 3588 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_71_34
timestamp 1676037725
transform 1 0 4232 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_71_38
timestamp 1676037725
transform 1 0 4600 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_50
timestamp 1676037725
transform 1 0 5704 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_71_57
timestamp 1676037725
transform 1 0 6348 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_79
timestamp 1676037725
transform 1 0 8372 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_71_83
timestamp 1676037725
transform 1 0 8740 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_89
timestamp 1676037725
transform 1 0 9292 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_71_110
timestamp 1676037725
transform 1 0 11224 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_113
timestamp 1676037725
transform 1 0 11500 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_124
timestamp 1676037725
transform 1 0 12512 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_128
timestamp 1676037725
transform 1 0 12880 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_132
timestamp 1676037725
transform 1 0 13248 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_71_153
timestamp 1676037725
transform 1 0 15180 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_71_157
timestamp 1676037725
transform 1 0 15548 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_71_165
timestamp 1676037725
transform 1 0 16284 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_71_169
timestamp 1676037725
transform 1 0 16652 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_180
timestamp 1676037725
transform 1 0 17664 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_184
timestamp 1676037725
transform 1 0 18032 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_208
timestamp 1676037725
transform 1 0 20240 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_71_212
timestamp 1676037725
transform 1 0 20608 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_218
timestamp 1676037725
transform 1 0 21160 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_71_222
timestamp 1676037725
transform 1 0 21528 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_225
timestamp 1676037725
transform 1 0 21804 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_236
timestamp 1676037725
transform 1 0 22816 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_260
timestamp 1676037725
transform 1 0 25024 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_72_3
timestamp 1676037725
transform 1 0 1380 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_72_9
timestamp 1676037725
transform 1 0 1932 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_13
timestamp 1676037725
transform 1 0 2300 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_72_25
timestamp 1676037725
transform 1 0 3404 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_72_29
timestamp 1676037725
transform 1 0 3772 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_72_39
timestamp 1676037725
transform 1 0 4692 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_72_43
timestamp 1676037725
transform 1 0 5060 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_72_49
timestamp 1676037725
transform 1 0 5612 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_53
timestamp 1676037725
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_65
timestamp 1676037725
transform 1 0 7084 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_72_82
timestamp 1676037725
transform 1 0 8648 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_85
timestamp 1676037725
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_97
timestamp 1676037725
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_109
timestamp 1676037725
transform 1 0 11132 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_72_130
timestamp 1676037725
transform 1 0 13064 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_72_134
timestamp 1676037725
transform 1 0 13432 0 1 41344
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_72_141
timestamp 1676037725
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_72_173
timestamp 1676037725
transform 1 0 17020 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_72_177
timestamp 1676037725
transform 1 0 17388 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_72_181
timestamp 1676037725
transform 1 0 17756 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_72_194
timestamp 1676037725
transform 1 0 18952 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_72_197
timestamp 1676037725
transform 1 0 19228 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_208
timestamp 1676037725
transform 1 0 20240 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_212
timestamp 1676037725
transform 1 0 20608 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_222
timestamp 1676037725
transform 1 0 21528 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_226
timestamp 1676037725
transform 1 0 21896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_236
timestamp 1676037725
transform 1 0 22816 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_72_250
timestamp 1676037725
transform 1 0 24104 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_72_253
timestamp 1676037725
transform 1 0 24380 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_72_264
timestamp 1676037725
transform 1 0 25392 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_3
timestamp 1676037725
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_15
timestamp 1676037725
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_27
timestamp 1676037725
transform 1 0 3588 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_32
timestamp 1676037725
transform 1 0 4048 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_36
timestamp 1676037725
transform 1 0 4416 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_48
timestamp 1676037725
transform 1 0 5520 0 -1 42432
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_73_57
timestamp 1676037725
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_69
timestamp 1676037725
transform 1 0 7452 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_93
timestamp 1676037725
transform 1 0 9660 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_97
timestamp 1676037725
transform 1 0 10028 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_73_109
timestamp 1676037725
transform 1 0 11132 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_73_113
timestamp 1676037725
transform 1 0 11500 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_73_125
timestamp 1676037725
transform 1 0 12604 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_73_133
timestamp 1676037725
transform 1 0 13340 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_73_156
timestamp 1676037725
transform 1 0 15456 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_73_160
timestamp 1676037725
transform 1 0 15824 0 -1 42432
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_73_169
timestamp 1676037725
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_181
timestamp 1676037725
transform 1 0 17756 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_202
timestamp 1676037725
transform 1 0 19688 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_73_206
timestamp 1676037725
transform 1 0 20056 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_209
timestamp 1676037725
transform 1 0 20332 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_222
timestamp 1676037725
transform 1 0 21528 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_225
timestamp 1676037725
transform 1 0 21804 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_236
timestamp 1676037725
transform 1 0 22816 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_240
timestamp 1676037725
transform 1 0 23184 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_261
timestamp 1676037725
transform 1 0 25116 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_73_265
timestamp 1676037725
transform 1 0 25484 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_3
timestamp 1676037725
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_15
timestamp 1676037725
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1676037725
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_29
timestamp 1676037725
transform 1 0 3772 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_74_37
timestamp 1676037725
transform 1 0 4508 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_74_41
timestamp 1676037725
transform 1 0 4876 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_74_49
timestamp 1676037725
transform 1 0 5612 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_74_54
timestamp 1676037725
transform 1 0 6072 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_60
timestamp 1676037725
transform 1 0 6624 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_67
timestamp 1676037725
transform 1 0 7268 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_74
timestamp 1676037725
transform 1 0 7912 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_74_82
timestamp 1676037725
transform 1 0 8648 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_74_85
timestamp 1676037725
transform 1 0 8924 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_74_88
timestamp 1676037725
transform 1 0 9200 0 1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_74_99
timestamp 1676037725
transform 1 0 10212 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_111
timestamp 1676037725
transform 1 0 11316 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_117
timestamp 1676037725
transform 1 0 11868 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_127
timestamp 1676037725
transform 1 0 12788 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1676037725
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_74_141
timestamp 1676037725
transform 1 0 14076 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_74_163
timestamp 1676037725
transform 1 0 16100 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_74_167
timestamp 1676037725
transform 1 0 16468 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_74_175
timestamp 1676037725
transform 1 0 17204 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_74_187
timestamp 1676037725
transform 1 0 18308 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_191
timestamp 1676037725
transform 1 0 18676 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1676037725
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_74_197
timestamp 1676037725
transform 1 0 19228 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_74_219
timestamp 1676037725
transform 1 0 21252 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_74_226
timestamp 1676037725
transform 1 0 21896 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_74_250
timestamp 1676037725
transform 1 0 24104 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_74_253
timestamp 1676037725
transform 1 0 24380 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_74_258
timestamp 1676037725
transform 1 0 24840 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_74_262
timestamp 1676037725
transform 1 0 25208 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_75_3
timestamp 1676037725
transform 1 0 1380 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_9
timestamp 1676037725
transform 1 0 1932 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_75_13
timestamp 1676037725
transform 1 0 2300 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_17
timestamp 1676037725
transform 1 0 2668 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_29
timestamp 1676037725
transform 1 0 3772 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_41
timestamp 1676037725
transform 1 0 4876 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_47
timestamp 1676037725
transform 1 0 5428 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_51
timestamp 1676037725
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1676037725
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1676037725
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_69
timestamp 1676037725
transform 1 0 7452 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_75
timestamp 1676037725
transform 1 0 8004 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_75_78
timestamp 1676037725
transform 1 0 8280 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_75_102
timestamp 1676037725
transform 1 0 10488 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_75_106
timestamp 1676037725
transform 1 0 10856 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_75_113
timestamp 1676037725
transform 1 0 11500 0 -1 43520
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_75_130
timestamp 1676037725
transform 1 0 13064 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_142
timestamp 1676037725
transform 1 0 14168 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_154
timestamp 1676037725
transform 1 0 15272 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_75_166
timestamp 1676037725
transform 1 0 16376 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_75_169
timestamp 1676037725
transform 1 0 16652 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_75_180
timestamp 1676037725
transform 1 0 17664 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_184
timestamp 1676037725
transform 1 0 18032 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_196
timestamp 1676037725
transform 1 0 19136 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_208
timestamp 1676037725
transform 1 0 20240 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_220
timestamp 1676037725
transform 1 0 21344 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_75_225
timestamp 1676037725
transform 1 0 21804 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_75_247
timestamp 1676037725
transform 1 0 23828 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_75_254
timestamp 1676037725
transform 1 0 24472 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_260
timestamp 1676037725
transform 1 0 25024 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_75_264
timestamp 1676037725
transform 1 0 25392 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_3
timestamp 1676037725
transform 1 0 1380 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_8
timestamp 1676037725
transform 1 0 1840 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_12
timestamp 1676037725
transform 1 0 2208 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_24
timestamp 1676037725
transform 1 0 3312 0 1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_76_29
timestamp 1676037725
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_41
timestamp 1676037725
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_53
timestamp 1676037725
transform 1 0 5980 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_76_61
timestamp 1676037725
transform 1 0 6716 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_65
timestamp 1676037725
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_77
timestamp 1676037725
transform 1 0 8188 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_76_82
timestamp 1676037725
transform 1 0 8648 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_87
timestamp 1676037725
transform 1 0 9108 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_91
timestamp 1676037725
transform 1 0 9476 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_97
timestamp 1676037725
transform 1 0 10028 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_76_105
timestamp 1676037725
transform 1 0 10764 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_76_109
timestamp 1676037725
transform 1 0 11132 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_112
timestamp 1676037725
transform 1 0 11408 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_76_137
timestamp 1676037725
transform 1 0 13708 0 1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_76_143
timestamp 1676037725
transform 1 0 14260 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_155
timestamp 1676037725
transform 1 0 15364 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_159
timestamp 1676037725
transform 1 0 15732 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_76_180
timestamp 1676037725
transform 1 0 17664 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_184
timestamp 1676037725
transform 1 0 18032 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_76_197
timestamp 1676037725
transform 1 0 19228 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_219
timestamp 1676037725
transform 1 0 21252 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_223
timestamp 1676037725
transform 1 0 21620 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_76_247
timestamp 1676037725
transform 1 0 23828 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1676037725
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_76_253
timestamp 1676037725
transform 1 0 24380 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_258
timestamp 1676037725
transform 1 0 24840 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_262
timestamp 1676037725
transform 1 0 25208 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_77_3
timestamp 1676037725
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_15
timestamp 1676037725
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_27
timestamp 1676037725
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_39
timestamp 1676037725
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1676037725
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1676037725
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_57
timestamp 1676037725
transform 1 0 6348 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_77_63
timestamp 1676037725
transform 1 0 6900 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_69
timestamp 1676037725
transform 1 0 7452 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_76
timestamp 1676037725
transform 1 0 8096 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_77_84
timestamp 1676037725
transform 1 0 8832 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_88
timestamp 1676037725
transform 1 0 9200 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_110
timestamp 1676037725
transform 1 0 11224 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_113
timestamp 1676037725
transform 1 0 11500 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_124
timestamp 1676037725
transform 1 0 12512 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_77_132
timestamp 1676037725
transform 1 0 13248 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_77_136
timestamp 1676037725
transform 1 0 13616 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_77_151
timestamp 1676037725
transform 1 0 14996 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_77_155
timestamp 1676037725
transform 1 0 15364 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1676037725
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_77_169
timestamp 1676037725
transform 1 0 16652 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_77_177
timestamp 1676037725
transform 1 0 17388 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_77_200
timestamp 1676037725
transform 1 0 19504 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_77_204
timestamp 1676037725
transform 1 0 19872 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_77_216
timestamp 1676037725
transform 1 0 20976 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1676037725
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_77_225
timestamp 1676037725
transform 1 0 21804 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_247
timestamp 1676037725
transform 1 0 23828 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_77_251
timestamp 1676037725
transform 1 0 24196 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_77_264
timestamp 1676037725
transform 1 0 25392 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_78_3
timestamp 1676037725
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_15
timestamp 1676037725
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1676037725
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_29
timestamp 1676037725
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_41
timestamp 1676037725
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_53
timestamp 1676037725
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_78_65
timestamp 1676037725
transform 1 0 7084 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_78_72
timestamp 1676037725
transform 1 0 7728 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_78_76
timestamp 1676037725
transform 1 0 8096 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_80
timestamp 1676037725
transform 1 0 8464 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_78_85
timestamp 1676037725
transform 1 0 8924 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_91
timestamp 1676037725
transform 1 0 9476 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_78_94
timestamp 1676037725
transform 1 0 9752 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_100
timestamp 1676037725
transform 1 0 10304 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_78_124
timestamp 1676037725
transform 1 0 12512 0 1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_78_128
timestamp 1676037725
transform 1 0 12880 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_78_141
timestamp 1676037725
transform 1 0 14076 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_78_163
timestamp 1676037725
transform 1 0 16100 0 1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_78_167
timestamp 1676037725
transform 1 0 16468 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_179
timestamp 1676037725
transform 1 0 17572 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_191
timestamp 1676037725
transform 1 0 18676 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1676037725
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_78_197
timestamp 1676037725
transform 1 0 19228 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_219
timestamp 1676037725
transform 1 0 21252 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_232
timestamp 1676037725
transform 1 0 22448 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_78_245
timestamp 1676037725
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1676037725
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_253
timestamp 1676037725
transform 1 0 24380 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_78_259
timestamp 1676037725
transform 1 0 24932 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_78_264
timestamp 1676037725
transform 1 0 25392 0 1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_79_5
timestamp 1676037725
transform 1 0 1564 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_17
timestamp 1676037725
transform 1 0 2668 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_29
timestamp 1676037725
transform 1 0 3772 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_41
timestamp 1676037725
transform 1 0 4876 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_53
timestamp 1676037725
transform 1 0 5980 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_79_57
timestamp 1676037725
transform 1 0 6348 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_79_65
timestamp 1676037725
transform 1 0 7084 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_79_68
timestamp 1676037725
transform 1 0 7360 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_79_74
timestamp 1676037725
transform 1 0 7912 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_78
timestamp 1676037725
transform 1 0 8280 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_82
timestamp 1676037725
transform 1 0 8648 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_97
timestamp 1676037725
transform 1 0 10028 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_79_105
timestamp 1676037725
transform 1 0 10764 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_79_110
timestamp 1676037725
transform 1 0 11224 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_79_113
timestamp 1676037725
transform 1 0 11500 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_79_119
timestamp 1676037725
transform 1 0 12052 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_79_123
timestamp 1676037725
transform 1 0 12420 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_79_131
timestamp 1676037725
transform 1 0 13156 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_79_153
timestamp 1676037725
transform 1 0 15180 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_79_157
timestamp 1676037725
transform 1 0 15548 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_79_165
timestamp 1676037725
transform 1 0 16284 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_79_169
timestamp 1676037725
transform 1 0 16652 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_79_191
timestamp 1676037725
transform 1 0 18676 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_79_195
timestamp 1676037725
transform 1 0 19044 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_79_200
timestamp 1676037725
transform 1 0 19504 0 -1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_79_211
timestamp 1676037725
transform 1 0 20516 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1676037725
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_225
timestamp 1676037725
transform 1 0 21804 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_79_233
timestamp 1676037725
transform 1 0 22540 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_236
timestamp 1676037725
transform 1 0 22816 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_79_264
timestamp 1676037725
transform 1 0 25392 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_3
timestamp 1676037725
transform 1 0 1380 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_80_15
timestamp 1676037725
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1676037725
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_29
timestamp 1676037725
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_41
timestamp 1676037725
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_53
timestamp 1676037725
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_65
timestamp 1676037725
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_77
timestamp 1676037725
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1676037725
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_85
timestamp 1676037725
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_97
timestamp 1676037725
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_109
timestamp 1676037725
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_121
timestamp 1676037725
transform 1 0 12236 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_133
timestamp 1676037725
transform 1 0 13340 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_139
timestamp 1676037725
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_141
timestamp 1676037725
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_153
timestamp 1676037725
transform 1 0 15180 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_159
timestamp 1676037725
transform 1 0 15732 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_80_180
timestamp 1676037725
transform 1 0 17664 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_80_186
timestamp 1676037725
transform 1 0 18216 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_80_194
timestamp 1676037725
transform 1 0 18952 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_197
timestamp 1676037725
transform 1 0 19228 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_208
timestamp 1676037725
transform 1 0 20240 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_212
timestamp 1676037725
transform 1 0 20608 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_222
timestamp 1676037725
transform 1 0 21528 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_234
timestamp 1676037725
transform 1 0 22632 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_246
timestamp 1676037725
transform 1 0 23736 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_80_250
timestamp 1676037725
transform 1 0 24104 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_253
timestamp 1676037725
transform 1 0 24380 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_258
timestamp 1676037725
transform 1 0 24840 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_262
timestamp 1676037725
transform 1 0 25208 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_81_3
timestamp 1676037725
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_15
timestamp 1676037725
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_27
timestamp 1676037725
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_39
timestamp 1676037725
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_51
timestamp 1676037725
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1676037725
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_57
timestamp 1676037725
transform 1 0 6348 0 -1 46784
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_81_68
timestamp 1676037725
transform 1 0 7360 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_80
timestamp 1676037725
transform 1 0 8464 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_92
timestamp 1676037725
transform 1 0 9568 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_104
timestamp 1676037725
transform 1 0 10672 0 -1 46784
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_81_113
timestamp 1676037725
transform 1 0 11500 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_125
timestamp 1676037725
transform 1 0 12604 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_81_157
timestamp 1676037725
transform 1 0 15548 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_81_161
timestamp 1676037725
transform 1 0 15916 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_167
timestamp 1676037725
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_81_169
timestamp 1676037725
transform 1 0 16652 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_180
timestamp 1676037725
transform 1 0 17664 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_193
timestamp 1676037725
transform 1 0 18860 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_81_197
timestamp 1676037725
transform 1 0 19228 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_81_205
timestamp 1676037725
transform 1 0 19964 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_81_210
timestamp 1676037725
transform 1 0 20424 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_213
timestamp 1676037725
transform 1 0 20700 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_81_221
timestamp 1676037725
transform 1 0 21436 0 -1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_81_225
timestamp 1676037725
transform 1 0 21804 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_237
timestamp 1676037725
transform 1 0 22908 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_244
timestamp 1676037725
transform 1 0 23552 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_248
timestamp 1676037725
transform 1 0 23920 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_252
timestamp 1676037725
transform 1 0 24288 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_264
timestamp 1676037725
transform 1 0 25392 0 -1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_3
timestamp 1676037725
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_15
timestamp 1676037725
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1676037725
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_29
timestamp 1676037725
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_41
timestamp 1676037725
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_53
timestamp 1676037725
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_65
timestamp 1676037725
transform 1 0 7084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_77
timestamp 1676037725
transform 1 0 8188 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1676037725
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_85
timestamp 1676037725
transform 1 0 8924 0 1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_90
timestamp 1676037725
transform 1 0 9384 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_102
timestamp 1676037725
transform 1 0 10488 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_110
timestamp 1676037725
transform 1 0 11224 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_82_116
timestamp 1676037725
transform 1 0 11776 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_128
timestamp 1676037725
transform 1 0 12880 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_141
timestamp 1676037725
transform 1 0 14076 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_149
timestamp 1676037725
transform 1 0 14812 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_172
timestamp 1676037725
transform 1 0 16928 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_185
timestamp 1676037725
transform 1 0 18124 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_82_189
timestamp 1676037725
transform 1 0 18492 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_195
timestamp 1676037725
transform 1 0 19044 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_197
timestamp 1676037725
transform 1 0 19228 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_209
timestamp 1676037725
transform 1 0 20332 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_221
timestamp 1676037725
transform 1 0 21436 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_233
timestamp 1676037725
transform 1 0 22540 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_241
timestamp 1676037725
transform 1 0 23276 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_245
timestamp 1676037725
transform 1 0 23644 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_250
timestamp 1676037725
transform 1 0 24104 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_253
timestamp 1676037725
transform 1 0 24380 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_259
timestamp 1676037725
transform 1 0 24932 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_82_263
timestamp 1676037725
transform 1 0 25300 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_83_3
timestamp 1676037725
transform 1 0 1380 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_15
timestamp 1676037725
transform 1 0 2484 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_27
timestamp 1676037725
transform 1 0 3588 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_39
timestamp 1676037725
transform 1 0 4692 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_51
timestamp 1676037725
transform 1 0 5796 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_55
timestamp 1676037725
transform 1 0 6164 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_57
timestamp 1676037725
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_69
timestamp 1676037725
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_81
timestamp 1676037725
transform 1 0 8556 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_93
timestamp 1676037725
transform 1 0 9660 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_105
timestamp 1676037725
transform 1 0 10764 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_111
timestamp 1676037725
transform 1 0 11316 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_113
timestamp 1676037725
transform 1 0 11500 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_125
timestamp 1676037725
transform 1 0 12604 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_137
timestamp 1676037725
transform 1 0 13708 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_149
timestamp 1676037725
transform 1 0 14812 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_161
timestamp 1676037725
transform 1 0 15916 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_167
timestamp 1676037725
transform 1 0 16468 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_83_169
timestamp 1676037725
transform 1 0 16652 0 -1 47872
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_83_174
timestamp 1676037725
transform 1 0 17112 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_186
timestamp 1676037725
transform 1 0 18216 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_198
timestamp 1676037725
transform 1 0 19320 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_210
timestamp 1676037725
transform 1 0 20424 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_83_222
timestamp 1676037725
transform 1 0 21528 0 -1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_83_225
timestamp 1676037725
transform 1 0 21804 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_237
timestamp 1676037725
transform 1 0 22908 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_244
timestamp 1676037725
transform 1 0 23552 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_251
timestamp 1676037725
transform 1 0 24196 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_83_259
timestamp 1676037725
transform 1 0 24932 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_83_263
timestamp 1676037725
transform 1 0 25300 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_84_3
timestamp 1676037725
transform 1 0 1380 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_84_9
timestamp 1676037725
transform 1 0 1932 0 1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_84_13
timestamp 1676037725
transform 1 0 2300 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_84_25
timestamp 1676037725
transform 1 0 3404 0 1 47872
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_84_29
timestamp 1676037725
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_41
timestamp 1676037725
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_53
timestamp 1676037725
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_65
timestamp 1676037725
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_77
timestamp 1676037725
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_83
timestamp 1676037725
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_85
timestamp 1676037725
transform 1 0 8924 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_97
timestamp 1676037725
transform 1 0 10028 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_109
timestamp 1676037725
transform 1 0 11132 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_121
timestamp 1676037725
transform 1 0 12236 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_133
timestamp 1676037725
transform 1 0 13340 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_139
timestamp 1676037725
transform 1 0 13892 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_141
timestamp 1676037725
transform 1 0 14076 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_153
timestamp 1676037725
transform 1 0 15180 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_165
timestamp 1676037725
transform 1 0 16284 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_177
timestamp 1676037725
transform 1 0 17388 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_189
timestamp 1676037725
transform 1 0 18492 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_195
timestamp 1676037725
transform 1 0 19044 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_197
timestamp 1676037725
transform 1 0 19228 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_209
timestamp 1676037725
transform 1 0 20332 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_221
timestamp 1676037725
transform 1 0 21436 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_233
timestamp 1676037725
transform 1 0 22540 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_84_241
timestamp 1676037725
transform 1 0 23276 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_84_246
timestamp 1676037725
transform 1 0 23736 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_84_255
timestamp 1676037725
transform 1 0 24564 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_84_259
timestamp 1676037725
transform 1 0 24932 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_84_264
timestamp 1676037725
transform 1 0 25392 0 1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_85_3
timestamp 1676037725
transform 1 0 1380 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_15
timestamp 1676037725
transform 1 0 2484 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_27
timestamp 1676037725
transform 1 0 3588 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_39
timestamp 1676037725
transform 1 0 4692 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_51
timestamp 1676037725
transform 1 0 5796 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_55
timestamp 1676037725
transform 1 0 6164 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_57
timestamp 1676037725
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_69
timestamp 1676037725
transform 1 0 7452 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_81
timestamp 1676037725
transform 1 0 8556 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_93
timestamp 1676037725
transform 1 0 9660 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_105
timestamp 1676037725
transform 1 0 10764 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_111
timestamp 1676037725
transform 1 0 11316 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_85_113
timestamp 1676037725
transform 1 0 11500 0 -1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_85_118
timestamp 1676037725
transform 1 0 11960 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_130
timestamp 1676037725
transform 1 0 13064 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_142
timestamp 1676037725
transform 1 0 14168 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_154
timestamp 1676037725
transform 1 0 15272 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_85_166
timestamp 1676037725
transform 1 0 16376 0 -1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_85_169
timestamp 1676037725
transform 1 0 16652 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_181
timestamp 1676037725
transform 1 0 17756 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_193
timestamp 1676037725
transform 1 0 18860 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_205
timestamp 1676037725
transform 1 0 19964 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_217
timestamp 1676037725
transform 1 0 21068 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_223
timestamp 1676037725
transform 1 0 21620 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_225
timestamp 1676037725
transform 1 0 21804 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_237
timestamp 1676037725
transform 1 0 22908 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_249
timestamp 1676037725
transform 1 0 24012 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_255
timestamp 1676037725
transform 1 0 24564 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_85_258
timestamp 1676037725
transform 1 0 24840 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_85_264
timestamp 1676037725
transform 1 0 25392 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_86_3
timestamp 1676037725
transform 1 0 1380 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_86_21
timestamp 1676037725
transform 1 0 3036 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_27
timestamp 1676037725
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_86_29
timestamp 1676037725
transform 1 0 3772 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_35
timestamp 1676037725
transform 1 0 4324 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_86_59
timestamp 1676037725
transform 1 0 6532 0 1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_86_63
timestamp 1676037725
transform 1 0 6900 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_75
timestamp 1676037725
transform 1 0 8004 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_86_83
timestamp 1676037725
transform 1 0 8740 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_85
timestamp 1676037725
transform 1 0 8924 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_97
timestamp 1676037725
transform 1 0 10028 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_109
timestamp 1676037725
transform 1 0 11132 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_121
timestamp 1676037725
transform 1 0 12236 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_133
timestamp 1676037725
transform 1 0 13340 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_139
timestamp 1676037725
transform 1 0 13892 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_141
timestamp 1676037725
transform 1 0 14076 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_153
timestamp 1676037725
transform 1 0 15180 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_165
timestamp 1676037725
transform 1 0 16284 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_177
timestamp 1676037725
transform 1 0 17388 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_189
timestamp 1676037725
transform 1 0 18492 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_195
timestamp 1676037725
transform 1 0 19044 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_197
timestamp 1676037725
transform 1 0 19228 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_209
timestamp 1676037725
transform 1 0 20332 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_221
timestamp 1676037725
transform 1 0 21436 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_233
timestamp 1676037725
transform 1 0 22540 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_245
timestamp 1676037725
transform 1 0 23644 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_251
timestamp 1676037725
transform 1 0 24196 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_86_253
timestamp 1676037725
transform 1 0 24380 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_86_258
timestamp 1676037725
transform 1 0 24840 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_86_264
timestamp 1676037725
transform 1 0 25392 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_87_3
timestamp 1676037725
transform 1 0 1380 0 -1 50048
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_87_23
timestamp 1676037725
transform 1 0 3220 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_35
timestamp 1676037725
transform 1 0 4324 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_87_47
timestamp 1676037725
transform 1 0 5428 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_87_55
timestamp 1676037725
transform 1 0 6164 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_87_57
timestamp 1676037725
transform 1 0 6348 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_87_62
timestamp 1676037725
transform 1 0 6808 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_87_70
timestamp 1676037725
transform 1 0 7544 0 -1 50048
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_87_76
timestamp 1676037725
transform 1 0 8096 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_87_88
timestamp 1676037725
transform 1 0 9200 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_93
timestamp 1676037725
transform 1 0 9660 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_105
timestamp 1676037725
transform 1 0 10764 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_111
timestamp 1676037725
transform 1 0 11316 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_113
timestamp 1676037725
transform 1 0 11500 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_125
timestamp 1676037725
transform 1 0 12604 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_137
timestamp 1676037725
transform 1 0 13708 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_149
timestamp 1676037725
transform 1 0 14812 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_161
timestamp 1676037725
transform 1 0 15916 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_167
timestamp 1676037725
transform 1 0 16468 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_169
timestamp 1676037725
transform 1 0 16652 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_181
timestamp 1676037725
transform 1 0 17756 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_193
timestamp 1676037725
transform 1 0 18860 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_205
timestamp 1676037725
transform 1 0 19964 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_217
timestamp 1676037725
transform 1 0 21068 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_223
timestamp 1676037725
transform 1 0 21620 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_225
timestamp 1676037725
transform 1 0 21804 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_237
timestamp 1676037725
transform 1 0 22908 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_249
timestamp 1676037725
transform 1 0 24012 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_255
timestamp 1676037725
transform 1 0 24564 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_87_258
timestamp 1676037725
transform 1 0 24840 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_87_264
timestamp 1676037725
transform 1 0 25392 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_88_5
timestamp 1676037725
transform 1 0 1564 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_9
timestamp 1676037725
transform 1 0 1932 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_88_26
timestamp 1676037725
transform 1 0 3496 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_88_29
timestamp 1676037725
transform 1 0 3772 0 1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_88_47
timestamp 1676037725
transform 1 0 5428 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_59
timestamp 1676037725
transform 1 0 6532 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_71
timestamp 1676037725
transform 1 0 7636 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_83
timestamp 1676037725
transform 1 0 8740 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_88_85
timestamp 1676037725
transform 1 0 8924 0 1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_88_91
timestamp 1676037725
transform 1 0 9476 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_103
timestamp 1676037725
transform 1 0 10580 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_115
timestamp 1676037725
transform 1 0 11684 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_127
timestamp 1676037725
transform 1 0 12788 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_139
timestamp 1676037725
transform 1 0 13892 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_141
timestamp 1676037725
transform 1 0 14076 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_153
timestamp 1676037725
transform 1 0 15180 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_165
timestamp 1676037725
transform 1 0 16284 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_177
timestamp 1676037725
transform 1 0 17388 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_189
timestamp 1676037725
transform 1 0 18492 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_195
timestamp 1676037725
transform 1 0 19044 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_197
timestamp 1676037725
transform 1 0 19228 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_209
timestamp 1676037725
transform 1 0 20332 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_221
timestamp 1676037725
transform 1 0 21436 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_233
timestamp 1676037725
transform 1 0 22540 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_245
timestamp 1676037725
transform 1 0 23644 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_251
timestamp 1676037725
transform 1 0 24196 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_88_253
timestamp 1676037725
transform 1 0 24380 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_88_258
timestamp 1676037725
transform 1 0 24840 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_88_264
timestamp 1676037725
transform 1 0 25392 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_89_3
timestamp 1676037725
transform 1 0 1380 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_89_15
timestamp 1676037725
transform 1 0 2484 0 -1 51136
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_89_35
timestamp 1676037725
transform 1 0 4324 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_89_47
timestamp 1676037725
transform 1 0 5428 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_89_55
timestamp 1676037725
transform 1 0 6164 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_89_57
timestamp 1676037725
transform 1 0 6348 0 -1 51136
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_89_65
timestamp 1676037725
transform 1 0 7084 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_77
timestamp 1676037725
transform 1 0 8188 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_89
timestamp 1676037725
transform 1 0 9292 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_89_97
timestamp 1676037725
transform 1 0 10028 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_101
timestamp 1676037725
transform 1 0 10396 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_89_105
timestamp 1676037725
transform 1 0 10764 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_111
timestamp 1676037725
transform 1 0 11316 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_113
timestamp 1676037725
transform 1 0 11500 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_125
timestamp 1676037725
transform 1 0 12604 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_137
timestamp 1676037725
transform 1 0 13708 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_149
timestamp 1676037725
transform 1 0 14812 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_161
timestamp 1676037725
transform 1 0 15916 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_167
timestamp 1676037725
transform 1 0 16468 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_169
timestamp 1676037725
transform 1 0 16652 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_181
timestamp 1676037725
transform 1 0 17756 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_193
timestamp 1676037725
transform 1 0 18860 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_205
timestamp 1676037725
transform 1 0 19964 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_217
timestamp 1676037725
transform 1 0 21068 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_223
timestamp 1676037725
transform 1 0 21620 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_225
timestamp 1676037725
transform 1 0 21804 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_237
timestamp 1676037725
transform 1 0 22908 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_249
timestamp 1676037725
transform 1 0 24012 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_255
timestamp 1676037725
transform 1 0 24564 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_89_258
timestamp 1676037725
transform 1 0 24840 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_89_264
timestamp 1676037725
transform 1 0 25392 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_90_3
timestamp 1676037725
transform 1 0 1380 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_9
timestamp 1676037725
transform 1 0 1932 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_90_26
timestamp 1676037725
transform 1 0 3496 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_90_29
timestamp 1676037725
transform 1 0 3772 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_90_47
timestamp 1676037725
transform 1 0 5428 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_90_51
timestamp 1676037725
transform 1 0 5796 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_90_55
timestamp 1676037725
transform 1 0 6164 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_90_75
timestamp 1676037725
transform 1 0 8004 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_90_83
timestamp 1676037725
transform 1 0 8740 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_85
timestamp 1676037725
transform 1 0 8924 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_97
timestamp 1676037725
transform 1 0 10028 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_109
timestamp 1676037725
transform 1 0 11132 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_121
timestamp 1676037725
transform 1 0 12236 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_133
timestamp 1676037725
transform 1 0 13340 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_139
timestamp 1676037725
transform 1 0 13892 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_141
timestamp 1676037725
transform 1 0 14076 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_153
timestamp 1676037725
transform 1 0 15180 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_165
timestamp 1676037725
transform 1 0 16284 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_177
timestamp 1676037725
transform 1 0 17388 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_189
timestamp 1676037725
transform 1 0 18492 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_195
timestamp 1676037725
transform 1 0 19044 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_197
timestamp 1676037725
transform 1 0 19228 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_209
timestamp 1676037725
transform 1 0 20332 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_221
timestamp 1676037725
transform 1 0 21436 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_233
timestamp 1676037725
transform 1 0 22540 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_90_245
timestamp 1676037725
transform 1 0 23644 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_90_250
timestamp 1676037725
transform 1 0 24104 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_90_255
timestamp 1676037725
transform 1 0 24564 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_90_258
timestamp 1676037725
transform 1 0 24840 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_90_264
timestamp 1676037725
transform 1 0 25392 0 1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_91_3
timestamp 1676037725
transform 1 0 1380 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_91_15
timestamp 1676037725
transform 1 0 2484 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_91_34
timestamp 1676037725
transform 1 0 4232 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_91_54
timestamp 1676037725
transform 1 0 6072 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_91_57
timestamp 1676037725
transform 1 0 6348 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_91_79
timestamp 1676037725
transform 1 0 8372 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_91_103
timestamp 1676037725
transform 1 0 10580 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_91_111
timestamp 1676037725
transform 1 0 11316 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_91_113
timestamp 1676037725
transform 1 0 11500 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_91_118
timestamp 1676037725
transform 1 0 11960 0 -1 52224
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_91_123
timestamp 1676037725
transform 1 0 12420 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_135
timestamp 1676037725
transform 1 0 13524 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_147
timestamp 1676037725
transform 1 0 14628 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_159
timestamp 1676037725
transform 1 0 15732 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_91_167
timestamp 1676037725
transform 1 0 16468 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_169
timestamp 1676037725
transform 1 0 16652 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_181
timestamp 1676037725
transform 1 0 17756 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_193
timestamp 1676037725
transform 1 0 18860 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_205
timestamp 1676037725
transform 1 0 19964 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_217
timestamp 1676037725
transform 1 0 21068 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_223
timestamp 1676037725
transform 1 0 21620 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_225
timestamp 1676037725
transform 1 0 21804 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_91_237
timestamp 1676037725
transform 1 0 22908 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_91_244
timestamp 1676037725
transform 1 0 23552 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_91_249
timestamp 1676037725
transform 1 0 24012 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_91_256
timestamp 1676037725
transform 1 0 24656 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_91_264
timestamp 1676037725
transform 1 0 25392 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_92_3
timestamp 1676037725
transform 1 0 1380 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_9
timestamp 1676037725
transform 1 0 1932 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_92_26
timestamp 1676037725
transform 1 0 3496 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_92_29
timestamp 1676037725
transform 1 0 3772 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_92_41
timestamp 1676037725
transform 1 0 4876 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_45
timestamp 1676037725
transform 1 0 5244 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_92_62
timestamp 1676037725
transform 1 0 6808 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_92_82
timestamp 1676037725
transform 1 0 8648 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_92_85
timestamp 1676037725
transform 1 0 8924 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_92_93
timestamp 1676037725
transform 1 0 9660 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_92_111
timestamp 1676037725
transform 1 0 11316 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_115
timestamp 1676037725
transform 1 0 11684 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_92_119
timestamp 1676037725
transform 1 0 12052 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_126
timestamp 1676037725
transform 1 0 12696 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_130
timestamp 1676037725
transform 1 0 13064 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_92_135
timestamp 1676037725
transform 1 0 13524 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_92_139
timestamp 1676037725
transform 1 0 13892 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_143
timestamp 1676037725
transform 1 0 14260 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_155
timestamp 1676037725
transform 1 0 15364 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_167
timestamp 1676037725
transform 1 0 16468 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_179
timestamp 1676037725
transform 1 0 17572 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_191
timestamp 1676037725
transform 1 0 18676 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_195
timestamp 1676037725
transform 1 0 19044 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_197
timestamp 1676037725
transform 1 0 19228 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_209
timestamp 1676037725
transform 1 0 20332 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_221
timestamp 1676037725
transform 1 0 21436 0 1 52224
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_92_227
timestamp 1676037725
transform 1 0 21988 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_242
timestamp 1676037725
transform 1 0 23368 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_92_249
timestamp 1676037725
transform 1 0 24012 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_92_253
timestamp 1676037725
transform 1 0 24380 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_92_258
timestamp 1676037725
transform 1 0 24840 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_93_3
timestamp 1676037725
transform 1 0 1380 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_93_8
timestamp 1676037725
transform 1 0 1840 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_93_12
timestamp 1676037725
transform 1 0 2208 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_93_34
timestamp 1676037725
transform 1 0 4232 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_93_54
timestamp 1676037725
transform 1 0 6072 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_93_57
timestamp 1676037725
transform 1 0 6348 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_93_63
timestamp 1676037725
transform 1 0 6900 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_93_71
timestamp 1676037725
transform 1 0 7636 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_93_90
timestamp 1676037725
transform 1 0 9384 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_93_110
timestamp 1676037725
transform 1 0 11224 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_93_113
timestamp 1676037725
transform 1 0 11500 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_93_131
timestamp 1676037725
transform 1 0 13156 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_139
timestamp 1676037725
transform 1 0 13892 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_93_147
timestamp 1676037725
transform 1 0 14628 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_93_151
timestamp 1676037725
transform 1 0 14996 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_93_159
timestamp 1676037725
transform 1 0 15732 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_93_163
timestamp 1676037725
transform 1 0 16100 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_93_167
timestamp 1676037725
transform 1 0 16468 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_93_171
timestamp 1676037725
transform 1 0 16836 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_93_175
timestamp 1676037725
transform 1 0 17204 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_93_183
timestamp 1676037725
transform 1 0 17940 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_93_187
timestamp 1676037725
transform 1 0 18308 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_93_191
timestamp 1676037725
transform 1 0 18676 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_93_199
timestamp 1676037725
transform 1 0 19412 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_93_206
timestamp 1676037725
transform 1 0 20056 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_93_210
timestamp 1676037725
transform 1 0 20424 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_93_215
timestamp 1676037725
transform 1 0 20884 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_93_219
timestamp 1676037725
transform 1 0 21252 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_93_225
timestamp 1676037725
transform 1 0 21804 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_93_231
timestamp 1676037725
transform 1 0 22356 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_93_238
timestamp 1676037725
transform 1 0 23000 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_93_242
timestamp 1676037725
transform 1 0 23368 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_93_264
timestamp 1676037725
transform 1 0 25392 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_94_3
timestamp 1676037725
transform 1 0 1380 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_9
timestamp 1676037725
transform 1 0 1932 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_94_26
timestamp 1676037725
transform 1 0 3496 0 1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_94_31
timestamp 1676037725
transform 1 0 3956 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_94_43
timestamp 1676037725
transform 1 0 5060 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_94_62
timestamp 1676037725
transform 1 0 6808 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_94_82
timestamp 1676037725
transform 1 0 8648 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_94_85
timestamp 1676037725
transform 1 0 8924 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_94_93
timestamp 1676037725
transform 1 0 9660 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_94_111
timestamp 1676037725
transform 1 0 11316 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_131
timestamp 1676037725
transform 1 0 13156 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_94_138
timestamp 1676037725
transform 1 0 13800 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_141
timestamp 1676037725
transform 1 0 14076 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_147
timestamp 1676037725
transform 1 0 14628 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_151
timestamp 1676037725
transform 1 0 14996 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_157
timestamp 1676037725
transform 1 0 15548 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_94_163
timestamp 1676037725
transform 1 0 16100 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_171
timestamp 1676037725
transform 1 0 16836 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_178
timestamp 1676037725
transform 1 0 17480 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_182
timestamp 1676037725
transform 1 0 17848 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_187
timestamp 1676037725
transform 1 0 18308 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_94_194
timestamp 1676037725
transform 1 0 18952 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_197
timestamp 1676037725
transform 1 0 19228 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_203
timestamp 1676037725
transform 1 0 19780 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_209
timestamp 1676037725
transform 1 0 20332 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_94_215
timestamp 1676037725
transform 1 0 20884 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_223
timestamp 1676037725
transform 1 0 21620 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_230
timestamp 1676037725
transform 1 0 22264 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_94_250
timestamp 1676037725
transform 1 0 24104 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_253
timestamp 1676037725
transform 1 0 24380 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_258
timestamp 1676037725
transform 1 0 24840 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_262
timestamp 1676037725
transform 1 0 25208 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_95_3
timestamp 1676037725
transform 1 0 1380 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_9
timestamp 1676037725
transform 1 0 1932 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_26
timestamp 1676037725
transform 1 0 3496 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_29
timestamp 1676037725
transform 1 0 3772 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_37
timestamp 1676037725
transform 1 0 4508 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_54
timestamp 1676037725
transform 1 0 6072 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_57
timestamp 1676037725
transform 1 0 6348 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_65
timestamp 1676037725
transform 1 0 7084 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_82
timestamp 1676037725
transform 1 0 8648 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_85
timestamp 1676037725
transform 1 0 8924 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_93
timestamp 1676037725
transform 1 0 9660 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_110
timestamp 1676037725
transform 1 0 11224 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_95_113
timestamp 1676037725
transform 1 0 11500 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_95_135
timestamp 1676037725
transform 1 0 13524 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_95_141
timestamp 1676037725
transform 1 0 14076 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_145
timestamp 1676037725
transform 1 0 14444 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_151
timestamp 1676037725
transform 1 0 14996 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_159
timestamp 1676037725
transform 1 0 15732 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_166
timestamp 1676037725
transform 1 0 16376 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_169
timestamp 1676037725
transform 1 0 16652 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_175
timestamp 1676037725
transform 1 0 17204 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_183
timestamp 1676037725
transform 1 0 17940 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_191
timestamp 1676037725
transform 1 0 18676 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_95_195
timestamp 1676037725
transform 1 0 19044 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_197
timestamp 1676037725
transform 1 0 19228 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_203
timestamp 1676037725
transform 1 0 19780 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_211
timestamp 1676037725
transform 1 0 20516 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_219
timestamp 1676037725
transform 1 0 21252 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_95_223
timestamp 1676037725
transform 1 0 21620 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_225
timestamp 1676037725
transform 1 0 21804 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_230
timestamp 1676037725
transform 1 0 22264 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_250
timestamp 1676037725
transform 1 0 24104 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_253
timestamp 1676037725
transform 1 0 24380 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_258
timestamp 1676037725
transform 1 0 24840 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_262
timestamp 1676037725
transform 1 0 25208 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1676037725
transform -1 0 1840 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1676037725
transform -1 0 2576 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1676037725
transform 1 0 25116 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1676037725
transform 1 0 25116 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1676037725
transform 1 0 25116 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1676037725
transform 1 0 25116 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1676037725
transform 1 0 25116 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1676037725
transform 1 0 25116 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1676037725
transform 1 0 25116 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1676037725
transform 1 0 25116 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1676037725
transform 1 0 23828 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1676037725
transform 1 0 25116 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1676037725
transform 1 0 25116 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1676037725
transform 1 0 21252 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input15
timestamp 1676037725
transform -1 0 25392 0 -1 40256
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input16
timestamp 1676037725
transform -1 0 24104 0 -1 40256
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1676037725
transform 1 0 23828 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input18
timestamp 1676037725
transform -1 0 24104 0 1 41344
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1676037725
transform 1 0 25116 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1676037725
transform 1 0 25116 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input21
timestamp 1676037725
transform -1 0 25392 0 -1 44608
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input22
timestamp 1676037725
transform -1 0 25392 0 -1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1676037725
transform 1 0 24564 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1676037725
transform 1 0 23276 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1676037725
transform 1 0 23276 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1676037725
transform 1 0 23828 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1676037725
transform 1 0 23828 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1676037725
transform 1 0 23920 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1676037725
transform 1 0 25116 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1676037725
transform 1 0 25116 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1676037725
transform 1 0 25116 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input32
timestamp 1676037725
transform -1 0 25392 0 -1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1676037725
transform -1 0 1840 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input34 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4876 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input35
timestamp 1676037725
transform -1 0 5336 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1676037725
transform -1 0 5888 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input37
timestamp 1676037725
transform 1 0 5704 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input38
timestamp 1676037725
transform 1 0 6348 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input39
timestamp 1676037725
transform -1 0 6072 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input40
timestamp 1676037725
transform 1 0 7084 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input41
timestamp 1676037725
transform 1 0 7452 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input42
timestamp 1676037725
transform 1 0 6992 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input43
timestamp 1676037725
transform 1 0 8188 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input44
timestamp 1676037725
transform 1 0 1564 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input45
timestamp 1676037725
transform 1 0 8556 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input46
timestamp 1676037725
transform -1 0 8188 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input47
timestamp 1676037725
transform 1 0 9292 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input48
timestamp 1676037725
transform -1 0 9660 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input49
timestamp 1676037725
transform 1 0 10028 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input50
timestamp 1676037725
transform -1 0 11224 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input51
timestamp 1676037725
transform 1 0 11316 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input52
timestamp 1676037725
transform -1 0 8648 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1676037725
transform -1 0 11960 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input54
timestamp 1676037725
transform -1 0 12604 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input55
timestamp 1676037725
transform 1 0 1932 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input56
timestamp 1676037725
transform 1 0 1840 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input57
timestamp 1676037725
transform -1 0 3496 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input58
timestamp 1676037725
transform 1 0 3036 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input59
timestamp 1676037725
transform 1 0 2760 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input60
timestamp 1676037725
transform -1 0 3864 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input61
timestamp 1676037725
transform 1 0 4140 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input62
timestamp 1676037725
transform 1 0 4232 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1676037725
transform -1 0 12696 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input64
timestamp 1676037725
transform 1 0 16836 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input65
timestamp 1676037725
transform 1 0 16468 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1676037725
transform -1 0 17480 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input67
timestamp 1676037725
transform -1 0 17940 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input68
timestamp 1676037725
transform 1 0 18308 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input69
timestamp 1676037725
transform 1 0 17940 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input70
timestamp 1676037725
transform 1 0 18676 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input71
timestamp 1676037725
transform 1 0 19412 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input72
timestamp 1676037725
transform -1 0 19780 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input73
timestamp 1676037725
transform -1 0 20516 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input74
timestamp 1676037725
transform -1 0 14628 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input75
timestamp 1676037725
transform 1 0 19780 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input76
timestamp 1676037725
transform 1 0 20884 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input77
timestamp 1676037725
transform 1 0 20516 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input78
timestamp 1676037725
transform 1 0 21252 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input79
timestamp 1676037725
transform 1 0 21988 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input80
timestamp 1676037725
transform 1 0 21988 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input81
timestamp 1676037725
transform 1 0 21988 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input82
timestamp 1676037725
transform 1 0 22724 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input83
timestamp 1676037725
transform 1 0 24564 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input84
timestamp 1676037725
transform 1 0 24564 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input85
timestamp 1676037725
transform 1 0 13156 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input86
timestamp 1676037725
transform -1 0 13892 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input87
timestamp 1676037725
transform -1 0 13800 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input88
timestamp 1676037725
transform -1 0 14628 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input89
timestamp 1676037725
transform 1 0 14628 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input90
timestamp 1676037725
transform 1 0 15364 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input91
timestamp 1676037725
transform -1 0 16376 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input92
timestamp 1676037725
transform 1 0 15732 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input93
timestamp 1676037725
transform -1 0 1840 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input94
timestamp 1676037725
transform -1 0 1840 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input95
timestamp 1676037725
transform -1 0 1840 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input96
timestamp 1676037725
transform -1 0 1840 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input97
timestamp 1676037725
transform 1 0 1564 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  input98
timestamp 1676037725
transform -1 0 25392 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  input99
timestamp 1676037725
transform -1 0 1840 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input100
timestamp 1676037725
transform -1 0 24012 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input101
timestamp 1676037725
transform -1 0 24932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input102
timestamp 1676037725
transform -1 0 24104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input103
timestamp 1676037725
transform -1 0 23368 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input104
timestamp 1676037725
transform -1 0 25392 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input105
timestamp 1676037725
transform -1 0 25392 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input106
timestamp 1676037725
transform -1 0 25392 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input107
timestamp 1676037725
transform -1 0 25392 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input108
timestamp 1676037725
transform -1 0 25392 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input109
timestamp 1676037725
transform -1 0 25392 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input110
timestamp 1676037725
transform -1 0 25392 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input111
timestamp 1676037725
transform -1 0 25392 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input112
timestamp 1676037725
transform 1 0 25024 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input113
timestamp 1676037725
transform 1 0 24380 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input114
timestamp 1676037725
transform 1 0 23828 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input115
timestamp 1676037725
transform 1 0 1564 0 1 45696
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input116
timestamp 1676037725
transform 1 0 1564 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input117
timestamp 1676037725
transform 1 0 1564 0 -1 51136
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input118
timestamp 1676037725
transform 1 0 3956 0 1 52224
box -38 -48 958 592
use sky130_fd_sc_hd__conb_1  left_tile_225
timestamp 1676037725
transform 1 0 25116 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  output119 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20056 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output120
timestamp 1676037725
transform -1 0 5428 0 1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output121
timestamp 1676037725
transform 1 0 22632 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output122
timestamp 1676037725
transform 1 0 22080 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output123
timestamp 1676037725
transform 1 0 23920 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output124
timestamp 1676037725
transform 1 0 23920 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output125
timestamp 1676037725
transform 1 0 22080 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output126
timestamp 1676037725
transform 1 0 23920 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output127
timestamp 1676037725
transform 1 0 22632 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output128
timestamp 1676037725
transform -1 0 23552 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output129
timestamp 1676037725
transform 1 0 23920 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output130
timestamp 1676037725
transform 1 0 23920 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output131
timestamp 1676037725
transform 1 0 23920 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output132
timestamp 1676037725
transform -1 0 24104 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output133
timestamp 1676037725
transform -1 0 21528 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output134
timestamp 1676037725
transform -1 0 23552 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output135
timestamp 1676037725
transform -1 0 24104 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output136
timestamp 1676037725
transform -1 0 25392 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output137
timestamp 1676037725
transform -1 0 24104 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output138
timestamp 1676037725
transform -1 0 24104 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output139
timestamp 1676037725
transform -1 0 23552 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output140
timestamp 1676037725
transform -1 0 24104 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output141
timestamp 1676037725
transform 1 0 23920 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output142
timestamp 1676037725
transform -1 0 24104 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output143
timestamp 1676037725
transform 1 0 23920 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output144
timestamp 1676037725
transform -1 0 24104 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output145
timestamp 1676037725
transform 1 0 23920 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output146
timestamp 1676037725
transform 1 0 23920 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output147
timestamp 1676037725
transform -1 0 24104 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output148
timestamp 1676037725
transform 1 0 23920 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output149
timestamp 1676037725
transform 1 0 23920 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output150
timestamp 1676037725
transform -1 0 11224 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output151
timestamp 1676037725
transform 1 0 16836 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output152
timestamp 1676037725
transform 1 0 16836 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output153
timestamp 1676037725
transform 1 0 18676 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output154
timestamp 1676037725
transform 1 0 19412 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output155
timestamp 1676037725
transform 1 0 17388 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output156
timestamp 1676037725
transform 1 0 19412 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output157
timestamp 1676037725
transform 1 0 18676 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output158
timestamp 1676037725
transform 1 0 21988 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output159
timestamp 1676037725
transform 1 0 19412 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output160
timestamp 1676037725
transform 1 0 21252 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output161
timestamp 1676037725
transform -1 0 13800 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output162
timestamp 1676037725
transform 1 0 19596 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output163
timestamp 1676037725
transform 1 0 21252 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output164
timestamp 1676037725
transform 1 0 21988 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output165
timestamp 1676037725
transform 1 0 20700 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output166
timestamp 1676037725
transform 1 0 21988 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output167
timestamp 1676037725
transform 1 0 23828 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output168
timestamp 1676037725
transform 1 0 22540 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output169
timestamp 1676037725
transform 1 0 22080 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output170
timestamp 1676037725
transform 1 0 22080 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output171
timestamp 1676037725
transform 1 0 20792 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output172
timestamp 1676037725
transform 1 0 12972 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output173
timestamp 1676037725
transform 1 0 12328 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output174
timestamp 1676037725
transform -1 0 14444 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output175
timestamp 1676037725
transform 1 0 14260 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output176
timestamp 1676037725
transform -1 0 15916 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output177
timestamp 1676037725
transform -1 0 16284 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output178
timestamp 1676037725
transform 1 0 16836 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output179
timestamp 1676037725
transform 1 0 16100 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output180
timestamp 1676037725
transform -1 0 3036 0 1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output181
timestamp 1676037725
transform -1 0 6072 0 -1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output182
timestamp 1676037725
transform -1 0 3496 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output183
timestamp 1676037725
transform -1 0 6072 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output184
timestamp 1676037725
transform -1 0 6808 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output185
timestamp 1676037725
transform -1 0 8004 0 1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output186
timestamp 1676037725
transform 1 0 6900 0 -1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output187
timestamp 1676037725
transform -1 0 6072 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output188
timestamp 1676037725
transform -1 0 6808 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output189
timestamp 1676037725
transform -1 0 8648 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output190
timestamp 1676037725
transform 1 0 7176 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output191
timestamp 1676037725
transform -1 0 3220 0 -1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output192
timestamp 1676037725
transform -1 0 9384 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output193
timestamp 1676037725
transform -1 0 10580 0 -1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output194
timestamp 1676037725
transform -1 0 8648 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output195
timestamp 1676037725
transform 1 0 9844 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output196
timestamp 1676037725
transform 1 0 9752 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output197
timestamp 1676037725
transform -1 0 11316 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output198
timestamp 1676037725
transform 1 0 9752 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output199
timestamp 1676037725
transform 1 0 11684 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output200
timestamp 1676037725
transform 1 0 11684 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output201
timestamp 1676037725
transform 1 0 12052 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output202
timestamp 1676037725
transform -1 0 3496 0 1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output203
timestamp 1676037725
transform -1 0 3496 0 1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output204
timestamp 1676037725
transform -1 0 4324 0 -1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output205
timestamp 1676037725
transform -1 0 3496 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output206
timestamp 1676037725
transform -1 0 4232 0 -1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output207
timestamp 1676037725
transform -1 0 5428 0 1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output208
timestamp 1676037725
transform -1 0 4232 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output209
timestamp 1676037725
transform -1 0 3496 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output210
timestamp 1676037725
transform -1 0 3036 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output211
timestamp 1676037725
transform 1 0 1564 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output212
timestamp 1676037725
transform 1 0 1564 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output213
timestamp 1676037725
transform 1 0 1564 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output214
timestamp 1676037725
transform -1 0 3036 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output215
timestamp 1676037725
transform 1 0 1564 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output216
timestamp 1676037725
transform 1 0 1564 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output217
timestamp 1676037725
transform 1 0 1564 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output218
timestamp 1676037725
transform -1 0 19228 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output219
timestamp 1676037725
transform 1 0 23920 0 -1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output220
timestamp 1676037725
transform -1 0 24104 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output221
timestamp 1676037725
transform -1 0 23552 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output222
timestamp 1676037725
transform -1 0 25392 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output223
timestamp 1676037725
transform -1 0 21528 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output224
timestamp 1676037725
transform -1 0 24104 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 25852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 25852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 25852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 25852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 25852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 25852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 25852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 25852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 25852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 25852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 25852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1676037725
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1676037725
transform -1 0 25852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1676037725
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1676037725
transform -1 0 25852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1676037725
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1676037725
transform -1 0 25852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1676037725
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1676037725
transform -1 0 25852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1676037725
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1676037725
transform -1 0 25852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1676037725
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1676037725
transform -1 0 25852 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1676037725
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1676037725
transform -1 0 25852 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1676037725
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1676037725
transform -1 0 25852 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1676037725
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1676037725
transform -1 0 25852 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1676037725
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1676037725
transform -1 0 25852 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1676037725
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1676037725
transform -1 0 25852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1676037725
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1676037725
transform -1 0 25852 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1676037725
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1676037725
transform -1 0 25852 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1676037725
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1676037725
transform -1 0 25852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1676037725
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1676037725
transform -1 0 25852 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1676037725
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1676037725
transform -1 0 25852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1676037725
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1676037725
transform -1 0 25852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1676037725
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1676037725
transform -1 0 25852 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1676037725
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1676037725
transform -1 0 25852 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1676037725
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1676037725
transform -1 0 25852 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1676037725
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1676037725
transform -1 0 25852 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1676037725
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1676037725
transform -1 0 25852 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1676037725
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1676037725
transform -1 0 25852 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1676037725
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1676037725
transform -1 0 25852 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1676037725
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1676037725
transform -1 0 25852 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1676037725
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1676037725
transform -1 0 25852 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1676037725
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1676037725
transform -1 0 25852 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1676037725
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1676037725
transform -1 0 25852 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1676037725
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1676037725
transform -1 0 25852 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1676037725
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1676037725
transform -1 0 25852 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1676037725
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1676037725
transform -1 0 25852 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1676037725
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1676037725
transform -1 0 25852 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1676037725
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1676037725
transform -1 0 25852 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1676037725
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1676037725
transform -1 0 25852 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1676037725
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1676037725
transform -1 0 25852 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1676037725
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1676037725
transform -1 0 25852 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1676037725
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1676037725
transform -1 0 25852 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1676037725
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1676037725
transform -1 0 25852 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1676037725
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1676037725
transform -1 0 25852 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1676037725
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1676037725
transform -1 0 25852 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1676037725
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1676037725
transform -1 0 25852 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1676037725
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1676037725
transform -1 0 25852 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1676037725
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1676037725
transform -1 0 25852 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1676037725
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1676037725
transform -1 0 25852 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1676037725
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1676037725
transform -1 0 25852 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1676037725
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1676037725
transform -1 0 25852 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1676037725
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1676037725
transform -1 0 25852 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1676037725
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1676037725
transform -1 0 25852 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1676037725
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1676037725
transform -1 0 25852 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1676037725
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1676037725
transform -1 0 25852 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1676037725
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1676037725
transform -1 0 25852 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1676037725
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1676037725
transform -1 0 25852 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1676037725
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1676037725
transform -1 0 25852 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1676037725
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1676037725
transform -1 0 25852 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1676037725
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1676037725
transform -1 0 25852 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1676037725
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1676037725
transform -1 0 25852 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1676037725
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1676037725
transform -1 0 25852 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1676037725
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1676037725
transform -1 0 25852 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1676037725
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1676037725
transform -1 0 25852 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1676037725
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1676037725
transform -1 0 25852 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1676037725
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1676037725
transform -1 0 25852 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1676037725
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1676037725
transform -1 0 25852 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1676037725
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1676037725
transform -1 0 25852 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1676037725
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1676037725
transform -1 0 25852 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1676037725
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1676037725
transform -1 0 25852 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1676037725
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1676037725
transform -1 0 25852 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1676037725
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1676037725
transform -1 0 25852 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1676037725
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1676037725
transform -1 0 25852 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1676037725
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1676037725
transform -1 0 25852 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1676037725
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1676037725
transform -1 0 25852 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1676037725
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1676037725
transform -1 0 25852 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1676037725
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1676037725
transform -1 0 25852 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1676037725
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1676037725
transform -1 0 25852 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1676037725
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1676037725
transform -1 0 25852 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1676037725
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1676037725
transform -1 0 25852 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1676037725
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1676037725
transform -1 0 25852 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1676037725
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1676037725
transform -1 0 25852 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1676037725
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1676037725
transform -1 0 25852 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1676037725
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1676037725
transform -1 0 25852 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1676037725
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1676037725
transform -1 0 25852 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1676037725
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1676037725
transform -1 0 25852 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1676037725
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1676037725
transform -1 0 25852 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1676037725
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1676037725
transform -1 0 25852 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1676037725
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1676037725
transform -1 0 25852 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1676037725
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1676037725
transform -1 0 25852 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 17848 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 13340 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 14260 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 15640 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 17112 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 18676 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 20516 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22908 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform -1 0 25116 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_0__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 24748 0 -1 21760
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 21988 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform -1 0 21436 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_0__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 21160 0 -1 22848
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 14536 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 14536 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 16928 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 21252 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 20424 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21436 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22264 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 23184 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 24012 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 19596 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 14536 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 17020 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 16284 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 14260 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 16836 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 20792 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform -1 0 22264 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 18676 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 10488 0 -1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 18676 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22264 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform -1 0 25300 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 23460 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 25024 0 -1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 22264 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 25116 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 23000 0 1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 21436 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22724 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 23184 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform -1 0 25392 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 25300 0 -1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 21988 0 -1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform -1 0 23828 0 1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 23828 0 -1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 21252 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 18400 0 -1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19412 0 1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 21252 0 1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 17848 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 19504 0 -1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 18676 0 -1 45696
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 15824 0 1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 17664 0 1 45696
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 16928 0 1 46784
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 14260 0 1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 15548 0 -1 46784
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 15180 0 -1 45696
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 14260 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 15456 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 15180 0 -1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform -1 0 13800 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11868 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 13524 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 10672 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11224 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 13616 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 13524 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 11040 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 10028 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 8096 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 6532 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 8096 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 6256 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 6348 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 7912 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 10948 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 10488 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 8648 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 6808 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 9292 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 11224 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 12604 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 14168 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 16836 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 15916 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 17296 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19412 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 21528 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 21988 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22632 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 23920 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 23460 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 22632 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 21528 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 19872 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 18952 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 16836 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 4416 0 1 48960
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 9384 0 -1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 10672 0 1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11776 0 1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 12144 0 -1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 9384 0 -1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 12236 0 1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 11224 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 7544 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 9752 0 -1 38080
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 7912 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform -1 0 6716 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_0__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 5244 0 1 36992
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 7084 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 4232 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 6716 0 -1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 10948 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 7728 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 9108 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 9476 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform -1 0 6992 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 5520 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 6716 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform -1 0 5336 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 4232 0 -1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 6348 0 1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 6532 0 -1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 7820 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 11224 0 1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 15180 0 1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 19504 0 -1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 17020 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_1.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15548 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_1.mux_l1_in_1_
timestamp 1676037725
transform 1 0 17664 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_1.mux_l1_in_2_
timestamp 1676037725
transform -1 0 12696 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_1.mux_l2_in_0_
timestamp 1676037725
transform 1 0 15088 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_1.mux_l2_in_1_
timestamp 1676037725
transform -1 0 13524 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_1.mux_l2_in_1__275
timestamp 1676037725
transform 1 0 13524 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_1.mux_l3_in_0_
timestamp 1676037725
transform 1 0 14352 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 14628 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_3.mux_l1_in_0_
timestamp 1676037725
transform -1 0 18216 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_3.mux_l1_in_1_
timestamp 1676037725
transform 1 0 19412 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_3.mux_l2_in_0_
timestamp 1676037725
transform 1 0 17940 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_3.mux_l2_in_1_
timestamp 1676037725
transform -1 0 17664 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_3.mux_l2_in_1__226
timestamp 1676037725
transform -1 0 16928 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_3.mux_l3_in_0_
timestamp 1676037725
transform 1 0 17848 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 17296 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_5.mux_l1_in_0_
timestamp 1676037725
transform -1 0 21436 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_5.mux_l1_in_1_
timestamp 1676037725
transform -1 0 22816 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_5.mux_l1_in_2_
timestamp 1676037725
transform 1 0 20700 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_5.mux_l2_in_0_
timestamp 1676037725
transform -1 0 22816 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_5.mux_l2_in_1_
timestamp 1676037725
transform -1 0 20240 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_5.mux_l2_in_1__229
timestamp 1676037725
transform 1 0 21988 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_5.mux_l3_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 20332 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_7.mux_l1_in_0_
timestamp 1676037725
transform -1 0 18768 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_7.mux_l1_in_1_
timestamp 1676037725
transform 1 0 20424 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_7.mux_l1_in_2_
timestamp 1676037725
transform -1 0 18584 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_7.mux_l1_in_3__231
timestamp 1676037725
transform 1 0 18032 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_7.mux_l1_in_3_
timestamp 1676037725
transform -1 0 17664 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_7.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19228 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_7.mux_l2_in_1_
timestamp 1676037725
transform -1 0 18952 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_7.mux_l3_in_0_
timestamp 1676037725
transform 1 0 18124 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 17296 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_11.mux_l1_in_0_
timestamp 1676037725
transform -1 0 17296 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_11.mux_l1_in_1_
timestamp 1676037725
transform 1 0 19228 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_11.mux_l1_in_2_
timestamp 1676037725
transform 1 0 16284 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_11.mux_l1_in_3__276
timestamp 1676037725
transform 1 0 13524 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_11.mux_l1_in_3_
timestamp 1676037725
transform -1 0 13800 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_11.mux_l2_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_11.mux_l2_in_1_
timestamp 1676037725
transform -1 0 16284 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_11.mux_l3_in_0_
timestamp 1676037725
transform 1 0 15548 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 16008 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_13.mux_l1_in_0_
timestamp 1676037725
transform -1 0 17940 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_13.mux_l1_in_1_
timestamp 1676037725
transform 1 0 20608 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_13.mux_l1_in_2_
timestamp 1676037725
transform -1 0 18216 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_13.mux_l2_in_0_
timestamp 1676037725
transform -1 0 20240 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_13.mux_l2_in_1__277
timestamp 1676037725
transform 1 0 20424 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_13.mux_l2_in_1_
timestamp 1676037725
transform -1 0 20056 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_13.mux_l3_in_0_
timestamp 1676037725
transform 1 0 19504 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18584 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_21.mux_l1_in_0_
timestamp 1676037725
transform -1 0 20516 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_21.mux_l1_in_1_
timestamp 1676037725
transform 1 0 22632 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_21.mux_l1_in_2_
timestamp 1676037725
transform -1 0 20608 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_21.mux_l2_in_0_
timestamp 1676037725
transform -1 0 22816 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_21.mux_l2_in_1__278
timestamp 1676037725
transform 1 0 23828 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_21.mux_l2_in_1_
timestamp 1676037725
transform -1 0 23460 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_21.mux_l3_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 21252 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_29.mux_l1_in_0_
timestamp 1676037725
transform -1 0 17664 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_29.mux_l1_in_1_
timestamp 1676037725
transform 1 0 19964 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_29.mux_l1_in_2_
timestamp 1676037725
transform 1 0 18032 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_29.mux_l2_in_0_
timestamp 1676037725
transform 1 0 17204 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_29.mux_l2_in_1__279
timestamp 1676037725
transform 1 0 18216 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_29.mux_l2_in_1_
timestamp 1676037725
transform 1 0 17020 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_29.mux_l3_in_0_
timestamp 1676037725
transform 1 0 16744 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 15548 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_37.mux_l1_in_0_
timestamp 1676037725
transform -1 0 18860 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_37.mux_l1_in_1_
timestamp 1676037725
transform 1 0 19044 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_37.mux_l2_in_0_
timestamp 1676037725
transform 1 0 18032 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_37.mux_l2_in_1__227
timestamp 1676037725
transform 1 0 13156 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_37.mux_l2_in_1_
timestamp 1676037725
transform -1 0 13524 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_37.mux_l3_in_0_
timestamp 1676037725
transform 1 0 14260 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 13156 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_45.mux_l1_in_0_
timestamp 1676037725
transform -1 0 21068 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_45.mux_l2_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_45.mux_l2_in_1_
timestamp 1676037725
transform 1 0 22632 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_45.mux_l2_in_1__228
timestamp 1676037725
transform 1 0 23092 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_45.mux_l3_in_0_
timestamp 1676037725
transform 1 0 20792 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19412 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_53.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14996 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_53.mux_l1_in_1__230
timestamp 1676037725
transform -1 0 14904 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_53.mux_l1_in_1_
timestamp 1676037725
transform 1 0 15272 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_53.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11316 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_0__1_.mux_bottom_track_53.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 9844 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_0.mux_l1_in_0_
timestamp 1676037725
transform -1 0 21528 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_0.mux_l1_in_1_
timestamp 1676037725
transform -1 0 22724 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_0.mux_l2_in_0_
timestamp 1676037725
transform -1 0 22816 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_0.mux_l2_in_1__232
timestamp 1676037725
transform -1 0 22264 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_0.mux_l2_in_1_
timestamp 1676037725
transform -1 0 22632 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_0.mux_l3_in_0_
timestamp 1676037725
transform -1 0 24012 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 24196 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_2.mux_l1_in_0_
timestamp 1676037725
transform 1 0 22816 0 1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_2.mux_l1_in_1_
timestamp 1676037725
transform 1 0 21988 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_2.mux_l1_in_2_
timestamp 1676037725
transform -1 0 20792 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_2.mux_l2_in_0_
timestamp 1676037725
transform -1 0 22816 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_2.mux_l2_in_1_
timestamp 1676037725
transform -1 0 22816 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_2.mux_l2_in_1__238
timestamp 1676037725
transform 1 0 23368 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_2.mux_l3_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 24840 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_4.mux_l1_in_0_
timestamp 1676037725
transform -1 0 22448 0 1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_4.mux_l1_in_1_
timestamp 1676037725
transform -1 0 21528 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_4.mux_l2_in_0_
timestamp 1676037725
transform 1 0 21896 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_4.mux_l2_in_1__249
timestamp 1676037725
transform 1 0 20240 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_4.mux_l2_in_1_
timestamp 1676037725
transform -1 0 20240 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_4.mux_l3_in_0_
timestamp 1676037725
transform -1 0 22356 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 23644 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_6.mux_l1_in_0_
timestamp 1676037725
transform -1 0 21528 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_6.mux_l1_in_1_
timestamp 1676037725
transform -1 0 22264 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_6.mux_l1_in_2_
timestamp 1676037725
transform -1 0 20332 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_6.mux_l2_in_0_
timestamp 1676037725
transform -1 0 23828 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_6.mux_l2_in_1__258
timestamp 1676037725
transform 1 0 23184 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_6.mux_l2_in_1_
timestamp 1676037725
transform -1 0 23552 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_6.mux_l3_in_0_
timestamp 1676037725
transform -1 0 24104 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 24840 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_8.mux_l1_in_0_
timestamp 1676037725
transform -1 0 21528 0 1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_8.mux_l1_in_1_
timestamp 1676037725
transform -1 0 21528 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_8.mux_l1_in_2_
timestamp 1676037725
transform -1 0 18952 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_8.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_8.mux_l2_in_1__259
timestamp 1676037725
transform -1 0 21528 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_8.mux_l2_in_1_
timestamp 1676037725
transform -1 0 22816 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_8.mux_l3_in_0_
timestamp 1676037725
transform -1 0 22816 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 23828 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_10.mux_l1_in_0_
timestamp 1676037725
transform 1 0 19688 0 -1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_10.mux_l1_in_1_
timestamp 1676037725
transform 1 0 19504 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_10.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19412 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_10.mux_l2_in_1__233
timestamp 1676037725
transform 1 0 16836 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_10.mux_l2_in_1_
timestamp 1676037725
transform -1 0 16744 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_10.mux_l3_in_0_
timestamp 1676037725
transform -1 0 20240 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 24104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_12.mux_l1_in_0_
timestamp 1676037725
transform -1 0 20240 0 1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_12.mux_l2_in_0_
timestamp 1676037725
transform -1 0 20240 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_12.mux_l2_in_1__234
timestamp 1676037725
transform 1 0 19412 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_12.mux_l2_in_1_
timestamp 1676037725
transform -1 0 17296 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_12.mux_l3_in_0_
timestamp 1676037725
transform -1 0 20700 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 22264 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_14.mux_l1_in_0_
timestamp 1676037725
transform 1 0 18032 0 -1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_14.mux_l2_in_0_
timestamp 1676037725
transform 1 0 17480 0 1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_14.mux_l2_in_1_
timestamp 1676037725
transform -1 0 16468 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_14.mux_l2_in_1__235
timestamp 1676037725
transform 1 0 16100 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_14.mux_l3_in_0_
timestamp 1676037725
transform -1 0 18216 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 22264 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_16.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_16.mux_l2_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_16.mux_l2_in_1__236
timestamp 1676037725
transform 1 0 14352 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_16.mux_l2_in_1_
timestamp 1676037725
transform -1 0 14536 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_16.mux_l3_in_0_
timestamp 1676037725
transform -1 0 16652 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 19780 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_18.mux_l1_in_0_
timestamp 1676037725
transform 1 0 17296 0 1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_18.mux_l2_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_18.mux_l2_in_1__237
timestamp 1676037725
transform 1 0 14076 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_18.mux_l2_in_1_
timestamp 1676037725
transform -1 0 13708 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_18.mux_l3_in_0_
timestamp 1676037725
transform -1 0 16284 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 19688 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_20.mux_l1_in_0_
timestamp 1676037725
transform -1 0 14996 0 -1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_20.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14904 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_20.mux_l2_in_1_
timestamp 1676037725
transform -1 0 13708 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_20.mux_l2_in_1__239
timestamp 1676037725
transform 1 0 13340 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_20.mux_l3_in_0_
timestamp 1676037725
transform -1 0 15456 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 19504 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_22.mux_l1_in_0_
timestamp 1676037725
transform -1 0 13708 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_22.mux_l2_in_0_
timestamp 1676037725
transform 1 0 13432 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_22.mux_l2_in_1__240
timestamp 1676037725
transform 1 0 11684 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_22.mux_l2_in_1_
timestamp 1676037725
transform -1 0 11408 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_22.mux_l3_in_0_
timestamp 1676037725
transform -1 0 13800 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 18216 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_24.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14628 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_24.mux_l1_in_1__241
timestamp 1676037725
transform 1 0 12604 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_24.mux_l1_in_1_
timestamp 1676037725
transform -1 0 12972 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_24.mux_l2_in_0_
timestamp 1676037725
transform -1 0 15088 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 19688 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_26.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14812 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_26.mux_l1_in_1__242
timestamp 1676037725
transform 1 0 10672 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_26.mux_l1_in_1_
timestamp 1676037725
transform -1 0 11040 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_26.mux_l2_in_0_
timestamp 1676037725
transform -1 0 13616 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 17756 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_28.mux_l1_in_0_
timestamp 1676037725
transform 1 0 11776 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_28.mux_l1_in_1__243
timestamp 1676037725
transform 1 0 8740 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_28.mux_l1_in_1_
timestamp 1676037725
transform -1 0 8280 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_28.mux_l2_in_0_
timestamp 1676037725
transform -1 0 10856 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 15824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_30.mux_l1_in_0_
timestamp 1676037725
transform 1 0 11776 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_30.mux_l1_in_1_
timestamp 1676037725
transform -1 0 8372 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_30.mux_l1_in_1__244
timestamp 1676037725
transform 1 0 8648 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_30.mux_l2_in_0_
timestamp 1676037725
transform -1 0 10764 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 15732 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_32.mux_l1_in_0_
timestamp 1676037725
transform 1 0 11868 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_32.mux_l1_in_1__245
timestamp 1676037725
transform -1 0 7544 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_32.mux_l1_in_1_
timestamp 1676037725
transform -1 0 8648 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_32.mux_l2_in_0_
timestamp 1676037725
transform -1 0 11224 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 16192 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_34.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14260 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_34.mux_l1_in_1__246
timestamp 1676037725
transform 1 0 10856 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_34.mux_l1_in_1_
timestamp 1676037725
transform -1 0 10488 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_34.mux_l2_in_0_
timestamp 1676037725
transform -1 0 13156 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 18216 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_36.mux_l1_in_0_
timestamp 1676037725
transform 1 0 11408 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_36.mux_l2_in_0_
timestamp 1676037725
transform -1 0 8372 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_36.mux_l2_in_1__247
timestamp 1676037725
transform -1 0 6072 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_36.mux_l2_in_1_
timestamp 1676037725
transform -1 0 7360 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_36.mux_l3_in_0_
timestamp 1676037725
transform -1 0 9660 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 16468 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_38.mux_l1_in_0_
timestamp 1676037725
transform -1 0 12880 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_38.mux_l2_in_0__248
timestamp 1676037725
transform 1 0 16100 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_38.mux_l2_in_0_
timestamp 1676037725
transform -1 0 15088 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_38.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 18400 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_40.mux_l1_in_0_
timestamp 1676037725
transform -1 0 14720 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_40.mux_l2_in_0_
timestamp 1676037725
transform -1 0 17664 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_40.mux_l2_in_0__250
timestamp 1676037725
transform -1 0 16928 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_40.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 19872 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_44.mux_l1_in_0_
timestamp 1676037725
transform -1 0 16376 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_44.mux_l2_in_0_
timestamp 1676037725
transform -1 0 18952 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_44.mux_l2_in_0__251
timestamp 1676037725
transform 1 0 18492 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_44.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 22264 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_46.mux_l1_in_0_
timestamp 1676037725
transform -1 0 17940 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_46.mux_l2_in_0_
timestamp 1676037725
transform -1 0 20700 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_46.mux_l2_in_0__252
timestamp 1676037725
transform 1 0 20608 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_46.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 22908 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_48.mux_l1_in_0_
timestamp 1676037725
transform -1 0 20240 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_48.mux_l2_in_0__253
timestamp 1676037725
transform 1 0 23828 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_48.mux_l2_in_0_
timestamp 1676037725
transform -1 0 22264 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_48.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 23920 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_50.mux_l1_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_50.mux_l1_in_1__254
timestamp 1676037725
transform 1 0 19504 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_50.mux_l1_in_1_
timestamp 1676037725
transform -1 0 19964 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_50.mux_l2_in_0_
timestamp 1676037725
transform -1 0 21528 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_50.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 23368 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_52.mux_l1_in_0_
timestamp 1676037725
transform -1 0 20240 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_52.mux_l2_in_0_
timestamp 1676037725
transform -1 0 21528 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_52.mux_l2_in_0__255
timestamp 1676037725
transform 1 0 23000 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_52.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 23000 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_54.mux_l1_in_0_
timestamp 1676037725
transform -1 0 18860 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_54.mux_l2_in_0__256
timestamp 1676037725
transform 1 0 20608 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_54.mux_l2_in_0_
timestamp 1676037725
transform -1 0 20240 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_54.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 22264 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_56.mux_l1_in_0_
timestamp 1676037725
transform -1 0 17848 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_56.mux_l2_in_0__257
timestamp 1676037725
transform 1 0 19044 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_56.mux_l2_in_0_
timestamp 1676037725
transform -1 0 18952 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_56.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 21344 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_0.mux_l1_in_0_
timestamp 1676037725
transform -1 0 10212 0 1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_0.mux_l1_in_1_
timestamp 1676037725
transform 1 0 17388 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_0.mux_l1_in_2_
timestamp 1676037725
transform 1 0 15180 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_0.mux_l1_in_3_
timestamp 1676037725
transform -1 0 10948 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_0.mux_l1_in_3__260
timestamp 1676037725
transform 1 0 10948 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_0.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12236 0 -1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_0.mux_l2_in_1_
timestamp 1676037725
transform -1 0 12512 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_0.mux_l3_in_0_
timestamp 1676037725
transform 1 0 11684 0 -1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 11960 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_2.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15180 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_2.mux_l1_in_1_
timestamp 1676037725
transform 1 0 18124 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_2.mux_l1_in_2_
timestamp 1676037725
transform 1 0 11868 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_2.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14260 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_2.mux_l2_in_1_
timestamp 1676037725
transform -1 0 12604 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_2.mux_l2_in_1__263
timestamp 1676037725
transform 1 0 12236 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_2.mux_l3_in_0_
timestamp 1676037725
transform 1 0 11776 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 11776 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_4.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14444 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_4.mux_l1_in_1_
timestamp 1676037725
transform 1 0 18216 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_4.mux_l1_in_2_
timestamp 1676037725
transform 1 0 10120 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_4.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12972 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_4.mux_l2_in_1__267
timestamp 1676037725
transform 1 0 10488 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_4.mux_l2_in_1_
timestamp 1676037725
transform -1 0 10396 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_4.mux_l3_in_0_
timestamp 1676037725
transform 1 0 9752 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 10028 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_6.mux_l1_in_0_
timestamp 1676037725
transform -1 0 9936 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_6.mux_l1_in_1_
timestamp 1676037725
transform 1 0 17112 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_6.mux_l1_in_2_
timestamp 1676037725
transform 1 0 12972 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_6.mux_l1_in_3__270
timestamp 1676037725
transform 1 0 7452 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_6.mux_l1_in_3_
timestamp 1676037725
transform -1 0 7912 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_6.mux_l2_in_0_
timestamp 1676037725
transform 1 0 9476 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_6.mux_l2_in_1_
timestamp 1676037725
transform 1 0 9016 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_6.mux_l3_in_0_
timestamp 1676037725
transform -1 0 8464 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 8648 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_10.mux_l1_in_0_
timestamp 1676037725
transform -1 0 8556 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_10.mux_l1_in_1_
timestamp 1676037725
transform 1 0 16836 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_10.mux_l1_in_2_
timestamp 1676037725
transform 1 0 12604 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_10.mux_l1_in_3__261
timestamp 1676037725
transform 1 0 8832 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_10.mux_l1_in_3_
timestamp 1676037725
transform -1 0 7820 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_10.mux_l2_in_0_
timestamp 1676037725
transform 1 0 9752 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_10.mux_l2_in_1_
timestamp 1676037725
transform 1 0 9936 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_10.mux_l3_in_0_
timestamp 1676037725
transform 1 0 7728 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 8096 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_12.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14260 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_12.mux_l1_in_1_
timestamp 1676037725
transform 1 0 17296 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_12.mux_l1_in_2_
timestamp 1676037725
transform -1 0 9936 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_12.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12236 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_12.mux_l2_in_1_
timestamp 1676037725
transform -1 0 9936 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_12.mux_l2_in_1__262
timestamp 1676037725
transform -1 0 8740 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_12.mux_l3_in_0_
timestamp 1676037725
transform 1 0 9752 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 7912 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_20.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14076 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_20.mux_l1_in_1_
timestamp 1676037725
transform 1 0 18492 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_20.mux_l1_in_2_
timestamp 1676037725
transform 1 0 9108 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_20.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11684 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_20.mux_l2_in_1_
timestamp 1676037725
transform -1 0 8280 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_20.mux_l2_in_1__264
timestamp 1676037725
transform 1 0 8188 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_20.mux_l3_in_0_
timestamp 1676037725
transform 1 0 7636 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 7268 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_28.mux_l1_in_0_
timestamp 1676037725
transform 1 0 11684 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_28.mux_l1_in_1_
timestamp 1676037725
transform 1 0 12328 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_28.mux_l2_in_0_
timestamp 1676037725
transform 1 0 9108 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_28.mux_l2_in_1__265
timestamp 1676037725
transform 1 0 4968 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_28.mux_l2_in_1_
timestamp 1676037725
transform -1 0 5336 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_28.mux_l3_in_0_
timestamp 1676037725
transform 1 0 5152 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 5796 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_36.mux_l1_in_0_
timestamp 1676037725
transform 1 0 12604 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_36.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11960 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_36.mux_l2_in_1_
timestamp 1676037725
transform -1 0 8648 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_36.mux_l2_in_1__266
timestamp 1676037725
transform 1 0 8556 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_36.mux_l3_in_0_
timestamp 1676037725
transform 1 0 7820 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 7084 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_44.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16836 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_44.mux_l1_in_1__268
timestamp 1676037725
transform 1 0 10948 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_44.mux_l1_in_1_
timestamp 1676037725
transform -1 0 11500 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_44.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11960 0 1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_44.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 9108 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_52.mux_l1_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_52.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19688 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_52.mux_l2_in_1__269
timestamp 1676037725
transform -1 0 14812 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_52.mux_l2_in_1_
timestamp 1676037725
transform -1 0 15640 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_52.mux_l3_in_0_
timestamp 1676037725
transform 1 0 15732 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 10948 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1676037725
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1676037725
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1676037725
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1676037725
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1676037725
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1676037725
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1676037725
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1676037725
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1676037725
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1676037725
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1676037725
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1676037725
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1676037725
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1676037725
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1676037725
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1676037725
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1676037725
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1676037725
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1676037725
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1676037725
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1676037725
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1676037725
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1676037725
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1676037725
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1676037725
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1676037725
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1676037725
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1676037725
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1676037725
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1676037725
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1676037725
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1676037725
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1676037725
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1676037725
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1676037725
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1676037725
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1676037725
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1676037725
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1676037725
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1676037725
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1676037725
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1676037725
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1676037725
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1676037725
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1676037725
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1676037725
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1676037725
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1676037725
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1676037725
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1676037725
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1676037725
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1676037725
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1676037725
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1676037725
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1676037725
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1676037725
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1676037725
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1676037725
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1676037725
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1676037725
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1676037725
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1676037725
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1676037725
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1676037725
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1676037725
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1676037725
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1676037725
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1676037725
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1676037725
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1676037725
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1676037725
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1676037725
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1676037725
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1676037725
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1676037725
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1676037725
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1676037725
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1676037725
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1676037725
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1676037725
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1676037725
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1676037725
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1676037725
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1676037725
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1676037725
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1676037725
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1676037725
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1676037725
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1676037725
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1676037725
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1676037725
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1676037725
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1676037725
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1676037725
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1676037725
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1676037725
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1676037725
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1676037725
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1676037725
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1676037725
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1676037725
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1676037725
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1676037725
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1676037725
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1676037725
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1676037725
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1676037725
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1676037725
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1676037725
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1676037725
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1676037725
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1676037725
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1676037725
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1676037725
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1676037725
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1676037725
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1676037725
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1676037725
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1676037725
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1676037725
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1676037725
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1676037725
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1676037725
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1676037725
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1676037725
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1676037725
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1676037725
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1676037725
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1676037725
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1676037725
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1676037725
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1676037725
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1676037725
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1676037725
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1676037725
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1676037725
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1676037725
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1676037725
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1676037725
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1676037725
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1676037725
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1676037725
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1676037725
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1676037725
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1676037725
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1676037725
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1676037725
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1676037725
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1676037725
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1676037725
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1676037725
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1676037725
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1676037725
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1676037725
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1676037725
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1676037725
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1676037725
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1676037725
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1676037725
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1676037725
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1676037725
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1676037725
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1676037725
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1676037725
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1676037725
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1676037725
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1676037725
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1676037725
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1676037725
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1676037725
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1676037725
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1676037725
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1676037725
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1676037725
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1676037725
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1676037725
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1676037725
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1676037725
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1676037725
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1676037725
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1676037725
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1676037725
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1676037725
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1676037725
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1676037725
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1676037725
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1676037725
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1676037725
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1676037725
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1676037725
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1676037725
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1676037725
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1676037725
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1676037725
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1676037725
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1676037725
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1676037725
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1676037725
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1676037725
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1676037725
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1676037725
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1676037725
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1676037725
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1676037725
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1676037725
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1676037725
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1676037725
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1676037725
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1676037725
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1676037725
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1676037725
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1676037725
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1676037725
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1676037725
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1676037725
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1676037725
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1676037725
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1676037725
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1676037725
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1676037725
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1676037725
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1676037725
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1676037725
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1676037725
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1676037725
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1676037725
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1676037725
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1676037725
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1676037725
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1676037725
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1676037725
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1676037725
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1676037725
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1676037725
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1676037725
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1676037725
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1676037725
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1676037725
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1676037725
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1676037725
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1676037725
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1676037725
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1676037725
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1676037725
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1676037725
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1676037725
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1676037725
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1676037725
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1676037725
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1676037725
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1676037725
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1676037725
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1676037725
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1676037725
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1676037725
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1676037725
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1676037725
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1676037725
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1676037725
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1676037725
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1676037725
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1676037725
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1676037725
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1676037725
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1676037725
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1676037725
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1676037725
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1676037725
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1676037725
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1676037725
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1676037725
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1676037725
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1676037725
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1676037725
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1676037725
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1676037725
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1676037725
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1676037725
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1676037725
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1676037725
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1676037725
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1676037725
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1676037725
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1676037725
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1676037725
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1676037725
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1676037725
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1676037725
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1676037725
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1676037725
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1676037725
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1676037725
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1676037725
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1676037725
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1676037725
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1676037725
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1676037725
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1676037725
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1676037725
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1676037725
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1676037725
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1676037725
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1676037725
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1676037725
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1676037725
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1676037725
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1676037725
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1676037725
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1676037725
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1676037725
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1676037725
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1676037725
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1676037725
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1676037725
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1676037725
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1676037725
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1676037725
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1676037725
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1676037725
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1676037725
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1676037725
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1676037725
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1676037725
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1676037725
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1676037725
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1676037725
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1676037725
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1676037725
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1676037725
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1676037725
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1676037725
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1676037725
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1676037725
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1676037725
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1676037725
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1676037725
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1676037725
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1676037725
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1676037725
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1676037725
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1676037725
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1676037725
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1676037725
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1676037725
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1676037725
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1676037725
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1676037725
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1676037725
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1676037725
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1676037725
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1676037725
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1676037725
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1676037725
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1676037725
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1676037725
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1676037725
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1676037725
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1676037725
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1676037725
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1676037725
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1676037725
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1676037725
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1676037725
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1676037725
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1676037725
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1676037725
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1676037725
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1676037725
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1676037725
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1676037725
transform 1 0 19136 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1676037725
transform 1 0 24288 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1676037725
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1676037725
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1676037725
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1676037725
transform 1 0 21712 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1676037725
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1676037725
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1676037725
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1676037725
transform 1 0 19136 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1676037725
transform 1 0 24288 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1676037725
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1676037725
transform 1 0 11408 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1676037725
transform 1 0 16560 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1676037725
transform 1 0 21712 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1676037725
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1676037725
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1676037725
transform 1 0 13984 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1676037725
transform 1 0 19136 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1676037725
transform 1 0 24288 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1676037725
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1676037725
transform 1 0 11408 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1676037725
transform 1 0 16560 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1676037725
transform 1 0 21712 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1676037725
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1676037725
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1676037725
transform 1 0 13984 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1676037725
transform 1 0 19136 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1676037725
transform 1 0 24288 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1676037725
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1676037725
transform 1 0 11408 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1676037725
transform 1 0 16560 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1676037725
transform 1 0 21712 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1676037725
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1676037725
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1676037725
transform 1 0 13984 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1676037725
transform 1 0 19136 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1676037725
transform 1 0 24288 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1676037725
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1676037725
transform 1 0 11408 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1676037725
transform 1 0 16560 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1676037725
transform 1 0 21712 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1676037725
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1676037725
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1676037725
transform 1 0 13984 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1676037725
transform 1 0 19136 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1676037725
transform 1 0 24288 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1676037725
transform 1 0 3680 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1676037725
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1676037725
transform 1 0 8832 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1676037725
transform 1 0 11408 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1676037725
transform 1 0 13984 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1676037725
transform 1 0 16560 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1676037725
transform 1 0 19136 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1676037725
transform 1 0 21712 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1676037725
transform 1 0 24288 0 -1 54400
box -38 -48 130 592
<< labels >>
flabel metal4 s 7944 2128 8264 54448 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 17944 2128 18264 54448 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2944 2128 3264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 12944 2128 13264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 22944 2128 23264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 54952 800 55072 0 FreeSans 480 0 0 0 ccff_head
port 2 nsew signal input
flabel metal3 s 0 1776 800 1896 0 FreeSans 480 0 0 0 ccff_head_0
port 3 nsew signal input
flabel metal3 s 26200 4224 27000 4344 0 FreeSans 480 0 0 0 ccff_tail
port 4 nsew signal tristate
flabel metal2 s 938 56200 994 57000 0 FreeSans 224 90 0 0 ccff_tail_0
port 5 nsew signal tristate
flabel metal3 s 26200 25304 27000 25424 0 FreeSans 480 0 0 0 chanx_right_in[0]
port 6 nsew signal input
flabel metal3 s 26200 32104 27000 32224 0 FreeSans 480 0 0 0 chanx_right_in[10]
port 7 nsew signal input
flabel metal3 s 26200 32784 27000 32904 0 FreeSans 480 0 0 0 chanx_right_in[11]
port 8 nsew signal input
flabel metal3 s 26200 33464 27000 33584 0 FreeSans 480 0 0 0 chanx_right_in[12]
port 9 nsew signal input
flabel metal3 s 26200 34144 27000 34264 0 FreeSans 480 0 0 0 chanx_right_in[13]
port 10 nsew signal input
flabel metal3 s 26200 34824 27000 34944 0 FreeSans 480 0 0 0 chanx_right_in[14]
port 11 nsew signal input
flabel metal3 s 26200 35504 27000 35624 0 FreeSans 480 0 0 0 chanx_right_in[15]
port 12 nsew signal input
flabel metal3 s 26200 36184 27000 36304 0 FreeSans 480 0 0 0 chanx_right_in[16]
port 13 nsew signal input
flabel metal3 s 26200 36864 27000 36984 0 FreeSans 480 0 0 0 chanx_right_in[17]
port 14 nsew signal input
flabel metal3 s 26200 37544 27000 37664 0 FreeSans 480 0 0 0 chanx_right_in[18]
port 15 nsew signal input
flabel metal3 s 26200 38224 27000 38344 0 FreeSans 480 0 0 0 chanx_right_in[19]
port 16 nsew signal input
flabel metal3 s 26200 25984 27000 26104 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 17 nsew signal input
flabel metal3 s 26200 38904 27000 39024 0 FreeSans 480 0 0 0 chanx_right_in[20]
port 18 nsew signal input
flabel metal3 s 26200 39584 27000 39704 0 FreeSans 480 0 0 0 chanx_right_in[21]
port 19 nsew signal input
flabel metal3 s 26200 40264 27000 40384 0 FreeSans 480 0 0 0 chanx_right_in[22]
port 20 nsew signal input
flabel metal3 s 26200 40944 27000 41064 0 FreeSans 480 0 0 0 chanx_right_in[23]
port 21 nsew signal input
flabel metal3 s 26200 41624 27000 41744 0 FreeSans 480 0 0 0 chanx_right_in[24]
port 22 nsew signal input
flabel metal3 s 26200 42304 27000 42424 0 FreeSans 480 0 0 0 chanx_right_in[25]
port 23 nsew signal input
flabel metal3 s 26200 42984 27000 43104 0 FreeSans 480 0 0 0 chanx_right_in[26]
port 24 nsew signal input
flabel metal3 s 26200 43664 27000 43784 0 FreeSans 480 0 0 0 chanx_right_in[27]
port 25 nsew signal input
flabel metal3 s 26200 44344 27000 44464 0 FreeSans 480 0 0 0 chanx_right_in[28]
port 26 nsew signal input
flabel metal3 s 26200 45024 27000 45144 0 FreeSans 480 0 0 0 chanx_right_in[29]
port 27 nsew signal input
flabel metal3 s 26200 26664 27000 26784 0 FreeSans 480 0 0 0 chanx_right_in[2]
port 28 nsew signal input
flabel metal3 s 26200 27344 27000 27464 0 FreeSans 480 0 0 0 chanx_right_in[3]
port 29 nsew signal input
flabel metal3 s 26200 28024 27000 28144 0 FreeSans 480 0 0 0 chanx_right_in[4]
port 30 nsew signal input
flabel metal3 s 26200 28704 27000 28824 0 FreeSans 480 0 0 0 chanx_right_in[5]
port 31 nsew signal input
flabel metal3 s 26200 29384 27000 29504 0 FreeSans 480 0 0 0 chanx_right_in[6]
port 32 nsew signal input
flabel metal3 s 26200 30064 27000 30184 0 FreeSans 480 0 0 0 chanx_right_in[7]
port 33 nsew signal input
flabel metal3 s 26200 30744 27000 30864 0 FreeSans 480 0 0 0 chanx_right_in[8]
port 34 nsew signal input
flabel metal3 s 26200 31424 27000 31544 0 FreeSans 480 0 0 0 chanx_right_in[9]
port 35 nsew signal input
flabel metal3 s 26200 4904 27000 5024 0 FreeSans 480 0 0 0 chanx_right_out[0]
port 36 nsew signal tristate
flabel metal3 s 26200 11704 27000 11824 0 FreeSans 480 0 0 0 chanx_right_out[10]
port 37 nsew signal tristate
flabel metal3 s 26200 12384 27000 12504 0 FreeSans 480 0 0 0 chanx_right_out[11]
port 38 nsew signal tristate
flabel metal3 s 26200 13064 27000 13184 0 FreeSans 480 0 0 0 chanx_right_out[12]
port 39 nsew signal tristate
flabel metal3 s 26200 13744 27000 13864 0 FreeSans 480 0 0 0 chanx_right_out[13]
port 40 nsew signal tristate
flabel metal3 s 26200 14424 27000 14544 0 FreeSans 480 0 0 0 chanx_right_out[14]
port 41 nsew signal tristate
flabel metal3 s 26200 15104 27000 15224 0 FreeSans 480 0 0 0 chanx_right_out[15]
port 42 nsew signal tristate
flabel metal3 s 26200 15784 27000 15904 0 FreeSans 480 0 0 0 chanx_right_out[16]
port 43 nsew signal tristate
flabel metal3 s 26200 16464 27000 16584 0 FreeSans 480 0 0 0 chanx_right_out[17]
port 44 nsew signal tristate
flabel metal3 s 26200 17144 27000 17264 0 FreeSans 480 0 0 0 chanx_right_out[18]
port 45 nsew signal tristate
flabel metal3 s 26200 17824 27000 17944 0 FreeSans 480 0 0 0 chanx_right_out[19]
port 46 nsew signal tristate
flabel metal3 s 26200 5584 27000 5704 0 FreeSans 480 0 0 0 chanx_right_out[1]
port 47 nsew signal tristate
flabel metal3 s 26200 18504 27000 18624 0 FreeSans 480 0 0 0 chanx_right_out[20]
port 48 nsew signal tristate
flabel metal3 s 26200 19184 27000 19304 0 FreeSans 480 0 0 0 chanx_right_out[21]
port 49 nsew signal tristate
flabel metal3 s 26200 19864 27000 19984 0 FreeSans 480 0 0 0 chanx_right_out[22]
port 50 nsew signal tristate
flabel metal3 s 26200 20544 27000 20664 0 FreeSans 480 0 0 0 chanx_right_out[23]
port 51 nsew signal tristate
flabel metal3 s 26200 21224 27000 21344 0 FreeSans 480 0 0 0 chanx_right_out[24]
port 52 nsew signal tristate
flabel metal3 s 26200 21904 27000 22024 0 FreeSans 480 0 0 0 chanx_right_out[25]
port 53 nsew signal tristate
flabel metal3 s 26200 22584 27000 22704 0 FreeSans 480 0 0 0 chanx_right_out[26]
port 54 nsew signal tristate
flabel metal3 s 26200 23264 27000 23384 0 FreeSans 480 0 0 0 chanx_right_out[27]
port 55 nsew signal tristate
flabel metal3 s 26200 23944 27000 24064 0 FreeSans 480 0 0 0 chanx_right_out[28]
port 56 nsew signal tristate
flabel metal3 s 26200 24624 27000 24744 0 FreeSans 480 0 0 0 chanx_right_out[29]
port 57 nsew signal tristate
flabel metal3 s 26200 6264 27000 6384 0 FreeSans 480 0 0 0 chanx_right_out[2]
port 58 nsew signal tristate
flabel metal3 s 26200 6944 27000 7064 0 FreeSans 480 0 0 0 chanx_right_out[3]
port 59 nsew signal tristate
flabel metal3 s 26200 7624 27000 7744 0 FreeSans 480 0 0 0 chanx_right_out[4]
port 60 nsew signal tristate
flabel metal3 s 26200 8304 27000 8424 0 FreeSans 480 0 0 0 chanx_right_out[5]
port 61 nsew signal tristate
flabel metal3 s 26200 8984 27000 9104 0 FreeSans 480 0 0 0 chanx_right_out[6]
port 62 nsew signal tristate
flabel metal3 s 26200 9664 27000 9784 0 FreeSans 480 0 0 0 chanx_right_out[7]
port 63 nsew signal tristate
flabel metal3 s 26200 10344 27000 10464 0 FreeSans 480 0 0 0 chanx_right_out[8]
port 64 nsew signal tristate
flabel metal3 s 26200 11024 27000 11144 0 FreeSans 480 0 0 0 chanx_right_out[9]
port 65 nsew signal tristate
flabel metal2 s 1122 0 1178 800 0 FreeSans 224 90 0 0 chany_bottom_in[0]
port 66 nsew signal input
flabel metal2 s 4802 0 4858 800 0 FreeSans 224 90 0 0 chany_bottom_in[10]
port 67 nsew signal input
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 chany_bottom_in[11]
port 68 nsew signal input
flabel metal2 s 5538 0 5594 800 0 FreeSans 224 90 0 0 chany_bottom_in[12]
port 69 nsew signal input
flabel metal2 s 5906 0 5962 800 0 FreeSans 224 90 0 0 chany_bottom_in[13]
port 70 nsew signal input
flabel metal2 s 6274 0 6330 800 0 FreeSans 224 90 0 0 chany_bottom_in[14]
port 71 nsew signal input
flabel metal2 s 6642 0 6698 800 0 FreeSans 224 90 0 0 chany_bottom_in[15]
port 72 nsew signal input
flabel metal2 s 7010 0 7066 800 0 FreeSans 224 90 0 0 chany_bottom_in[16]
port 73 nsew signal input
flabel metal2 s 7378 0 7434 800 0 FreeSans 224 90 0 0 chany_bottom_in[17]
port 74 nsew signal input
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 chany_bottom_in[18]
port 75 nsew signal input
flabel metal2 s 8114 0 8170 800 0 FreeSans 224 90 0 0 chany_bottom_in[19]
port 76 nsew signal input
flabel metal2 s 1490 0 1546 800 0 FreeSans 224 90 0 0 chany_bottom_in[1]
port 77 nsew signal input
flabel metal2 s 8482 0 8538 800 0 FreeSans 224 90 0 0 chany_bottom_in[20]
port 78 nsew signal input
flabel metal2 s 8850 0 8906 800 0 FreeSans 224 90 0 0 chany_bottom_in[21]
port 79 nsew signal input
flabel metal2 s 9218 0 9274 800 0 FreeSans 224 90 0 0 chany_bottom_in[22]
port 80 nsew signal input
flabel metal2 s 9586 0 9642 800 0 FreeSans 224 90 0 0 chany_bottom_in[23]
port 81 nsew signal input
flabel metal2 s 9954 0 10010 800 0 FreeSans 224 90 0 0 chany_bottom_in[24]
port 82 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 chany_bottom_in[25]
port 83 nsew signal input
flabel metal2 s 10690 0 10746 800 0 FreeSans 224 90 0 0 chany_bottom_in[26]
port 84 nsew signal input
flabel metal2 s 11058 0 11114 800 0 FreeSans 224 90 0 0 chany_bottom_in[27]
port 85 nsew signal input
flabel metal2 s 11426 0 11482 800 0 FreeSans 224 90 0 0 chany_bottom_in[28]
port 86 nsew signal input
flabel metal2 s 11794 0 11850 800 0 FreeSans 224 90 0 0 chany_bottom_in[29]
port 87 nsew signal input
flabel metal2 s 1858 0 1914 800 0 FreeSans 224 90 0 0 chany_bottom_in[2]
port 88 nsew signal input
flabel metal2 s 2226 0 2282 800 0 FreeSans 224 90 0 0 chany_bottom_in[3]
port 89 nsew signal input
flabel metal2 s 2594 0 2650 800 0 FreeSans 224 90 0 0 chany_bottom_in[4]
port 90 nsew signal input
flabel metal2 s 2962 0 3018 800 0 FreeSans 224 90 0 0 chany_bottom_in[5]
port 91 nsew signal input
flabel metal2 s 3330 0 3386 800 0 FreeSans 224 90 0 0 chany_bottom_in[6]
port 92 nsew signal input
flabel metal2 s 3698 0 3754 800 0 FreeSans 224 90 0 0 chany_bottom_in[7]
port 93 nsew signal input
flabel metal2 s 4066 0 4122 800 0 FreeSans 224 90 0 0 chany_bottom_in[8]
port 94 nsew signal input
flabel metal2 s 4434 0 4490 800 0 FreeSans 224 90 0 0 chany_bottom_in[9]
port 95 nsew signal input
flabel metal2 s 12162 0 12218 800 0 FreeSans 224 90 0 0 chany_bottom_out[0]
port 96 nsew signal tristate
flabel metal2 s 15842 0 15898 800 0 FreeSans 224 90 0 0 chany_bottom_out[10]
port 97 nsew signal tristate
flabel metal2 s 16210 0 16266 800 0 FreeSans 224 90 0 0 chany_bottom_out[11]
port 98 nsew signal tristate
flabel metal2 s 16578 0 16634 800 0 FreeSans 224 90 0 0 chany_bottom_out[12]
port 99 nsew signal tristate
flabel metal2 s 16946 0 17002 800 0 FreeSans 224 90 0 0 chany_bottom_out[13]
port 100 nsew signal tristate
flabel metal2 s 17314 0 17370 800 0 FreeSans 224 90 0 0 chany_bottom_out[14]
port 101 nsew signal tristate
flabel metal2 s 17682 0 17738 800 0 FreeSans 224 90 0 0 chany_bottom_out[15]
port 102 nsew signal tristate
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 chany_bottom_out[16]
port 103 nsew signal tristate
flabel metal2 s 18418 0 18474 800 0 FreeSans 224 90 0 0 chany_bottom_out[17]
port 104 nsew signal tristate
flabel metal2 s 18786 0 18842 800 0 FreeSans 224 90 0 0 chany_bottom_out[18]
port 105 nsew signal tristate
flabel metal2 s 19154 0 19210 800 0 FreeSans 224 90 0 0 chany_bottom_out[19]
port 106 nsew signal tristate
flabel metal2 s 12530 0 12586 800 0 FreeSans 224 90 0 0 chany_bottom_out[1]
port 107 nsew signal tristate
flabel metal2 s 19522 0 19578 800 0 FreeSans 224 90 0 0 chany_bottom_out[20]
port 108 nsew signal tristate
flabel metal2 s 19890 0 19946 800 0 FreeSans 224 90 0 0 chany_bottom_out[21]
port 109 nsew signal tristate
flabel metal2 s 20258 0 20314 800 0 FreeSans 224 90 0 0 chany_bottom_out[22]
port 110 nsew signal tristate
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 chany_bottom_out[23]
port 111 nsew signal tristate
flabel metal2 s 20994 0 21050 800 0 FreeSans 224 90 0 0 chany_bottom_out[24]
port 112 nsew signal tristate
flabel metal2 s 21362 0 21418 800 0 FreeSans 224 90 0 0 chany_bottom_out[25]
port 113 nsew signal tristate
flabel metal2 s 21730 0 21786 800 0 FreeSans 224 90 0 0 chany_bottom_out[26]
port 114 nsew signal tristate
flabel metal2 s 22098 0 22154 800 0 FreeSans 224 90 0 0 chany_bottom_out[27]
port 115 nsew signal tristate
flabel metal2 s 22466 0 22522 800 0 FreeSans 224 90 0 0 chany_bottom_out[28]
port 116 nsew signal tristate
flabel metal2 s 22834 0 22890 800 0 FreeSans 224 90 0 0 chany_bottom_out[29]
port 117 nsew signal tristate
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 chany_bottom_out[2]
port 118 nsew signal tristate
flabel metal2 s 13266 0 13322 800 0 FreeSans 224 90 0 0 chany_bottom_out[3]
port 119 nsew signal tristate
flabel metal2 s 13634 0 13690 800 0 FreeSans 224 90 0 0 chany_bottom_out[4]
port 120 nsew signal tristate
flabel metal2 s 14002 0 14058 800 0 FreeSans 224 90 0 0 chany_bottom_out[5]
port 121 nsew signal tristate
flabel metal2 s 14370 0 14426 800 0 FreeSans 224 90 0 0 chany_bottom_out[6]
port 122 nsew signal tristate
flabel metal2 s 14738 0 14794 800 0 FreeSans 224 90 0 0 chany_bottom_out[7]
port 123 nsew signal tristate
flabel metal2 s 15106 0 15162 800 0 FreeSans 224 90 0 0 chany_bottom_out[8]
port 124 nsew signal tristate
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 chany_bottom_out[9]
port 125 nsew signal tristate
flabel metal2 s 12346 56200 12402 57000 0 FreeSans 224 90 0 0 chany_top_in_0[0]
port 126 nsew signal input
flabel metal2 s 16026 56200 16082 57000 0 FreeSans 224 90 0 0 chany_top_in_0[10]
port 127 nsew signal input
flabel metal2 s 16394 56200 16450 57000 0 FreeSans 224 90 0 0 chany_top_in_0[11]
port 128 nsew signal input
flabel metal2 s 16762 56200 16818 57000 0 FreeSans 224 90 0 0 chany_top_in_0[12]
port 129 nsew signal input
flabel metal2 s 17130 56200 17186 57000 0 FreeSans 224 90 0 0 chany_top_in_0[13]
port 130 nsew signal input
flabel metal2 s 17498 56200 17554 57000 0 FreeSans 224 90 0 0 chany_top_in_0[14]
port 131 nsew signal input
flabel metal2 s 17866 56200 17922 57000 0 FreeSans 224 90 0 0 chany_top_in_0[15]
port 132 nsew signal input
flabel metal2 s 18234 56200 18290 57000 0 FreeSans 224 90 0 0 chany_top_in_0[16]
port 133 nsew signal input
flabel metal2 s 18602 56200 18658 57000 0 FreeSans 224 90 0 0 chany_top_in_0[17]
port 134 nsew signal input
flabel metal2 s 18970 56200 19026 57000 0 FreeSans 224 90 0 0 chany_top_in_0[18]
port 135 nsew signal input
flabel metal2 s 19338 56200 19394 57000 0 FreeSans 224 90 0 0 chany_top_in_0[19]
port 136 nsew signal input
flabel metal2 s 12714 56200 12770 57000 0 FreeSans 224 90 0 0 chany_top_in_0[1]
port 137 nsew signal input
flabel metal2 s 19706 56200 19762 57000 0 FreeSans 224 90 0 0 chany_top_in_0[20]
port 138 nsew signal input
flabel metal2 s 20074 56200 20130 57000 0 FreeSans 224 90 0 0 chany_top_in_0[21]
port 139 nsew signal input
flabel metal2 s 20442 56200 20498 57000 0 FreeSans 224 90 0 0 chany_top_in_0[22]
port 140 nsew signal input
flabel metal2 s 20810 56200 20866 57000 0 FreeSans 224 90 0 0 chany_top_in_0[23]
port 141 nsew signal input
flabel metal2 s 21178 56200 21234 57000 0 FreeSans 224 90 0 0 chany_top_in_0[24]
port 142 nsew signal input
flabel metal2 s 21546 56200 21602 57000 0 FreeSans 224 90 0 0 chany_top_in_0[25]
port 143 nsew signal input
flabel metal2 s 21914 56200 21970 57000 0 FreeSans 224 90 0 0 chany_top_in_0[26]
port 144 nsew signal input
flabel metal2 s 22282 56200 22338 57000 0 FreeSans 224 90 0 0 chany_top_in_0[27]
port 145 nsew signal input
flabel metal2 s 22650 56200 22706 57000 0 FreeSans 224 90 0 0 chany_top_in_0[28]
port 146 nsew signal input
flabel metal2 s 23018 56200 23074 57000 0 FreeSans 224 90 0 0 chany_top_in_0[29]
port 147 nsew signal input
flabel metal2 s 13082 56200 13138 57000 0 FreeSans 224 90 0 0 chany_top_in_0[2]
port 148 nsew signal input
flabel metal2 s 13450 56200 13506 57000 0 FreeSans 224 90 0 0 chany_top_in_0[3]
port 149 nsew signal input
flabel metal2 s 13818 56200 13874 57000 0 FreeSans 224 90 0 0 chany_top_in_0[4]
port 150 nsew signal input
flabel metal2 s 14186 56200 14242 57000 0 FreeSans 224 90 0 0 chany_top_in_0[5]
port 151 nsew signal input
flabel metal2 s 14554 56200 14610 57000 0 FreeSans 224 90 0 0 chany_top_in_0[6]
port 152 nsew signal input
flabel metal2 s 14922 56200 14978 57000 0 FreeSans 224 90 0 0 chany_top_in_0[7]
port 153 nsew signal input
flabel metal2 s 15290 56200 15346 57000 0 FreeSans 224 90 0 0 chany_top_in_0[8]
port 154 nsew signal input
flabel metal2 s 15658 56200 15714 57000 0 FreeSans 224 90 0 0 chany_top_in_0[9]
port 155 nsew signal input
flabel metal2 s 1306 56200 1362 57000 0 FreeSans 224 90 0 0 chany_top_out_0[0]
port 156 nsew signal tristate
flabel metal2 s 4986 56200 5042 57000 0 FreeSans 224 90 0 0 chany_top_out_0[10]
port 157 nsew signal tristate
flabel metal2 s 5354 56200 5410 57000 0 FreeSans 224 90 0 0 chany_top_out_0[11]
port 158 nsew signal tristate
flabel metal2 s 5722 56200 5778 57000 0 FreeSans 224 90 0 0 chany_top_out_0[12]
port 159 nsew signal tristate
flabel metal2 s 6090 56200 6146 57000 0 FreeSans 224 90 0 0 chany_top_out_0[13]
port 160 nsew signal tristate
flabel metal2 s 6458 56200 6514 57000 0 FreeSans 224 90 0 0 chany_top_out_0[14]
port 161 nsew signal tristate
flabel metal2 s 6826 56200 6882 57000 0 FreeSans 224 90 0 0 chany_top_out_0[15]
port 162 nsew signal tristate
flabel metal2 s 7194 56200 7250 57000 0 FreeSans 224 90 0 0 chany_top_out_0[16]
port 163 nsew signal tristate
flabel metal2 s 7562 56200 7618 57000 0 FreeSans 224 90 0 0 chany_top_out_0[17]
port 164 nsew signal tristate
flabel metal2 s 7930 56200 7986 57000 0 FreeSans 224 90 0 0 chany_top_out_0[18]
port 165 nsew signal tristate
flabel metal2 s 8298 56200 8354 57000 0 FreeSans 224 90 0 0 chany_top_out_0[19]
port 166 nsew signal tristate
flabel metal2 s 1674 56200 1730 57000 0 FreeSans 224 90 0 0 chany_top_out_0[1]
port 167 nsew signal tristate
flabel metal2 s 8666 56200 8722 57000 0 FreeSans 224 90 0 0 chany_top_out_0[20]
port 168 nsew signal tristate
flabel metal2 s 9034 56200 9090 57000 0 FreeSans 224 90 0 0 chany_top_out_0[21]
port 169 nsew signal tristate
flabel metal2 s 9402 56200 9458 57000 0 FreeSans 224 90 0 0 chany_top_out_0[22]
port 170 nsew signal tristate
flabel metal2 s 9770 56200 9826 57000 0 FreeSans 224 90 0 0 chany_top_out_0[23]
port 171 nsew signal tristate
flabel metal2 s 10138 56200 10194 57000 0 FreeSans 224 90 0 0 chany_top_out_0[24]
port 172 nsew signal tristate
flabel metal2 s 10506 56200 10562 57000 0 FreeSans 224 90 0 0 chany_top_out_0[25]
port 173 nsew signal tristate
flabel metal2 s 10874 56200 10930 57000 0 FreeSans 224 90 0 0 chany_top_out_0[26]
port 174 nsew signal tristate
flabel metal2 s 11242 56200 11298 57000 0 FreeSans 224 90 0 0 chany_top_out_0[27]
port 175 nsew signal tristate
flabel metal2 s 11610 56200 11666 57000 0 FreeSans 224 90 0 0 chany_top_out_0[28]
port 176 nsew signal tristate
flabel metal2 s 11978 56200 12034 57000 0 FreeSans 224 90 0 0 chany_top_out_0[29]
port 177 nsew signal tristate
flabel metal2 s 2042 56200 2098 57000 0 FreeSans 224 90 0 0 chany_top_out_0[2]
port 178 nsew signal tristate
flabel metal2 s 2410 56200 2466 57000 0 FreeSans 224 90 0 0 chany_top_out_0[3]
port 179 nsew signal tristate
flabel metal2 s 2778 56200 2834 57000 0 FreeSans 224 90 0 0 chany_top_out_0[4]
port 180 nsew signal tristate
flabel metal2 s 3146 56200 3202 57000 0 FreeSans 224 90 0 0 chany_top_out_0[5]
port 181 nsew signal tristate
flabel metal2 s 3514 56200 3570 57000 0 FreeSans 224 90 0 0 chany_top_out_0[6]
port 182 nsew signal tristate
flabel metal2 s 3882 56200 3938 57000 0 FreeSans 224 90 0 0 chany_top_out_0[7]
port 183 nsew signal tristate
flabel metal2 s 4250 56200 4306 57000 0 FreeSans 224 90 0 0 chany_top_out_0[8]
port 184 nsew signal tristate
flabel metal2 s 4618 56200 4674 57000 0 FreeSans 224 90 0 0 chany_top_out_0[9]
port 185 nsew signal tristate
flabel metal3 s 0 13336 800 13456 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_dir[0]
port 186 nsew signal tristate
flabel metal3 s 0 15648 800 15768 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_dir[1]
port 187 nsew signal tristate
flabel metal3 s 0 17960 800 18080 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_dir[2]
port 188 nsew signal tristate
flabel metal3 s 0 20272 800 20392 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_dir[3]
port 189 nsew signal tristate
flabel metal3 s 0 31832 800 31952 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_in[0]
port 190 nsew signal input
flabel metal3 s 0 34144 800 34264 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_in[1]
port 191 nsew signal input
flabel metal3 s 0 36456 800 36576 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_in[2]
port 192 nsew signal input
flabel metal3 s 0 38768 800 38888 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_in[3]
port 193 nsew signal input
flabel metal3 s 0 22584 800 22704 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_out[0]
port 194 nsew signal tristate
flabel metal3 s 0 24896 800 25016 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_out[1]
port 195 nsew signal tristate
flabel metal3 s 0 27208 800 27328 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_out[2]
port 196 nsew signal tristate
flabel metal3 s 0 29520 800 29640 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_out[3]
port 197 nsew signal tristate
flabel metal3 s 0 41080 800 41200 0 FreeSans 480 0 0 0 isol_n
port 198 nsew signal input
flabel metal2 s 23202 0 23258 800 0 FreeSans 224 90 0 0 prog_clk
port 199 nsew signal input
flabel metal2 s 23570 0 23626 800 0 FreeSans 224 90 0 0 prog_reset_bottom_in
port 200 nsew signal input
flabel metal2 s 23938 0 23994 800 0 FreeSans 224 90 0 0 prog_reset_bottom_out
port 201 nsew signal tristate
flabel metal3 s 0 43392 800 43512 0 FreeSans 480 0 0 0 prog_reset_left_in
port 202 nsew signal input
flabel metal3 s 26200 45704 27000 45824 0 FreeSans 480 0 0 0 prog_reset_right_out
port 203 nsew signal tristate
flabel metal2 s 24490 56200 24546 57000 0 FreeSans 224 90 0 0 prog_reset_top_in
port 204 nsew signal input
flabel metal2 s 24122 56200 24178 57000 0 FreeSans 224 90 0 0 prog_reset_top_out
port 205 nsew signal tristate
flabel metal2 s 24306 0 24362 800 0 FreeSans 224 90 0 0 reset_bottom_in
port 206 nsew signal input
flabel metal2 s 24674 0 24730 800 0 FreeSans 224 90 0 0 reset_bottom_out
port 207 nsew signal tristate
flabel metal3 s 26200 46384 27000 46504 0 FreeSans 480 0 0 0 reset_right_in
port 208 nsew signal input
flabel metal2 s 25226 56200 25282 57000 0 FreeSans 224 90 0 0 reset_top_in
port 209 nsew signal input
flabel metal2 s 24858 56200 24914 57000 0 FreeSans 224 90 0 0 reset_top_out
port 210 nsew signal tristate
flabel metal3 s 26200 47064 27000 47184 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
port 211 nsew signal input
flabel metal3 s 26200 47744 27000 47864 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_
port 212 nsew signal input
flabel metal3 s 26200 48424 27000 48544 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
port 213 nsew signal input
flabel metal3 s 26200 49104 27000 49224 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_
port 214 nsew signal input
flabel metal3 s 26200 49784 27000 49904 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
port 215 nsew signal input
flabel metal3 s 26200 50464 27000 50584 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_
port 216 nsew signal input
flabel metal3 s 26200 51144 27000 51264 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_
port 217 nsew signal input
flabel metal3 s 26200 51824 27000 51944 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_
port 218 nsew signal input
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_0__pin_inpad_0_
port 219 nsew signal tristate
flabel metal3 s 0 6400 800 6520 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_1__pin_inpad_0_
port 220 nsew signal tristate
flabel metal3 s 0 8712 800 8832 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_2__pin_inpad_0_
port 221 nsew signal tristate
flabel metal3 s 0 11024 800 11144 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_3__pin_inpad_0_
port 222 nsew signal tristate
flabel metal2 s 25042 0 25098 800 0 FreeSans 224 90 0 0 test_enable_bottom_in
port 223 nsew signal input
flabel metal2 s 25410 0 25466 800 0 FreeSans 224 90 0 0 test_enable_bottom_out
port 224 nsew signal tristate
flabel metal3 s 26200 52504 27000 52624 0 FreeSans 480 0 0 0 test_enable_right_in
port 225 nsew signal input
flabel metal2 s 25962 56200 26018 57000 0 FreeSans 224 90 0 0 test_enable_top_in
port 226 nsew signal input
flabel metal2 s 25594 56200 25650 57000 0 FreeSans 224 90 0 0 test_enable_top_out
port 227 nsew signal tristate
flabel metal3 s 0 45704 800 45824 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
port 228 nsew signal input
flabel metal3 s 0 48016 800 48136 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
port 229 nsew signal input
flabel metal3 s 0 50328 800 50448 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
port 230 nsew signal input
flabel metal3 s 0 52640 800 52760 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
port 231 nsew signal input
rlabel metal1 13478 54400 13478 54400 0 VGND
rlabel metal1 13478 53856 13478 53856 0 VPWR
rlabel metal1 5014 23494 5014 23494 0 cby_0__1_.cby_0__1_.ccff_tail
rlabel metal1 4232 23290 4232 23290 0 cby_0__1_.cby_0__1_.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_
rlabel metal1 4094 22542 4094 22542 0 cby_0__1_.cby_0__1_.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_
rlabel metal2 4002 20196 4002 20196 0 cby_0__1_.cby_0__1_.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_
rlabel metal2 3450 21148 3450 21148 0 cby_0__1_.cby_0__1_.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_
rlabel metal1 6854 20774 6854 20774 0 cby_0__1_.cby_0__1_.mem_right_ipin_0.ccff_tail
rlabel metal2 12604 12036 12604 12036 0 cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[0\]
rlabel metal1 10074 18054 10074 18054 0 cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[1\]
rlabel metal1 5428 20026 5428 20026 0 cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[2\]
rlabel metal1 6900 14246 6900 14246 0 cby_0__1_.cby_0__1_.mem_right_ipin_1.ccff_tail
rlabel metal1 15226 17714 15226 17714 0 cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[0\]
rlabel metal1 13662 14858 13662 14858 0 cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[1\]
rlabel metal2 8878 14620 8878 14620 0 cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[2\]
rlabel metal1 5842 17136 5842 17136 0 cby_0__1_.cby_0__1_.mem_right_ipin_2.ccff_tail
rlabel metal1 15042 12274 15042 12274 0 cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[0\]
rlabel metal1 7544 15402 7544 15402 0 cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[1\]
rlabel metal1 6440 17578 6440 17578 0 cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[2\]
rlabel metal1 13248 18190 13248 18190 0 cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[0\]
rlabel metal1 8234 21012 8234 21012 0 cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[1\]
rlabel metal1 7544 21590 7544 21590 0 cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[2\]
rlabel metal2 12742 15606 12742 15606 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 7406 21760 7406 21760 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 6532 21658 6532 21658 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 10534 17102 10534 17102 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 13662 19414 13662 19414 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 12558 22950 12558 22950 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 9522 18938 9522 18938 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 9890 17306 9890 17306 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 9982 19822 9982 19822 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 8004 20298 8004 20298 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 8694 21998 8694 21998 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal2 9154 20672 9154 20672 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 14260 14994 14260 14994 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 8556 16218 8556 16218 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 7038 16218 7038 16218 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 14168 15130 14168 15130 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 14306 19754 14306 19754 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 13616 17578 13616 17578 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 10488 21862 10488 21862 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 10902 15572 10902 15572 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 12558 16864 12558 16864 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 9430 14586 9430 14586 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 10028 16490 10028 16490 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 9246 15946 9246 15946 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 14766 11322 14766 11322 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 6348 17306 6348 17306 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 4738 17306 4738 17306 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 13892 12410 13892 12410 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 13202 21352 13202 21352 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 12098 18088 12098 18088 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 8418 19822 8418 19822 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 11822 14960 11822 14960 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 11086 17306 11086 17306 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 7682 17306 7682 17306 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal2 8786 16524 8786 16524 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 7268 17034 7268 17034 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal2 11638 17000 11638 17000 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 5888 22202 5888 22202 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 4048 21522 4048 21522 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal2 12466 18870 12466 18870 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 13110 19618 13110 19618 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 11178 20842 11178 20842 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 9798 16422 9798 16422 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 9936 19482 9936 19482 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 9246 21114 9246 21114 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 7498 21114 7498 21114 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 7544 23494 7544 23494 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 6716 22610 6716 22610 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 3634 24718 3634 24718 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.ccff_tail
rlabel metal1 2254 22032 2254 22032 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
rlabel metal1 2438 26010 2438 26010 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_out
rlabel via1 3519 27098 3519 27098 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 4232 20502 4232 20502 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.ccff_tail
rlabel metal1 2806 19822 2806 19822 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
rlabel metal2 2254 23766 2254 23766 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_out
rlabel metal1 3979 26010 3979 26010 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 5704 20230 5704 20230 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.ccff_tail
rlabel metal1 2898 21454 2898 21454 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
rlabel metal2 2162 22134 2162 22134 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_out
rlabel metal1 4071 24038 4071 24038 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal2 4094 16762 4094 16762 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
rlabel metal2 2898 21556 2898 21556 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_out
rlabel metal1 3979 22746 3979 22746 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 2438 53210 2438 53210 0 ccff_head
rlabel metal1 2576 3502 2576 3502 0 ccff_head_0
rlabel metal2 23414 5321 23414 5321 0 ccff_tail
rlabel metal1 2668 52666 2668 52666 0 ccff_tail_0
rlabel metal2 25346 23987 25346 23987 0 chanx_right_in[0]
rlabel metal2 25346 32283 25346 32283 0 chanx_right_in[10]
rlabel via2 25346 32861 25346 32861 0 chanx_right_in[11]
rlabel metal2 25346 33677 25346 33677 0 chanx_right_in[12]
rlabel metal1 25392 35054 25392 35054 0 chanx_right_in[13]
rlabel metal2 25346 35513 25346 35513 0 chanx_right_in[14]
rlabel metal1 25070 36754 25070 36754 0 chanx_right_in[15]
rlabel metal2 25346 36737 25346 36737 0 chanx_right_in[16]
rlabel metal1 24748 37162 24748 37162 0 chanx_right_in[17]
rlabel metal1 25392 38318 25392 38318 0 chanx_right_in[18]
rlabel metal1 24840 40358 24840 40358 0 chanx_right_in[19]
rlabel metal1 21252 25874 21252 25874 0 chanx_right_in[1]
rlabel metal2 25346 39457 25346 39457 0 chanx_right_in[20]
rlabel metal1 24518 39950 24518 39950 0 chanx_right_in[21]
rlabel metal1 23506 39610 23506 39610 0 chanx_right_in[22]
rlabel metal3 25584 41004 25584 41004 0 chanx_right_in[23]
rlabel metal2 25530 42109 25530 42109 0 chanx_right_in[24]
rlabel metal2 25346 43605 25346 43605 0 chanx_right_in[25]
rlabel metal2 25530 43333 25530 43333 0 chanx_right_in[26]
rlabel metal1 25070 45866 25070 45866 0 chanx_right_in[27]
rlabel metal1 24932 43962 24932 43962 0 chanx_right_in[28]
rlabel metal2 23874 45713 23874 45713 0 chanx_right_in[29]
rlabel metal1 24610 28594 24610 28594 0 chanx_right_in[2]
rlabel metal2 25438 27251 25438 27251 0 chanx_right_in[3]
rlabel metal1 24794 28390 24794 28390 0 chanx_right_in[4]
rlabel metal2 24150 28951 24150 28951 0 chanx_right_in[5]
rlabel metal1 25392 28526 25392 28526 0 chanx_right_in[6]
rlabel metal2 25346 29869 25346 29869 0 chanx_right_in[7]
rlabel metal1 25116 31790 25116 31790 0 chanx_right_in[8]
rlabel metal2 25346 31399 25346 31399 0 chanx_right_in[9]
rlabel metal3 25676 11764 25676 11764 0 chanx_right_out[10]
rlabel metal1 24104 12886 24104 12886 0 chanx_right_out[11]
rlabel metal3 25538 13124 25538 13124 0 chanx_right_out[12]
rlabel metal2 24794 13277 24794 13277 0 chanx_right_out[13]
rlabel metal1 24104 15062 24104 15062 0 chanx_right_out[14]
rlabel metal2 25162 14569 25162 14569 0 chanx_right_out[15]
rlabel metal1 24380 15538 24380 15538 0 chanx_right_out[16]
rlabel metal1 23552 16014 23552 16014 0 chanx_right_out[17]
rlabel metal3 25538 17204 25538 17204 0 chanx_right_out[18]
rlabel metal3 25584 17884 25584 17884 0 chanx_right_out[19]
rlabel metal2 24794 5389 24794 5389 0 chanx_right_out[1]
rlabel metal2 23414 18139 23414 18139 0 chanx_right_out[20]
rlabel metal2 22126 19329 22126 19329 0 chanx_right_out[21]
rlabel metal1 23736 19414 23736 19414 0 chanx_right_out[22]
rlabel metal1 24288 19890 24288 19890 0 chanx_right_out[23]
rlabel metal1 24472 19346 24472 19346 0 chanx_right_out[24]
rlabel metal1 24150 22066 24150 22066 0 chanx_right_out[25]
rlabel metal1 24150 23154 24150 23154 0 chanx_right_out[26]
rlabel metal1 23230 23630 23230 23630 0 chanx_right_out[27]
rlabel metal1 24150 24242 24150 24242 0 chanx_right_out[28]
rlabel metal2 25162 24225 25162 24225 0 chanx_right_out[29]
rlabel metal1 24150 6834 24150 6834 0 chanx_right_out[2]
rlabel metal2 24794 6613 24794 6613 0 chanx_right_out[3]
rlabel metal1 24196 7922 24196 7922 0 chanx_right_out[4]
rlabel metal2 24794 7837 24794 7837 0 chanx_right_out[5]
rlabel metal2 25162 8789 25162 8789 0 chanx_right_out[6]
rlabel metal1 24150 10098 24150 10098 0 chanx_right_out[7]
rlabel metal2 24794 9945 24794 9945 0 chanx_right_out[8]
rlabel metal2 24794 10829 24794 10829 0 chanx_right_out[9]
rlabel metal1 1380 4114 1380 4114 0 chany_bottom_in[0]
rlabel metal1 4738 3366 4738 3366 0 chany_bottom_in[10]
rlabel metal1 5290 2278 5290 2278 0 chany_bottom_in[11]
rlabel metal1 5612 3502 5612 3502 0 chany_bottom_in[12]
rlabel metal1 5888 3026 5888 3026 0 chany_bottom_in[13]
rlabel metal1 6348 3502 6348 3502 0 chany_bottom_in[14]
rlabel metal1 6578 2278 6578 2278 0 chany_bottom_in[15]
rlabel metal2 7038 1792 7038 1792 0 chany_bottom_in[16]
rlabel metal1 7314 3366 7314 3366 0 chany_bottom_in[17]
rlabel metal2 7774 1554 7774 1554 0 chany_bottom_in[18]
rlabel metal1 8050 2822 8050 2822 0 chany_bottom_in[19]
rlabel metal2 1518 1792 1518 1792 0 chany_bottom_in[1]
rlabel metal1 8740 2278 8740 2278 0 chany_bottom_in[20]
rlabel metal1 8648 3910 8648 3910 0 chany_bottom_in[21]
rlabel metal1 9292 4114 9292 4114 0 chany_bottom_in[22]
rlabel metal1 9660 2822 9660 2822 0 chany_bottom_in[23]
rlabel metal2 9982 1792 9982 1792 0 chany_bottom_in[24]
rlabel metal1 10764 3026 10764 3026 0 chany_bottom_in[25]
rlabel metal1 11040 3502 11040 3502 0 chany_bottom_in[26]
rlabel metal1 10120 2278 10120 2278 0 chany_bottom_in[27]
rlabel metal1 12006 2414 12006 2414 0 chany_bottom_in[28]
rlabel metal1 12190 2958 12190 2958 0 chany_bottom_in[29]
rlabel metal1 1794 2822 1794 2822 0 chany_bottom_in[2]
rlabel metal1 2070 2414 2070 2414 0 chany_bottom_in[3]
rlabel metal1 3036 2482 3036 2482 0 chany_bottom_in[4]
rlabel metal1 2990 3502 2990 3502 0 chany_bottom_in[5]
rlabel metal1 3128 3026 3128 3026 0 chany_bottom_in[6]
rlabel metal1 3772 3026 3772 3026 0 chany_bottom_in[7]
rlabel metal1 4002 2278 4002 2278 0 chany_bottom_in[8]
rlabel metal1 4370 3026 4370 3026 0 chany_bottom_in[9]
rlabel metal2 12190 1622 12190 1622 0 chany_bottom_out[0]
rlabel metal2 15870 1860 15870 1860 0 chany_bottom_out[10]
rlabel metal2 16238 2404 16238 2404 0 chany_bottom_out[11]
rlabel metal2 16606 1826 16606 1826 0 chany_bottom_out[12]
rlabel metal2 16974 1588 16974 1588 0 chany_bottom_out[13]
rlabel metal2 17342 1792 17342 1792 0 chany_bottom_out[14]
rlabel metal2 17710 2166 17710 2166 0 chany_bottom_out[15]
rlabel metal2 18078 823 18078 823 0 chany_bottom_out[16]
rlabel metal2 18446 823 18446 823 0 chany_bottom_out[17]
rlabel metal2 18814 1792 18814 1792 0 chany_bottom_out[18]
rlabel metal2 19182 2098 19182 2098 0 chany_bottom_out[19]
rlabel metal2 12558 2098 12558 2098 0 chany_bottom_out[1]
rlabel metal2 19550 2948 19550 2948 0 chany_bottom_out[20]
rlabel metal2 19918 1503 19918 1503 0 chany_bottom_out[21]
rlabel metal2 20286 2404 20286 2404 0 chany_bottom_out[22]
rlabel metal2 20654 3254 20654 3254 0 chany_bottom_out[23]
rlabel metal2 21022 1792 21022 1792 0 chany_bottom_out[24]
rlabel metal2 21390 2370 21390 2370 0 chany_bottom_out[25]
rlabel metal2 21758 1775 21758 1775 0 chany_bottom_out[26]
rlabel metal1 22126 6188 22126 6188 0 chany_bottom_out[27]
rlabel metal1 22540 7310 22540 7310 0 chany_bottom_out[28]
rlabel metal2 22034 4862 22034 4862 0 chany_bottom_out[29]
rlabel metal2 12926 1435 12926 1435 0 chany_bottom_out[2]
rlabel metal2 13294 1554 13294 1554 0 chany_bottom_out[3]
rlabel metal2 13662 1860 13662 1860 0 chany_bottom_out[4]
rlabel metal2 14030 2166 14030 2166 0 chany_bottom_out[5]
rlabel metal2 14398 1554 14398 1554 0 chany_bottom_out[6]
rlabel metal2 14766 1860 14766 1860 0 chany_bottom_out[7]
rlabel metal2 15134 1622 15134 1622 0 chany_bottom_out[8]
rlabel metal2 15502 2166 15502 2166 0 chany_bottom_out[9]
rlabel metal2 12374 52292 12374 52292 0 chany_top_in_0[0]
rlabel metal1 16882 54196 16882 54196 0 chany_top_in_0[10]
rlabel metal1 16468 53550 16468 53550 0 chany_top_in_0[11]
rlabel metal1 17020 53550 17020 53550 0 chany_top_in_0[12]
rlabel metal1 17480 54162 17480 54162 0 chany_top_in_0[13]
rlabel metal1 17986 54230 17986 54230 0 chany_top_in_0[14]
rlabel metal1 17940 53550 17940 53550 0 chany_top_in_0[15]
rlabel metal1 18446 53210 18446 53210 0 chany_top_in_0[16]
rlabel metal1 19044 54162 19044 54162 0 chany_top_in_0[17]
rlabel metal1 19366 53550 19366 53550 0 chany_top_in_0[18]
rlabel metal1 20194 54162 20194 54162 0 chany_top_in_0[19]
rlabel metal1 13616 53142 13616 53142 0 chany_top_in_0[1]
rlabel metal1 19872 53074 19872 53074 0 chany_top_in_0[20]
rlabel metal1 20930 54196 20930 54196 0 chany_top_in_0[21]
rlabel metal1 20378 53754 20378 53754 0 chany_top_in_0[22]
rlabel metal1 21068 53550 21068 53550 0 chany_top_in_0[23]
rlabel metal2 21206 55192 21206 55192 0 chany_top_in_0[24]
rlabel metal2 21574 54886 21574 54886 0 chany_top_in_0[25]
rlabel metal1 21988 53074 21988 53074 0 chany_top_in_0[26]
rlabel metal1 22632 53074 22632 53074 0 chany_top_in_0[27]
rlabel metal1 24794 54196 24794 54196 0 chany_top_in_0[28]
rlabel metal2 23230 56236 23230 56236 0 chany_top_in_0[29]
rlabel metal1 13018 52394 13018 52394 0 chany_top_in_0[2]
rlabel metal1 13662 53074 13662 53074 0 chany_top_in_0[3]
rlabel metal2 13846 55260 13846 55260 0 chany_top_in_0[4]
rlabel metal1 14398 53550 14398 53550 0 chany_top_in_0[5]
rlabel metal1 14490 54298 14490 54298 0 chany_top_in_0[6]
rlabel metal1 15226 54230 15226 54230 0 chany_top_in_0[7]
rlabel metal1 15732 54162 15732 54162 0 chany_top_in_0[8]
rlabel metal1 15548 53754 15548 53754 0 chany_top_in_0[9]
rlabel metal1 1564 49266 1564 49266 0 chany_top_out_0[0]
rlabel metal2 5014 54138 5014 54138 0 chany_top_out_0[10]
rlabel metal1 4186 54094 4186 54094 0 chany_top_out_0[11]
rlabel metal1 5658 53006 5658 53006 0 chany_top_out_0[12]
rlabel metal2 6118 54376 6118 54376 0 chany_top_out_0[13]
rlabel metal2 6486 54376 6486 54376 0 chany_top_out_0[14]
rlabel metal2 6854 54461 6854 54461 0 chany_top_out_0[15]
rlabel metal1 6394 54094 6394 54094 0 chany_top_out_0[16]
rlabel metal1 6946 53618 6946 53618 0 chany_top_out_0[17]
rlabel metal2 7958 55711 7958 55711 0 chany_top_out_0[18]
rlabel metal2 8326 54920 8326 54920 0 chany_top_out_0[19]
rlabel metal1 1840 49878 1840 49878 0 chany_top_out_0[1]
rlabel metal2 8694 54614 8694 54614 0 chany_top_out_0[20]
rlabel metal1 9384 53550 9384 53550 0 chany_top_out_0[21]
rlabel metal1 8786 54094 8786 54094 0 chany_top_out_0[22]
rlabel metal1 10074 52530 10074 52530 0 chany_top_out_0[23]
rlabel metal1 10212 53006 10212 53006 0 chany_top_out_0[24]
rlabel metal2 10534 54920 10534 54920 0 chany_top_out_0[25]
rlabel metal2 10902 55226 10902 55226 0 chany_top_out_0[26]
rlabel metal1 11730 53006 11730 53006 0 chany_top_out_0[27]
rlabel metal1 11914 53618 11914 53618 0 chany_top_out_0[28]
rlabel metal2 12006 55158 12006 55158 0 chany_top_out_0[29]
rlabel metal1 2162 50354 2162 50354 0 chany_top_out_0[2]
rlabel metal2 2438 53832 2438 53832 0 chany_top_out_0[3]
rlabel metal2 2806 55711 2806 55711 0 chany_top_out_0[4]
rlabel metal2 3174 55711 3174 55711 0 chany_top_out_0[5]
rlabel metal2 3542 54070 3542 54070 0 chany_top_out_0[6]
rlabel metal2 4048 53244 4048 53244 0 chany_top_out_0[7]
rlabel metal1 4002 53006 4002 53006 0 chany_top_out_0[8]
rlabel metal1 3818 53618 3818 53618 0 chany_top_out_0[9]
rlabel metal1 19412 41582 19412 41582 0 clknet_0_prog_clk
rlabel metal1 5382 8602 5382 8602 0 clknet_4_0_0_prog_clk
rlabel metal1 6302 38386 6302 38386 0 clknet_4_10_0_prog_clk
rlabel metal2 14306 43792 14306 43792 0 clknet_4_11_0_prog_clk
rlabel metal2 19550 38046 19550 38046 0 clknet_4_12_0_prog_clk
rlabel metal1 23230 37876 23230 37876 0 clknet_4_13_0_prog_clk
rlabel metal1 18584 41650 18584 41650 0 clknet_4_14_0_prog_clk
rlabel metal2 22034 42942 22034 42942 0 clknet_4_15_0_prog_clk
rlabel metal2 11270 11424 11270 11424 0 clknet_4_1_0_prog_clk
rlabel metal2 5014 20740 5014 20740 0 clknet_4_2_0_prog_clk
rlabel metal1 13846 20978 13846 20978 0 clknet_4_3_0_prog_clk
rlabel metal1 17894 12274 17894 12274 0 clknet_4_4_0_prog_clk
rlabel metal1 22678 18292 22678 18292 0 clknet_4_5_0_prog_clk
rlabel metal1 16330 22066 16330 22066 0 clknet_4_6_0_prog_clk
rlabel metal1 24886 21454 24886 21454 0 clknet_4_7_0_prog_clk
rlabel metal2 7774 32878 7774 32878 0 clknet_4_8_0_prog_clk
rlabel metal1 13478 34646 13478 34646 0 clknet_4_9_0_prog_clk
rlabel metal3 1234 13396 1234 13396 0 gfpga_pad_io_soc_dir[0]
rlabel metal3 1004 15708 1004 15708 0 gfpga_pad_io_soc_dir[1]
rlabel metal3 1004 18020 1004 18020 0 gfpga_pad_io_soc_dir[2]
rlabel metal3 1004 20332 1004 20332 0 gfpga_pad_io_soc_dir[3]
rlabel metal1 1472 32402 1472 32402 0 gfpga_pad_io_soc_in[0]
rlabel metal2 1610 34391 1610 34391 0 gfpga_pad_io_soc_in[1]
rlabel metal1 1472 36754 1472 36754 0 gfpga_pad_io_soc_in[2]
rlabel metal1 1426 38930 1426 38930 0 gfpga_pad_io_soc_in[3]
rlabel metal3 820 22644 820 22644 0 gfpga_pad_io_soc_out[0]
rlabel metal3 1004 24956 1004 24956 0 gfpga_pad_io_soc_out[1]
rlabel metal3 1004 27268 1004 27268 0 gfpga_pad_io_soc_out[2]
rlabel metal3 1004 29580 1004 29580 0 gfpga_pad_io_soc_out[3]
rlabel metal2 1702 41327 1702 41327 0 isol_n
rlabel metal1 2944 52870 2944 52870 0 net1
rlabel metal1 18630 34952 18630 34952 0 net10
rlabel metal1 24288 52122 24288 52122 0 net100
rlabel metal1 24840 2618 24840 2618 0 net101
rlabel metal2 24610 44302 24610 44302 0 net102
rlabel metal1 23598 47226 23598 47226 0 net103
rlabel metal1 16284 17306 16284 17306 0 net104
rlabel metal1 17526 18802 17526 18802 0 net105
rlabel metal1 18952 43418 18952 43418 0 net106
rlabel metal2 21482 45356 21482 45356 0 net107
rlabel metal1 18768 15470 18768 15470 0 net108
rlabel metal1 13662 13362 13662 13362 0 net109
rlabel metal1 19504 34510 19504 34510 0 net11
rlabel metal1 25392 51238 25392 51238 0 net110
rlabel metal1 25438 51782 25438 51782 0 net111
rlabel metal2 25254 6256 25254 6256 0 net112
rlabel metal1 24288 47770 24288 47770 0 net113
rlabel metal1 23690 47770 23690 47770 0 net114
rlabel metal2 14766 37502 14766 37502 0 net115
rlabel metal1 14076 34646 14076 34646 0 net116
rlabel metal1 14536 38250 14536 38250 0 net117
rlabel metal1 4416 52462 4416 52462 0 net118
rlabel metal1 20102 6324 20102 6324 0 net119
rlabel metal1 22402 38896 22402 38896 0 net12
rlabel metal1 11684 37298 11684 37298 0 net120
rlabel metal2 22678 12036 22678 12036 0 net121
rlabel metal1 21574 12410 21574 12410 0 net122
rlabel metal1 21482 15912 21482 15912 0 net123
rlabel metal2 23966 14382 23966 14382 0 net124
rlabel metal2 22126 16286 22126 16286 0 net125
rlabel metal2 22954 14110 22954 14110 0 net126
rlabel metal1 22448 19754 22448 19754 0 net127
rlabel metal1 24150 18666 24150 18666 0 net128
rlabel metal1 23460 20842 23460 20842 0 net129
rlabel metal1 17434 38250 17434 38250 0 net13
rlabel metal1 23184 22406 23184 22406 0 net130
rlabel metal1 24426 5202 24426 5202 0 net131
rlabel metal1 24380 17646 24380 17646 0 net132
rlabel metal1 21896 19346 21896 19346 0 net133
rlabel metal2 23414 20713 23414 20713 0 net134
rlabel metal1 24426 19822 24426 19822 0 net135
rlabel metal1 25070 26282 25070 26282 0 net136
rlabel metal1 24150 21998 24150 21998 0 net137
rlabel metal1 24196 23086 24196 23086 0 net138
rlabel metal1 23644 23698 23644 23698 0 net139
rlabel metal1 18308 24242 18308 24242 0 net14
rlabel metal1 24288 24174 24288 24174 0 net140
rlabel metal2 24150 24412 24150 24412 0 net141
rlabel metal1 24058 6732 24058 6732 0 net142
rlabel metal1 23644 6290 23644 6290 0 net143
rlabel metal1 24150 7854 24150 7854 0 net144
rlabel metal2 24150 8636 24150 8636 0 net145
rlabel metal2 24058 9724 24058 9724 0 net146
rlabel metal1 24334 10030 24334 10030 0 net147
rlabel metal2 16238 5678 16238 5678 0 net148
rlabel metal2 23966 11084 23966 11084 0 net149
rlabel metal1 16146 39440 16146 39440 0 net15
rlabel metal1 11730 14858 11730 14858 0 net150
rlabel metal2 16882 4182 16882 4182 0 net151
rlabel metal1 16054 4114 16054 4114 0 net152
rlabel metal1 17848 4998 17848 4998 0 net153
rlabel metal1 17756 2346 17756 2346 0 net154
rlabel metal1 16928 4590 16928 4590 0 net155
rlabel metal1 18630 3502 18630 3502 0 net156
rlabel metal1 18676 4114 18676 4114 0 net157
rlabel metal1 20516 2550 20516 2550 0 net158
rlabel metal1 19136 5746 19136 5746 0 net159
rlabel via2 19918 29699 19918 29699 0 net16
rlabel metal1 21206 3502 21206 3502 0 net160
rlabel metal2 13754 3842 13754 3842 0 net161
rlabel metal1 19550 5202 19550 5202 0 net162
rlabel metal1 21252 4590 21252 4590 0 net163
rlabel metal1 20976 13906 20976 13906 0 net164
rlabel metal1 19734 8874 19734 8874 0 net165
rlabel metal1 19090 6698 19090 6698 0 net166
rlabel metal2 23506 7854 23506 7854 0 net167
rlabel metal1 19596 7786 19596 7786 0 net168
rlabel metal2 20194 6086 20194 6086 0 net169
rlabel metal1 15272 34714 15272 34714 0 net17
rlabel metal1 20562 6426 20562 6426 0 net170
rlabel metal1 20240 6630 20240 6630 0 net171
rlabel metal1 12880 4114 12880 4114 0 net172
rlabel metal1 12098 9962 12098 9962 0 net173
rlabel metal1 13984 12138 13984 12138 0 net174
rlabel metal1 13984 12614 13984 12614 0 net175
rlabel via3 15709 2652 15709 2652 0 net176
rlabel metal1 16376 3026 16376 3026 0 net177
rlabel metal2 15732 4692 15732 4692 0 net178
rlabel metal1 15594 3502 15594 3502 0 net179
rlabel metal2 14582 36397 14582 36397 0 net18
rlabel metal1 3174 40630 3174 40630 0 net180
rlabel metal1 6026 52020 6026 52020 0 net181
rlabel metal2 5934 52870 5934 52870 0 net182
rlabel metal1 6624 44982 6624 44982 0 net183
rlabel metal1 7130 45526 7130 45526 0 net184
rlabel metal2 7774 51217 7774 51217 0 net185
rlabel metal1 6900 49946 6900 49946 0 net186
rlabel metal1 6463 54162 6463 54162 0 net187
rlabel metal2 8326 43520 8326 43520 0 net188
rlabel metal1 9062 52462 9062 52462 0 net189
rlabel metal1 18814 35564 18814 35564 0 net19
rlabel metal1 7636 49946 7636 49946 0 net190
rlabel metal2 3726 46036 3726 46036 0 net191
rlabel metal1 9844 43962 9844 43962 0 net192
rlabel metal1 10258 51986 10258 51986 0 net193
rlabel metal1 9200 54162 9200 54162 0 net194
rlabel metal1 9752 52462 9752 52462 0 net195
rlabel metal1 9614 53074 9614 53074 0 net196
rlabel metal2 11086 48994 11086 48994 0 net197
rlabel metal2 9890 52598 9890 52598 0 net198
rlabel metal1 11224 53074 11224 53074 0 net199
rlabel metal1 2668 3706 2668 3706 0 net2
rlabel metal2 17618 36193 17618 36193 0 net20
rlabel metal2 11914 52836 11914 52836 0 net200
rlabel metal1 12052 52666 12052 52666 0 net201
rlabel metal1 3726 50286 3726 50286 0 net202
rlabel metal1 5106 51306 5106 51306 0 net203
rlabel metal2 4186 46818 4186 46818 0 net204
rlabel metal1 3772 52462 3772 52462 0 net205
rlabel metal1 4738 51986 4738 51986 0 net206
rlabel metal1 5704 51374 5704 51374 0 net207
rlabel metal1 4094 53108 4094 53108 0 net208
rlabel metal1 4830 53550 4830 53550 0 net209
rlabel metal1 16652 38318 16652 38318 0 net21
rlabel metal2 2806 15266 2806 15266 0 net210
rlabel metal1 1932 18598 1932 18598 0 net211
rlabel metal1 1840 18258 1840 18258 0 net212
rlabel metal2 1794 21148 1794 21148 0 net213
rlabel metal1 2760 21862 2760 21862 0 net214
rlabel metal1 1886 22746 1886 22746 0 net215
rlabel metal1 2024 24650 2024 24650 0 net216
rlabel metal1 1932 27098 1932 27098 0 net217
rlabel metal1 19182 5236 19182 5236 0 net218
rlabel metal2 24150 45628 24150 45628 0 net219
rlabel metal2 20562 40528 20562 40528 0 net22
rlabel metal2 23966 53414 23966 53414 0 net220
rlabel metal1 23506 8500 23506 8500 0 net221
rlabel metal1 25070 53074 25070 53074 0 net222
rlabel metal1 21482 7412 21482 7412 0 net223
rlabel metal1 24334 47702 24334 47702 0 net224
rlabel metal2 25346 4879 25346 4879 0 net225
rlabel metal1 17066 20570 17066 20570 0 net226
rlabel metal1 13248 27438 13248 27438 0 net227
rlabel metal1 23230 31858 23230 31858 0 net228
rlabel metal1 20930 21658 20930 21658 0 net229
rlabel metal1 18124 40358 18124 40358 0 net23
rlabel metal1 15272 36754 15272 36754 0 net230
rlabel metal1 17664 22610 17664 22610 0 net231
rlabel metal2 22218 28798 22218 28798 0 net232
rlabel metal2 16330 36414 16330 36414 0 net233
rlabel metal1 18170 37230 18170 37230 0 net234
rlabel metal2 16146 38080 16146 38080 0 net235
rlabel metal1 14260 39066 14260 39066 0 net236
rlabel metal1 13708 37842 13708 37842 0 net237
rlabel metal2 23414 40800 23414 40800 0 net238
rlabel metal2 13386 32640 13386 32640 0 net239
rlabel metal1 22586 38998 22586 38998 0 net24
rlabel metal2 10994 29886 10994 29886 0 net240
rlabel metal2 12558 25024 12558 25024 0 net241
rlabel metal2 10626 26826 10626 26826 0 net242
rlabel metal1 8096 26010 8096 26010 0 net243
rlabel metal2 8694 26486 8694 26486 0 net244
rlabel metal1 7866 24174 7866 24174 0 net245
rlabel metal1 10488 23698 10488 23698 0 net246
rlabel metal1 6486 9554 6486 9554 0 net247
rlabel metal1 15134 11118 15134 11118 0 net248
rlabel metal1 20056 33966 20056 33966 0 net249
rlabel metal1 16698 25330 16698 25330 0 net25
rlabel metal2 17250 13056 17250 13056 0 net250
rlabel metal2 18538 15232 18538 15232 0 net251
rlabel metal1 20470 15538 20470 15538 0 net252
rlabel metal2 21850 15946 21850 15946 0 net253
rlabel metal2 19550 15572 19550 15572 0 net254
rlabel metal1 22954 13362 22954 13362 0 net255
rlabel metal1 20240 11050 20240 11050 0 net256
rlabel metal1 18814 13294 18814 13294 0 net257
rlabel metal2 23230 34816 23230 34816 0 net258
rlabel metal2 21758 40596 21758 40596 0 net259
rlabel metal1 17618 26350 17618 26350 0 net26
rlabel metal1 10764 36890 10764 36890 0 net260
rlabel metal1 8142 31314 8142 31314 0 net261
rlabel metal1 9108 32538 9108 32538 0 net262
rlabel metal1 12236 37978 12236 37978 0 net263
rlabel metal1 8050 31450 8050 31450 0 net264
rlabel metal1 4968 31450 4968 31450 0 net265
rlabel metal1 8418 38318 8418 38318 0 net266
rlabel metal1 10258 35054 10258 35054 0 net267
rlabel metal2 11086 38590 11086 38590 0 net268
rlabel metal1 14996 35054 14996 35054 0 net269
rlabel metal1 19136 33626 19136 33626 0 net27
rlabel metal2 7498 31518 7498 31518 0 net270
rlabel metal1 10396 23018 10396 23018 0 net271
rlabel metal2 11730 20094 11730 20094 0 net272
rlabel metal1 9154 16116 9154 16116 0 net273
rlabel metal1 9016 23834 9016 23834 0 net274
rlabel metal2 13570 21216 13570 21216 0 net275
rlabel metal2 13570 23936 13570 23936 0 net276
rlabel metal1 20056 24922 20056 24922 0 net277
rlabel metal1 23460 25194 23460 25194 0 net278
rlabel metal1 17848 28458 17848 28458 0 net279
rlabel metal1 18584 35054 18584 35054 0 net28
rlabel metal1 19228 34714 19228 34714 0 net29
rlabel metal1 20056 24106 20056 24106 0 net3
rlabel metal1 22770 32334 22770 32334 0 net30
rlabel metal1 17020 36890 17020 36890 0 net31
rlabel metal1 17296 30702 17296 30702 0 net32
rlabel metal1 3772 3978 3772 3978 0 net33
rlabel metal2 5106 3944 5106 3944 0 net34
rlabel metal1 5152 3162 5152 3162 0 net35
rlabel metal2 16054 4420 16054 4420 0 net36
rlabel metal2 12834 37587 12834 37587 0 net37
rlabel metal1 6624 3706 6624 3706 0 net38
rlabel metal1 7130 2482 7130 2482 0 net39
rlabel metal1 17526 31858 17526 31858 0 net4
rlabel metal1 10764 5542 10764 5542 0 net40
rlabel metal1 7728 3706 7728 3706 0 net41
rlabel metal1 8418 2550 8418 2550 0 net42
rlabel metal2 8418 3978 8418 3978 0 net43
rlabel metal1 3404 3638 3404 3638 0 net44
rlabel metal2 8878 4963 8878 4963 0 net45
rlabel metal1 7912 3978 7912 3978 0 net46
rlabel metal1 10810 3978 10810 3978 0 net47
rlabel metal1 10672 3366 10672 3366 0 net48
rlabel metal1 14352 3434 14352 3434 0 net49
rlabel metal1 24426 32742 24426 32742 0 net5
rlabel metal1 13386 5746 13386 5746 0 net50
rlabel metal1 12604 3706 12604 3706 0 net51
rlabel metal1 12144 2006 12144 2006 0 net52
rlabel metal1 13662 2618 13662 2618 0 net53
rlabel metal2 12282 4963 12282 4963 0 net54
rlabel metal2 2162 10608 2162 10608 0 net55
rlabel metal1 4554 2448 4554 2448 0 net56
rlabel metal2 3174 2244 3174 2244 0 net57
rlabel metal1 3358 3706 3358 3706 0 net58
rlabel metal1 3910 2958 3910 2958 0 net59
rlabel metal2 20838 30362 20838 30362 0 net6
rlabel metal1 4140 2890 4140 2890 0 net60
rlabel metal1 4462 2550 4462 2550 0 net61
rlabel metal1 4462 3128 4462 3128 0 net62
rlabel metal1 13340 40494 13340 40494 0 net63
rlabel metal1 15548 13498 15548 13498 0 net64
rlabel metal1 16813 44506 16813 44506 0 net65
rlabel metal1 17342 46682 17342 46682 0 net66
rlabel metal1 18078 47022 18078 47022 0 net67
rlabel metal2 18492 42364 18492 42364 0 net68
rlabel metal1 16054 15062 16054 15062 0 net69
rlabel metal1 19688 32538 19688 32538 0 net7
rlabel metal1 18630 46682 18630 46682 0 net70
rlabel metal1 19964 46682 19964 46682 0 net71
rlabel metal3 19481 44268 19481 44268 0 net72
rlabel metal1 20838 45866 20838 45866 0 net73
rlabel metal2 12834 15827 12834 15827 0 net74
rlabel metal1 19780 46002 19780 46002 0 net75
rlabel metal1 21160 41446 21160 41446 0 net76
rlabel via2 21482 44285 21482 44285 0 net77
rlabel via3 21459 45492 21459 45492 0 net78
rlabel metal1 21114 45526 21114 45526 0 net79
rlabel metal1 20102 36142 20102 36142 0 net8
rlabel metal1 21298 46002 21298 46002 0 net80
rlabel metal1 20608 11730 20608 11730 0 net81
rlabel metal2 22770 52054 22770 52054 0 net82
rlabel metal2 21942 45227 21942 45227 0 net83
rlabel metal1 24564 53414 24564 53414 0 net84
rlabel metal1 14674 15470 14674 15470 0 net85
rlabel metal1 13340 12954 13340 12954 0 net86
rlabel metal1 14122 44506 14122 44506 0 net87
rlabel metal1 13110 12138 13110 12138 0 net88
rlabel metal1 13156 13498 13156 13498 0 net89
rlabel metal1 18722 33388 18722 33388 0 net9
rlabel metal2 16238 17187 16238 17187 0 net90
rlabel metal1 17710 47056 17710 47056 0 net91
rlabel metal1 15502 12206 15502 12206 0 net92
rlabel metal2 2622 29308 2622 29308 0 net93
rlabel metal2 2714 31110 2714 31110 0 net94
rlabel metal1 1886 36550 1886 36550 0 net95
rlabel metal1 2898 38726 2898 38726 0 net96
rlabel metal1 9752 17646 9752 17646 0 net97
rlabel metal2 25070 21862 25070 21862 0 net98
rlabel metal1 1932 43418 1932 43418 0 net99
rlabel metal2 23230 1639 23230 1639 0 prog_clk
rlabel metal1 24518 2890 24518 2890 0 prog_reset_bottom_in
rlabel metal2 20562 4012 20562 4012 0 prog_reset_bottom_out
rlabel metal1 1472 43758 1472 43758 0 prog_reset_left_in
rlabel metal2 24794 45577 24794 45577 0 prog_reset_right_out
rlabel metal2 24518 55711 24518 55711 0 prog_reset_top_in
rlabel metal1 23874 54094 23874 54094 0 prog_reset_top_out
rlabel metal1 24610 2414 24610 2414 0 reset_bottom_in
rlabel metal2 24702 1761 24702 1761 0 reset_bottom_out
rlabel metal1 24564 46410 24564 46410 0 reset_right_in
rlabel metal2 23506 52496 23506 52496 0 reset_top_in
rlabel metal2 24886 54614 24886 54614 0 reset_top_out
rlabel metal2 25530 47277 25530 47277 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
rlabel metal2 24794 48263 24794 48263 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_
rlabel metal2 25346 48841 25346 48841 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
rlabel metal2 24794 49487 24794 49487 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_
rlabel metal2 25346 50065 25346 50065 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
rlabel metal2 25346 50711 25346 50711 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_
rlabel metal2 25346 51289 25346 51289 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_
rlabel metal2 25254 51935 25254 51935 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_
rlabel metal3 1970 4148 1970 4148 0 right_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal3 1924 6460 1924 6460 0 right_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal3 1786 8772 1786 8772 0 right_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal3 2016 11084 2016 11084 0 right_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal2 18630 15844 18630 15844 0 sb_0__1_.mem_bottom_track_1.ccff_head
rlabel metal2 16054 20570 16054 20570 0 sb_0__1_.mem_bottom_track_1.ccff_tail
rlabel metal1 15686 17850 15686 17850 0 sb_0__1_.mem_bottom_track_1.mem_out\[0\]
rlabel metal1 15410 22746 15410 22746 0 sb_0__1_.mem_bottom_track_1.mem_out\[1\]
rlabel metal1 20194 21318 20194 21318 0 sb_0__1_.mem_bottom_track_11.ccff_head
rlabel metal1 16790 24718 16790 24718 0 sb_0__1_.mem_bottom_track_11.ccff_tail
rlabel metal1 17526 32266 17526 32266 0 sb_0__1_.mem_bottom_track_11.mem_out\[0\]
rlabel metal1 16192 26554 16192 26554 0 sb_0__1_.mem_bottom_track_11.mem_out\[1\]
rlabel metal2 21114 24684 21114 24684 0 sb_0__1_.mem_bottom_track_13.ccff_tail
rlabel metal2 21206 32037 21206 32037 0 sb_0__1_.mem_bottom_track_13.mem_out\[0\]
rlabel metal1 19504 27642 19504 27642 0 sb_0__1_.mem_bottom_track_13.mem_out\[1\]
rlabel metal1 24932 24718 24932 24718 0 sb_0__1_.mem_bottom_track_21.ccff_tail
rlabel metal1 20056 26418 20056 26418 0 sb_0__1_.mem_bottom_track_21.mem_out\[0\]
rlabel metal1 24012 27574 24012 27574 0 sb_0__1_.mem_bottom_track_21.mem_out\[1\]
rlabel metal1 16514 28730 16514 28730 0 sb_0__1_.mem_bottom_track_29.ccff_tail
rlabel metal1 17066 32368 17066 32368 0 sb_0__1_.mem_bottom_track_29.mem_out\[0\]
rlabel metal1 16238 28594 16238 28594 0 sb_0__1_.mem_bottom_track_29.mem_out\[1\]
rlabel metal1 20608 20366 20608 20366 0 sb_0__1_.mem_bottom_track_3.ccff_tail
rlabel metal1 17618 26860 17618 26860 0 sb_0__1_.mem_bottom_track_3.mem_out\[0\]
rlabel metal1 18952 20502 18952 20502 0 sb_0__1_.mem_bottom_track_3.mem_out\[1\]
rlabel metal1 16652 32810 16652 32810 0 sb_0__1_.mem_bottom_track_37.ccff_tail
rlabel metal2 15962 32164 15962 32164 0 sb_0__1_.mem_bottom_track_37.mem_out\[0\]
rlabel metal1 15870 32198 15870 32198 0 sb_0__1_.mem_bottom_track_37.mem_out\[1\]
rlabel metal1 20332 33014 20332 33014 0 sb_0__1_.mem_bottom_track_45.ccff_tail
rlabel metal1 20332 33898 20332 33898 0 sb_0__1_.mem_bottom_track_45.mem_out\[0\]
rlabel metal2 23230 32572 23230 32572 0 sb_0__1_.mem_bottom_track_45.mem_out\[1\]
rlabel metal1 23874 20570 23874 20570 0 sb_0__1_.mem_bottom_track_5.ccff_tail
rlabel metal1 22264 21046 22264 21046 0 sb_0__1_.mem_bottom_track_5.mem_out\[0\]
rlabel metal2 24288 21828 24288 21828 0 sb_0__1_.mem_bottom_track_5.mem_out\[1\]
rlabel metal1 10488 43214 10488 43214 0 sb_0__1_.mem_bottom_track_53.mem_out\[0\]
rlabel metal1 22172 21590 22172 21590 0 sb_0__1_.mem_bottom_track_7.mem_out\[0\]
rlabel metal1 19734 21454 19734 21454 0 sb_0__1_.mem_bottom_track_7.mem_out\[1\]
rlabel metal2 18814 38590 18814 38590 0 sb_0__1_.mem_right_track_0.ccff_head
rlabel metal1 23644 30158 23644 30158 0 sb_0__1_.mem_right_track_0.ccff_tail
rlabel metal1 20608 31858 20608 31858 0 sb_0__1_.mem_right_track_0.mem_out\[0\]
rlabel metal2 22218 29801 22218 29801 0 sb_0__1_.mem_right_track_0.mem_out\[1\]
rlabel metal2 22126 42806 22126 42806 0 sb_0__1_.mem_right_track_10.ccff_head
rlabel metal1 19872 43690 19872 43690 0 sb_0__1_.mem_right_track_10.ccff_tail
rlabel metal1 21436 44234 21436 44234 0 sb_0__1_.mem_right_track_10.mem_out\[0\]
rlabel metal1 20010 41684 20010 41684 0 sb_0__1_.mem_right_track_10.mem_out\[1\]
rlabel metal1 19412 44438 19412 44438 0 sb_0__1_.mem_right_track_12.ccff_tail
rlabel metal2 20930 44370 20930 44370 0 sb_0__1_.mem_right_track_12.mem_out\[0\]
rlabel metal1 18676 42126 18676 42126 0 sb_0__1_.mem_right_track_12.mem_out\[1\]
rlabel metal1 17480 45866 17480 45866 0 sb_0__1_.mem_right_track_14.ccff_tail
rlabel metal1 18124 44506 18124 44506 0 sb_0__1_.mem_right_track_14.mem_out\[0\]
rlabel metal2 16882 44030 16882 44030 0 sb_0__1_.mem_right_track_14.mem_out\[1\]
rlabel metal1 15640 46614 15640 46614 0 sb_0__1_.mem_right_track_16.ccff_tail
rlabel via1 16606 46546 16606 46546 0 sb_0__1_.mem_right_track_16.mem_out\[0\]
rlabel metal1 17434 43180 17434 43180 0 sb_0__1_.mem_right_track_16.mem_out\[1\]
rlabel metal1 15364 42126 15364 42126 0 sb_0__1_.mem_right_track_18.ccff_tail
rlabel metal1 17894 47158 17894 47158 0 sb_0__1_.mem_right_track_18.mem_out\[0\]
rlabel metal1 13652 42874 13652 42874 0 sb_0__1_.mem_right_track_18.mem_out\[1\]
rlabel metal1 24932 39474 24932 39474 0 sb_0__1_.mem_right_track_2.ccff_tail
rlabel metal1 20516 36210 20516 36210 0 sb_0__1_.mem_right_track_2.mem_out\[0\]
rlabel metal1 22218 41004 22218 41004 0 sb_0__1_.mem_right_track_2.mem_out\[1\]
rlabel metal1 13064 35122 13064 35122 0 sb_0__1_.mem_right_track_20.ccff_tail
rlabel metal1 14122 41990 14122 41990 0 sb_0__1_.mem_right_track_20.mem_out\[0\]
rlabel metal1 14444 37774 14444 37774 0 sb_0__1_.mem_right_track_20.mem_out\[1\]
rlabel metal1 13064 29682 13064 29682 0 sb_0__1_.mem_right_track_22.ccff_tail
rlabel metal1 13570 35598 13570 35598 0 sb_0__1_.mem_right_track_22.mem_out\[0\]
rlabel metal1 14030 33490 14030 33490 0 sb_0__1_.mem_right_track_22.mem_out\[1\]
rlabel metal2 13478 24956 13478 24956 0 sb_0__1_.mem_right_track_24.ccff_tail
rlabel metal1 12972 25806 12972 25806 0 sb_0__1_.mem_right_track_24.mem_out\[0\]
rlabel metal2 12650 27234 12650 27234 0 sb_0__1_.mem_right_track_26.ccff_tail
rlabel metal2 15410 28628 15410 28628 0 sb_0__1_.mem_right_track_26.mem_out\[0\]
rlabel metal1 7084 27982 7084 27982 0 sb_0__1_.mem_right_track_28.ccff_tail
rlabel metal1 9568 29274 9568 29274 0 sb_0__1_.mem_right_track_28.mem_out\[0\]
rlabel metal1 7222 26418 7222 26418 0 sb_0__1_.mem_right_track_30.ccff_tail
rlabel metal1 9200 27982 9200 27982 0 sb_0__1_.mem_right_track_30.mem_out\[0\]
rlabel metal1 9384 24718 9384 24718 0 sb_0__1_.mem_right_track_32.ccff_tail
rlabel metal2 12466 27829 12466 27829 0 sb_0__1_.mem_right_track_32.mem_out\[0\]
rlabel metal1 12466 23596 12466 23596 0 sb_0__1_.mem_right_track_34.ccff_tail
rlabel metal1 13570 27880 13570 27880 0 sb_0__1_.mem_right_track_34.mem_out\[0\]
rlabel metal1 9246 12138 9246 12138 0 sb_0__1_.mem_right_track_36.ccff_tail
rlabel metal1 8510 18802 8510 18802 0 sb_0__1_.mem_right_track_36.mem_out\[0\]
rlabel metal1 6762 9452 6762 9452 0 sb_0__1_.mem_right_track_36.mem_out\[1\]
rlabel metal1 13708 11186 13708 11186 0 sb_0__1_.mem_right_track_38.ccff_tail
rlabel metal1 11776 12410 11776 12410 0 sb_0__1_.mem_right_track_38.mem_out\[0\]
rlabel metal2 21758 35904 21758 35904 0 sb_0__1_.mem_right_track_4.ccff_tail
rlabel metal1 21850 44948 21850 44948 0 sb_0__1_.mem_right_track_4.mem_out\[0\]
rlabel metal1 21712 37162 21712 37162 0 sb_0__1_.mem_right_track_4.mem_out\[1\]
rlabel metal1 16238 12750 16238 12750 0 sb_0__1_.mem_right_track_40.ccff_tail
rlabel metal2 14490 13328 14490 13328 0 sb_0__1_.mem_right_track_40.mem_out\[0\]
rlabel metal1 17664 15674 17664 15674 0 sb_0__1_.mem_right_track_44.ccff_tail
rlabel metal1 16192 15402 16192 15402 0 sb_0__1_.mem_right_track_44.mem_out\[0\]
rlabel metal2 21206 16864 21206 16864 0 sb_0__1_.mem_right_track_46.ccff_tail
rlabel metal2 19090 18122 19090 18122 0 sb_0__1_.mem_right_track_46.mem_out\[0\]
rlabel metal1 23552 17306 23552 17306 0 sb_0__1_.mem_right_track_48.ccff_tail
rlabel metal1 22310 17272 22310 17272 0 sb_0__1_.mem_right_track_48.mem_out\[0\]
rlabel metal1 22356 18598 22356 18598 0 sb_0__1_.mem_right_track_50.ccff_tail
rlabel metal1 23098 18938 23098 18938 0 sb_0__1_.mem_right_track_50.mem_out\[0\]
rlabel metal1 20884 13158 20884 13158 0 sb_0__1_.mem_right_track_52.ccff_tail
rlabel metal2 21666 14790 21666 14790 0 sb_0__1_.mem_right_track_52.mem_out\[0\]
rlabel metal1 19412 11186 19412 11186 0 sb_0__1_.mem_right_track_54.ccff_tail
rlabel metal2 19550 11565 19550 11565 0 sb_0__1_.mem_right_track_54.mem_out\[0\]
rlabel metal2 17158 14382 17158 14382 0 sb_0__1_.mem_right_track_56.mem_out\[0\]
rlabel metal1 23506 36244 23506 36244 0 sb_0__1_.mem_right_track_6.ccff_tail
rlabel metal1 21344 36210 21344 36210 0 sb_0__1_.mem_right_track_6.mem_out\[0\]
rlabel metal2 25070 35360 25070 35360 0 sb_0__1_.mem_right_track_6.mem_out\[1\]
rlabel metal1 20838 46036 20838 46036 0 sb_0__1_.mem_right_track_8.mem_out\[0\]
rlabel metal1 22218 39984 22218 39984 0 sb_0__1_.mem_right_track_8.mem_out\[1\]
rlabel metal2 12374 43996 12374 43996 0 sb_0__1_.mem_top_track_0.ccff_tail
rlabel metal1 17572 40562 17572 40562 0 sb_0__1_.mem_top_track_0.mem_out\[0\]
rlabel metal1 12834 43180 12834 43180 0 sb_0__1_.mem_top_track_0.mem_out\[1\]
rlabel metal1 5934 38522 5934 38522 0 sb_0__1_.mem_top_track_10.ccff_head
rlabel metal1 6624 35802 6624 35802 0 sb_0__1_.mem_top_track_10.ccff_tail
rlabel metal1 13754 35530 13754 35530 0 sb_0__1_.mem_top_track_10.mem_out\[0\]
rlabel metal1 10626 37298 10626 37298 0 sb_0__1_.mem_top_track_10.mem_out\[1\]
rlabel metal2 9522 35156 9522 35156 0 sb_0__1_.mem_top_track_12.ccff_tail
rlabel metal1 8510 34510 8510 34510 0 sb_0__1_.mem_top_track_12.mem_out\[0\]
rlabel metal1 12627 34034 12627 34034 0 sb_0__1_.mem_top_track_12.mem_out\[1\]
rlabel metal1 11546 40902 11546 40902 0 sb_0__1_.mem_top_track_2.ccff_tail
rlabel metal1 13616 43622 13616 43622 0 sb_0__1_.mem_top_track_2.mem_out\[0\]
rlabel metal1 14398 39474 14398 39474 0 sb_0__1_.mem_top_track_2.mem_out\[1\]
rlabel metal1 5980 32810 5980 32810 0 sb_0__1_.mem_top_track_20.ccff_tail
rlabel metal1 14858 32878 14858 32878 0 sb_0__1_.mem_top_track_20.mem_out\[0\]
rlabel metal1 12282 32912 12282 32912 0 sb_0__1_.mem_top_track_20.mem_out\[1\]
rlabel metal1 5750 36652 5750 36652 0 sb_0__1_.mem_top_track_28.ccff_tail
rlabel metal2 11638 34272 11638 34272 0 sb_0__1_.mem_top_track_28.mem_out\[0\]
rlabel metal1 5750 34034 5750 34034 0 sb_0__1_.mem_top_track_28.mem_out\[1\]
rlabel metal1 8418 41242 8418 41242 0 sb_0__1_.mem_top_track_36.ccff_tail
rlabel metal1 12811 39474 12811 39474 0 sb_0__1_.mem_top_track_36.mem_out\[0\]
rlabel metal1 12489 38386 12489 38386 0 sb_0__1_.mem_top_track_36.mem_out\[1\]
rlabel metal1 9936 37910 9936 37910 0 sb_0__1_.mem_top_track_4.ccff_tail
rlabel metal1 15364 38386 15364 38386 0 sb_0__1_.mem_top_track_4.mem_out\[0\]
rlabel metal1 13570 36652 13570 36652 0 sb_0__1_.mem_top_track_4.mem_out\[1\]
rlabel metal1 13018 41480 13018 41480 0 sb_0__1_.mem_top_track_44.ccff_tail
rlabel metal1 17434 38420 17434 38420 0 sb_0__1_.mem_top_track_44.mem_out\[0\]
rlabel metal1 18032 41718 18032 41718 0 sb_0__1_.mem_top_track_52.mem_out\[0\]
rlabel metal2 17342 36448 17342 36448 0 sb_0__1_.mem_top_track_52.mem_out\[1\]
rlabel metal1 12834 36040 12834 36040 0 sb_0__1_.mem_top_track_6.mem_out\[0\]
rlabel metal2 10166 37655 10166 37655 0 sb_0__1_.mem_top_track_6.mem_out\[1\]
rlabel metal1 19642 6766 19642 6766 0 sb_0__1_.mux_bottom_track_1.out
rlabel metal2 15594 26316 15594 26316 0 sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 16606 25262 16606 25262 0 sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 12650 21352 12650 21352 0 sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 14996 20570 14996 20570 0 sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 14766 20944 14766 20944 0 sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 14582 17238 14582 17238 0 sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 16790 6766 16790 6766 0 sb_0__1_.mux_bottom_track_11.out
rlabel metal2 17342 29376 17342 29376 0 sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18584 32266 18584 32266 0 sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 16054 24242 16054 24242 0 sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 14812 24106 14812 24106 0 sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 16468 23834 16468 23834 0 sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 15962 23936 15962 23936 0 sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 15686 23494 15686 23494 0 sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 18584 8942 18584 8942 0 sb_0__1_.mux_bottom_track_13.out
rlabel metal1 19504 28526 19504 28526 0 sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20240 28526 20240 28526 0 sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 19550 25636 19550 25636 0 sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 20010 26316 20010 26316 0 sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 19918 24378 19918 24378 0 sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 19182 24038 19182 24038 0 sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 20838 7854 20838 7854 0 sb_0__1_.mux_bottom_track_21.out
rlabel metal2 20470 29104 20470 29104 0 sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22540 28186 22540 28186 0 sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 22908 25330 22908 25330 0 sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 25300 22950 25300 22950 0 sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 25024 23086 25024 23086 0 sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 21482 15062 21482 15062 0 sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 16054 8942 16054 8942 0 sb_0__1_.mux_bottom_track_29.out
rlabel metal1 17664 31450 17664 31450 0 sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19366 34918 19366 34918 0 sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 17802 28186 17802 28186 0 sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 17250 29206 17250 29206 0 sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 17112 27438 17112 27438 0 sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 16284 20434 16284 20434 0 sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 18400 6290 18400 6290 0 sb_0__1_.mux_bottom_track_3.out
rlabel metal2 18446 25415 18446 25415 0 sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18906 24922 18906 24922 0 sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 18170 24582 18170 24582 0 sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 18262 20026 18262 20026 0 sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 17526 17034 17526 17034 0 sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 13984 9622 13984 9622 0 sb_0__1_.mux_bottom_track_37.out
rlabel metal2 18538 34510 18538 34510 0 sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18768 32538 18768 32538 0 sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 16514 32538 16514 32538 0 sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 14076 27370 14076 27370 0 sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 13846 21998 13846 21998 0 sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 18492 10030 18492 10030 0 sb_0__1_.mux_bottom_track_45.out
rlabel metal2 22494 36210 22494 36210 0 sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21666 29614 21666 29614 0 sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 22402 32538 22402 32538 0 sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 20332 19822 20332 19822 0 sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 20010 8636 20010 8636 0 sb_0__1_.mux_bottom_track_5.out
rlabel metal2 21390 26588 21390 26588 0 sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22586 24922 22586 24922 0 sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20240 21998 20240 21998 0 sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 22632 20570 22632 20570 0 sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 22402 21250 22402 21250 0 sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 20608 14994 20608 14994 0 sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 10534 10030 10534 10030 0 sb_0__1_.mux_bottom_track_53.out
rlabel metal1 15042 37128 15042 37128 0 sb_0__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 15318 37060 15318 37060 0 sb_0__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 10304 36074 10304 36074 0 sb_0__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 18768 7854 18768 7854 0 sb_0__1_.mux_bottom_track_7.out
rlabel metal1 19228 26010 19228 26010 0 sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 19642 28254 19642 28254 0 sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 18492 21522 18492 21522 0 sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 18492 21658 18492 21658 0 sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 18676 23188 18676 23188 0 sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 18538 21114 18538 21114 0 sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 17158 19550 17158 19550 0 sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 24472 25262 24472 25262 0 sb_0__1_.mux_right_track_0.out
rlabel metal1 21896 31926 21896 31926 0 sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22540 31926 22540 31926 0 sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 23460 29682 23460 29682 0 sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 23092 28730 23092 28730 0 sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 23966 28764 23966 28764 0 sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 24288 32198 24288 32198 0 sb_0__1_.mux_right_track_10.out
rlabel metal1 19826 41650 19826 41650 0 sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19688 41446 19688 41446 0 sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19596 38318 19596 38318 0 sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 18032 36346 18032 36346 0 sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 22770 37383 22770 37383 0 sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 25070 28526 25070 28526 0 sb_0__1_.mux_right_track_12.out
rlabel metal1 20148 45798 20148 45798 0 sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 20194 39712 20194 39712 0 sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 17986 37094 17986 37094 0 sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 20608 38726 20608 38726 0 sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 23092 32198 23092 32198 0 sb_0__1_.mux_right_track_14.out
rlabel metal1 18170 42670 18170 42670 0 sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17618 42534 17618 42534 0 sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 16514 38522 16514 38522 0 sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 22034 32436 22034 32436 0 sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 20746 33082 20746 33082 0 sb_0__1_.mux_right_track_16.out
rlabel metal1 17250 43418 17250 43418 0 sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 16790 43078 16790 43078 0 sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14996 39066 14996 39066 0 sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 19550 32912 19550 32912 0 sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 21298 27642 21298 27642 0 sb_0__1_.mux_right_track_18.out
rlabel metal2 17342 44064 17342 44064 0 sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 16330 39066 16330 39066 0 sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14444 37978 14444 37978 0 sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 16836 38726 16836 38726 0 sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 24748 33830 24748 33830 0 sb_0__1_.mux_right_track_2.out
rlabel metal1 22586 42330 22586 42330 0 sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 22218 38624 22218 38624 0 sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 22586 38658 22586 38658 0 sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 25116 39338 25116 39338 0 sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 24104 39338 24104 39338 0 sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 24656 33966 24656 33966 0 sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 21666 25296 21666 25296 0 sb_0__1_.mux_right_track_20.out
rlabel metal1 15180 44234 15180 44234 0 sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 14950 35632 14950 35632 0 sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14352 33082 14352 33082 0 sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 15732 33286 15732 33286 0 sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 22954 20808 22954 20808 0 sb_0__1_.mux_right_track_22.out
rlabel metal2 13938 34867 13938 34867 0 sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13386 29682 13386 29682 0 sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 13156 29614 13156 29614 0 sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 17986 25330 17986 25330 0 sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 24564 18734 24564 18734 0 sb_0__1_.mux_right_track_24.out
rlabel metal1 14628 24242 14628 24242 0 sb_0__1_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 14260 24038 14260 24038 0 sb_0__1_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 18354 20842 18354 20842 0 sb_0__1_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 21252 19754 21252 19754 0 sb_0__1_.mux_right_track_26.out
rlabel metal1 13800 26282 13800 26282 0 sb_0__1_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13202 26418 13202 26418 0 sb_0__1_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 15640 23698 15640 23698 0 sb_0__1_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 21206 19822 21206 19822 0 sb_0__1_.mux_right_track_28.out
rlabel metal1 10626 27098 10626 27098 0 sb_0__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 8556 25738 8556 25738 0 sb_0__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 13478 22440 13478 22440 0 sb_0__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 21390 17578 21390 17578 0 sb_0__1_.mux_right_track_30.out
rlabel metal1 10350 25942 10350 25942 0 sb_0__1_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 10350 26384 10350 26384 0 sb_0__1_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_1_X
rlabel via2 15502 21539 15502 21539 0 sb_0__1_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 20562 16082 20562 16082 0 sb_0__1_.mux_right_track_32.out
rlabel metal2 10718 26316 10718 26316 0 sb_0__1_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 9706 24378 9706 24378 0 sb_0__1_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 15088 19822 15088 19822 0 sb_0__1_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 19918 16150 19918 16150 0 sb_0__1_.mux_right_track_34.out
rlabel metal1 13340 23766 13340 23766 0 sb_0__1_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 11592 23834 11592 23834 0 sb_0__1_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 16422 19346 16422 19346 0 sb_0__1_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 17618 12376 17618 12376 0 sb_0__1_.mux_right_track_36.out
rlabel metal1 8050 17646 8050 17646 0 sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 8740 12954 8740 12954 0 sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 8280 12818 8280 12818 0 sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 16238 12274 16238 12274 0 sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 22494 11526 22494 11526 0 sb_0__1_.mux_right_track_38.out
rlabel metal1 13708 13430 13708 13430 0 sb_0__1_.mux_right_track_38.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17365 11118 17365 11118 0 sb_0__1_.mux_right_track_38.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24564 27438 24564 27438 0 sb_0__1_.mux_right_track_4.out
rlabel metal1 22448 39338 22448 39338 0 sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21482 39304 21482 39304 0 sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21896 35122 21896 35122 0 sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 20470 34170 20470 34170 0 sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 23414 31620 23414 31620 0 sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 19826 11832 19826 11832 0 sb_0__1_.mux_right_track_40.out
rlabel metal1 17112 12954 17112 12954 0 sb_0__1_.mux_right_track_40.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 19596 12580 19596 12580 0 sb_0__1_.mux_right_track_40.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 22494 14042 22494 14042 0 sb_0__1_.mux_right_track_44.out
rlabel metal1 18400 15538 18400 15538 0 sb_0__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20010 15402 20010 15402 0 sb_0__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 23138 13838 23138 13838 0 sb_0__1_.mux_right_track_46.out
rlabel metal1 20102 16558 20102 16558 0 sb_0__1_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22678 13872 22678 13872 0 sb_0__1_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24334 9962 24334 9962 0 sb_0__1_.mux_right_track_48.out
rlabel metal1 21160 15470 21160 15470 0 sb_0__1_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 23506 13294 23506 13294 0 sb_0__1_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 22954 14246 22954 14246 0 sb_0__1_.mux_right_track_50.out
rlabel metal1 21298 18734 21298 18734 0 sb_0__1_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20148 15130 20148 15130 0 sb_0__1_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 21482 16490 21482 16490 0 sb_0__1_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 23000 8942 23000 8942 0 sb_0__1_.mux_right_track_52.out
rlabel metal2 21022 14688 21022 14688 0 sb_0__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21712 14042 21712 14042 0 sb_0__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24656 6766 24656 6766 0 sb_0__1_.mux_right_track_54.out
rlabel metal1 19734 12648 19734 12648 0 sb_0__1_.mux_right_track_54.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 22034 10404 22034 10404 0 sb_0__1_.mux_right_track_54.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 24334 9146 24334 9146 0 sb_0__1_.mux_right_track_56.out
rlabel metal2 18446 14110 18446 14110 0 sb_0__1_.mux_right_track_56.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20010 13498 20010 13498 0 sb_0__1_.mux_right_track_56.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 24794 28798 24794 28798 0 sb_0__1_.mux_right_track_6.out
rlabel metal2 23322 39893 23322 39893 0 sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22540 36346 22540 36346 0 sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20378 31994 20378 31994 0 sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 23690 36210 23690 36210 0 sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 23598 35258 23598 35258 0 sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 24334 36006 24334 36006 0 sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 24104 33830 24104 33830 0 sb_0__1_.mux_right_track_8.out
rlabel metal1 25024 41446 25024 41446 0 sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21482 40120 21482 40120 0 sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19688 37094 19688 37094 0 sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 23460 41514 23460 41514 0 sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 22724 40154 22724 40154 0 sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 23552 38726 23552 38726 0 sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 11868 48858 11868 48858 0 sb_0__1_.mux_top_track_0.out
rlabel metal1 10626 42534 10626 42534 0 sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 14168 43282 14168 43282 0 sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 15042 35530 15042 35530 0 sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 10902 39508 10902 39508 0 sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 12236 43418 12236 43418 0 sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 12558 41242 12558 41242 0 sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 11730 46614 11730 46614 0 sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 7912 44506 7912 44506 0 sb_0__1_.mux_top_track_10.out
rlabel metal1 10166 37230 10166 37230 0 sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 16882 36176 16882 36176 0 sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 10442 31756 10442 31756 0 sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 7636 31892 7636 31892 0 sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 9016 37162 9016 37162 0 sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 9982 35428 9982 35428 0 sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 7820 44370 7820 44370 0 sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 7774 42534 7774 42534 0 sb_0__1_.mux_top_track_12.out
rlabel metal1 13064 33966 13064 33966 0 sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 14168 33898 14168 33898 0 sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 9614 32810 9614 32810 0 sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 11638 34170 11638 34170 0 sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 10028 33082 10028 33082 0 sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 9660 36890 9660 36890 0 sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 11684 51986 11684 51986 0 sb_0__1_.mux_top_track_2.out
rlabel metal1 14996 39406 14996 39406 0 sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 16422 35190 16422 35190 0 sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 11960 33626 11960 33626 0 sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 14398 39610 14398 39610 0 sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 12466 39066 12466 39066 0 sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 11684 42330 11684 42330 0 sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 7314 42534 7314 42534 0 sb_0__1_.mux_top_track_20.out
rlabel metal1 14076 34714 14076 34714 0 sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17664 30090 17664 30090 0 sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 8418 31790 8418 31790 0 sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 10764 33014 10764 33014 0 sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 8050 31926 8050 31926 0 sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 7682 38329 7682 38329 0 sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 6164 43418 6164 43418 0 sb_0__1_.mux_top_track_28.out
rlabel metal2 9614 35292 9614 35292 0 sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 12374 32912 12374 32912 0 sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 9154 35530 9154 35530 0 sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 5474 36754 5474 36754 0 sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 5382 43282 5382 43282 0 sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 6624 51374 6624 51374 0 sb_0__1_.mux_top_track_36.out
rlabel metal1 12558 38182 12558 38182 0 sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 10902 38454 10902 38454 0 sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 8464 38522 8464 38522 0 sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 7590 41786 7590 41786 0 sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 9982 48110 9982 48110 0 sb_0__1_.mux_top_track_4.out
rlabel metal1 13984 36890 13984 36890 0 sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 15916 33354 15916 33354 0 sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 10028 31450 10028 31450 0 sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 12742 36890 12742 36890 0 sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 10350 37128 10350 37128 0 sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 9798 42262 9798 42262 0 sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 6808 51442 6808 51442 0 sb_0__1_.mux_top_track_44.out
rlabel metal2 12466 42432 12466 42432 0 sb_0__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 11776 38522 11776 38522 0 sb_0__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 12006 42568 12006 42568 0 sb_0__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 9660 45254 9660 45254 0 sb_0__1_.mux_top_track_52.out
rlabel metal1 21114 36890 21114 36890 0 sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19504 36890 19504 36890 0 sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 15778 35258 15778 35258 0 sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 14720 39542 14720 39542 0 sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 8602 48110 8602 48110 0 sb_0__1_.mux_top_track_6.out
rlabel metal1 9936 38386 9936 38386 0 sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 17158 36601 17158 36601 0 sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 12926 30906 12926 30906 0 sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 7728 32198 7728 32198 0 sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 9430 38522 9430 38522 0 sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 8786 34714 8786 34714 0 sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 8418 42534 8418 42534 0 sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 24932 3502 24932 3502 0 test_enable_bottom_in
rlabel metal2 25438 1639 25438 1639 0 test_enable_bottom_out
rlabel metal1 24656 51986 24656 51986 0 test_enable_right_in
rlabel metal1 24656 51510 24656 51510 0 test_enable_top_in
rlabel metal1 24426 53686 24426 53686 0 test_enable_top_out
rlabel metal1 1334 45594 1334 45594 0 top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal1 1518 48042 1518 48042 0 top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal1 1288 50422 1288 50422 0 top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal1 4002 52564 4002 52564 0 top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
<< properties >>
string FIXED_BBOX 0 0 27000 57000
<< end >>
