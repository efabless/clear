* NGSPICE file created from cbx_1__0_.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_1 abstract view
.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_4 abstract view
.subckt sky130_fd_sc_hd__or2b_4 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_4 abstract view
.subckt sky130_fd_sc_hd__ebufn_4 A TE_B VGND VNB VPB VPWR Z
.ends

.subckt cbx_1__0_ IO_ISOL_N SC_IN_BOT SC_IN_TOP SC_OUT_BOT SC_OUT_TOP VGND VPWR bottom_grid_pin_0_
+ bottom_grid_pin_10_ bottom_grid_pin_12_ bottom_grid_pin_14_ bottom_grid_pin_16_
+ bottom_grid_pin_2_ bottom_grid_pin_4_ bottom_grid_pin_6_ bottom_grid_pin_8_ ccff_head
+ ccff_tail chanx_left_in[0] chanx_left_in[10] chanx_left_in[11] chanx_left_in[12]
+ chanx_left_in[13] chanx_left_in[14] chanx_left_in[15] chanx_left_in[16] chanx_left_in[17]
+ chanx_left_in[18] chanx_left_in[19] chanx_left_in[1] chanx_left_in[2] chanx_left_in[3]
+ chanx_left_in[4] chanx_left_in[5] chanx_left_in[6] chanx_left_in[7] chanx_left_in[8]
+ chanx_left_in[9] chanx_left_out[0] chanx_left_out[10] chanx_left_out[11] chanx_left_out[12]
+ chanx_left_out[13] chanx_left_out[14] chanx_left_out[15] chanx_left_out[16] chanx_left_out[17]
+ chanx_left_out[18] chanx_left_out[19] chanx_left_out[1] chanx_left_out[2] chanx_left_out[3]
+ chanx_left_out[4] chanx_left_out[5] chanx_left_out[6] chanx_left_out[7] chanx_left_out[8]
+ chanx_left_out[9] chanx_right_in[0] chanx_right_in[10] chanx_right_in[11] chanx_right_in[12]
+ chanx_right_in[13] chanx_right_in[14] chanx_right_in[15] chanx_right_in[16] chanx_right_in[17]
+ chanx_right_in[18] chanx_right_in[19] chanx_right_in[1] chanx_right_in[2] chanx_right_in[3]
+ chanx_right_in[4] chanx_right_in[5] chanx_right_in[6] chanx_right_in[7] chanx_right_in[8]
+ chanx_right_in[9] chanx_right_out[0] chanx_right_out[10] chanx_right_out[11] chanx_right_out[12]
+ chanx_right_out[13] chanx_right_out[14] chanx_right_out[15] chanx_right_out[16]
+ chanx_right_out[17] chanx_right_out[18] chanx_right_out[19] chanx_right_out[1] chanx_right_out[2]
+ chanx_right_out[3] chanx_right_out[4] chanx_right_out[5] chanx_right_out[6] chanx_right_out[7]
+ chanx_right_out[8] chanx_right_out[9] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[0] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[1]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[2] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[3] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[4]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[5] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[6] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[7]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[8] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[0] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[1]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[2] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[3] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[4]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[5] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[6] gfpga_pad_EMBEDDED_IO_HD_SOC_IN[7]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[8] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[0] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[1]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[2] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[3] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[4]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[5] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[6] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[7]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[8] prog_clk_0_N_in prog_clk_0_W_out top_width_0_height_0__pin_0_
+ top_width_0_height_0__pin_10_ top_width_0_height_0__pin_11_lower top_width_0_height_0__pin_11_upper
+ top_width_0_height_0__pin_12_ top_width_0_height_0__pin_13_lower top_width_0_height_0__pin_13_upper
+ top_width_0_height_0__pin_14_ top_width_0_height_0__pin_15_lower top_width_0_height_0__pin_15_upper
+ top_width_0_height_0__pin_16_ top_width_0_height_0__pin_17_lower top_width_0_height_0__pin_17_upper
+ top_width_0_height_0__pin_1_lower top_width_0_height_0__pin_1_upper top_width_0_height_0__pin_2_
+ top_width_0_height_0__pin_3_lower top_width_0_height_0__pin_3_upper top_width_0_height_0__pin_4_
+ top_width_0_height_0__pin_5_lower top_width_0_height_0__pin_5_upper top_width_0_height_0__pin_6_
+ top_width_0_height_0__pin_7_lower top_width_0_height_0__pin_7_upper top_width_0_height_0__pin_8_
+ top_width_0_height_0__pin_9_lower top_width_0_height_0__pin_9_upper
XANTENNA_mux_top_ipin_7.mux_l1_in_0__A1 chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_1.mux_l1_in_1_ chanx_right_in[3] chanx_left_in[3] mux_top_ipin_1.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_1.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_top_ipin_7.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_8.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
X_83_ SC_IN_BOT VGND VGND VPWR VPWR SC_OUT_TOP sky130_fd_sc_hd__buf_2
XFILLER_13_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE_A
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_5.mux_l1_in_2__A1 chanx_left_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_158 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_66_ _66_/A VGND VGND VPWR VPWR gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[2] sky130_fd_sc_hd__buf_2
Xmux_top_ipin_6.mux_l2_in_0_ mux_top_ipin_6.mux_l1_in_1_/X mux_top_ipin_6.mux_l1_in_0_/X
+ mux_top_ipin_6.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_top_ipin_6.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_49_ chanx_left_in[14] VGND VGND VPWR VPWR chanx_right_out[14] sky130_fd_sc_hd__buf_2
XFILLER_18_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_6.mux_l1_in_1_ chanx_right_in[2] chanx_left_in[2] mux_top_ipin_6.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_6.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_3.mux_l2_in_3__A1 chanx_right_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_2.mux_l1_in_0__A0 chanx_right_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_150 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE_A
+ top_width_0_height_0__pin_10_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_ipin_0.mux_l1_in_2__A0 chanx_right_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_ipin_1.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_top_ipin_1.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_1.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XTAP_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_156 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_24 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_82_ SC_IN_TOP VGND VGND VPWR VPWR SC_OUT_BOT sky130_fd_sc_hd__buf_2
XANTENNA_mux_top_ipin_0.mux_l2_in_1__A0 chanx_left_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_65_ _65_/A VGND VGND VPWR VPWR gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[1] sky130_fd_sc_hd__buf_2
XFILLER_5_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_prog_clk_0_W_FTB01_A prog_clk_0_N_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_48_ chanx_left_in[13] VGND VGND VPWR VPWR chanx_right_out[13] sky130_fd_sc_hd__buf_2
XANTENNA_logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE_B_N
+ IO_ISOL_N VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_6.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_top_ipin_6.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_6.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_top_ipin_2.mux_l1_in_0__A1 chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_ipin_0.mux_l1_in_2__A1 chanx_left_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_ipin_7.mux_l2_in_2__A0 chanx_left_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_81_ top_width_0_height_0__pin_9_lower VGND VGND VPWR VPWR top_width_0_height_0__pin_9_upper
+ sky130_fd_sc_hd__buf_2
XFILLER_8_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_36 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_64_ _64_/A VGND VGND VPWR VPWR gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[0] sky130_fd_sc_hd__buf_2
Xlogical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR _60_/A
+ VGND VGND VPWR VPWR logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y
+ sky130_fd_sc_hd__inv_1
XFILLER_5_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_4.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_4.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR bottom_grid_pin_8_ sky130_fd_sc_hd__buf_4
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_47_ chanx_left_in[12] VGND VGND VPWR VPWR chanx_right_out[12] sky130_fd_sc_hd__buf_2
XFILLER_15_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_80_ top_width_0_height_0__pin_7_lower VGND VGND VPWR VPWR top_width_0_height_0__pin_7_upper
+ sky130_fd_sc_hd__buf_2
XANTENNA_mux_top_ipin_7.mux_l2_in_2__A1 chanx_right_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_59 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_63_ _63_/A VGND VGND VPWR VPWR gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[8] sky130_fd_sc_hd__buf_2
Xprog_clk_0_FTB00 prog_clk_0_N_in VGND VGND VPWR VPWR prog_clk_0_FTB00/X sky130_fd_sc_hd__buf_8
XANTENNA_mux_top_ipin_4.mux_l1_in_1__A0 chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE_B_N
+ IO_ISOL_N VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_46_ chanx_left_in[11] VGND VGND VPWR VPWR chanx_right_out[11] sky130_fd_sc_hd__buf_2
XFILLER_18_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29_ chanx_right_in[14] VGND VGND VPWR VPWR chanx_left_out[14] sky130_fd_sc_hd__buf_2
XFILLER_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_ipin_2.mux_l2_in_2__A0 chanx_left_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20__A chanx_right_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xlogical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
+ prog_clk_0_FTB00/X logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A
+ VGND VGND VPWR VPWR logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A
+ sky130_fd_sc_hd__dfxtp_1
XTAP_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xlogical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A
+ IO_ISOL_N VGND VGND VPWR VPWR _60_/A sky130_fd_sc_hd__or2b_4
XFILLER_21_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_ipin_2.mux_l2_in_3_ _11_/HI chanx_right_in[18] mux_top_ipin_2.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_2.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_62_ _62_/A VGND VGND VPWR VPWR gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[7] sky130_fd_sc_hd__buf_2
XFILLER_2_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_4.mux_l1_in_1__A1 chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE_A
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_45_ chanx_left_in[10] VGND VGND VPWR VPWR chanx_right_out[10] sky130_fd_sc_hd__buf_2
Xmux_top_ipin_2.mux_l4_in_0_ mux_top_ipin_2.mux_l3_in_1_/X mux_top_ipin_2.mux_l3_in_0_/X
+ mux_top_ipin_2.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_2.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA__23__A chanx_right_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE_A
+ top_width_0_height_0__pin_8_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_28_ chanx_right_in[13] VGND VGND VPWR VPWR chanx_left_out[13] sky130_fd_sc_hd__buf_2
XANTENNA_logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE_A
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_7.mux_l2_in_3_ _16_/HI chanx_right_in[17] mux_top_ipin_7.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_7.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XANTENNA__18__A chanx_right_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_2.mux_l3_in_1_ mux_top_ipin_2.mux_l2_in_3_/X mux_top_ipin_2.mux_l2_in_2_/X
+ mux_top_ipin_2.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_2.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_2.mux_l2_in_2__A1 chanx_right_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_ipin_2.mux_l2_in_2_ chanx_left_in[18] chanx_right_in[12] mux_top_ipin_2.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_2.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XANTENNA__31__A chanx_right_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_7.mux_l4_in_0_ mux_top_ipin_7.mux_l3_in_1_/X mux_top_ipin_7.mux_l3_in_0_/X
+ mux_top_ipin_7.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_7.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__26__A chanx_right_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_61_ _61_/A VGND VGND VPWR VPWR gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[6] sky130_fd_sc_hd__buf_2
XFILLER_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_7.mux_l3_in_1_ mux_top_ipin_7.mux_l2_in_3_/X mux_top_ipin_7.mux_l2_in_2_/X
+ mux_top_ipin_7.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_7.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_44_ chanx_left_in[9] VGND VGND VPWR VPWR chanx_right_out[9] sky130_fd_sc_hd__buf_2
XFILLER_1_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27_ chanx_right_in[12] VGND VGND VPWR VPWR chanx_left_out[12] sky130_fd_sc_hd__buf_2
Xmux_top_ipin_7.mux_l2_in_2_ chanx_left_in[17] chanx_right_in[11] mux_top_ipin_7.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_7.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xlogical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
+ prog_clk_0_FTB00/X logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A
+ VGND VGND VPWR VPWR ccff_tail sky130_fd_sc_hd__dfxtp_1
XFILLER_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__34__A chanx_right_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_2.mux_l3_in_0_ mux_top_ipin_2.mux_l2_in_1_/X mux_top_ipin_2.mux_l2_in_0_/X
+ mux_top_ipin_2.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_2.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_8.mux_l1_in_0__A0 chanx_right_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__29__A chanx_right_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_6.mux_l1_in_2__A0 chanx_right_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_2.mux_l2_in_1_ chanx_left_in[12] mux_top_ipin_2.mux_l1_in_2_/X mux_top_ipin_2.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_2.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__42__A chanx_left_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_60_ _60_/A VGND VGND VPWR VPWR gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[5] sky130_fd_sc_hd__buf_2
XFILLER_4_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_2.mux_l1_in_2_ chanx_right_in[6] chanx_left_in[6] mux_top_ipin_2.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_2.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_6.mux_l2_in_1__A0 chanx_left_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_7.mux_l3_in_0_ mux_top_ipin_7.mux_l2_in_1_/X mux_top_ipin_7.mux_l2_in_0_/X
+ mux_top_ipin_7.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_7.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA__37__A chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_7.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_7.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR bottom_grid_pin_14_ sky130_fd_sc_hd__buf_4
X_43_ chanx_left_in[8] VGND VGND VPWR VPWR chanx_right_out[8] sky130_fd_sc_hd__buf_2
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_7.mux_l2_in_1_ chanx_left_in[11] mux_top_ipin_7.mux_l1_in_2_/X mux_top_ipin_7.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_7.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
X_26_ chanx_right_in[11] VGND VGND VPWR VPWR chanx_left_out[11] sky130_fd_sc_hd__buf_2
XFILLER_1_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__50__A chanx_left_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09_ VGND VGND VPWR VPWR _09_/HI _09_/LO sky130_fd_sc_hd__conb_1
XANTENNA_mux_top_ipin_8.mux_l1_in_0__A1 chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__45__A chanx_left_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_ipin_7.mux_l1_in_2_ chanx_right_in[7] chanx_left_in[7] mux_top_ipin_7.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_7.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_6.mux_l1_in_2__A1 chanx_left_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_2.mux_l2_in_0_ mux_top_ipin_2.mux_l1_in_1_/X mux_top_ipin_2.mux_l1_in_0_/X
+ mux_top_ipin_2.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_top_ipin_2.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xlogical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR _55_/A
+ VGND VGND VPWR VPWR logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y
+ sky130_fd_sc_hd__inv_1
XFILLER_4_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_2.mux_l1_in_1_ chanx_right_in[2] chanx_left_in[2] mux_top_ipin_2.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_2.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_top_ipin_1.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_top_ipin_1.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA__53__A chanx_left_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_42_ chanx_left_in[7] VGND VGND VPWR VPWR chanx_right_out[7] sky130_fd_sc_hd__buf_2
XANTENNA_mux_top_ipin_4.mux_l2_in_3__A1 chanx_right_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_3.mux_l1_in_0__A0 chanx_right_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__48__A chanx_left_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_7.mux_l2_in_0_ mux_top_ipin_7.mux_l1_in_1_/X mux_top_ipin_7.mux_l1_in_0_/X
+ mux_top_ipin_7.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_top_ipin_7.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_25_ chanx_right_in[10] VGND VGND VPWR VPWR chanx_left_out[10] sky130_fd_sc_hd__buf_2
XFILLER_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_1.mux_l1_in_2__A0 chanx_right_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_ipin_7.mux_l1_in_1_ chanx_right_in[3] chanx_left_in[3] mux_top_ipin_7.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_7.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xlogical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A
+ IO_ISOL_N VGND VGND VPWR VPWR _58_/A sky130_fd_sc_hd__or2b_4
XANTENNA_mux_top_ipin_1.mux_l2_in_1__A0 chanx_left_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_top_ipin_4.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_top_ipin_4.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_8_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE_A
+ top_width_0_height_0__pin_6_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_top_ipin_1.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_1.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_2.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_top_ipin_2.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_2.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
X_41_ chanx_left_in[6] VGND VGND VPWR VPWR chanx_right_out[6] sky130_fd_sc_hd__buf_2
XANTENNA_mux_top_ipin_3.mux_l1_in_0__A1 chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_24_ chanx_right_in[9] VGND VGND VPWR VPWR chanx_left_out[9] sky130_fd_sc_hd__buf_2
XFILLER_19_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_1.mux_l1_in_2__A1 chanx_left_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_top_ipin_7.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_top_ipin_7.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_0.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR bottom_grid_pin_0_ sky130_fd_sc_hd__buf_4
XFILLER_21_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_7.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_top_ipin_7.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_7.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XTAP_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_8.mux_l2_in_2__A0 chanx_left_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE_A
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xlogical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE gfpga_pad_EMBEDDED_IO_HD_SOC_IN[6]
+ logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y VGND
+ VGND VPWR VPWR top_width_0_height_0__pin_13_lower sky130_fd_sc_hd__ebufn_4
Xmem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_top_ipin_4.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_4.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_12_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_top_ipin_1.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_1.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
X_40_ chanx_left_in[5] VGND VGND VPWR VPWR chanx_right_out[5] sky130_fd_sc_hd__buf_2
XANTENNA__80__A top_width_0_height_0__pin_7_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23_ chanx_right_in[8] VGND VGND VPWR VPWR chanx_left_out[8] sky130_fd_sc_hd__buf_2
Xmem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_top_ipin_7.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_7.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_21_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_8.mux_l2_in_2__A1 chanx_right_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xlogical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE gfpga_pad_EMBEDDED_IO_HD_SOC_IN[3]
+ logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y VGND
+ VGND VPWR VPWR top_width_0_height_0__pin_7_lower sky130_fd_sc_hd__ebufn_4
XFILLER_7_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_154 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_top_ipin_4.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_4.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA__83__A SC_IN_BOT VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_5.mux_l1_in_1__A0 chanx_right_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xlogical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
+ prog_clk_0_FTB00/X logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A
+ VGND VGND VPWR VPWR logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__78__A top_width_0_height_0__pin_3_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_top_ipin_0.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_1.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
Xlogical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR _59_/A
+ VGND VGND VPWR VPWR logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y
+ sky130_fd_sc_hd__inv_1
X_22_ chanx_right_in[7] VGND VGND VPWR VPWR chanx_left_out[7] sky130_fd_sc_hd__buf_2
XANTENNA_mux_top_ipin_3.mux_l2_in_2__A0 chanx_left_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_top_ipin_7.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_7.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_10_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xlogical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE gfpga_pad_EMBEDDED_IO_HD_SOC_IN[0]
+ logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y VGND
+ VGND VPWR VPWR top_width_0_height_0__pin_1_lower sky130_fd_sc_hd__ebufn_4
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__86__A chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_top_ipin_3.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_4.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_12_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_5.mux_l1_in_1__A1 chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_top_ipin_3.mux_l2_in_3_ _12_/HI chanx_right_in[19] mux_top_ipin_3.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_3.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21_ chanx_right_in[6] VGND VGND VPWR VPWR chanx_left_out[6] sky130_fd_sc_hd__buf_2
XFILLER_1_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_3.mux_l2_in_2__A1 chanx_right_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_top_ipin_6.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_7.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_18_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_3.mux_l4_in_0_ mux_top_ipin_3.mux_l3_in_1_/X mux_top_ipin_3.mux_l3_in_0_/X
+ mux_top_ipin_3.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_3.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE_A
+ top_width_0_height_0__pin_4_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_0.mux_l1_in_1__A0 chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_top_ipin_8.mux_l2_in_3_ _17_/HI chanx_right_in[18] mux_top_ipin_8.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_8.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
Xlogical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A
+ IO_ISOL_N VGND VGND VPWR VPWR _56_/A sky130_fd_sc_hd__or2b_4
Xmux_top_ipin_3.mux_l3_in_1_ mux_top_ipin_3.mux_l2_in_3_/X mux_top_ipin_3.mux_l2_in_2_/X
+ mux_top_ipin_3.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_3.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_3.mux_l2_in_2_ chanx_left_in[19] chanx_right_in[13] mux_top_ipin_3.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_3.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_21 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_top_ipin_8.mux_l4_in_0_ mux_top_ipin_8.mux_l3_in_1_/X mux_top_ipin_8.mux_l3_in_0_/X
+ mux_top_ipin_8.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_8.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20_ chanx_right_in[5] VGND VGND VPWR VPWR chanx_left_out[5] sky130_fd_sc_hd__buf_2
XFILLER_19_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_8.mux_l3_in_1_ mux_top_ipin_8.mux_l2_in_3_/X mux_top_ipin_8.mux_l2_in_2_/X
+ mux_top_ipin_8.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_8.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XTAP_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_ipin_7.mux_l1_in_2__A0 chanx_right_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_8.mux_l2_in_2_ chanx_left_in[18] chanx_right_in[12] mux_top_ipin_8.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_8.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_3.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR bottom_grid_pin_6_ sky130_fd_sc_hd__buf_4
XANTENNA_mux_top_ipin_0.mux_l1_in_1__A1 chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_3.mux_l3_in_0_ mux_top_ipin_3.mux_l2_in_1_/X mux_top_ipin_3.mux_l2_in_0_/X
+ mux_top_ipin_3.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_3.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_98 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_7.mux_l2_in_1__A0 chanx_left_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_3.mux_l2_in_1_ chanx_left_in[13] mux_top_ipin_3.mux_l1_in_2_/X mux_top_ipin_3.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_3.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE_A
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_3.mux_l1_in_2_ chanx_right_in[7] chanx_left_in[7] mux_top_ipin_3.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_3.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xlogical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR _63_/A
+ VGND VGND VPWR VPWR logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y
+ sky130_fd_sc_hd__inv_1
X_79_ top_width_0_height_0__pin_5_lower VGND VGND VPWR VPWR top_width_0_height_0__pin_5_upper
+ sky130_fd_sc_hd__buf_2
XTAP_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_8.mux_l3_in_0_ mux_top_ipin_8.mux_l2_in_1_/X mux_top_ipin_8.mux_l2_in_0_/X
+ mux_top_ipin_8.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_8.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_19_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_top_ipin_7.mux_l1_in_2__A1 chanx_left_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_8.mux_l2_in_1_ chanx_left_in[12] mux_top_ipin_8.mux_l1_in_2_/X mux_top_ipin_8.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_8.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_ipin_8.mux_l1_in_2_ chanx_right_in[8] chanx_left_in[8] mux_top_ipin_8.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_8.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_5.mux_l2_in_3__A1 chanx_right_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_3.mux_l2_in_0_ mux_top_ipin_3.mux_l1_in_1_/X mux_top_ipin_3.mux_l1_in_0_/X
+ mux_top_ipin_3.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_top_ipin_3.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_ipin_4.mux_l1_in_0__A0 chanx_right_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_2.mux_l1_in_2__A0 chanx_right_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_78_ top_width_0_height_0__pin_3_lower VGND VGND VPWR VPWR top_width_0_height_0__pin_3_upper
+ sky130_fd_sc_hd__buf_2
Xmux_top_ipin_3.mux_l1_in_1_ chanx_right_in[3] chanx_left_in[3] mux_top_ipin_3.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_3.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XTAP_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_ipin_2.mux_l2_in_1__A0 chanx_left_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_ipin_8.mux_l2_in_0_ mux_top_ipin_8.mux_l1_in_1_/X mux_top_ipin_8.mux_l1_in_0_/X
+ mux_top_ipin_8.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_top_ipin_8.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xlogical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
+ prog_clk_0_FTB00/X logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A
+ VGND VGND VPWR VPWR logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A
+ sky130_fd_sc_hd__dfxtp_1
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_prog_clk_0_FTB00_A prog_clk_0_N_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_8.mux_l1_in_1_ chanx_right_in[2] chanx_left_in[2] mux_top_ipin_8.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_8.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_ipin_4.mux_l1_in_0__A1 chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE_A
+ top_width_0_height_0__pin_2_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_2.mux_l1_in_2__A1 chanx_left_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_77_ top_width_0_height_0__pin_1_lower VGND VGND VPWR VPWR top_width_0_height_0__pin_1_upper
+ sky130_fd_sc_hd__buf_2
Xmux_top_ipin_3.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_top_ipin_3.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_3.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XTAP_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xlogical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE ccff_tail
+ IO_ISOL_N VGND VGND VPWR VPWR _63_/A sky130_fd_sc_hd__or2b_4
XANTENNA_mux_top_ipin_0.mux_l2_in_3__A1 chanx_right_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21__A chanx_right_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_8.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_top_ipin_8.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_8.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_76_ top_width_0_height_0__pin_17_lower VGND VGND VPWR VPWR top_width_0_height_0__pin_17_upper
+ sky130_fd_sc_hd__buf_2
XTAP_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24__A chanx_right_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_59_ _59_/A VGND VGND VPWR VPWR gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[4] sky130_fd_sc_hd__buf_2
XANTENNA__19__A chanx_right_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_6.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_6.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR bottom_grid_pin_12_ sky130_fd_sc_hd__buf_4
XANTENNA_mux_top_ipin_6.mux_l1_in_1__A0 chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__32__A chanx_right_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__27__A chanx_right_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_4.mux_l2_in_2__A0 chanx_left_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_75_ top_width_0_height_0__pin_15_lower VGND VGND VPWR VPWR top_width_0_height_0__pin_15_upper
+ sky130_fd_sc_hd__buf_2
XTAP_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_156 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__40__A chanx_left_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_58_ _58_/A VGND VGND VPWR VPWR gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[3] sky130_fd_sc_hd__buf_2
XFILLER_21_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__35__A chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE_A
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_6.mux_l1_in_1__A1 chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_100 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__43__A chanx_left_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_4.mux_l2_in_2__A1 chanx_right_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__38__A chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xlogical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR _58_/A
+ VGND VGND VPWR VPWR logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y
+ sky130_fd_sc_hd__inv_1
X_74_ top_width_0_height_0__pin_13_lower VGND VGND VPWR VPWR top_width_0_height_0__pin_13_upper
+ sky130_fd_sc_hd__buf_2
XTAP_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_ipin_4.mux_l2_in_3_ _13_/HI chanx_right_in[14] mux_top_ipin_4.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_4.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XTAP_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_ipin_1.mux_l1_in_1__A0 chanx_right_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_57_ _57_/A VGND VGND VPWR VPWR gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[2] sky130_fd_sc_hd__buf_2
XANTENNA__51__A chanx_left_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__46__A chanx_left_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_top_ipin_0.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_top_ipin_0.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xlogical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE top_width_0_height_0__pin_0_
+ _55_/A VGND VGND VPWR VPWR _64_/A sky130_fd_sc_hd__ebufn_4
Xmux_top_ipin_4.mux_l4_in_0_ mux_top_ipin_4.mux_l3_in_1_/X mux_top_ipin_4.mux_l3_in_0_/X
+ mux_top_ipin_4.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_4.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE_A
+ top_width_0_height_0__pin_0_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_4.mux_l3_in_1_ mux_top_ipin_4.mux_l2_in_3_/X mux_top_ipin_4.mux_l2_in_2_/X
+ mux_top_ipin_4.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_4.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xlogical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
+ prog_clk_0_FTB00/X logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A
+ VGND VGND VPWR VPWR logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__54__A chanx_left_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_73_ top_width_0_height_0__pin_11_lower VGND VGND VPWR VPWR top_width_0_height_0__pin_11_upper
+ sky130_fd_sc_hd__buf_2
XTAP_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_ipin_4.mux_l2_in_2_ chanx_left_in[14] chanx_right_in[8] mux_top_ipin_4.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_4.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XTAP_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_8.mux_l1_in_2__A0 chanx_right_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_1.mux_l1_in_1__A1 chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_top_ipin_3.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_top_ipin_3.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xprog_clk_0_W_FTB01 prog_clk_0_N_in VGND VGND VPWR VPWR prog_clk_0_W_out sky130_fd_sc_hd__buf_4
XANTENNA__49__A chanx_left_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_56_ _56_/A VGND VGND VPWR VPWR gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[1] sky130_fd_sc_hd__buf_2
XFILLER_2_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_52 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xlogical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A
+ IO_ISOL_N VGND VGND VPWR VPWR _61_/A sky130_fd_sc_hd__or2b_4
X_39_ chanx_left_in[4] VGND VGND VPWR VPWR chanx_right_out[4] sky130_fd_sc_hd__buf_2
XANTENNA_mux_top_ipin_8.mux_l2_in_1__A0 chanx_left_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_top_ipin_0.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_0.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_ipin_4.mux_l3_in_0_ mux_top_ipin_4.mux_l2_in_1_/X mux_top_ipin_4.mux_l2_in_0_/X
+ mux_top_ipin_4.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_4.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xlogical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE gfpga_pad_EMBEDDED_IO_HD_SOC_IN[8]
+ logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y VGND
+ VGND VPWR VPWR top_width_0_height_0__pin_17_lower sky130_fd_sc_hd__ebufn_4
Xmem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_top_ipin_6.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_top_ipin_6.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_5_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_72_ _72_/A VGND VGND VPWR VPWR gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[8] sky130_fd_sc_hd__buf_2
XTAP_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_ipin_8.mux_l1_in_2__A1 chanx_left_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_4.mux_l2_in_1_ chanx_left_in[8] mux_top_ipin_4.mux_l1_in_2_/X mux_top_ipin_4.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_4.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_top_ipin_3.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_3.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
X_55_ _55_/A VGND VGND VPWR VPWR gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[0] sky130_fd_sc_hd__buf_2
XFILLER_2_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_73 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xlogical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE top_width_0_height_0__pin_2_
+ _56_/A VGND VGND VPWR VPWR _65_/A sky130_fd_sc_hd__ebufn_4
Xmux_top_ipin_4.mux_l1_in_2_ chanx_right_in[4] chanx_left_in[4] mux_top_ipin_4.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_4.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_38_ chanx_left_in[3] VGND VGND VPWR VPWR chanx_right_out[3] sky130_fd_sc_hd__buf_2
XFILLER_11_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_top_ipin_0.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_0.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_8_52 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_ipin_6.mux_l2_in_3__A1 chanx_right_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__73__A top_width_0_height_0__pin_11_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_5.mux_l1_in_0__A0 chanx_right_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xlogical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE gfpga_pad_EMBEDDED_IO_HD_SOC_IN[5]
+ logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y VGND
+ VGND VPWR VPWR top_width_0_height_0__pin_11_lower sky130_fd_sc_hd__ebufn_4
XANTENNA_mux_top_ipin_3.mux_l1_in_2__A0 chanx_right_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_top_ipin_6.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_6.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
X_71_ _71_/A VGND VGND VPWR VPWR gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[7] sky130_fd_sc_hd__buf_2
XTAP_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_ipin_4.mux_l2_in_0_ mux_top_ipin_4.mux_l1_in_1_/X mux_top_ipin_4.mux_l1_in_0_/X
+ mux_top_ipin_4.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_top_ipin_4.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XTAP_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__81__A top_width_0_height_0__pin_9_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_3.mux_l2_in_1__A0 chanx_left_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_54_ chanx_left_in[19] VGND VGND VPWR VPWR chanx_right_out[19] sky130_fd_sc_hd__buf_2
Xmem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_top_ipin_3.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_3.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
Xlogical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR _62_/A
+ VGND VGND VPWR VPWR logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y
+ sky130_fd_sc_hd__inv_1
XFILLER_14_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_4.mux_l1_in_1_ chanx_right_in[2] chanx_left_in[2] mux_top_ipin_4.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_4.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_37_ chanx_left_in[2] VGND VGND VPWR VPWR chanx_right_out[2] sky130_fd_sc_hd__buf_2
XFILLER_11_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X ccff_head VGND VGND
+ VPWR VPWR mux_top_ipin_0.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_8_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_ipin_5.mux_l1_in_0__A1 chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xlogical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE gfpga_pad_EMBEDDED_IO_HD_SOC_IN[2]
+ logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y VGND
+ VGND VPWR VPWR top_width_0_height_0__pin_5_lower sky130_fd_sc_hd__ebufn_4
XANTENNA_mux_top_ipin_3.mux_l1_in_2__A1 chanx_left_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__84__A chanx_right_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_top_ipin_6.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_6.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE_A
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__79__A top_width_0_height_0__pin_5_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_70_ _70_/A VGND VGND VPWR VPWR gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[6] sky130_fd_sc_hd__buf_2
XTAP_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_53_ chanx_left_in[18] VGND VGND VPWR VPWR chanx_right_out[18] sky130_fd_sc_hd__buf_2
Xmem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_top_ipin_2.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_3.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
Xlogical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE top_width_0_height_0__pin_4_
+ _57_/A VGND VGND VPWR VPWR _66_/A sky130_fd_sc_hd__ebufn_4
XANTENNA_mux_top_ipin_1.mux_l2_in_3__A1 chanx_right_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_top_ipin_4.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_top_ipin_4.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_4.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36_ chanx_left_in[1] VGND VGND VPWR VPWR chanx_right_out[1] sky130_fd_sc_hd__buf_2
XANTENNA_mux_top_ipin_0.mux_l1_in_0__A0 chanx_right_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19_ chanx_right_in[4] VGND VGND VPWR VPWR chanx_left_out[4] sky130_fd_sc_hd__buf_2
XFILLER_4_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_top_ipin_5.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_6.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_2.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR bottom_grid_pin_4_ sky130_fd_sc_hd__buf_4
XTAP_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_52_ chanx_left_in[17] VGND VGND VPWR VPWR chanx_right_out[17] sky130_fd_sc_hd__buf_2
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_7.mux_l1_in_1__A0 chanx_right_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xlogical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A
+ IO_ISOL_N VGND VGND VPWR VPWR _59_/A sky130_fd_sc_hd__or2b_4
XFILLER_14_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_0.mux_l1_in_0__A1 chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_35_ chanx_left_in[0] VGND VGND VPWR VPWR chanx_right_out[0] sky130_fd_sc_hd__buf_2
XFILLER_22_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xlogical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
+ prog_clk_0_FTB00/X mux_top_ipin_8.mux_l4_in_0_/S VGND VGND VPWR VPWR logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A
+ sky130_fd_sc_hd__dfxtp_1
X_18_ chanx_right_in[3] VGND VGND VPWR VPWR chanx_left_out[3] sky130_fd_sc_hd__buf_2
XANTENNA_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE_B_N
+ IO_ISOL_N VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_5.mux_l2_in_2__A0 chanx_left_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xlogical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE top_width_0_height_0__pin_6_
+ _58_/A VGND VGND VPWR VPWR _67_/A sky130_fd_sc_hd__ebufn_4
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_51_ chanx_left_in[16] VGND VGND VPWR VPWR chanx_right_out[16] sky130_fd_sc_hd__buf_2
XANTENNA_mux_top_ipin_7.mux_l1_in_1__A1 chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34_ chanx_right_in[19] VGND VGND VPWR VPWR chanx_left_out[19] sky130_fd_sc_hd__buf_2
XFILLER_20_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17_ VGND VGND VPWR VPWR _17_/HI _17_/LO sky130_fd_sc_hd__conb_1
XFILLER_3_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_0.mux_l2_in_3_ _09_/HI chanx_right_in[16] mux_top_ipin_0.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_0.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_5.mux_l2_in_2__A1 chanx_right_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_ipin_2.mux_l1_in_1__A0 chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_0.mux_l4_in_0_ mux_top_ipin_0.mux_l3_in_1_/X mux_top_ipin_0.mux_l3_in_0_/X
+ mux_top_ipin_0.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_0.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE_A
+ top_width_0_height_0__pin_16_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_50_ chanx_left_in[15] VGND VGND VPWR VPWR chanx_right_out[15] sky130_fd_sc_hd__buf_2
Xmux_top_ipin_5.mux_l2_in_3_ _14_/HI chanx_right_in[15] mux_top_ipin_5.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_5.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
X_33_ chanx_right_in[18] VGND VGND VPWR VPWR chanx_left_out[18] sky130_fd_sc_hd__buf_2
Xlogical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
+ prog_clk_0_FTB00/X logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A
+ VGND VGND VPWR VPWR logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A
+ sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_0.mux_l3_in_1_ mux_top_ipin_0.mux_l2_in_3_/X mux_top_ipin_0.mux_l2_in_2_/X
+ mux_top_ipin_0.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_0.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_0.mux_l2_in_2__A0 chanx_left_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16_ VGND VGND VPWR VPWR _16_/HI _16_/LO sky130_fd_sc_hd__conb_1
XFILLER_10_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE_B_N
+ IO_ISOL_N VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_5.mux_l4_in_0_ mux_top_ipin_5.mux_l3_in_1_/X mux_top_ipin_5.mux_l3_in_0_/X
+ mux_top_ipin_5.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_5.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_0.mux_l2_in_2_ chanx_left_in[16] chanx_right_in[10] mux_top_ipin_0.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_0.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xlogical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE top_width_0_height_0__pin_8_
+ _59_/A VGND VGND VPWR VPWR _68_/A sky130_fd_sc_hd__ebufn_4
XANTENNA_mux_top_ipin_2.mux_l1_in_1__A1 chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_5.mux_l3_in_1_ mux_top_ipin_5.mux_l2_in_3_/X mux_top_ipin_5.mux_l2_in_2_/X
+ mux_top_ipin_5.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_5.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xlogical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR _57_/A
+ VGND VGND VPWR VPWR logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y
+ sky130_fd_sc_hd__inv_1
XFILLER_14_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32_ chanx_right_in[17] VGND VGND VPWR VPWR chanx_left_out[17] sky130_fd_sc_hd__buf_2
Xmux_top_ipin_5.mux_l2_in_2_ chanx_left_in[15] chanx_right_in[9] mux_top_ipin_5.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_5.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XANTENNA_logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE_A
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_0.mux_l2_in_2__A1 chanx_right_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_0.mux_l3_in_0_ mux_top_ipin_0.mux_l2_in_1_/X mux_top_ipin_0.mux_l2_in_0_/X
+ mux_top_ipin_0.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_0.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15_ VGND VGND VPWR VPWR _15_/HI _15_/LO sky130_fd_sc_hd__conb_1
XFILLER_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_0.mux_l2_in_1_ chanx_left_in[10] mux_top_ipin_0.mux_l1_in_2_/X mux_top_ipin_0.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_0.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_0.mux_l1_in_2_ chanx_right_in[4] chanx_left_in[4] mux_top_ipin_0.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_0.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_5.mux_l3_in_0_ mux_top_ipin_5.mux_l2_in_1_/X mux_top_ipin_5.mux_l2_in_0_/X
+ mux_top_ipin_5.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_5.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_5.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_5.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR bottom_grid_pin_10_ sky130_fd_sc_hd__buf_4
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xlogical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A
+ IO_ISOL_N VGND VGND VPWR VPWR _57_/A sky130_fd_sc_hd__or2b_4
XFILLER_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_7.mux_l2_in_3__A1 chanx_right_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_5.mux_l2_in_1_ chanx_left_in[9] mux_top_ipin_5.mux_l1_in_2_/X mux_top_ipin_5.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_5.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
X_31_ chanx_right_in[16] VGND VGND VPWR VPWR chanx_left_out[16] sky130_fd_sc_hd__buf_2
XFILLER_22_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE_B_N
+ IO_ISOL_N VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_6.mux_l1_in_0__A0 chanx_right_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14_ VGND VGND VPWR VPWR _14_/HI _14_/LO sky130_fd_sc_hd__conb_1
Xmux_top_ipin_5.mux_l1_in_2_ chanx_right_in[5] chanx_left_in[5] mux_top_ipin_5.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_5.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22__A chanx_right_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_4.mux_l1_in_2__A0 chanx_right_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_0.mux_l2_in_0_ mux_top_ipin_0.mux_l1_in_1_/X mux_top_ipin_0.mux_l1_in_0_/X
+ mux_top_ipin_0.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_top_ipin_0.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xlogical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE top_width_0_height_0__pin_10_
+ _60_/A VGND VGND VPWR VPWR _69_/A sky130_fd_sc_hd__ebufn_4
XFILLER_14_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_4.mux_l2_in_1__A0 chanx_left_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_0.mux_l1_in_1_ chanx_right_in[2] chanx_left_in[2] mux_top_ipin_0.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_0.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA__30__A chanx_right_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25__A chanx_right_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30_ chanx_right_in[15] VGND VGND VPWR VPWR chanx_left_out[15] sky130_fd_sc_hd__buf_2
Xmux_top_ipin_5.mux_l2_in_0_ mux_top_ipin_5.mux_l1_in_1_/X mux_top_ipin_5.mux_l1_in_0_/X
+ mux_top_ipin_5.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_top_ipin_5.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_6.mux_l1_in_0__A1 chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13_ VGND VGND VPWR VPWR _13_/HI _13_/LO sky130_fd_sc_hd__conb_1
XFILLER_17_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_5.mux_l1_in_1_ chanx_right_in[3] chanx_left_in[3] mux_top_ipin_5.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_5.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_ipin_4.mux_l1_in_2__A1 chanx_left_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE_A
+ top_width_0_height_0__pin_14_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__33__A chanx_right_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__28__A chanx_right_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_0.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_top_ipin_0.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_0.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_2.mux_l2_in_3__A1 chanx_right_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_1.mux_l1_in_0__A0 chanx_right_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE_B_N
+ IO_ISOL_N VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xlogical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR _61_/A
+ VGND VGND VPWR VPWR logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y
+ sky130_fd_sc_hd__inv_1
XANTENNA__41__A chanx_left_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__36__A chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12_ VGND VGND VPWR VPWR _12_/HI _12_/LO sky130_fd_sc_hd__conb_1
XFILLER_6_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_5.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_top_ipin_5.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_5.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xlogical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE top_width_0_height_0__pin_12_
+ _61_/A VGND VGND VPWR VPWR _70_/A sky130_fd_sc_hd__ebufn_4
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__44__A chanx_left_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xlogical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
+ prog_clk_0_FTB00/X logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A
+ VGND VGND VPWR VPWR logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_8.mux_l1_in_1__A0 chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_1.mux_l1_in_0__A1 chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__39__A chanx_left_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_128 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__52__A chanx_left_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11_ VGND VGND VPWR VPWR _11_/HI _11_/LO sky130_fd_sc_hd__conb_1
XFILLER_6_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_6.mux_l2_in_2__A0 chanx_left_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__47__A chanx_left_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_top_ipin_2.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_top_ipin_2.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE_A
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_8.mux_l1_in_1__A1 chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_8.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_8.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR bottom_grid_pin_16_ sky130_fd_sc_hd__buf_4
XANTENNA_logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE_B_N
+ IO_ISOL_N VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xlogical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A
+ IO_ISOL_N VGND VGND VPWR VPWR _55_/A sky130_fd_sc_hd__or2b_4
X_10_ VGND VGND VPWR VPWR _10_/HI _10_/LO sky130_fd_sc_hd__conb_1
XANTENNA_mux_top_ipin_6.mux_l2_in_2__A1 chanx_right_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xlogical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE top_width_0_height_0__pin_14_
+ _62_/A VGND VGND VPWR VPWR _71_/A sky130_fd_sc_hd__ebufn_4
Xmem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_top_ipin_5.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_top_ipin_5.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0__D ccff_head VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_3.mux_l1_in_1__A0 chanx_right_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_top_ipin_2.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_2.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_1.mux_l2_in_3_ _10_/HI chanx_right_in[17] mux_top_ipin_1.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_1.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xlogical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE gfpga_pad_EMBEDDED_IO_HD_SOC_IN[7]
+ logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y VGND
+ VGND VPWR VPWR top_width_0_height_0__pin_15_lower sky130_fd_sc_hd__ebufn_4
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_top_ipin_1.mux_l2_in_2__A0 chanx_left_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_top_ipin_8.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_top_ipin_8.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_22_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_86_ chanx_right_in[2] VGND VGND VPWR VPWR chanx_left_out[2] sky130_fd_sc_hd__buf_2
Xmux_top_ipin_1.mux_l4_in_0_ mux_top_ipin_1.mux_l3_in_1_/X mux_top_ipin_1.mux_l3_in_0_/X
+ mux_top_ipin_1.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_1.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE_A
+ top_width_0_height_0__pin_12_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_top_ipin_5.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_5.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
X_69_ _69_/A VGND VGND VPWR VPWR gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[5] sky130_fd_sc_hd__buf_2
XFILLER_0_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_6.mux_l2_in_3_ _15_/HI chanx_right_in[16] mux_top_ipin_6.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_6.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_1.mux_l3_in_1_ mux_top_ipin_1.mux_l2_in_3_/X mux_top_ipin_1.mux_l2_in_2_/X
+ mux_top_ipin_1.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_1.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_3.mux_l1_in_1__A1 chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_top_ipin_2.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_2.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_20_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xlogical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE gfpga_pad_EMBEDDED_IO_HD_SOC_IN[4]
+ logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y VGND
+ VGND VPWR VPWR top_width_0_height_0__pin_9_lower sky130_fd_sc_hd__ebufn_4
Xmux_top_ipin_1.mux_l2_in_2_ chanx_left_in[17] chanx_right_in[11] mux_top_ipin_1.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_1.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XANTENNA_logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE_B_N
+ IO_ISOL_N VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_6.mux_l4_in_0_ mux_top_ipin_6.mux_l3_in_1_/X mux_top_ipin_6.mux_l3_in_0_/X
+ mux_top_ipin_6.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_6.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XTAP_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__82__A SC_IN_TOP VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_1.mux_l2_in_2__A1 chanx_right_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_top_ipin_8.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_8.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_9_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_85_ chanx_right_in[1] VGND VGND VPWR VPWR chanx_left_out[1] sky130_fd_sc_hd__buf_2
Xmux_top_ipin_6.mux_l3_in_1_ mux_top_ipin_6.mux_l2_in_3_/X mux_top_ipin_6.mux_l2_in_2_/X
+ mux_top_ipin_6.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_6.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xlogical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE top_width_0_height_0__pin_16_
+ _63_/A VGND VGND VPWR VPWR _72_/A sky130_fd_sc_hd__ebufn_4
XFILLER_6_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__77__A top_width_0_height_0__pin_1_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_1.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR bottom_grid_pin_2_ sky130_fd_sc_hd__buf_4
XFILLER_17_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_top_ipin_5.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_5.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
X_68_ _68_/A VGND VGND VPWR VPWR gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[4] sky130_fd_sc_hd__buf_2
Xmux_top_ipin_6.mux_l2_in_2_ chanx_left_in[16] chanx_right_in[10] mux_top_ipin_6.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_6.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_174 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_top_ipin_1.mux_l3_in_0_ mux_top_ipin_1.mux_l2_in_1_/X mux_top_ipin_1.mux_l2_in_0_/X
+ mux_top_ipin_1.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_1.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_top_ipin_1.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_2.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
Xlogical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE gfpga_pad_EMBEDDED_IO_HD_SOC_IN[1]
+ logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y VGND
+ VGND VPWR VPWR top_width_0_height_0__pin_3_lower sky130_fd_sc_hd__ebufn_4
XFILLER_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_1.mux_l2_in_1_ chanx_left_in[11] mux_top_ipin_1.mux_l1_in_2_/X mux_top_ipin_1.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_1.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA__85__A chanx_right_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_ipin_8.mux_l2_in_3__A1 chanx_right_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_7.mux_l1_in_0__A0 chanx_right_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_1.mux_l1_in_2_ chanx_right_in[5] chanx_left_in[5] mux_top_ipin_1.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_1.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xmem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_top_ipin_8.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_8.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
Xlogical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR _56_/A
+ VGND VGND VPWR VPWR logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y
+ sky130_fd_sc_hd__inv_1
X_84_ chanx_right_in[0] VGND VGND VPWR VPWR chanx_left_out[0] sky130_fd_sc_hd__buf_2
Xmux_top_ipin_6.mux_l3_in_0_ mux_top_ipin_6.mux_l2_in_1_/X mux_top_ipin_6.mux_l2_in_0_/X
+ mux_top_ipin_6.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_6.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_ipin_5.mux_l1_in_2__A0 chanx_right_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_top_ipin_4.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_5.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
Xlogical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
+ prog_clk_0_FTB00/X logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A
+ VGND VGND VPWR VPWR logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A
+ sky130_fd_sc_hd__dfxtp_1
X_67_ _67_/A VGND VGND VPWR VPWR gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[3] sky130_fd_sc_hd__buf_2
XFILLER_2_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_6.mux_l2_in_1_ chanx_left_in[10] mux_top_ipin_6.mux_l1_in_2_/X mux_top_ipin_6.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_6.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_5.mux_l2_in_1__A0 chanx_left_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE_B_N
+ IO_ISOL_N VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_6.mux_l1_in_2_ chanx_right_in[6] chanx_left_in[6] mux_top_ipin_6.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_6.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_1.mux_l2_in_0_ mux_top_ipin_1.mux_l1_in_1_/X mux_top_ipin_1.mux_l1_in_0_/X
+ mux_top_ipin_1.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_top_ipin_1.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xlogical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE/A
+ IO_ISOL_N VGND VGND VPWR VPWR _62_/A sky130_fd_sc_hd__or2b_4
.ends

