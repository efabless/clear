magic
tech sky130A
magscale 1 2
timestamp 1656943069
<< obsli1 >>
rect 1104 2159 18860 14705
<< obsm1 >>
rect 934 1504 19398 15360
<< metal2 >>
rect 1122 16400 1178 17200
rect 3330 16400 3386 17200
rect 5538 16400 5594 17200
rect 7746 16400 7802 17200
rect 9954 16400 10010 17200
rect 12162 16400 12218 17200
rect 14370 16400 14426 17200
rect 16578 16400 16634 17200
rect 18786 16400 18842 17200
rect 1214 0 1270 800
rect 2042 0 2098 800
rect 2870 0 2926 800
rect 3698 0 3754 800
rect 4526 0 4582 800
rect 5354 0 5410 800
rect 6182 0 6238 800
rect 7010 0 7066 800
rect 7838 0 7894 800
rect 8666 0 8722 800
rect 9494 0 9550 800
rect 10322 0 10378 800
rect 11150 0 11206 800
rect 11978 0 12034 800
rect 12806 0 12862 800
rect 13634 0 13690 800
rect 14462 0 14518 800
rect 15290 0 15346 800
rect 16118 0 16174 800
rect 16946 0 17002 800
rect 17774 0 17830 800
rect 18602 0 18658 800
<< obsm2 >>
rect 938 16344 1066 16697
rect 1234 16344 3274 16697
rect 3442 16344 5482 16697
rect 5650 16344 7690 16697
rect 7858 16344 9898 16697
rect 10066 16344 12106 16697
rect 12274 16344 14314 16697
rect 14482 16344 16522 16697
rect 16690 16344 18730 16697
rect 18898 16344 19392 16697
rect 938 856 19392 16344
rect 938 303 1158 856
rect 1326 303 1986 856
rect 2154 303 2814 856
rect 2982 303 3642 856
rect 3810 303 4470 856
rect 4638 303 5298 856
rect 5466 303 6126 856
rect 6294 303 6954 856
rect 7122 303 7782 856
rect 7950 303 8610 856
rect 8778 303 9438 856
rect 9606 303 10266 856
rect 10434 303 11094 856
rect 11262 303 11922 856
rect 12090 303 12750 856
rect 12918 303 13578 856
rect 13746 303 14406 856
rect 14574 303 15234 856
rect 15402 303 16062 856
rect 16230 303 16890 856
rect 17058 303 17718 856
rect 17886 303 18546 856
rect 18714 303 19392 856
<< metal3 >>
rect 0 16600 800 16720
rect 19200 16464 20000 16584
rect 0 16192 800 16312
rect 19200 16056 20000 16176
rect 0 15784 800 15904
rect 19200 15648 20000 15768
rect 0 15376 800 15496
rect 19200 15240 20000 15360
rect 0 14968 800 15088
rect 19200 14832 20000 14952
rect 0 14560 800 14680
rect 19200 14424 20000 14544
rect 0 14152 800 14272
rect 19200 14016 20000 14136
rect 0 13744 800 13864
rect 19200 13608 20000 13728
rect 0 13336 800 13456
rect 19200 13200 20000 13320
rect 0 12928 800 13048
rect 19200 12792 20000 12912
rect 0 12520 800 12640
rect 19200 12384 20000 12504
rect 0 12112 800 12232
rect 19200 11976 20000 12096
rect 0 11704 800 11824
rect 19200 11568 20000 11688
rect 0 11296 800 11416
rect 19200 11160 20000 11280
rect 0 10888 800 11008
rect 19200 10752 20000 10872
rect 0 10480 800 10600
rect 19200 10344 20000 10464
rect 0 10072 800 10192
rect 19200 9936 20000 10056
rect 0 9664 800 9784
rect 19200 9528 20000 9648
rect 0 9256 800 9376
rect 19200 9120 20000 9240
rect 0 8848 800 8968
rect 19200 8712 20000 8832
rect 0 8440 800 8560
rect 19200 8304 20000 8424
rect 0 8032 800 8152
rect 19200 7896 20000 8016
rect 0 7624 800 7744
rect 19200 7488 20000 7608
rect 0 7216 800 7336
rect 19200 7080 20000 7200
rect 0 6808 800 6928
rect 19200 6672 20000 6792
rect 0 6400 800 6520
rect 19200 6264 20000 6384
rect 0 5992 800 6112
rect 19200 5856 20000 5976
rect 0 5584 800 5704
rect 19200 5448 20000 5568
rect 0 5176 800 5296
rect 19200 5040 20000 5160
rect 0 4768 800 4888
rect 19200 4632 20000 4752
rect 0 4360 800 4480
rect 19200 4224 20000 4344
rect 0 3952 800 4072
rect 19200 3816 20000 3936
rect 0 3544 800 3664
rect 19200 3408 20000 3528
rect 0 3136 800 3256
rect 19200 3000 20000 3120
rect 0 2728 800 2848
rect 19200 2592 20000 2712
rect 0 2320 800 2440
rect 19200 2184 20000 2304
rect 0 1912 800 2032
rect 19200 1776 20000 1896
rect 0 1504 800 1624
rect 19200 1368 20000 1488
rect 0 1096 800 1216
rect 19200 960 20000 1080
rect 0 688 800 808
rect 19200 552 20000 672
rect 0 280 800 400
<< obsm3 >>
rect 880 16664 19200 16693
rect 880 16520 19120 16664
rect 800 16392 19120 16520
rect 880 16384 19120 16392
rect 880 16256 19200 16384
rect 880 16112 19120 16256
rect 800 15984 19120 16112
rect 880 15976 19120 15984
rect 880 15848 19200 15976
rect 880 15704 19120 15848
rect 800 15576 19120 15704
rect 880 15568 19120 15576
rect 880 15440 19200 15568
rect 880 15296 19120 15440
rect 800 15168 19120 15296
rect 880 15160 19120 15168
rect 880 15032 19200 15160
rect 880 14888 19120 15032
rect 800 14760 19120 14888
rect 880 14752 19120 14760
rect 880 14624 19200 14752
rect 880 14480 19120 14624
rect 800 14352 19120 14480
rect 880 14344 19120 14352
rect 880 14216 19200 14344
rect 880 14072 19120 14216
rect 800 13944 19120 14072
rect 880 13936 19120 13944
rect 880 13808 19200 13936
rect 880 13664 19120 13808
rect 800 13536 19120 13664
rect 880 13528 19120 13536
rect 880 13400 19200 13528
rect 880 13256 19120 13400
rect 800 13128 19120 13256
rect 880 13120 19120 13128
rect 880 12992 19200 13120
rect 880 12848 19120 12992
rect 800 12720 19120 12848
rect 880 12712 19120 12720
rect 880 12584 19200 12712
rect 880 12440 19120 12584
rect 800 12312 19120 12440
rect 880 12304 19120 12312
rect 880 12176 19200 12304
rect 880 12032 19120 12176
rect 800 11904 19120 12032
rect 880 11896 19120 11904
rect 880 11768 19200 11896
rect 880 11624 19120 11768
rect 800 11496 19120 11624
rect 880 11488 19120 11496
rect 880 11360 19200 11488
rect 880 11216 19120 11360
rect 800 11088 19120 11216
rect 880 11080 19120 11088
rect 880 10952 19200 11080
rect 880 10808 19120 10952
rect 800 10680 19120 10808
rect 880 10672 19120 10680
rect 880 10544 19200 10672
rect 880 10400 19120 10544
rect 800 10272 19120 10400
rect 880 10264 19120 10272
rect 880 10136 19200 10264
rect 880 9992 19120 10136
rect 800 9864 19120 9992
rect 880 9856 19120 9864
rect 880 9728 19200 9856
rect 880 9584 19120 9728
rect 800 9456 19120 9584
rect 880 9448 19120 9456
rect 880 9320 19200 9448
rect 880 9176 19120 9320
rect 800 9048 19120 9176
rect 880 9040 19120 9048
rect 880 8912 19200 9040
rect 880 8768 19120 8912
rect 800 8640 19120 8768
rect 880 8632 19120 8640
rect 880 8504 19200 8632
rect 880 8360 19120 8504
rect 800 8232 19120 8360
rect 880 8224 19120 8232
rect 880 8096 19200 8224
rect 880 7952 19120 8096
rect 800 7824 19120 7952
rect 880 7816 19120 7824
rect 880 7688 19200 7816
rect 880 7544 19120 7688
rect 800 7416 19120 7544
rect 880 7408 19120 7416
rect 880 7280 19200 7408
rect 880 7136 19120 7280
rect 800 7008 19120 7136
rect 880 7000 19120 7008
rect 880 6872 19200 7000
rect 880 6728 19120 6872
rect 800 6600 19120 6728
rect 880 6592 19120 6600
rect 880 6464 19200 6592
rect 880 6320 19120 6464
rect 800 6192 19120 6320
rect 880 6184 19120 6192
rect 880 6056 19200 6184
rect 880 5912 19120 6056
rect 800 5784 19120 5912
rect 880 5776 19120 5784
rect 880 5648 19200 5776
rect 880 5504 19120 5648
rect 800 5376 19120 5504
rect 880 5368 19120 5376
rect 880 5240 19200 5368
rect 880 5096 19120 5240
rect 800 4968 19120 5096
rect 880 4960 19120 4968
rect 880 4832 19200 4960
rect 880 4688 19120 4832
rect 800 4560 19120 4688
rect 880 4552 19120 4560
rect 880 4424 19200 4552
rect 880 4280 19120 4424
rect 800 4152 19120 4280
rect 880 4144 19120 4152
rect 880 4016 19200 4144
rect 880 3872 19120 4016
rect 800 3744 19120 3872
rect 880 3736 19120 3744
rect 880 3608 19200 3736
rect 880 3464 19120 3608
rect 800 3336 19120 3464
rect 880 3328 19120 3336
rect 880 3200 19200 3328
rect 880 3056 19120 3200
rect 800 2928 19120 3056
rect 880 2920 19120 2928
rect 880 2792 19200 2920
rect 880 2648 19120 2792
rect 800 2520 19120 2648
rect 880 2512 19120 2520
rect 880 2384 19200 2512
rect 880 2240 19120 2384
rect 800 2112 19120 2240
rect 880 2104 19120 2112
rect 880 1976 19200 2104
rect 880 1832 19120 1976
rect 800 1704 19120 1832
rect 880 1696 19120 1704
rect 880 1568 19200 1696
rect 880 1424 19120 1568
rect 800 1296 19120 1424
rect 880 1288 19120 1296
rect 880 1160 19200 1288
rect 880 1016 19120 1160
rect 800 888 19120 1016
rect 880 880 19120 888
rect 880 752 19200 880
rect 880 608 19120 752
rect 800 480 19120 608
rect 880 472 19120 480
rect 880 307 19200 472
<< metal4 >>
rect 3168 2128 3488 14736
rect 5392 2128 5712 14736
rect 7616 2128 7936 14736
rect 9840 2128 10160 14736
rect 12064 2128 12384 14736
rect 14288 2128 14608 14736
rect 16512 2128 16832 14736
<< obsm4 >>
rect 2451 14816 17789 16149
rect 2451 2347 3088 14816
rect 3568 2347 5312 14816
rect 5792 2347 7536 14816
rect 8016 2347 9760 14816
rect 10240 2347 11984 14816
rect 12464 2347 14208 14816
rect 14688 2347 16432 14816
rect 16912 2347 17789 14816
<< labels >>
rlabel metal2 s 1122 16400 1178 17200 6 IO_ISOL_N
port 1 nsew signal input
rlabel metal2 s 16946 0 17002 800 6 SC_IN_BOT
port 2 nsew signal input
rlabel metal2 s 3330 16400 3386 17200 6 SC_IN_TOP
port 3 nsew signal input
rlabel metal2 s 17774 0 17830 800 6 SC_OUT_BOT
port 4 nsew signal output
rlabel metal2 s 5538 16400 5594 17200 6 SC_OUT_TOP
port 5 nsew signal output
rlabel metal4 s 5392 2128 5712 14736 6 VGND
port 6 nsew ground bidirectional
rlabel metal4 s 9840 2128 10160 14736 6 VGND
port 6 nsew ground bidirectional
rlabel metal4 s 14288 2128 14608 14736 6 VGND
port 6 nsew ground bidirectional
rlabel metal4 s 3168 2128 3488 14736 6 VPWR
port 7 nsew power bidirectional
rlabel metal4 s 7616 2128 7936 14736 6 VPWR
port 7 nsew power bidirectional
rlabel metal4 s 12064 2128 12384 14736 6 VPWR
port 7 nsew power bidirectional
rlabel metal4 s 16512 2128 16832 14736 6 VPWR
port 7 nsew power bidirectional
rlabel metal2 s 2042 0 2098 800 6 bottom_grid_pin_0_
port 8 nsew signal output
rlabel metal2 s 10322 0 10378 800 6 bottom_grid_pin_10_
port 9 nsew signal output
rlabel metal2 s 11150 0 11206 800 6 bottom_grid_pin_11_
port 10 nsew signal output
rlabel metal2 s 11978 0 12034 800 6 bottom_grid_pin_12_
port 11 nsew signal output
rlabel metal2 s 12806 0 12862 800 6 bottom_grid_pin_13_
port 12 nsew signal output
rlabel metal2 s 13634 0 13690 800 6 bottom_grid_pin_14_
port 13 nsew signal output
rlabel metal2 s 14462 0 14518 800 6 bottom_grid_pin_15_
port 14 nsew signal output
rlabel metal2 s 2870 0 2926 800 6 bottom_grid_pin_1_
port 15 nsew signal output
rlabel metal2 s 3698 0 3754 800 6 bottom_grid_pin_2_
port 16 nsew signal output
rlabel metal2 s 4526 0 4582 800 6 bottom_grid_pin_3_
port 17 nsew signal output
rlabel metal2 s 5354 0 5410 800 6 bottom_grid_pin_4_
port 18 nsew signal output
rlabel metal2 s 6182 0 6238 800 6 bottom_grid_pin_5_
port 19 nsew signal output
rlabel metal2 s 7010 0 7066 800 6 bottom_grid_pin_6_
port 20 nsew signal output
rlabel metal2 s 7838 0 7894 800 6 bottom_grid_pin_7_
port 21 nsew signal output
rlabel metal2 s 8666 0 8722 800 6 bottom_grid_pin_8_
port 22 nsew signal output
rlabel metal2 s 9494 0 9550 800 6 bottom_grid_pin_9_
port 23 nsew signal output
rlabel metal2 s 15290 0 15346 800 6 bottom_width_0_height_0__pin_0_
port 24 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 bottom_width_0_height_0__pin_1_lower
port 25 nsew signal output
rlabel metal2 s 1214 0 1270 800 6 bottom_width_0_height_0__pin_1_upper
port 26 nsew signal output
rlabel metal2 s 7746 16400 7802 17200 6 ccff_head
port 27 nsew signal input
rlabel metal2 s 9954 16400 10010 17200 6 ccff_tail
port 28 nsew signal output
rlabel metal3 s 0 8848 800 8968 6 chanx_left_in[0]
port 29 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 chanx_left_in[10]
port 30 nsew signal input
rlabel metal3 s 0 13336 800 13456 6 chanx_left_in[11]
port 31 nsew signal input
rlabel metal3 s 0 13744 800 13864 6 chanx_left_in[12]
port 32 nsew signal input
rlabel metal3 s 0 14152 800 14272 6 chanx_left_in[13]
port 33 nsew signal input
rlabel metal3 s 0 14560 800 14680 6 chanx_left_in[14]
port 34 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 chanx_left_in[15]
port 35 nsew signal input
rlabel metal3 s 0 15376 800 15496 6 chanx_left_in[16]
port 36 nsew signal input
rlabel metal3 s 0 15784 800 15904 6 chanx_left_in[17]
port 37 nsew signal input
rlabel metal3 s 0 16192 800 16312 6 chanx_left_in[18]
port 38 nsew signal input
rlabel metal3 s 0 16600 800 16720 6 chanx_left_in[19]
port 39 nsew signal input
rlabel metal3 s 0 9256 800 9376 6 chanx_left_in[1]
port 40 nsew signal input
rlabel metal3 s 0 9664 800 9784 6 chanx_left_in[2]
port 41 nsew signal input
rlabel metal3 s 0 10072 800 10192 6 chanx_left_in[3]
port 42 nsew signal input
rlabel metal3 s 0 10480 800 10600 6 chanx_left_in[4]
port 43 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 chanx_left_in[5]
port 44 nsew signal input
rlabel metal3 s 0 11296 800 11416 6 chanx_left_in[6]
port 45 nsew signal input
rlabel metal3 s 0 11704 800 11824 6 chanx_left_in[7]
port 46 nsew signal input
rlabel metal3 s 0 12112 800 12232 6 chanx_left_in[8]
port 47 nsew signal input
rlabel metal3 s 0 12520 800 12640 6 chanx_left_in[9]
port 48 nsew signal input
rlabel metal3 s 0 688 800 808 6 chanx_left_out[0]
port 49 nsew signal output
rlabel metal3 s 0 4768 800 4888 6 chanx_left_out[10]
port 50 nsew signal output
rlabel metal3 s 0 5176 800 5296 6 chanx_left_out[11]
port 51 nsew signal output
rlabel metal3 s 0 5584 800 5704 6 chanx_left_out[12]
port 52 nsew signal output
rlabel metal3 s 0 5992 800 6112 6 chanx_left_out[13]
port 53 nsew signal output
rlabel metal3 s 0 6400 800 6520 6 chanx_left_out[14]
port 54 nsew signal output
rlabel metal3 s 0 6808 800 6928 6 chanx_left_out[15]
port 55 nsew signal output
rlabel metal3 s 0 7216 800 7336 6 chanx_left_out[16]
port 56 nsew signal output
rlabel metal3 s 0 7624 800 7744 6 chanx_left_out[17]
port 57 nsew signal output
rlabel metal3 s 0 8032 800 8152 6 chanx_left_out[18]
port 58 nsew signal output
rlabel metal3 s 0 8440 800 8560 6 chanx_left_out[19]
port 59 nsew signal output
rlabel metal3 s 0 1096 800 1216 6 chanx_left_out[1]
port 60 nsew signal output
rlabel metal3 s 0 1504 800 1624 6 chanx_left_out[2]
port 61 nsew signal output
rlabel metal3 s 0 1912 800 2032 6 chanx_left_out[3]
port 62 nsew signal output
rlabel metal3 s 0 2320 800 2440 6 chanx_left_out[4]
port 63 nsew signal output
rlabel metal3 s 0 2728 800 2848 6 chanx_left_out[5]
port 64 nsew signal output
rlabel metal3 s 0 3136 800 3256 6 chanx_left_out[6]
port 65 nsew signal output
rlabel metal3 s 0 3544 800 3664 6 chanx_left_out[7]
port 66 nsew signal output
rlabel metal3 s 0 3952 800 4072 6 chanx_left_out[8]
port 67 nsew signal output
rlabel metal3 s 0 4360 800 4480 6 chanx_left_out[9]
port 68 nsew signal output
rlabel metal3 s 19200 8712 20000 8832 6 chanx_right_in[0]
port 69 nsew signal input
rlabel metal3 s 19200 12792 20000 12912 6 chanx_right_in[10]
port 70 nsew signal input
rlabel metal3 s 19200 13200 20000 13320 6 chanx_right_in[11]
port 71 nsew signal input
rlabel metal3 s 19200 13608 20000 13728 6 chanx_right_in[12]
port 72 nsew signal input
rlabel metal3 s 19200 14016 20000 14136 6 chanx_right_in[13]
port 73 nsew signal input
rlabel metal3 s 19200 14424 20000 14544 6 chanx_right_in[14]
port 74 nsew signal input
rlabel metal3 s 19200 14832 20000 14952 6 chanx_right_in[15]
port 75 nsew signal input
rlabel metal3 s 19200 15240 20000 15360 6 chanx_right_in[16]
port 76 nsew signal input
rlabel metal3 s 19200 15648 20000 15768 6 chanx_right_in[17]
port 77 nsew signal input
rlabel metal3 s 19200 16056 20000 16176 6 chanx_right_in[18]
port 78 nsew signal input
rlabel metal3 s 19200 16464 20000 16584 6 chanx_right_in[19]
port 79 nsew signal input
rlabel metal3 s 19200 9120 20000 9240 6 chanx_right_in[1]
port 80 nsew signal input
rlabel metal3 s 19200 9528 20000 9648 6 chanx_right_in[2]
port 81 nsew signal input
rlabel metal3 s 19200 9936 20000 10056 6 chanx_right_in[3]
port 82 nsew signal input
rlabel metal3 s 19200 10344 20000 10464 6 chanx_right_in[4]
port 83 nsew signal input
rlabel metal3 s 19200 10752 20000 10872 6 chanx_right_in[5]
port 84 nsew signal input
rlabel metal3 s 19200 11160 20000 11280 6 chanx_right_in[6]
port 85 nsew signal input
rlabel metal3 s 19200 11568 20000 11688 6 chanx_right_in[7]
port 86 nsew signal input
rlabel metal3 s 19200 11976 20000 12096 6 chanx_right_in[8]
port 87 nsew signal input
rlabel metal3 s 19200 12384 20000 12504 6 chanx_right_in[9]
port 88 nsew signal input
rlabel metal3 s 19200 552 20000 672 6 chanx_right_out[0]
port 89 nsew signal output
rlabel metal3 s 19200 4632 20000 4752 6 chanx_right_out[10]
port 90 nsew signal output
rlabel metal3 s 19200 5040 20000 5160 6 chanx_right_out[11]
port 91 nsew signal output
rlabel metal3 s 19200 5448 20000 5568 6 chanx_right_out[12]
port 92 nsew signal output
rlabel metal3 s 19200 5856 20000 5976 6 chanx_right_out[13]
port 93 nsew signal output
rlabel metal3 s 19200 6264 20000 6384 6 chanx_right_out[14]
port 94 nsew signal output
rlabel metal3 s 19200 6672 20000 6792 6 chanx_right_out[15]
port 95 nsew signal output
rlabel metal3 s 19200 7080 20000 7200 6 chanx_right_out[16]
port 96 nsew signal output
rlabel metal3 s 19200 7488 20000 7608 6 chanx_right_out[17]
port 97 nsew signal output
rlabel metal3 s 19200 7896 20000 8016 6 chanx_right_out[18]
port 98 nsew signal output
rlabel metal3 s 19200 8304 20000 8424 6 chanx_right_out[19]
port 99 nsew signal output
rlabel metal3 s 19200 960 20000 1080 6 chanx_right_out[1]
port 100 nsew signal output
rlabel metal3 s 19200 1368 20000 1488 6 chanx_right_out[2]
port 101 nsew signal output
rlabel metal3 s 19200 1776 20000 1896 6 chanx_right_out[3]
port 102 nsew signal output
rlabel metal3 s 19200 2184 20000 2304 6 chanx_right_out[4]
port 103 nsew signal output
rlabel metal3 s 19200 2592 20000 2712 6 chanx_right_out[5]
port 104 nsew signal output
rlabel metal3 s 19200 3000 20000 3120 6 chanx_right_out[6]
port 105 nsew signal output
rlabel metal3 s 19200 3408 20000 3528 6 chanx_right_out[7]
port 106 nsew signal output
rlabel metal3 s 19200 3816 20000 3936 6 chanx_right_out[8]
port 107 nsew signal output
rlabel metal3 s 19200 4224 20000 4344 6 chanx_right_out[9]
port 108 nsew signal output
rlabel metal2 s 14370 16400 14426 17200 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR
port 109 nsew signal output
rlabel metal2 s 16578 16400 16634 17200 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN
port 110 nsew signal input
rlabel metal2 s 18786 16400 18842 17200 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT
port 111 nsew signal output
rlabel metal2 s 18602 0 18658 800 6 prog_clk_0_S_in
port 112 nsew signal input
rlabel metal3 s 0 280 800 400 6 prog_clk_0_W_out
port 113 nsew signal output
rlabel metal2 s 12162 16400 12218 17200 6 top_grid_pin_0_
port 114 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 20000 17200
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1196012
string GDS_FILE /home/marwan/clear_signoff_final/openlane/cbx_1__2_/runs/cbx_1__2_/results/signoff/cbx_1__2_.magic.gds
string GDS_START 84912
<< end >>

