magic
tech sky130A
magscale 1 2
timestamp 1656241648
<< viali >>
rect 8309 22185 8343 22219
rect 14289 22185 14323 22219
rect 10609 22117 10643 22151
rect 13645 22117 13679 22151
rect 5457 22049 5491 22083
rect 6009 22049 6043 22083
rect 6193 22049 6227 22083
rect 6745 22049 6779 22083
rect 8217 22049 8251 22083
rect 9689 22049 9723 22083
rect 10517 22049 10551 22083
rect 12449 22049 12483 22083
rect 12725 22049 12759 22083
rect 16957 22049 16991 22083
rect 17693 22049 17727 22083
rect 20637 22049 20671 22083
rect 1961 21981 1995 22015
rect 2605 21981 2639 22015
rect 3249 21981 3283 22015
rect 4077 21981 4111 22015
rect 4261 21981 4295 22015
rect 4813 21981 4847 22015
rect 5181 21981 5215 22015
rect 5733 21981 5767 22015
rect 6561 21981 6595 22015
rect 7021 21981 7055 22015
rect 7481 21981 7515 22015
rect 7757 21981 7791 22015
rect 8493 21981 8527 22015
rect 8769 21981 8803 22015
rect 10241 21981 10275 22015
rect 10793 21981 10827 22015
rect 11069 21981 11103 22015
rect 11345 21981 11379 22015
rect 11529 21981 11563 22015
rect 12081 21981 12115 22015
rect 12173 21981 12207 22015
rect 13461 21981 13495 22015
rect 13737 21981 13771 22015
rect 14473 21981 14507 22015
rect 15485 21981 15519 22015
rect 15761 21981 15795 22015
rect 16037 21981 16071 22015
rect 16313 21981 16347 22015
rect 18705 21981 18739 22015
rect 18981 21981 19015 22015
rect 19349 21981 19383 22015
rect 19717 21981 19751 22015
rect 20177 21981 20211 22015
rect 20913 21981 20947 22015
rect 21373 21981 21407 22015
rect 21833 21981 21867 22015
rect 22293 21981 22327 22015
rect 22845 21981 22879 22015
rect 7205 21913 7239 21947
rect 9045 21913 9079 21947
rect 14105 21913 14139 21947
rect 14657 21913 14691 21947
rect 14933 21913 14967 21947
rect 15117 21913 15151 21947
rect 17049 21913 17083 21947
rect 17877 21913 17911 21947
rect 22753 21913 22787 21947
rect 1777 21845 1811 21879
rect 2421 21845 2455 21879
rect 3065 21845 3099 21879
rect 3893 21845 3927 21879
rect 4445 21845 4479 21879
rect 4629 21845 4663 21879
rect 4997 21845 5031 21879
rect 5549 21845 5583 21879
rect 6377 21845 6411 21879
rect 6837 21845 6871 21879
rect 7297 21845 7331 21879
rect 7573 21845 7607 21879
rect 7849 21845 7883 21879
rect 8585 21845 8619 21879
rect 9137 21845 9171 21879
rect 9505 21845 9539 21879
rect 9597 21845 9631 21879
rect 10057 21845 10091 21879
rect 10885 21845 10919 21879
rect 11161 21845 11195 21879
rect 11713 21845 11747 21879
rect 11897 21845 11931 21879
rect 12357 21845 12391 21879
rect 12909 21845 12943 21879
rect 13001 21845 13035 21879
rect 13369 21845 13403 21879
rect 13921 21845 13955 21879
rect 14749 21845 14783 21879
rect 15301 21845 15335 21879
rect 15577 21845 15611 21879
rect 15853 21845 15887 21879
rect 16129 21845 16163 21879
rect 16405 21845 16439 21879
rect 17141 21845 17175 21879
rect 17509 21845 17543 21879
rect 17969 21845 18003 21879
rect 18337 21845 18371 21879
rect 18521 21845 18555 21879
rect 18797 21845 18831 21879
rect 19533 21845 19567 21879
rect 19901 21845 19935 21879
rect 20361 21845 20395 21879
rect 20821 21845 20855 21879
rect 21281 21845 21315 21879
rect 21557 21845 21591 21879
rect 22017 21845 22051 21879
rect 22477 21845 22511 21879
rect 23029 21845 23063 21879
rect 1501 21641 1535 21675
rect 2421 21641 2455 21675
rect 2973 21641 3007 21675
rect 3249 21641 3283 21675
rect 3709 21641 3743 21675
rect 4997 21641 5031 21675
rect 7757 21641 7791 21675
rect 8309 21641 8343 21675
rect 10333 21641 10367 21675
rect 10977 21641 11011 21675
rect 11713 21641 11747 21675
rect 12541 21641 12575 21675
rect 13093 21641 13127 21675
rect 13461 21641 13495 21675
rect 15478 21641 15512 21675
rect 17509 21641 17543 21675
rect 18889 21641 18923 21675
rect 19165 21641 19199 21675
rect 19533 21641 19567 21675
rect 20545 21641 20579 21675
rect 21465 21641 21499 21675
rect 22293 21641 22327 21675
rect 4445 21573 4479 21607
rect 5917 21573 5951 21607
rect 8769 21573 8803 21607
rect 10609 21573 10643 21607
rect 11345 21573 11379 21607
rect 13001 21573 13035 21607
rect 13921 21573 13955 21607
rect 16037 21573 16071 21607
rect 16221 21573 16255 21607
rect 16405 21573 16439 21607
rect 19993 21573 20027 21607
rect 1685 21505 1719 21539
rect 2053 21505 2087 21539
rect 2329 21505 2363 21539
rect 2605 21505 2639 21539
rect 2881 21505 2915 21539
rect 3157 21505 3191 21539
rect 3433 21505 3467 21539
rect 3525 21505 3559 21539
rect 3985 21505 4019 21539
rect 4905 21505 4939 21539
rect 5181 21505 5215 21539
rect 5547 21505 5581 21539
rect 6653 21505 6687 21539
rect 7021 21505 7055 21539
rect 9597 21505 9631 21539
rect 10057 21505 10091 21539
rect 11161 21505 11195 21539
rect 11529 21505 11563 21539
rect 12081 21505 12115 21539
rect 12173 21505 12207 21539
rect 15209 21505 15243 21539
rect 17325 21505 17359 21539
rect 17693 21505 17727 21539
rect 19073 21505 19107 21539
rect 19349 21505 19383 21539
rect 19901 21505 19935 21539
rect 20361 21505 20395 21539
rect 21097 21505 21131 21539
rect 22201 21505 22235 21539
rect 22845 21505 22879 21539
rect 3801 21437 3835 21471
rect 4261 21437 4295 21471
rect 7849 21437 7883 21471
rect 8033 21437 8067 21471
rect 8861 21437 8895 21471
rect 9045 21437 9079 21471
rect 9689 21437 9723 21471
rect 9873 21437 9907 21471
rect 11897 21437 11931 21471
rect 12817 21437 12851 21471
rect 15439 21437 15473 21471
rect 15945 21437 15979 21471
rect 16773 21437 16807 21471
rect 17969 21437 18003 21471
rect 18245 21437 18279 21471
rect 20085 21437 20119 21471
rect 20821 21437 20855 21471
rect 21005 21437 21039 21471
rect 22385 21437 22419 21471
rect 1869 21369 1903 21403
rect 2145 21369 2179 21403
rect 2697 21369 2731 21403
rect 5365 21369 5399 21403
rect 6837 21369 6871 21403
rect 13737 21369 13771 21403
rect 21649 21369 21683 21403
rect 4721 21301 4755 21335
rect 5825 21301 5859 21335
rect 6469 21301 6503 21335
rect 7389 21301 7423 21335
rect 8401 21301 8435 21335
rect 9229 21301 9263 21335
rect 13553 21301 13587 21335
rect 14105 21301 14139 21335
rect 17785 21301 17819 21335
rect 21833 21301 21867 21335
rect 22661 21301 22695 21335
rect 23029 21301 23063 21335
rect 3985 21097 4019 21131
rect 4353 21097 4387 21131
rect 8033 21097 8067 21131
rect 9781 21097 9815 21131
rect 9965 21097 9999 21131
rect 12817 21097 12851 21131
rect 13737 21097 13771 21131
rect 14473 21097 14507 21131
rect 17049 21097 17083 21131
rect 18061 21097 18095 21131
rect 18613 21097 18647 21131
rect 20085 21097 20119 21131
rect 22661 21097 22695 21131
rect 2789 21029 2823 21063
rect 14105 21029 14139 21063
rect 17233 21029 17267 21063
rect 4813 20961 4847 20995
rect 7297 20961 7331 20995
rect 8585 20961 8619 20995
rect 9137 20961 9171 20995
rect 10057 20961 10091 20995
rect 10520 20961 10554 20995
rect 12265 20961 12299 20995
rect 12357 20961 12391 20995
rect 13553 20961 13587 20995
rect 14565 20961 14599 20995
rect 15071 20961 15105 20995
rect 17877 20961 17911 20995
rect 19349 20961 19383 20995
rect 19533 20961 19567 20995
rect 20916 20961 20950 20995
rect 3617 20893 3651 20927
rect 4169 20893 4203 20927
rect 6837 20893 6871 20927
rect 10793 20893 10827 20927
rect 13921 20893 13955 20927
rect 14289 20893 14323 20927
rect 15301 20893 15335 20927
rect 18245 20893 18279 20927
rect 18521 20893 18555 20927
rect 18797 20893 18831 20927
rect 20269 20893 20303 20927
rect 20453 20893 20487 20927
rect 21189 20893 21223 20927
rect 22477 20893 22511 20927
rect 22845 20893 22879 20927
rect 3341 20825 3375 20859
rect 6570 20825 6604 20859
rect 7113 20825 7147 20859
rect 7573 20825 7607 20859
rect 9321 20825 9355 20859
rect 13277 20825 13311 20859
rect 19073 20825 19107 20859
rect 19625 20825 19659 20859
rect 3893 20757 3927 20791
rect 4905 20757 4939 20791
rect 4997 20757 5031 20791
rect 5365 20757 5399 20791
rect 5457 20757 5491 20791
rect 7481 20757 7515 20791
rect 7941 20757 7975 20791
rect 8401 20757 8435 20791
rect 8493 20757 8527 20791
rect 9413 20757 9447 20791
rect 10523 20757 10557 20791
rect 11897 20757 11931 20791
rect 12449 20757 12483 20791
rect 12909 20757 12943 20791
rect 13369 20757 13403 20791
rect 15031 20757 15065 20791
rect 16405 20757 16439 20791
rect 16497 20757 16531 20791
rect 16773 20757 16807 20791
rect 17601 20757 17635 20791
rect 17693 20757 17727 20791
rect 18337 20757 18371 20791
rect 19993 20757 20027 20791
rect 20919 20757 20953 20791
rect 22293 20757 22327 20791
rect 23029 20757 23063 20791
rect 4721 20553 4755 20587
rect 7389 20553 7423 20587
rect 8683 20553 8717 20587
rect 10057 20553 10091 20587
rect 10701 20553 10735 20587
rect 11161 20553 11195 20587
rect 11989 20553 12023 20587
rect 13645 20553 13679 20587
rect 13737 20553 13771 20587
rect 14197 20553 14231 20587
rect 14749 20553 14783 20587
rect 15577 20553 15611 20587
rect 15945 20553 15979 20587
rect 17601 20553 17635 20587
rect 18343 20553 18377 20587
rect 19993 20553 20027 20587
rect 20637 20553 20671 20587
rect 21097 20553 21131 20587
rect 21281 20553 21315 20587
rect 6377 20485 6411 20519
rect 6561 20485 6595 20519
rect 22201 20485 22235 20519
rect 4445 20417 4479 20451
rect 5926 20417 5960 20451
rect 6745 20417 6779 20451
rect 7757 20417 7791 20451
rect 8953 20417 8987 20451
rect 10609 20417 10643 20451
rect 11529 20417 11563 20451
rect 11805 20417 11839 20451
rect 12449 20417 12483 20451
rect 13277 20417 13311 20451
rect 14105 20417 14139 20451
rect 15117 20417 15151 20451
rect 16037 20417 16071 20451
rect 17049 20417 17083 20451
rect 18613 20417 18647 20451
rect 20085 20417 20119 20451
rect 20729 20417 20763 20451
rect 21373 20417 21407 20451
rect 22845 20417 22879 20451
rect 6193 20349 6227 20383
rect 7849 20349 7883 20383
rect 8033 20349 8067 20383
rect 8217 20349 8251 20383
rect 8680 20351 8714 20385
rect 10793 20349 10827 20383
rect 12541 20349 12575 20383
rect 12725 20349 12759 20383
rect 13001 20349 13035 20383
rect 13185 20349 13219 20383
rect 14289 20349 14323 20383
rect 15209 20349 15243 20383
rect 15301 20349 15335 20383
rect 16129 20349 16163 20383
rect 17141 20349 17175 20383
rect 17233 20349 17267 20383
rect 17877 20349 17911 20383
rect 18340 20349 18374 20383
rect 20453 20349 20487 20383
rect 22293 20349 22327 20383
rect 22477 20349 22511 20383
rect 11713 20281 11747 20315
rect 21557 20281 21591 20315
rect 4261 20213 4295 20247
rect 4813 20213 4847 20247
rect 6929 20213 6963 20247
rect 7113 20213 7147 20247
rect 10241 20213 10275 20247
rect 12081 20213 12115 20247
rect 14565 20213 14599 20247
rect 16405 20213 16439 20247
rect 16681 20213 16715 20247
rect 19717 20213 19751 20247
rect 20269 20213 20303 20247
rect 21833 20213 21867 20247
rect 22661 20213 22695 20247
rect 23029 20213 23063 20247
rect 3249 20009 3283 20043
rect 9873 20009 9907 20043
rect 10885 20009 10919 20043
rect 11069 20009 11103 20043
rect 12265 20009 12299 20043
rect 14381 20009 14415 20043
rect 15209 20009 15243 20043
rect 16865 20009 16899 20043
rect 17693 20009 17727 20043
rect 18797 20009 18831 20043
rect 20821 20009 20855 20043
rect 22753 20009 22787 20043
rect 4077 19941 4111 19975
rect 10701 19941 10735 19975
rect 11989 19941 12023 19975
rect 12173 19941 12207 19975
rect 13461 19941 13495 19975
rect 14289 19941 14323 19975
rect 9229 19873 9263 19907
rect 11621 19873 11655 19907
rect 12909 19873 12943 19907
rect 13921 19873 13955 19907
rect 14933 19873 14967 19907
rect 15761 19873 15795 19907
rect 16129 19873 16163 19907
rect 17509 19873 17543 19907
rect 18153 19873 18187 19907
rect 18245 19873 18279 19907
rect 21376 19873 21410 19907
rect 21649 19873 21683 19907
rect 3065 19805 3099 19839
rect 3525 19805 3559 19839
rect 5457 19805 5491 19839
rect 6929 19805 6963 19839
rect 8134 19805 8168 19839
rect 8401 19805 8435 19839
rect 9413 19805 9447 19839
rect 13277 19805 13311 19839
rect 14105 19805 14139 19839
rect 15577 19805 15611 19839
rect 16405 19805 16439 19839
rect 17233 19805 17267 19839
rect 18061 19805 18095 19839
rect 18613 19805 18647 19839
rect 18889 19805 18923 19839
rect 19257 19805 19291 19839
rect 20913 19805 20947 19839
rect 22845 19805 22879 19839
rect 5190 19737 5224 19771
rect 6684 19737 6718 19771
rect 9505 19737 9539 19771
rect 11437 19737 11471 19771
rect 16313 19737 16347 19771
rect 17325 19737 17359 19771
rect 19524 19737 19558 19771
rect 3341 19669 3375 19703
rect 3985 19669 4019 19703
rect 5549 19669 5583 19703
rect 7021 19669 7055 19703
rect 8493 19669 8527 19703
rect 11161 19669 11195 19703
rect 11713 19669 11747 19703
rect 12633 19669 12667 19703
rect 12725 19669 12759 19703
rect 13093 19669 13127 19703
rect 13645 19669 13679 19703
rect 14749 19669 14783 19703
rect 14841 19669 14875 19703
rect 15669 19669 15703 19703
rect 16773 19669 16807 19703
rect 19073 19669 19107 19703
rect 20637 19669 20671 19703
rect 21379 19669 21413 19703
rect 23029 19669 23063 19703
rect 2881 19465 2915 19499
rect 4077 19465 4111 19499
rect 4445 19465 4479 19499
rect 4721 19465 4755 19499
rect 7757 19465 7791 19499
rect 11529 19465 11563 19499
rect 13461 19465 13495 19499
rect 14381 19465 14415 19499
rect 15853 19465 15887 19499
rect 16221 19465 16255 19499
rect 16497 19465 16531 19499
rect 16681 19465 16715 19499
rect 17049 19465 17083 19499
rect 17509 19465 17543 19499
rect 20637 19465 20671 19499
rect 21189 19465 21223 19499
rect 21833 19465 21867 19499
rect 2145 19397 2179 19431
rect 3249 19397 3283 19431
rect 15494 19397 15528 19431
rect 17141 19397 17175 19431
rect 18644 19397 18678 19431
rect 2237 19329 2271 19363
rect 3341 19329 3375 19363
rect 5834 19329 5868 19363
rect 8861 19329 8895 19363
rect 9274 19329 9308 19363
rect 10802 19329 10836 19363
rect 12653 19329 12687 19363
rect 13369 19329 13403 19363
rect 14013 19329 14047 19363
rect 15761 19329 15795 19363
rect 20094 19329 20128 19363
rect 20545 19329 20579 19363
rect 20821 19329 20855 19363
rect 21281 19329 21315 19363
rect 22201 19329 22235 19363
rect 22845 19329 22879 19363
rect 1961 19261 1995 19295
rect 3433 19261 3467 19295
rect 3893 19261 3927 19295
rect 3985 19261 4019 19295
rect 6101 19261 6135 19295
rect 9091 19261 9125 19295
rect 9597 19261 9631 19295
rect 11069 19261 11103 19295
rect 12909 19261 12943 19295
rect 13553 19261 13587 19295
rect 13829 19261 13863 19295
rect 17233 19261 17267 19295
rect 18889 19261 18923 19295
rect 20361 19261 20395 19295
rect 21097 19261 21131 19295
rect 22293 19261 22327 19295
rect 22477 19261 22511 19295
rect 2605 19193 2639 19227
rect 9689 19193 9723 19227
rect 6377 19125 6411 19159
rect 6561 19125 6595 19159
rect 6745 19125 6779 19159
rect 7021 19125 7055 19159
rect 7389 19125 7423 19159
rect 11161 19125 11195 19159
rect 13001 19125 13035 19159
rect 14289 19125 14323 19159
rect 18981 19125 19015 19159
rect 21649 19125 21683 19159
rect 22753 19125 22787 19159
rect 23029 19125 23063 19159
rect 3985 18921 4019 18955
rect 5917 18921 5951 18955
rect 7389 18921 7423 18955
rect 11069 18921 11103 18955
rect 13001 18921 13035 18955
rect 15761 18921 15795 18955
rect 19073 18921 19107 18955
rect 22385 18921 22419 18955
rect 3617 18853 3651 18887
rect 18705 18853 18739 18887
rect 20913 18853 20947 18887
rect 2053 18785 2087 18819
rect 3065 18785 3099 18819
rect 13921 18785 13955 18819
rect 15853 18785 15887 18819
rect 22937 18785 22971 18819
rect 5558 18717 5592 18751
rect 5825 18717 5859 18751
rect 7297 18717 7331 18751
rect 8513 18717 8547 18751
rect 8769 18717 8803 18751
rect 9689 18717 9723 18751
rect 11161 18717 11195 18751
rect 11437 18717 11471 18751
rect 11621 18717 11655 18751
rect 13645 18717 13679 18751
rect 14197 18717 14231 18751
rect 14381 18717 14415 18751
rect 17325 18717 17359 18751
rect 18889 18717 18923 18751
rect 19349 18717 19383 18751
rect 20821 18717 20855 18751
rect 22293 18717 22327 18751
rect 22845 18717 22879 18751
rect 3157 18649 3191 18683
rect 4169 18649 4203 18683
rect 4353 18649 4387 18683
rect 7052 18649 7086 18683
rect 9934 18649 9968 18683
rect 11888 18649 11922 18683
rect 14648 18649 14682 18683
rect 16120 18649 16154 18683
rect 17592 18649 17626 18683
rect 20554 18649 20588 18683
rect 22037 18649 22071 18683
rect 2237 18581 2271 18615
rect 2329 18581 2363 18615
rect 2697 18581 2731 18615
rect 3249 18581 3283 18615
rect 4445 18581 4479 18615
rect 8953 18581 8987 18615
rect 17233 18581 17267 18615
rect 19441 18581 19475 18615
rect 22753 18581 22787 18615
rect 2053 18377 2087 18411
rect 2145 18377 2179 18411
rect 8125 18377 8159 18411
rect 9689 18377 9723 18411
rect 11345 18377 11379 18411
rect 15577 18377 15611 18411
rect 16405 18377 16439 18411
rect 18061 18377 18095 18411
rect 19533 18377 19567 18411
rect 21373 18377 21407 18411
rect 21649 18377 21683 18411
rect 22293 18377 22327 18411
rect 22753 18377 22787 18411
rect 23029 18377 23063 18411
rect 6990 18309 7024 18343
rect 8462 18309 8496 18343
rect 10210 18309 10244 18343
rect 12756 18309 12790 18343
rect 13645 18309 13679 18343
rect 14372 18309 14406 18343
rect 18420 18309 18454 18343
rect 22201 18309 22235 18343
rect 1869 18241 1903 18275
rect 2329 18241 2363 18275
rect 3249 18241 3283 18275
rect 4465 18241 4499 18275
rect 4721 18241 4755 18275
rect 4813 18241 4847 18275
rect 5069 18241 5103 18275
rect 8217 18241 8251 18275
rect 9965 18241 9999 18275
rect 13001 18241 13035 18275
rect 13185 18241 13219 18275
rect 14105 18241 14139 18275
rect 15945 18241 15979 18275
rect 16681 18241 16715 18275
rect 16948 18241 16982 18275
rect 18153 18241 18187 18275
rect 19625 18241 19659 18275
rect 19892 18241 19926 18275
rect 21189 18241 21223 18275
rect 21465 18241 21499 18275
rect 22845 18241 22879 18275
rect 2973 18173 3007 18207
rect 6377 18173 6411 18207
rect 6561 18173 6595 18207
rect 6745 18173 6779 18207
rect 13737 18173 13771 18207
rect 13829 18173 13863 18207
rect 16037 18173 16071 18207
rect 16129 18173 16163 18207
rect 22385 18173 22419 18207
rect 13277 18105 13311 18139
rect 3341 18037 3375 18071
rect 6193 18037 6227 18071
rect 9597 18037 9631 18071
rect 11621 18037 11655 18071
rect 15485 18037 15519 18071
rect 21005 18037 21039 18071
rect 21833 18037 21867 18071
rect 1961 17833 1995 17867
rect 2881 17833 2915 17867
rect 3801 17833 3835 17867
rect 7481 17833 7515 17867
rect 9505 17833 9539 17867
rect 10977 17833 11011 17867
rect 12725 17833 12759 17867
rect 13921 17833 13955 17867
rect 15485 17833 15519 17867
rect 16957 17833 16991 17867
rect 20637 17833 20671 17867
rect 13737 17765 13771 17799
rect 19073 17765 19107 17799
rect 21465 17765 21499 17799
rect 2605 17697 2639 17731
rect 3341 17697 3375 17731
rect 3525 17697 3559 17731
rect 4261 17697 4295 17731
rect 4445 17697 4479 17731
rect 13369 17697 13403 17731
rect 15577 17697 15611 17731
rect 18429 17697 18463 17731
rect 19257 17697 19291 17731
rect 20913 17697 20947 17731
rect 21649 17697 21683 17731
rect 22845 17697 22879 17731
rect 22937 17697 22971 17731
rect 1777 17629 1811 17663
rect 2421 17629 2455 17663
rect 3249 17629 3283 17663
rect 4629 17629 4663 17663
rect 6101 17629 6135 17663
rect 10629 17629 10663 17663
rect 10885 17629 10919 17663
rect 12357 17629 12391 17663
rect 14105 17629 14139 17663
rect 15844 17629 15878 17663
rect 18162 17629 18196 17663
rect 18613 17629 18647 17663
rect 18889 17629 18923 17663
rect 21097 17629 21131 17663
rect 21833 17629 21867 17663
rect 4874 17561 4908 17595
rect 6368 17561 6402 17595
rect 12090 17561 12124 17595
rect 14372 17561 14406 17595
rect 19524 17561 19558 17595
rect 21925 17561 21959 17595
rect 22753 17561 22787 17595
rect 2053 17493 2087 17527
rect 2513 17493 2547 17527
rect 4169 17493 4203 17527
rect 6009 17493 6043 17527
rect 7665 17493 7699 17527
rect 8217 17493 8251 17527
rect 8493 17493 8527 17527
rect 12541 17493 12575 17527
rect 13093 17493 13127 17527
rect 13185 17493 13219 17527
rect 17049 17493 17083 17527
rect 18797 17493 18831 17527
rect 21005 17493 21039 17527
rect 22293 17493 22327 17527
rect 22385 17493 22419 17527
rect 2237 17289 2271 17323
rect 2697 17289 2731 17323
rect 3157 17289 3191 17323
rect 3617 17289 3651 17323
rect 8401 17289 8435 17323
rect 9873 17289 9907 17323
rect 12357 17289 12391 17323
rect 12541 17289 12575 17323
rect 14197 17289 14231 17323
rect 14565 17289 14599 17323
rect 17325 17289 17359 17323
rect 17601 17289 17635 17323
rect 19441 17289 19475 17323
rect 21189 17289 21223 17323
rect 22753 17289 22787 17323
rect 7288 17221 7322 17255
rect 8760 17221 8794 17255
rect 10232 17221 10266 17255
rect 11989 17221 12023 17255
rect 12900 17221 12934 17255
rect 15792 17221 15826 17255
rect 16221 17221 16255 17255
rect 16405 17221 16439 17255
rect 20576 17221 20610 17255
rect 2881 17153 2915 17187
rect 2973 17153 3007 17187
rect 3709 17153 3743 17187
rect 5926 17153 5960 17187
rect 11897 17153 11931 17187
rect 12633 17153 12667 17187
rect 16037 17153 16071 17187
rect 16865 17153 16899 17187
rect 17141 17153 17175 17187
rect 17417 17153 17451 17187
rect 17693 17153 17727 17187
rect 17969 17153 18003 17187
rect 18236 17153 18270 17187
rect 21281 17153 21315 17187
rect 22201 17153 22235 17187
rect 22845 17153 22879 17187
rect 2329 17085 2363 17119
rect 2513 17085 2547 17119
rect 3525 17085 3559 17119
rect 6193 17085 6227 17119
rect 7021 17085 7055 17119
rect 8493 17085 8527 17119
rect 9965 17085 9999 17119
rect 11805 17085 11839 17119
rect 20821 17085 20855 17119
rect 21097 17085 21131 17119
rect 21925 17085 21959 17119
rect 22109 17085 22143 17119
rect 23029 17085 23063 17119
rect 4721 17017 4755 17051
rect 11345 17017 11379 17051
rect 14657 17017 14691 17051
rect 1869 16949 1903 16983
rect 4077 16949 4111 16983
rect 4813 16949 4847 16983
rect 6377 16949 6411 16983
rect 14013 16949 14047 16983
rect 16773 16949 16807 16983
rect 17049 16949 17083 16983
rect 17877 16949 17911 16983
rect 19349 16949 19383 16983
rect 21649 16949 21683 16983
rect 22569 16949 22603 16983
rect 3801 16745 3835 16779
rect 8769 16745 8803 16779
rect 16681 16745 16715 16779
rect 18245 16745 18279 16779
rect 22477 16745 22511 16779
rect 22753 16745 22787 16779
rect 4629 16677 4663 16711
rect 2697 16609 2731 16643
rect 2973 16609 3007 16643
rect 3157 16609 3191 16643
rect 4261 16609 4295 16643
rect 4445 16609 4479 16643
rect 5457 16609 5491 16643
rect 11621 16609 11655 16643
rect 18061 16609 18095 16643
rect 20637 16609 20671 16643
rect 20729 16609 20763 16643
rect 22109 16609 22143 16643
rect 22201 16609 22235 16643
rect 3249 16541 3283 16575
rect 4813 16541 4847 16575
rect 7389 16541 7423 16575
rect 8953 16541 8987 16575
rect 9597 16541 9631 16575
rect 9781 16541 9815 16575
rect 11345 16541 11379 16575
rect 12265 16541 12299 16575
rect 13737 16541 13771 16575
rect 14749 16541 14783 16575
rect 15016 16541 15050 16575
rect 17794 16541 17828 16575
rect 18613 16541 18647 16575
rect 18889 16541 18923 16575
rect 21005 16541 21039 16575
rect 22661 16541 22695 16575
rect 23121 16541 23155 16575
rect 2421 16473 2455 16507
rect 5702 16473 5736 16507
rect 6929 16473 6963 16507
rect 7656 16473 7690 16507
rect 11078 16473 11112 16507
rect 20370 16473 20404 16507
rect 2053 16405 2087 16439
rect 2513 16405 2547 16439
rect 3617 16405 3651 16439
rect 4169 16405 4203 16439
rect 6837 16405 6871 16439
rect 9965 16405 9999 16439
rect 11713 16405 11747 16439
rect 11805 16405 11839 16439
rect 12173 16405 12207 16439
rect 16129 16405 16163 16439
rect 16313 16405 16347 16439
rect 16497 16405 16531 16439
rect 18521 16405 18555 16439
rect 18797 16405 18831 16439
rect 19073 16405 19107 16439
rect 19257 16405 19291 16439
rect 21649 16405 21683 16439
rect 22017 16405 22051 16439
rect 22937 16405 22971 16439
rect 1685 16201 1719 16235
rect 1961 16201 1995 16235
rect 2421 16201 2455 16235
rect 2881 16201 2915 16235
rect 3709 16201 3743 16235
rect 4169 16201 4203 16235
rect 4813 16201 4847 16235
rect 9873 16201 9907 16235
rect 14013 16201 14047 16235
rect 15669 16201 15703 16235
rect 15853 16201 15887 16235
rect 16221 16201 16255 16235
rect 16865 16201 16899 16235
rect 17049 16201 17083 16235
rect 17233 16201 17267 16235
rect 17509 16201 17543 16235
rect 17693 16201 17727 16235
rect 18245 16201 18279 16235
rect 21189 16201 21223 16235
rect 22569 16201 22603 16235
rect 3249 16133 3283 16167
rect 5926 16133 5960 16167
rect 9514 16133 9548 16167
rect 11529 16133 11563 16167
rect 13921 16133 13955 16167
rect 17877 16133 17911 16167
rect 21557 16133 21591 16167
rect 1501 16065 1535 16099
rect 1777 16065 1811 16099
rect 4077 16065 4111 16099
rect 9781 16065 9815 16099
rect 10997 16065 11031 16099
rect 11253 16065 11287 16099
rect 12265 16065 12299 16099
rect 12532 16065 12566 16099
rect 15137 16065 15171 16099
rect 15393 16065 15427 16099
rect 16497 16065 16531 16099
rect 19461 16065 19495 16099
rect 19717 16065 19751 16099
rect 19809 16065 19843 16099
rect 20065 16065 20099 16099
rect 21373 16065 21407 16099
rect 22109 16065 22143 16099
rect 22201 16065 22235 16099
rect 22845 16065 22879 16099
rect 23121 16065 23155 16099
rect 2237 15997 2271 16031
rect 2329 15997 2363 16031
rect 3341 15997 3375 16031
rect 3525 15997 3559 16031
rect 4261 15997 4295 16031
rect 6193 15997 6227 16031
rect 18061 15997 18095 16031
rect 21925 15997 21959 16031
rect 2789 15929 2823 15963
rect 22661 15929 22695 15963
rect 6377 15861 6411 15895
rect 8401 15861 8435 15895
rect 13645 15861 13679 15895
rect 18337 15861 18371 15895
rect 22937 15861 22971 15895
rect 1961 15657 1995 15691
rect 4261 15657 4295 15691
rect 10425 15657 10459 15691
rect 11989 15657 12023 15691
rect 12173 15657 12207 15691
rect 15485 15657 15519 15691
rect 17049 15657 17083 15691
rect 18613 15657 18647 15691
rect 20637 15657 20671 15691
rect 21465 15657 21499 15691
rect 17141 15589 17175 15623
rect 22753 15589 22787 15623
rect 2697 15521 2731 15555
rect 3525 15521 3559 15555
rect 11897 15521 11931 15555
rect 12541 15521 12575 15555
rect 18521 15521 18555 15555
rect 19257 15521 19291 15555
rect 20821 15521 20855 15555
rect 21005 15521 21039 15555
rect 22201 15521 22235 15555
rect 1685 15453 1719 15487
rect 1777 15453 1811 15487
rect 3249 15453 3283 15487
rect 4169 15453 4203 15487
rect 5374 15453 5408 15487
rect 5641 15453 5675 15487
rect 7113 15453 7147 15487
rect 7297 15453 7331 15487
rect 9045 15453 9079 15487
rect 9312 15453 9346 15487
rect 11630 15453 11664 15487
rect 14105 15453 14139 15487
rect 15669 15453 15703 15487
rect 15936 15453 15970 15487
rect 18889 15453 18923 15487
rect 19513 15453 19547 15487
rect 21097 15453 21131 15487
rect 21557 15453 21591 15487
rect 21741 15453 21775 15487
rect 21925 15453 21959 15487
rect 23029 15453 23063 15487
rect 2513 15385 2547 15419
rect 3341 15385 3375 15419
rect 6846 15385 6880 15419
rect 7542 15385 7576 15419
rect 12808 15385 12842 15419
rect 14372 15385 14406 15419
rect 18254 15385 18288 15419
rect 1501 15317 1535 15351
rect 2053 15317 2087 15351
rect 2421 15317 2455 15351
rect 2881 15317 2915 15351
rect 3985 15317 4019 15351
rect 5733 15317 5767 15351
rect 8677 15317 8711 15351
rect 10517 15317 10551 15351
rect 13921 15317 13955 15351
rect 19073 15317 19107 15351
rect 22293 15317 22327 15351
rect 22385 15317 22419 15351
rect 22845 15317 22879 15351
rect 1961 15113 1995 15147
rect 2881 15113 2915 15147
rect 4813 15113 4847 15147
rect 11345 15113 11379 15147
rect 13185 15113 13219 15147
rect 16037 15113 16071 15147
rect 18245 15113 18279 15147
rect 19809 15113 19843 15147
rect 20637 15113 20671 15147
rect 21465 15113 21499 15147
rect 21649 15113 21683 15147
rect 22109 15113 22143 15147
rect 3249 15045 3283 15079
rect 8738 15045 8772 15079
rect 10232 15045 10266 15079
rect 14298 15045 14332 15079
rect 16129 15045 16163 15079
rect 16313 15045 16347 15079
rect 16948 15045 16982 15079
rect 20177 15045 20211 15079
rect 22845 15045 22879 15079
rect 1777 14977 1811 15011
rect 2421 14977 2455 15011
rect 4261 14977 4295 15011
rect 5926 14977 5960 15011
rect 14565 14977 14599 15011
rect 14657 14977 14691 15011
rect 14924 14977 14958 15011
rect 16681 14977 16715 15011
rect 18429 14977 18463 15011
rect 18696 14977 18730 15011
rect 20269 14977 20303 15011
rect 21097 14977 21131 15011
rect 22201 14977 22235 15011
rect 2145 14909 2179 14943
rect 2329 14909 2363 14943
rect 3341 14909 3375 14943
rect 3525 14909 3559 14943
rect 4537 14909 4571 14943
rect 6193 14909 6227 14943
rect 8493 14909 8527 14943
rect 9965 14909 9999 14943
rect 20085 14909 20119 14943
rect 20821 14909 20855 14943
rect 21005 14909 21039 14943
rect 22017 14909 22051 14943
rect 22661 14909 22695 14943
rect 2789 14841 2823 14875
rect 11529 14841 11563 14875
rect 18061 14841 18095 14875
rect 22569 14841 22603 14875
rect 6377 14773 6411 14807
rect 6561 14773 6595 14807
rect 7205 14773 7239 14807
rect 8309 14773 8343 14807
rect 9873 14773 9907 14807
rect 23121 14773 23155 14807
rect 1685 14569 1719 14603
rect 2881 14569 2915 14603
rect 12265 14569 12299 14603
rect 15485 14569 15519 14603
rect 17141 14569 17175 14603
rect 18797 14569 18831 14603
rect 18981 14569 19015 14603
rect 21465 14569 21499 14603
rect 23029 14569 23063 14603
rect 1961 14501 1995 14535
rect 4813 14501 4847 14535
rect 6377 14501 6411 14535
rect 9137 14501 9171 14535
rect 18705 14501 18739 14535
rect 2605 14433 2639 14467
rect 3525 14433 3559 14467
rect 4445 14433 4479 14467
rect 16957 14433 16991 14467
rect 19257 14433 19291 14467
rect 20913 14433 20947 14467
rect 22385 14433 22419 14467
rect 1501 14365 1535 14399
rect 1777 14365 1811 14399
rect 2513 14365 2547 14399
rect 3249 14365 3283 14399
rect 3341 14365 3375 14399
rect 6193 14365 6227 14399
rect 7757 14365 7791 14399
rect 7849 14365 7883 14399
rect 10517 14365 10551 14399
rect 13378 14365 13412 14399
rect 13645 14365 13679 14399
rect 13829 14365 13863 14399
rect 14105 14365 14139 14399
rect 19524 14365 19558 14399
rect 21649 14365 21683 14399
rect 21833 14365 21867 14399
rect 22109 14365 22143 14399
rect 2421 14297 2455 14331
rect 4169 14297 4203 14331
rect 4261 14297 4295 14331
rect 5948 14297 5982 14331
rect 7490 14297 7524 14331
rect 10250 14297 10284 14331
rect 14372 14297 14406 14331
rect 16690 14297 16724 14331
rect 18337 14297 18371 14331
rect 21097 14297 21131 14331
rect 2053 14229 2087 14263
rect 3801 14229 3835 14263
rect 10609 14229 10643 14263
rect 10793 14229 10827 14263
rect 10977 14229 11011 14263
rect 11437 14229 11471 14263
rect 15577 14229 15611 14263
rect 18521 14229 18555 14263
rect 20637 14229 20671 14263
rect 21005 14229 21039 14263
rect 22017 14229 22051 14263
rect 2329 14025 2363 14059
rect 2697 14025 2731 14059
rect 3157 14025 3191 14059
rect 3525 14025 3559 14059
rect 3985 14025 4019 14059
rect 4813 14025 4847 14059
rect 8493 14025 8527 14059
rect 9965 14025 9999 14059
rect 11529 14025 11563 14059
rect 14749 14025 14783 14059
rect 16773 14025 16807 14059
rect 17049 14025 17083 14059
rect 17785 14025 17819 14059
rect 21557 14025 21591 14059
rect 22937 14025 22971 14059
rect 2789 13957 2823 13991
rect 9606 13957 9640 13991
rect 12664 13957 12698 13991
rect 14933 13957 14967 13991
rect 21097 13957 21131 13991
rect 22109 13957 22143 13991
rect 3617 13889 3651 13923
rect 4353 13889 4387 13923
rect 5937 13889 5971 13923
rect 7858 13889 7892 13923
rect 8125 13889 8159 13923
rect 11078 13889 11112 13923
rect 11345 13889 11379 13923
rect 12909 13889 12943 13923
rect 13093 13889 13127 13923
rect 13369 13889 13403 13923
rect 13636 13889 13670 13923
rect 15117 13889 15151 13923
rect 15384 13889 15418 13923
rect 18909 13889 18943 13923
rect 19165 13889 19199 13923
rect 20381 13889 20415 13923
rect 20637 13889 20671 13923
rect 22201 13889 22235 13923
rect 22661 13889 22695 13923
rect 23121 13889 23155 13923
rect 2881 13821 2915 13855
rect 3801 13821 3835 13855
rect 4445 13821 4479 13855
rect 4629 13821 4663 13855
rect 6193 13821 6227 13855
rect 9873 13821 9907 13855
rect 20821 13821 20855 13855
rect 21005 13821 21039 13855
rect 22017 13821 22051 13855
rect 6745 13753 6779 13787
rect 16497 13753 16531 13787
rect 19257 13753 19291 13787
rect 21465 13753 21499 13787
rect 22569 13753 22603 13787
rect 6377 13685 6411 13719
rect 6561 13685 6595 13719
rect 8217 13685 8251 13719
rect 22845 13685 22879 13719
rect 1869 13481 1903 13515
rect 2605 13481 2639 13515
rect 6285 13481 6319 13515
rect 10517 13481 10551 13515
rect 11989 13481 12023 13515
rect 12173 13481 12207 13515
rect 19257 13481 19291 13515
rect 21557 13481 21591 13515
rect 22477 13481 22511 13515
rect 22845 13481 22879 13515
rect 6377 13413 6411 13447
rect 14105 13413 14139 13447
rect 18429 13413 18463 13447
rect 3157 13345 3191 13379
rect 11897 13345 11931 13379
rect 18613 13345 18647 13379
rect 18705 13345 18739 13379
rect 20637 13345 20671 13379
rect 20913 13345 20947 13379
rect 21925 13345 21959 13379
rect 2053 13277 2087 13311
rect 2973 13277 3007 13311
rect 4721 13277 4755 13311
rect 4905 13277 4939 13311
rect 5172 13277 5206 13311
rect 7757 13277 7791 13311
rect 8953 13277 8987 13311
rect 15485 13277 15519 13311
rect 15577 13277 15611 13311
rect 17049 13277 17083 13311
rect 18889 13277 18923 13311
rect 20381 13277 20415 13311
rect 22109 13277 22143 13311
rect 22569 13253 22603 13287
rect 23029 13277 23063 13311
rect 7490 13209 7524 13243
rect 9198 13209 9232 13243
rect 11630 13209 11664 13243
rect 15240 13209 15274 13243
rect 15844 13209 15878 13243
rect 17316 13209 17350 13243
rect 21097 13209 21131 13243
rect 2145 13141 2179 13175
rect 3065 13141 3099 13175
rect 4629 13141 4663 13175
rect 7849 13141 7883 13175
rect 10333 13141 10367 13175
rect 16957 13141 16991 13175
rect 19073 13141 19107 13175
rect 21005 13141 21039 13175
rect 21465 13141 21499 13175
rect 22017 13141 22051 13175
rect 22753 13141 22787 13175
rect 2513 12937 2547 12971
rect 3801 12937 3835 12971
rect 4169 12937 4203 12971
rect 6377 12937 6411 12971
rect 8401 12937 8435 12971
rect 13093 12937 13127 12971
rect 16313 12937 16347 12971
rect 16497 12937 16531 12971
rect 18245 12937 18279 12971
rect 21189 12937 21223 12971
rect 22109 12937 22143 12971
rect 22569 12937 22603 12971
rect 23121 12937 23155 12971
rect 5181 12869 5215 12903
rect 7266 12869 7300 12903
rect 17816 12869 17850 12903
rect 21465 12869 21499 12903
rect 2881 12801 2915 12835
rect 3709 12801 3743 12835
rect 4537 12801 4571 12835
rect 4629 12801 4663 12835
rect 7021 12801 7055 12835
rect 9606 12801 9640 12835
rect 11089 12801 11123 12835
rect 11345 12801 11379 12835
rect 12745 12801 12779 12835
rect 13001 12801 13035 12835
rect 13277 12801 13311 12835
rect 13544 12801 13578 12835
rect 14749 12801 14783 12835
rect 15016 12801 15050 12835
rect 18061 12801 18095 12835
rect 18337 12801 18371 12835
rect 18604 12801 18638 12835
rect 19809 12801 19843 12835
rect 20076 12801 20110 12835
rect 22201 12801 22235 12835
rect 22845 12801 22879 12835
rect 22937 12801 22971 12835
rect 2973 12733 3007 12767
rect 3157 12733 3191 12767
rect 3893 12733 3927 12767
rect 4813 12733 4847 12767
rect 9873 12733 9907 12767
rect 21281 12733 21315 12767
rect 21925 12733 21959 12767
rect 4997 12665 5031 12699
rect 8493 12665 8527 12699
rect 11621 12665 11655 12699
rect 14657 12665 14691 12699
rect 16129 12665 16163 12699
rect 3341 12597 3375 12631
rect 9965 12597 9999 12631
rect 16681 12597 16715 12631
rect 19717 12597 19751 12631
rect 22661 12597 22695 12631
rect 2053 12393 2087 12427
rect 3801 12393 3835 12427
rect 18521 12393 18555 12427
rect 17693 12325 17727 12359
rect 18797 12325 18831 12359
rect 19073 12325 19107 12359
rect 2697 12257 2731 12291
rect 3065 12257 3099 12291
rect 4721 12257 4755 12291
rect 14197 12257 14231 12291
rect 14841 12257 14875 12291
rect 16313 12257 16347 12291
rect 19257 12257 19291 12291
rect 20821 12257 20855 12291
rect 21649 12257 21683 12291
rect 22845 12257 22879 12291
rect 22937 12257 22971 12291
rect 3985 12189 4019 12223
rect 4905 12189 4939 12223
rect 6377 12189 6411 12223
rect 10057 12189 10091 12223
rect 12541 12189 12575 12223
rect 16580 12189 16614 12223
rect 18337 12189 18371 12223
rect 18613 12189 18647 12223
rect 18889 12189 18923 12223
rect 19513 12189 19547 12223
rect 21097 12189 21131 12223
rect 21925 12189 21959 12223
rect 22753 12189 22787 12223
rect 2421 12121 2455 12155
rect 3249 12121 3283 12155
rect 4537 12121 4571 12155
rect 5172 12121 5206 12155
rect 6622 12121 6656 12155
rect 10324 12121 10358 12155
rect 11529 12121 11563 12155
rect 11713 12121 11747 12155
rect 12808 12121 12842 12155
rect 17877 12121 17911 12155
rect 18153 12121 18187 12155
rect 21005 12121 21039 12155
rect 21833 12121 21867 12155
rect 2513 12053 2547 12087
rect 3157 12053 3191 12087
rect 3617 12053 3651 12087
rect 4077 12053 4111 12087
rect 4445 12053 4479 12087
rect 6285 12053 6319 12087
rect 7757 12053 7791 12087
rect 7849 12053 7883 12087
rect 8493 12053 8527 12087
rect 9229 12053 9263 12087
rect 9873 12053 9907 12087
rect 11437 12053 11471 12087
rect 13921 12053 13955 12087
rect 20637 12053 20671 12087
rect 21465 12053 21499 12087
rect 22293 12053 22327 12087
rect 22385 12053 22419 12087
rect 2605 11849 2639 11883
rect 2881 11849 2915 11883
rect 3617 11849 3651 11883
rect 3985 11849 4019 11883
rect 6377 11849 6411 11883
rect 10609 11849 10643 11883
rect 12909 11849 12943 11883
rect 17049 11849 17083 11883
rect 20453 11849 20487 11883
rect 20913 11849 20947 11883
rect 22201 11849 22235 11883
rect 3525 11781 3559 11815
rect 11774 11781 11808 11815
rect 16865 11781 16899 11815
rect 19340 11781 19374 11815
rect 20821 11781 20855 11815
rect 21557 11781 21591 11815
rect 2789 11713 2823 11747
rect 3065 11713 3099 11747
rect 4353 11713 4387 11747
rect 5926 11713 5960 11747
rect 6193 11713 6227 11747
rect 6561 11713 6595 11747
rect 8024 11713 8058 11747
rect 9229 11713 9263 11747
rect 9485 11713 9519 11747
rect 15770 11713 15804 11747
rect 18254 11713 18288 11747
rect 18797 11713 18831 11747
rect 22293 11713 22327 11747
rect 22845 11713 22879 11747
rect 23121 11713 23155 11747
rect 3709 11645 3743 11679
rect 4445 11645 4479 11679
rect 4629 11645 4663 11679
rect 7757 11645 7791 11679
rect 10701 11645 10735 11679
rect 11529 11645 11563 11679
rect 16037 11645 16071 11679
rect 18521 11645 18555 11679
rect 19073 11645 19107 11679
rect 20729 11645 20763 11679
rect 22385 11645 22419 11679
rect 3157 11577 3191 11611
rect 21373 11577 21407 11611
rect 22937 11577 22971 11611
rect 4813 11509 4847 11543
rect 9137 11509 9171 11543
rect 13093 11509 13127 11543
rect 13185 11509 13219 11543
rect 14657 11509 14691 11543
rect 16129 11509 16163 11543
rect 16497 11509 16531 11543
rect 17141 11509 17175 11543
rect 18705 11509 18739 11543
rect 18981 11509 19015 11543
rect 21281 11509 21315 11543
rect 21833 11509 21867 11543
rect 22661 11509 22695 11543
rect 3617 11305 3651 11339
rect 4261 11305 4295 11339
rect 5273 11305 5307 11339
rect 9045 11305 9079 11339
rect 12449 11305 12483 11339
rect 13921 11305 13955 11339
rect 19073 11305 19107 11339
rect 23029 11305 23063 11339
rect 6745 11237 6779 11271
rect 18429 11237 18463 11271
rect 20637 11237 20671 11271
rect 20729 11237 20763 11271
rect 22937 11237 22971 11271
rect 3065 11169 3099 11203
rect 4813 11169 4847 11203
rect 22109 11169 22143 11203
rect 22385 11169 22419 11203
rect 3249 11101 3283 11135
rect 4629 11101 4663 11135
rect 6653 11101 6687 11135
rect 8125 11101 8159 11135
rect 10425 11101 10459 11135
rect 11069 11101 11103 11135
rect 12541 11101 12575 11135
rect 14105 11101 14139 11135
rect 14841 11101 14875 11135
rect 15025 11101 15059 11135
rect 16497 11101 16531 11135
rect 16681 11101 16715 11135
rect 16865 11101 16899 11135
rect 17049 11101 17083 11135
rect 18889 11101 18923 11135
rect 19257 11101 19291 11135
rect 19524 11101 19558 11135
rect 22569 11101 22603 11135
rect 4721 11033 4755 11067
rect 6386 11033 6420 11067
rect 7858 11033 7892 11067
rect 10158 11033 10192 11067
rect 11336 11033 11370 11067
rect 12786 11033 12820 11067
rect 15292 11033 15326 11067
rect 17316 11033 17350 11067
rect 21842 11033 21876 11067
rect 22477 11033 22511 11067
rect 3157 10965 3191 10999
rect 8309 10965 8343 10999
rect 10517 10965 10551 10999
rect 16405 10965 16439 10999
rect 18705 10965 18739 10999
rect 3065 10761 3099 10795
rect 3893 10761 3927 10795
rect 5457 10761 5491 10795
rect 6193 10761 6227 10795
rect 6745 10761 6779 10795
rect 13553 10761 13587 10795
rect 22477 10761 22511 10795
rect 22569 10761 22603 10795
rect 4261 10693 4295 10727
rect 9606 10693 9640 10727
rect 11100 10693 11134 10727
rect 12440 10693 12474 10727
rect 14780 10693 14814 10727
rect 20821 10693 20855 10727
rect 21281 10693 21315 10727
rect 3249 10625 3283 10659
rect 4353 10625 4387 10659
rect 5549 10625 5583 10659
rect 8145 10625 8179 10659
rect 15025 10625 15059 10659
rect 16241 10625 16275 10659
rect 16497 10625 16531 10659
rect 16681 10625 16715 10659
rect 16937 10625 16971 10659
rect 18337 10625 18371 10659
rect 19156 10625 19190 10659
rect 20637 10625 20671 10659
rect 21833 10625 21867 10659
rect 23121 10625 23155 10659
rect 4537 10557 4571 10591
rect 4813 10557 4847 10591
rect 8401 10557 8435 10591
rect 9873 10557 9907 10591
rect 11345 10557 11379 10591
rect 12173 10557 12207 10591
rect 18797 10557 18831 10591
rect 18889 10557 18923 10591
rect 21373 10557 21407 10591
rect 21465 10557 21499 10591
rect 22661 10557 22695 10591
rect 8493 10489 8527 10523
rect 18061 10489 18095 10523
rect 18245 10489 18279 10523
rect 20453 10489 20487 10523
rect 7021 10421 7055 10455
rect 9965 10421 9999 10455
rect 11529 10421 11563 10455
rect 11713 10421 11747 10455
rect 13645 10421 13679 10455
rect 15117 10421 15151 10455
rect 18521 10421 18555 10455
rect 20269 10421 20303 10455
rect 20913 10421 20947 10455
rect 22017 10421 22051 10455
rect 22109 10421 22143 10455
rect 22937 10421 22971 10455
rect 2513 10217 2547 10251
rect 2789 10217 2823 10251
rect 5089 10217 5123 10251
rect 8953 10217 8987 10251
rect 17233 10217 17267 10251
rect 17417 10217 17451 10251
rect 17693 10217 17727 10251
rect 2881 10149 2915 10183
rect 5365 10149 5399 10183
rect 17049 10149 17083 10183
rect 17969 10149 18003 10183
rect 3433 10081 3467 10115
rect 4445 10081 4479 10115
rect 6745 10081 6779 10115
rect 6837 10081 6871 10115
rect 15577 10081 15611 10115
rect 15669 10081 15703 10115
rect 18889 10081 18923 10115
rect 20637 10081 20671 10115
rect 21281 10081 21315 10115
rect 21925 10081 21959 10115
rect 22201 10081 22235 10115
rect 22385 10081 22419 10115
rect 2329 10013 2363 10047
rect 2605 10013 2639 10047
rect 4261 10013 4295 10047
rect 4813 10013 4847 10047
rect 9505 10013 9539 10047
rect 11529 10013 11563 10047
rect 11621 10013 11655 10047
rect 13093 10013 13127 10047
rect 13645 10013 13679 10047
rect 15321 10013 15355 10047
rect 17785 10013 17819 10047
rect 18061 10013 18095 10047
rect 18613 10013 18647 10047
rect 22477 10013 22511 10047
rect 23121 10013 23155 10047
rect 4169 9945 4203 9979
rect 6478 9945 6512 9979
rect 7104 9945 7138 9979
rect 9965 9945 9999 9979
rect 11262 9945 11296 9979
rect 11866 9945 11900 9979
rect 15936 9945 15970 9979
rect 18521 9945 18555 9979
rect 20370 9945 20404 9979
rect 21557 9945 21591 9979
rect 21741 9945 21775 9979
rect 3249 9877 3283 9911
rect 3341 9877 3375 9911
rect 3801 9877 3835 9911
rect 4721 9877 4755 9911
rect 8217 9877 8251 9911
rect 8401 9877 8435 9911
rect 8493 9877 8527 9911
rect 10149 9877 10183 9911
rect 13001 9877 13035 9911
rect 14197 9877 14231 9911
rect 18245 9877 18279 9911
rect 19257 9877 19291 9911
rect 20729 9877 20763 9911
rect 21097 9877 21131 9911
rect 21189 9877 21223 9911
rect 22845 9877 22879 9911
rect 22937 9877 22971 9911
rect 4721 9673 4755 9707
rect 6377 9673 6411 9707
rect 6653 9673 6687 9707
rect 21373 9673 21407 9707
rect 22661 9673 22695 9707
rect 2973 9605 3007 9639
rect 10517 9605 10551 9639
rect 22293 9605 22327 9639
rect 1409 9537 1443 9571
rect 1685 9537 1719 9571
rect 2881 9537 2915 9571
rect 3597 9537 3631 9571
rect 4813 9537 4847 9571
rect 5069 9537 5103 9571
rect 7573 9537 7607 9571
rect 7840 9537 7874 9571
rect 9312 9537 9346 9571
rect 12642 9537 12676 9571
rect 12909 9537 12943 9571
rect 14114 9537 14148 9571
rect 14381 9537 14415 9571
rect 14473 9537 14507 9571
rect 15117 9537 15151 9571
rect 15384 9537 15418 9571
rect 17141 9537 17175 9571
rect 18530 9537 18564 9571
rect 19145 9537 19179 9571
rect 20821 9537 20855 9571
rect 20913 9537 20947 9571
rect 21557 9537 21591 9571
rect 22201 9537 22235 9571
rect 22845 9537 22879 9571
rect 23121 9537 23155 9571
rect 3065 9469 3099 9503
rect 3348 9469 3382 9503
rect 6929 9469 6963 9503
rect 9045 9469 9079 9503
rect 11345 9469 11379 9503
rect 18797 9469 18831 9503
rect 18889 9469 18923 9503
rect 20637 9469 20671 9503
rect 22477 9469 22511 9503
rect 1593 9401 1627 9435
rect 16681 9401 16715 9435
rect 16865 9401 16899 9435
rect 17233 9401 17267 9435
rect 21833 9401 21867 9435
rect 2513 9333 2547 9367
rect 6193 9333 6227 9367
rect 7481 9333 7515 9367
rect 8953 9333 8987 9367
rect 10425 9333 10459 9367
rect 10701 9333 10735 9367
rect 11529 9333 11563 9367
rect 13001 9333 13035 9367
rect 16497 9333 16531 9367
rect 17417 9333 17451 9367
rect 20269 9333 20303 9367
rect 20453 9333 20487 9367
rect 21281 9333 21315 9367
rect 22937 9333 22971 9367
rect 2789 9129 2823 9163
rect 5457 9129 5491 9163
rect 7021 9129 7055 9163
rect 7205 9129 7239 9163
rect 9045 9129 9079 9163
rect 13185 9129 13219 9163
rect 13369 9129 13403 9163
rect 19073 9129 19107 9163
rect 21465 9129 21499 9163
rect 22385 9129 22419 9163
rect 2881 9061 2915 9095
rect 2237 8993 2271 9027
rect 3433 8993 3467 9027
rect 6929 8993 6963 9027
rect 7389 8993 7423 9027
rect 10057 8993 10091 9027
rect 13093 8993 13127 9027
rect 17785 8993 17819 9027
rect 18705 8993 18739 9027
rect 20913 8993 20947 9027
rect 21649 8993 21683 9027
rect 22937 8993 22971 9027
rect 2421 8925 2455 8959
rect 4077 8925 4111 8959
rect 7645 8925 7679 8959
rect 9413 8925 9447 8959
rect 16313 8925 16347 8959
rect 18061 8925 18095 8959
rect 20637 8925 20671 8959
rect 21097 8925 21131 8959
rect 21925 8925 21959 8959
rect 22753 8925 22787 8959
rect 2329 8857 2363 8891
rect 3249 8857 3283 8891
rect 4344 8857 4378 8891
rect 6662 8857 6696 8891
rect 9965 8857 9999 8891
rect 10302 8857 10336 8891
rect 12826 8857 12860 8891
rect 16046 8857 16080 8891
rect 17518 8857 17552 8891
rect 20370 8857 20404 8891
rect 21833 8857 21867 8891
rect 22845 8857 22879 8891
rect 3341 8789 3375 8823
rect 5549 8789 5583 8823
rect 8769 8789 8803 8823
rect 11437 8789 11471 8823
rect 11529 8789 11563 8823
rect 11713 8789 11747 8823
rect 14933 8789 14967 8823
rect 16405 8789 16439 8823
rect 19257 8789 19291 8823
rect 21005 8789 21039 8823
rect 22293 8789 22327 8823
rect 1961 8585 1995 8619
rect 2513 8585 2547 8619
rect 3341 8585 3375 8619
rect 6193 8585 6227 8619
rect 14289 8585 14323 8619
rect 17509 8585 17543 8619
rect 21557 8585 21591 8619
rect 21833 8585 21867 8619
rect 2973 8517 3007 8551
rect 8156 8517 8190 8551
rect 11529 8517 11563 8551
rect 19524 8517 19558 8551
rect 22385 8517 22419 8551
rect 22937 8517 22971 8551
rect 2053 8449 2087 8483
rect 2881 8449 2915 8483
rect 4465 8449 4499 8483
rect 5069 8449 5103 8483
rect 9606 8449 9640 8483
rect 9873 8449 9907 8483
rect 9965 8449 9999 8483
rect 10232 8449 10266 8483
rect 12918 8449 12952 8483
rect 13185 8449 13219 8483
rect 13277 8449 13311 8483
rect 15413 8449 15447 8483
rect 18909 8449 18943 8483
rect 21097 8449 21131 8483
rect 21189 8449 21223 8483
rect 22661 8449 22695 8483
rect 1869 8381 1903 8415
rect 3157 8381 3191 8415
rect 4721 8381 4755 8415
rect 4813 8381 4847 8415
rect 8401 8381 8435 8415
rect 15669 8381 15703 8415
rect 19165 8381 19199 8415
rect 19257 8381 19291 8415
rect 21281 8381 21315 8415
rect 2421 8313 2455 8347
rect 6377 8313 6411 8347
rect 6561 8313 6595 8347
rect 6837 8313 6871 8347
rect 11805 8313 11839 8347
rect 15853 8313 15887 8347
rect 16037 8313 16071 8347
rect 16313 8313 16347 8347
rect 16497 8313 16531 8347
rect 16773 8313 16807 8347
rect 16957 8313 16991 8347
rect 17141 8313 17175 8347
rect 17325 8313 17359 8347
rect 17693 8313 17727 8347
rect 20729 8313 20763 8347
rect 22753 8313 22787 8347
rect 7021 8245 7055 8279
rect 8493 8245 8527 8279
rect 11345 8245 11379 8279
rect 17785 8245 17819 8279
rect 20637 8245 20671 8279
rect 2053 8041 2087 8075
rect 2881 8041 2915 8075
rect 5825 8041 5859 8075
rect 7389 8041 7423 8075
rect 18613 8041 18647 8075
rect 18429 7973 18463 8007
rect 22569 7973 22603 8007
rect 2697 7905 2731 7939
rect 3433 7905 3467 7939
rect 21192 7905 21226 7939
rect 21465 7905 21499 7939
rect 2513 7837 2547 7871
rect 4445 7837 4479 7871
rect 5917 7837 5951 7871
rect 8769 7837 8803 7871
rect 8953 7837 8987 7871
rect 9137 7837 9171 7871
rect 9321 7837 9355 7871
rect 9505 7837 9539 7871
rect 10977 7837 11011 7871
rect 12449 7837 12483 7871
rect 14105 7837 14139 7871
rect 15577 7837 15611 7871
rect 17049 7837 17083 7871
rect 18797 7837 18831 7871
rect 18889 7837 18923 7871
rect 20637 7837 20671 7871
rect 20729 7837 20763 7871
rect 23029 7837 23063 7871
rect 3249 7769 3283 7803
rect 4690 7769 4724 7803
rect 6184 7769 6218 7803
rect 8502 7769 8536 7803
rect 9772 7769 9806 7803
rect 11244 7769 11278 7803
rect 12694 7769 12728 7803
rect 14350 7769 14384 7803
rect 15822 7769 15856 7803
rect 17294 7769 17328 7803
rect 20370 7769 20404 7803
rect 2421 7701 2455 7735
rect 3341 7701 3375 7735
rect 7297 7701 7331 7735
rect 10885 7701 10919 7735
rect 12357 7701 12391 7735
rect 13829 7701 13863 7735
rect 15485 7701 15519 7735
rect 16957 7701 16991 7735
rect 19073 7701 19107 7735
rect 19257 7701 19291 7735
rect 21195 7701 21229 7735
rect 22661 7701 22695 7735
rect 22937 7701 22971 7735
rect 4813 7497 4847 7531
rect 9873 7497 9907 7531
rect 10333 7497 10367 7531
rect 10701 7497 10735 7531
rect 10977 7497 11011 7531
rect 11805 7497 11839 7531
rect 13369 7497 13403 7531
rect 16037 7497 16071 7531
rect 21097 7497 21131 7531
rect 23029 7497 23063 7531
rect 5926 7429 5960 7463
rect 10241 7429 10275 7463
rect 12234 7429 12268 7463
rect 14013 7429 14047 7463
rect 14197 7429 14231 7463
rect 16948 7429 16982 7463
rect 3341 7361 3375 7395
rect 3608 7361 3642 7395
rect 6193 7361 6227 7395
rect 6377 7361 6411 7395
rect 6561 7361 6595 7395
rect 6745 7361 6779 7395
rect 6929 7361 6963 7395
rect 7196 7361 7230 7395
rect 8401 7361 8435 7395
rect 8668 7361 8702 7395
rect 11989 7361 12023 7395
rect 13645 7361 13679 7395
rect 14473 7361 14507 7395
rect 14740 7361 14774 7395
rect 16313 7361 16347 7395
rect 18153 7361 18187 7395
rect 18409 7361 18443 7395
rect 19892 7361 19926 7395
rect 21557 7361 21591 7395
rect 22201 7361 22235 7395
rect 22845 7361 22879 7395
rect 10425 7293 10459 7327
rect 16681 7293 16715 7327
rect 19625 7293 19659 7327
rect 21925 7293 21959 7327
rect 22109 7293 22143 7327
rect 9781 7225 9815 7259
rect 21005 7225 21039 7259
rect 22569 7225 22603 7259
rect 4721 7157 4755 7191
rect 8309 7157 8343 7191
rect 13553 7157 13587 7191
rect 15853 7157 15887 7191
rect 16221 7157 16255 7191
rect 18061 7157 18095 7191
rect 19533 7157 19567 7191
rect 21373 7157 21407 7191
rect 22661 7157 22695 7191
rect 4813 6953 4847 6987
rect 5089 6953 5123 6987
rect 6653 6953 6687 6987
rect 7113 6953 7147 6987
rect 7297 6953 7331 6987
rect 8953 6953 8987 6987
rect 21465 6885 21499 6919
rect 6469 6817 6503 6851
rect 8677 6817 8711 6851
rect 10149 6817 10183 6851
rect 11069 6817 11103 6851
rect 11253 6817 11287 6851
rect 11529 6817 11563 6851
rect 12817 6817 12851 6851
rect 13001 6817 13035 6851
rect 13645 6817 13679 6851
rect 13737 6817 13771 6851
rect 16129 6817 16163 6851
rect 17785 6817 17819 6851
rect 19073 6817 19107 6851
rect 20637 6817 20671 6851
rect 20913 6817 20947 6851
rect 22201 6817 22235 6851
rect 6202 6749 6236 6783
rect 10793 6749 10827 6783
rect 10885 6749 10919 6783
rect 12725 6749 12759 6783
rect 14381 6749 14415 6783
rect 14565 6749 14599 6783
rect 14657 6749 14691 6783
rect 17877 6749 17911 6783
rect 22477 6749 22511 6783
rect 22845 6749 22879 6783
rect 8432 6681 8466 6715
rect 9413 6681 9447 6715
rect 13553 6681 13587 6715
rect 14924 6681 14958 6715
rect 16396 6681 16430 6715
rect 17969 6681 18003 6715
rect 20392 6681 20426 6715
rect 21097 6681 21131 6715
rect 22109 6681 22143 6715
rect 9321 6613 9355 6647
rect 9597 6613 9631 6647
rect 9965 6613 9999 6647
rect 10057 6613 10091 6647
rect 10425 6613 10459 6647
rect 12357 6613 12391 6647
rect 13185 6613 13219 6647
rect 16037 6613 16071 6647
rect 17509 6613 17543 6647
rect 18337 6613 18371 6647
rect 18429 6613 18463 6647
rect 18705 6613 18739 6647
rect 19257 6613 19291 6647
rect 21005 6613 21039 6647
rect 21649 6613 21683 6647
rect 22017 6613 22051 6647
rect 22661 6613 22695 6647
rect 23029 6613 23063 6647
rect 4813 6409 4847 6443
rect 6469 6409 6503 6443
rect 7573 6409 7607 6443
rect 8493 6409 8527 6443
rect 9321 6409 9355 6443
rect 10057 6409 10091 6443
rect 10885 6409 10919 6443
rect 12357 6409 12391 6443
rect 12725 6409 12759 6443
rect 12817 6409 12851 6443
rect 13277 6409 13311 6443
rect 16037 6409 16071 6443
rect 16405 6409 16439 6443
rect 17417 6409 17451 6443
rect 17969 6409 18003 6443
rect 18797 6409 18831 6443
rect 20637 6409 20671 6443
rect 21005 6409 21039 6443
rect 21465 6409 21499 6443
rect 21833 6409 21867 6443
rect 5926 6341 5960 6375
rect 8585 6341 8619 6375
rect 11805 6341 11839 6375
rect 15209 6341 15243 6375
rect 17049 6341 17083 6375
rect 18889 6341 18923 6375
rect 19524 6341 19558 6375
rect 6193 6273 6227 6307
rect 7665 6273 7699 6307
rect 9229 6273 9263 6307
rect 10149 6273 10183 6307
rect 10977 6273 11011 6307
rect 11897 6273 11931 6307
rect 14013 6273 14047 6307
rect 14473 6273 14507 6307
rect 15301 6273 15335 6307
rect 15945 6273 15979 6307
rect 17877 6273 17911 6307
rect 21097 6273 21131 6307
rect 22201 6273 22235 6307
rect 22845 6273 22879 6307
rect 7389 6205 7423 6239
rect 8769 6205 8803 6239
rect 9045 6205 9079 6239
rect 9965 6205 9999 6239
rect 10793 6205 10827 6239
rect 11621 6205 11655 6239
rect 13001 6205 13035 6239
rect 13829 6205 13863 6239
rect 13921 6205 13955 6239
rect 15393 6205 15427 6239
rect 15761 6205 15795 6239
rect 16773 6205 16807 6239
rect 16957 6205 16991 6239
rect 18061 6205 18095 6239
rect 18981 6205 19015 6239
rect 19257 6205 19291 6239
rect 20821 6205 20855 6239
rect 22293 6205 22327 6239
rect 22385 6205 22419 6239
rect 8033 6137 8067 6171
rect 12265 6137 12299 6171
rect 14381 6137 14415 6171
rect 21557 6137 21591 6171
rect 22661 6137 22695 6171
rect 8125 6069 8159 6103
rect 9689 6069 9723 6103
rect 10517 6069 10551 6103
rect 11345 6069 11379 6103
rect 14841 6069 14875 6103
rect 17509 6069 17543 6103
rect 18429 6069 18463 6103
rect 23029 6069 23063 6103
rect 9873 5865 9907 5899
rect 10057 5865 10091 5899
rect 12081 5865 12115 5899
rect 13921 5865 13955 5899
rect 17693 5865 17727 5899
rect 20913 5865 20947 5899
rect 21741 5865 21775 5899
rect 22661 5865 22695 5899
rect 7941 5797 7975 5831
rect 8769 5797 8803 5831
rect 16773 5797 16807 5831
rect 22293 5797 22327 5831
rect 7389 5729 7423 5763
rect 8217 5729 8251 5763
rect 9413 5729 9447 5763
rect 9505 5729 9539 5763
rect 10609 5729 10643 5763
rect 10701 5729 10735 5763
rect 11345 5729 11379 5763
rect 12725 5729 12759 5763
rect 14568 5729 14602 5763
rect 16129 5729 16163 5763
rect 16313 5729 16347 5763
rect 16957 5729 16991 5763
rect 18245 5729 18279 5763
rect 18521 5729 18555 5763
rect 19809 5729 19843 5763
rect 20177 5729 20211 5763
rect 21465 5729 21499 5763
rect 7573 5661 7607 5695
rect 8401 5661 8435 5695
rect 9321 5661 9355 5695
rect 10793 5661 10827 5695
rect 11621 5661 11655 5695
rect 13737 5661 13771 5695
rect 14105 5661 14139 5695
rect 14841 5661 14875 5695
rect 16405 5661 16439 5695
rect 17233 5661 17267 5695
rect 21373 5661 21407 5695
rect 21925 5661 21959 5695
rect 22845 5661 22879 5695
rect 7481 5593 7515 5627
rect 12449 5593 12483 5627
rect 12541 5593 12575 5627
rect 18061 5593 18095 5627
rect 19073 5593 19107 5627
rect 19625 5593 19659 5627
rect 20361 5593 20395 5627
rect 21281 5593 21315 5627
rect 22017 5593 22051 5627
rect 22477 5593 22511 5627
rect 8309 5525 8343 5559
rect 8953 5525 8987 5559
rect 11161 5525 11195 5559
rect 11529 5525 11563 5559
rect 11989 5525 12023 5559
rect 13645 5525 13679 5559
rect 14571 5525 14605 5559
rect 15945 5525 15979 5559
rect 17141 5525 17175 5559
rect 17601 5525 17635 5559
rect 18153 5525 18187 5559
rect 19257 5525 19291 5559
rect 19717 5525 19751 5559
rect 20453 5525 20487 5559
rect 20821 5525 20855 5559
rect 23029 5525 23063 5559
rect 8217 5321 8251 5355
rect 8769 5321 8803 5355
rect 9137 5321 9171 5355
rect 9689 5321 9723 5355
rect 12265 5321 12299 5355
rect 12357 5321 12391 5355
rect 15025 5321 15059 5355
rect 15393 5321 15427 5355
rect 15669 5321 15703 5355
rect 17049 5321 17083 5355
rect 17417 5321 17451 5355
rect 17969 5321 18003 5355
rect 19165 5321 19199 5355
rect 20085 5321 20119 5355
rect 22201 5321 22235 5355
rect 22753 5321 22787 5355
rect 8309 5253 8343 5287
rect 14381 5253 14415 5287
rect 14565 5253 14599 5287
rect 17877 5253 17911 5287
rect 22293 5253 22327 5287
rect 9229 5185 9263 5219
rect 14841 5185 14875 5219
rect 15117 5185 15151 5219
rect 16037 5185 16071 5219
rect 16129 5185 16163 5219
rect 18797 5185 18831 5219
rect 19625 5185 19659 5219
rect 20453 5185 20487 5219
rect 21281 5185 21315 5219
rect 22845 5185 22879 5219
rect 8125 5117 8159 5151
rect 9321 5117 9355 5151
rect 12081 5117 12115 5151
rect 16221 5117 16255 5151
rect 16773 5117 16807 5151
rect 16957 5117 16991 5151
rect 18061 5117 18095 5151
rect 18613 5117 18647 5151
rect 18705 5117 18739 5151
rect 19441 5117 19475 5151
rect 19533 5117 19567 5151
rect 20545 5117 20579 5151
rect 20637 5117 20671 5151
rect 21005 5117 21039 5151
rect 21189 5117 21223 5151
rect 22385 5117 22419 5151
rect 8677 5049 8711 5083
rect 21649 5049 21683 5083
rect 12725 4981 12759 5015
rect 14657 4981 14691 5015
rect 15301 4981 15335 5015
rect 17509 4981 17543 5015
rect 19993 4981 20027 5015
rect 21833 4981 21867 5015
rect 23029 4981 23063 5015
rect 8769 4777 8803 4811
rect 18337 4777 18371 4811
rect 19993 4777 20027 4811
rect 20729 4777 20763 4811
rect 9045 4709 9079 4743
rect 19073 4709 19107 4743
rect 8125 4641 8159 4675
rect 8309 4641 8343 4675
rect 17046 4641 17080 4675
rect 17509 4641 17543 4675
rect 17785 4641 17819 4675
rect 18705 4641 18739 4675
rect 19441 4641 19475 4675
rect 20269 4641 20303 4675
rect 21284 4641 21318 4675
rect 21557 4641 21591 4675
rect 8401 4573 8435 4607
rect 11713 4573 11747 4607
rect 12265 4573 12299 4607
rect 15393 4573 15427 4607
rect 16773 4573 16807 4607
rect 17969 4573 18003 4607
rect 18889 4573 18923 4607
rect 19533 4573 19567 4607
rect 20545 4573 20579 4607
rect 20821 4573 20855 4607
rect 22845 4573 22879 4607
rect 12449 4505 12483 4539
rect 17877 4505 17911 4539
rect 15577 4437 15611 4471
rect 15669 4437 15703 4471
rect 17042 4437 17076 4471
rect 19625 4437 19659 4471
rect 20361 4437 20395 4471
rect 21287 4437 21321 4471
rect 22661 4437 22695 4471
rect 23029 4437 23063 4471
rect 15761 4233 15795 4267
rect 16129 4233 16163 4267
rect 19073 4233 19107 4267
rect 19809 4233 19843 4267
rect 21281 4233 21315 4267
rect 22017 4233 22051 4267
rect 22293 4233 22327 4267
rect 15669 4165 15703 4199
rect 20637 4165 20671 4199
rect 18613 4097 18647 4131
rect 18889 4097 18923 4131
rect 19165 4097 19199 4131
rect 21373 4097 21407 4131
rect 21925 4097 21959 4131
rect 22477 4097 22511 4131
rect 22753 4097 22787 4131
rect 22845 4097 22879 4131
rect 15577 4029 15611 4063
rect 17785 4029 17819 4063
rect 18058 4029 18092 4063
rect 18198 4029 18232 4063
rect 18521 4029 18555 4063
rect 19625 4029 19659 4063
rect 19717 4029 19751 4063
rect 20729 4029 20763 4063
rect 20913 4029 20947 4063
rect 18797 3961 18831 3995
rect 21557 3961 21591 3995
rect 22569 3961 22603 3995
rect 16681 3893 16715 3927
rect 19349 3893 19383 3927
rect 20177 3893 20211 3927
rect 20269 3893 20303 3927
rect 23029 3893 23063 3927
rect 18061 3689 18095 3723
rect 19441 3689 19475 3723
rect 19625 3689 19659 3723
rect 17969 3621 18003 3655
rect 19073 3621 19107 3655
rect 19993 3621 20027 3655
rect 21005 3621 21039 3655
rect 22569 3621 22603 3655
rect 16865 3553 16899 3587
rect 17138 3553 17172 3587
rect 20453 3553 20487 3587
rect 20545 3553 20579 3587
rect 21833 3553 21867 3587
rect 22201 3553 22235 3587
rect 1593 3485 1627 3519
rect 17601 3485 17635 3519
rect 17785 3485 17819 3519
rect 18245 3485 18279 3519
rect 18797 3485 18831 3519
rect 18889 3485 18923 3519
rect 19257 3485 19291 3519
rect 19717 3485 19751 3519
rect 20821 3485 20855 3519
rect 21557 3485 21591 3519
rect 22293 3485 22327 3519
rect 22753 3485 22787 3519
rect 22845 3485 22879 3519
rect 20361 3417 20395 3451
rect 1409 3349 1443 3383
rect 15761 3349 15795 3383
rect 17134 3349 17168 3383
rect 18613 3349 18647 3383
rect 19901 3349 19935 3383
rect 21649 3349 21683 3383
rect 22477 3349 22511 3383
rect 23029 3349 23063 3383
rect 19986 3145 20020 3179
rect 22017 3145 22051 3179
rect 16221 3077 16255 3111
rect 8585 3009 8619 3043
rect 16497 3009 16531 3043
rect 19717 3009 19751 3043
rect 22109 3009 22143 3043
rect 22845 3009 22879 3043
rect 16681 2941 16715 2975
rect 17004 2941 17038 2975
rect 17144 2941 17178 2975
rect 17417 2941 17451 2975
rect 19990 2959 20024 2993
rect 20453 2941 20487 2975
rect 22385 2941 22419 2975
rect 22753 2941 22787 2975
rect 8401 2805 8435 2839
rect 8769 2805 8803 2839
rect 18521 2805 18555 2839
rect 18613 2805 18647 2839
rect 23029 2805 23063 2839
rect 10793 2601 10827 2635
rect 16773 2601 16807 2635
rect 22845 2601 22879 2635
rect 2513 2397 2547 2431
rect 6377 2397 6411 2431
rect 10609 2397 10643 2431
rect 22661 2397 22695 2431
rect 2329 2261 2363 2295
rect 10425 2261 10459 2295
rect 22477 2261 22511 2295
<< metal1 >>
rect 11974 22788 11980 22840
rect 12032 22828 12038 22840
rect 19058 22828 19064 22840
rect 12032 22800 19064 22828
rect 12032 22788 12038 22800
rect 19058 22788 19064 22800
rect 19116 22788 19122 22840
rect 9030 22720 9036 22772
rect 9088 22760 9094 22772
rect 20162 22760 20168 22772
rect 9088 22732 20168 22760
rect 9088 22720 9094 22732
rect 20162 22720 20168 22732
rect 20220 22720 20226 22772
rect 7466 22652 7472 22704
rect 7524 22692 7530 22704
rect 19702 22692 19708 22704
rect 7524 22664 19708 22692
rect 7524 22652 7530 22664
rect 19702 22652 19708 22664
rect 19760 22652 19766 22704
rect 5166 22584 5172 22636
rect 5224 22624 5230 22636
rect 19334 22624 19340 22636
rect 5224 22596 19340 22624
rect 5224 22584 5230 22596
rect 19334 22584 19340 22596
rect 19392 22584 19398 22636
rect 14550 22516 14556 22568
rect 14608 22556 14614 22568
rect 16298 22556 16304 22568
rect 14608 22528 16304 22556
rect 14608 22516 14614 22528
rect 16298 22516 16304 22528
rect 16356 22516 16362 22568
rect 14090 22448 14096 22500
rect 14148 22488 14154 22500
rect 20990 22488 20996 22500
rect 14148 22460 20996 22488
rect 14148 22448 14154 22460
rect 20990 22448 20996 22460
rect 21048 22448 21054 22500
rect 13814 22380 13820 22432
rect 13872 22420 13878 22432
rect 15562 22420 15568 22432
rect 13872 22392 15568 22420
rect 13872 22380 13878 22392
rect 15562 22380 15568 22392
rect 15620 22380 15626 22432
rect 1104 22330 23460 22352
rect 1104 22278 3749 22330
rect 3801 22278 3813 22330
rect 3865 22278 3877 22330
rect 3929 22278 3941 22330
rect 3993 22278 4005 22330
rect 4057 22278 9347 22330
rect 9399 22278 9411 22330
rect 9463 22278 9475 22330
rect 9527 22278 9539 22330
rect 9591 22278 9603 22330
rect 9655 22278 14945 22330
rect 14997 22278 15009 22330
rect 15061 22278 15073 22330
rect 15125 22278 15137 22330
rect 15189 22278 15201 22330
rect 15253 22278 20543 22330
rect 20595 22278 20607 22330
rect 20659 22278 20671 22330
rect 20723 22278 20735 22330
rect 20787 22278 20799 22330
rect 20851 22278 23460 22330
rect 1104 22256 23460 22278
rect 5718 22176 5724 22228
rect 5776 22216 5782 22228
rect 8297 22219 8355 22225
rect 8297 22216 8309 22219
rect 5776 22188 8309 22216
rect 5776 22176 5782 22188
rect 8297 22185 8309 22188
rect 8343 22185 8355 22219
rect 14277 22219 14335 22225
rect 14277 22216 14289 22219
rect 8297 22179 8355 22185
rect 12820 22188 14289 22216
rect 6656 22120 7604 22148
rect 5442 22080 5448 22092
rect 5403 22052 5448 22080
rect 5442 22040 5448 22052
rect 5500 22080 5506 22092
rect 5997 22083 6055 22089
rect 5500 22052 5764 22080
rect 5500 22040 5506 22052
rect 1949 22015 2007 22021
rect 1949 21981 1961 22015
rect 1995 22012 2007 22015
rect 2406 22012 2412 22024
rect 1995 21984 2412 22012
rect 1995 21981 2007 21984
rect 1949 21975 2007 21981
rect 2406 21972 2412 21984
rect 2464 21972 2470 22024
rect 2593 22015 2651 22021
rect 2593 21981 2605 22015
rect 2639 22012 2651 22015
rect 2958 22012 2964 22024
rect 2639 21984 2964 22012
rect 2639 21981 2651 21984
rect 2593 21975 2651 21981
rect 2958 21972 2964 21984
rect 3016 21972 3022 22024
rect 3234 22012 3240 22024
rect 3195 21984 3240 22012
rect 3234 21972 3240 21984
rect 3292 21972 3298 22024
rect 4065 22015 4123 22021
rect 4065 21981 4077 22015
rect 4111 22012 4123 22015
rect 4154 22012 4160 22024
rect 4111 21984 4160 22012
rect 4111 21981 4123 21984
rect 4065 21975 4123 21981
rect 4154 21972 4160 21984
rect 4212 21972 4218 22024
rect 4249 22015 4307 22021
rect 4249 21981 4261 22015
rect 4295 21981 4307 22015
rect 4249 21975 4307 21981
rect 4801 22015 4859 22021
rect 4801 21981 4813 22015
rect 4847 21981 4859 22015
rect 4801 21975 4859 21981
rect 3694 21904 3700 21956
rect 3752 21944 3758 21956
rect 4264 21944 4292 21975
rect 3752 21916 4292 21944
rect 4816 21944 4844 21975
rect 4982 21972 4988 22024
rect 5040 22012 5046 22024
rect 5736 22021 5764 22052
rect 5997 22049 6009 22083
rect 6043 22080 6055 22083
rect 6086 22080 6092 22092
rect 6043 22052 6092 22080
rect 6043 22049 6055 22052
rect 5997 22043 6055 22049
rect 6086 22040 6092 22052
rect 6144 22040 6150 22092
rect 6181 22083 6239 22089
rect 6181 22049 6193 22083
rect 6227 22080 6239 22083
rect 6454 22080 6460 22092
rect 6227 22052 6460 22080
rect 6227 22049 6239 22052
rect 6181 22043 6239 22049
rect 6454 22040 6460 22052
rect 6512 22040 6518 22092
rect 5169 22015 5227 22021
rect 5169 22012 5181 22015
rect 5040 21984 5181 22012
rect 5040 21972 5046 21984
rect 5169 21981 5181 21984
rect 5215 21981 5227 22015
rect 5169 21975 5227 21981
rect 5721 22015 5779 22021
rect 5721 21981 5733 22015
rect 5767 21981 5779 22015
rect 6104 22012 6132 22040
rect 6549 22015 6607 22021
rect 6549 22012 6561 22015
rect 6104 21984 6561 22012
rect 5721 21975 5779 21981
rect 6549 21981 6561 21984
rect 6595 21981 6607 22015
rect 6549 21975 6607 21981
rect 6656 21944 6684 22120
rect 6733 22083 6791 22089
rect 6733 22049 6745 22083
rect 6779 22080 6791 22083
rect 7374 22080 7380 22092
rect 6779 22052 7380 22080
rect 6779 22049 6791 22052
rect 6733 22043 6791 22049
rect 7374 22040 7380 22052
rect 7432 22080 7438 22092
rect 7576 22080 7604 22120
rect 7650 22108 7656 22160
rect 7708 22148 7714 22160
rect 7708 22120 9076 22148
rect 7708 22108 7714 22120
rect 8205 22083 8263 22089
rect 7432 22052 7512 22080
rect 7576 22052 8156 22080
rect 7432 22040 7438 22052
rect 6822 21972 6828 22024
rect 6880 22012 6886 22024
rect 7484 22021 7512 22052
rect 7009 22015 7067 22021
rect 7009 22012 7021 22015
rect 6880 21984 7021 22012
rect 6880 21972 6886 21984
rect 7009 21981 7021 21984
rect 7055 21981 7067 22015
rect 7009 21975 7067 21981
rect 7469 22015 7527 22021
rect 7469 21981 7481 22015
rect 7515 21981 7527 22015
rect 7745 22015 7803 22021
rect 7745 22012 7757 22015
rect 7469 21975 7527 21981
rect 7576 21984 7757 22012
rect 4816 21916 6684 21944
rect 7193 21947 7251 21953
rect 3752 21904 3758 21916
rect 7193 21913 7205 21947
rect 7239 21944 7251 21947
rect 7576 21944 7604 21984
rect 7745 21981 7757 21984
rect 7791 22012 7803 22015
rect 8018 22012 8024 22024
rect 7791 21984 8024 22012
rect 7791 21981 7803 21984
rect 7745 21975 7803 21981
rect 8018 21972 8024 21984
rect 8076 21972 8082 22024
rect 7239 21916 7604 21944
rect 8128 21944 8156 22052
rect 8205 22049 8217 22083
rect 8251 22080 8263 22083
rect 9048 22080 9076 22120
rect 9122 22108 9128 22160
rect 9180 22148 9186 22160
rect 10597 22151 10655 22157
rect 10597 22148 10609 22151
rect 9180 22120 9720 22148
rect 9180 22108 9186 22120
rect 9692 22094 9720 22120
rect 10428 22120 10609 22148
rect 9692 22089 9757 22094
rect 9677 22083 9757 22089
rect 8251 22052 8800 22080
rect 9048 22052 9352 22080
rect 8251 22049 8263 22052
rect 8205 22043 8263 22049
rect 8478 22012 8484 22024
rect 8439 21984 8484 22012
rect 8478 21972 8484 21984
rect 8536 21972 8542 22024
rect 8772 22021 8800 22052
rect 8757 22015 8815 22021
rect 8757 21981 8769 22015
rect 8803 22012 8815 22015
rect 9214 22012 9220 22024
rect 8803 21984 9220 22012
rect 8803 21981 8815 21984
rect 8757 21975 8815 21981
rect 9214 21972 9220 21984
rect 9272 21972 9278 22024
rect 9324 22012 9352 22052
rect 9677 22049 9689 22083
rect 9723 22066 9757 22083
rect 10428 22080 10456 22120
rect 10597 22117 10609 22120
rect 10643 22117 10655 22151
rect 10597 22111 10655 22117
rect 9723 22049 9735 22066
rect 9677 22043 9735 22049
rect 9876 22052 10456 22080
rect 10505 22083 10563 22089
rect 9876 22012 9904 22052
rect 10505 22049 10517 22083
rect 10551 22080 10563 22083
rect 11882 22080 11888 22092
rect 10551 22052 11888 22080
rect 10551 22049 10563 22052
rect 10505 22043 10563 22049
rect 9324 21984 9904 22012
rect 9950 21972 9956 22024
rect 10008 22012 10014 22024
rect 10226 22012 10232 22024
rect 10008 21984 10232 22012
rect 10008 21972 10014 21984
rect 10226 21972 10232 21984
rect 10284 21972 10290 22024
rect 10781 22015 10839 22021
rect 10781 21981 10793 22015
rect 10827 21981 10839 22015
rect 11054 22012 11060 22024
rect 11015 21984 11060 22012
rect 10781 21975 10839 21981
rect 9033 21947 9091 21953
rect 8128 21916 8616 21944
rect 7239 21913 7251 21916
rect 7193 21907 7251 21913
rect 1578 21836 1584 21888
rect 1636 21876 1642 21888
rect 1765 21879 1823 21885
rect 1765 21876 1777 21879
rect 1636 21848 1777 21876
rect 1636 21836 1642 21848
rect 1765 21845 1777 21848
rect 1811 21845 1823 21879
rect 1765 21839 1823 21845
rect 2222 21836 2228 21888
rect 2280 21876 2286 21888
rect 2409 21879 2467 21885
rect 2409 21876 2421 21879
rect 2280 21848 2421 21876
rect 2280 21836 2286 21848
rect 2409 21845 2421 21848
rect 2455 21845 2467 21879
rect 2409 21839 2467 21845
rect 2866 21836 2872 21888
rect 2924 21876 2930 21888
rect 3053 21879 3111 21885
rect 3053 21876 3065 21879
rect 2924 21848 3065 21876
rect 2924 21836 2930 21848
rect 3053 21845 3065 21848
rect 3099 21845 3111 21879
rect 3053 21839 3111 21845
rect 3510 21836 3516 21888
rect 3568 21876 3574 21888
rect 3881 21879 3939 21885
rect 3881 21876 3893 21879
rect 3568 21848 3893 21876
rect 3568 21836 3574 21848
rect 3881 21845 3893 21848
rect 3927 21845 3939 21879
rect 3881 21839 3939 21845
rect 4246 21836 4252 21888
rect 4304 21876 4310 21888
rect 4433 21879 4491 21885
rect 4433 21876 4445 21879
rect 4304 21848 4445 21876
rect 4304 21836 4310 21848
rect 4433 21845 4445 21848
rect 4479 21845 4491 21879
rect 4614 21876 4620 21888
rect 4575 21848 4620 21876
rect 4433 21839 4491 21845
rect 4614 21836 4620 21848
rect 4672 21836 4678 21888
rect 4798 21836 4804 21888
rect 4856 21876 4862 21888
rect 4985 21879 5043 21885
rect 4985 21876 4997 21879
rect 4856 21848 4997 21876
rect 4856 21836 4862 21848
rect 4985 21845 4997 21848
rect 5031 21845 5043 21879
rect 4985 21839 5043 21845
rect 5537 21879 5595 21885
rect 5537 21845 5549 21879
rect 5583 21876 5595 21879
rect 5810 21876 5816 21888
rect 5583 21848 5816 21876
rect 5583 21845 5595 21848
rect 5537 21839 5595 21845
rect 5810 21836 5816 21848
rect 5868 21836 5874 21888
rect 6362 21876 6368 21888
rect 6323 21848 6368 21876
rect 6362 21836 6368 21848
rect 6420 21836 6426 21888
rect 6454 21836 6460 21888
rect 6512 21876 6518 21888
rect 6825 21879 6883 21885
rect 6825 21876 6837 21879
rect 6512 21848 6837 21876
rect 6512 21836 6518 21848
rect 6825 21845 6837 21848
rect 6871 21845 6883 21879
rect 6825 21839 6883 21845
rect 6914 21836 6920 21888
rect 6972 21876 6978 21888
rect 7285 21879 7343 21885
rect 7285 21876 7297 21879
rect 6972 21848 7297 21876
rect 6972 21836 6978 21848
rect 7285 21845 7297 21848
rect 7331 21845 7343 21879
rect 7558 21876 7564 21888
rect 7519 21848 7564 21876
rect 7285 21839 7343 21845
rect 7558 21836 7564 21848
rect 7616 21836 7622 21888
rect 7834 21876 7840 21888
rect 7795 21848 7840 21876
rect 7834 21836 7840 21848
rect 7892 21836 7898 21888
rect 8588 21885 8616 21916
rect 9033 21913 9045 21947
rect 9079 21944 9091 21947
rect 10594 21944 10600 21956
rect 9079 21916 10600 21944
rect 9079 21913 9091 21916
rect 9033 21907 9091 21913
rect 10594 21904 10600 21916
rect 10652 21944 10658 21956
rect 10796 21944 10824 21975
rect 11054 21972 11060 21984
rect 11112 21972 11118 22024
rect 11348 22021 11376 22052
rect 11882 22040 11888 22052
rect 11940 22040 11946 22092
rect 12434 22080 12440 22092
rect 12084 22052 12440 22080
rect 11333 22015 11391 22021
rect 11333 21981 11345 22015
rect 11379 21981 11391 22015
rect 11514 22012 11520 22024
rect 11475 21984 11520 22012
rect 11333 21975 11391 21981
rect 11514 21972 11520 21984
rect 11572 21972 11578 22024
rect 12084 22021 12112 22052
rect 12434 22040 12440 22052
rect 12492 22080 12498 22092
rect 12710 22080 12716 22092
rect 12492 22052 12585 22080
rect 12671 22052 12716 22080
rect 12492 22040 12498 22052
rect 12710 22040 12716 22052
rect 12768 22080 12774 22092
rect 12820 22080 12848 22188
rect 14277 22185 14289 22188
rect 14323 22185 14335 22219
rect 14277 22179 14335 22185
rect 14458 22176 14464 22228
rect 14516 22216 14522 22228
rect 16022 22216 16028 22228
rect 14516 22188 16028 22216
rect 14516 22176 14522 22188
rect 16022 22176 16028 22188
rect 16080 22176 16086 22228
rect 16298 22176 16304 22228
rect 16356 22216 16362 22228
rect 22554 22216 22560 22228
rect 16356 22188 22560 22216
rect 16356 22176 16362 22188
rect 22554 22176 22560 22188
rect 22612 22176 22618 22228
rect 13630 22148 13636 22160
rect 13591 22120 13636 22148
rect 13630 22108 13636 22120
rect 13688 22108 13694 22160
rect 14826 22108 14832 22160
rect 14884 22148 14890 22160
rect 16114 22148 16120 22160
rect 14884 22120 16120 22148
rect 14884 22108 14890 22120
rect 16114 22108 16120 22120
rect 16172 22108 16178 22160
rect 16482 22108 16488 22160
rect 16540 22148 16546 22160
rect 16540 22120 16712 22148
rect 16540 22108 16546 22120
rect 12768 22052 12848 22080
rect 13096 22052 16620 22080
rect 12768 22040 12774 22052
rect 12069 22015 12127 22021
rect 12069 21981 12081 22015
rect 12115 21981 12127 22015
rect 12069 21975 12127 21981
rect 12161 22015 12219 22021
rect 12161 21981 12173 22015
rect 12207 22012 12219 22015
rect 12526 22012 12532 22024
rect 12207 21984 12532 22012
rect 12207 21981 12219 21984
rect 12161 21975 12219 21981
rect 12526 21972 12532 21984
rect 12584 21972 12590 22024
rect 10652 21916 10824 21944
rect 13096 21944 13124 22052
rect 13170 21972 13176 22024
rect 13228 22012 13234 22024
rect 13449 22015 13507 22021
rect 13449 22012 13461 22015
rect 13228 21984 13461 22012
rect 13228 21972 13234 21984
rect 13449 21981 13461 21984
rect 13495 21981 13507 22015
rect 13449 21975 13507 21981
rect 13464 21944 13492 21975
rect 13630 21972 13636 22024
rect 13688 22012 13694 22024
rect 13725 22015 13783 22021
rect 13725 22012 13737 22015
rect 13688 21984 13737 22012
rect 13688 21972 13694 21984
rect 13725 21981 13737 21984
rect 13771 21981 13783 22015
rect 13725 21975 13783 21981
rect 14461 22015 14519 22021
rect 14461 21981 14473 22015
rect 14507 22012 14519 22015
rect 14507 21984 15424 22012
rect 14507 21981 14519 21984
rect 14461 21975 14519 21981
rect 14093 21947 14151 21953
rect 14093 21944 14105 21947
rect 13096 21916 13400 21944
rect 13464 21916 14105 21944
rect 10652 21904 10658 21916
rect 8573 21879 8631 21885
rect 8573 21845 8585 21879
rect 8619 21845 8631 21879
rect 8573 21839 8631 21845
rect 9125 21879 9183 21885
rect 9125 21845 9137 21879
rect 9171 21876 9183 21879
rect 9214 21876 9220 21888
rect 9171 21848 9220 21876
rect 9171 21845 9183 21848
rect 9125 21839 9183 21845
rect 9214 21836 9220 21848
rect 9272 21836 9278 21888
rect 9490 21876 9496 21888
rect 9451 21848 9496 21876
rect 9490 21836 9496 21848
rect 9548 21836 9554 21888
rect 9585 21879 9643 21885
rect 9585 21845 9597 21879
rect 9631 21876 9643 21879
rect 9766 21876 9772 21888
rect 9631 21848 9772 21876
rect 9631 21845 9643 21848
rect 9585 21839 9643 21845
rect 9766 21836 9772 21848
rect 9824 21836 9830 21888
rect 10042 21876 10048 21888
rect 10003 21848 10048 21876
rect 10042 21836 10048 21848
rect 10100 21836 10106 21888
rect 10870 21876 10876 21888
rect 10831 21848 10876 21876
rect 10870 21836 10876 21848
rect 10928 21836 10934 21888
rect 11146 21876 11152 21888
rect 11107 21848 11152 21876
rect 11146 21836 11152 21848
rect 11204 21836 11210 21888
rect 11698 21876 11704 21888
rect 11659 21848 11704 21876
rect 11698 21836 11704 21848
rect 11756 21836 11762 21888
rect 11882 21876 11888 21888
rect 11843 21848 11888 21876
rect 11882 21836 11888 21848
rect 11940 21836 11946 21888
rect 12066 21836 12072 21888
rect 12124 21876 12130 21888
rect 12345 21879 12403 21885
rect 12345 21876 12357 21879
rect 12124 21848 12357 21876
rect 12124 21836 12130 21848
rect 12345 21845 12357 21848
rect 12391 21845 12403 21879
rect 12894 21876 12900 21888
rect 12855 21848 12900 21876
rect 12345 21839 12403 21845
rect 12894 21836 12900 21848
rect 12952 21836 12958 21888
rect 12986 21836 12992 21888
rect 13044 21876 13050 21888
rect 13372 21885 13400 21916
rect 14093 21913 14105 21916
rect 14139 21913 14151 21947
rect 14093 21907 14151 21913
rect 14366 21904 14372 21956
rect 14424 21944 14430 21956
rect 14645 21947 14703 21953
rect 14645 21944 14657 21947
rect 14424 21916 14657 21944
rect 14424 21904 14430 21916
rect 14645 21913 14657 21916
rect 14691 21944 14703 21947
rect 14921 21947 14979 21953
rect 14921 21944 14933 21947
rect 14691 21916 14933 21944
rect 14691 21913 14703 21916
rect 14645 21907 14703 21913
rect 14921 21913 14933 21916
rect 14967 21913 14979 21947
rect 14921 21907 14979 21913
rect 15010 21904 15016 21956
rect 15068 21944 15074 21956
rect 15105 21947 15163 21953
rect 15105 21944 15117 21947
rect 15068 21916 15117 21944
rect 15068 21904 15074 21916
rect 15105 21913 15117 21916
rect 15151 21913 15163 21947
rect 15396 21944 15424 21984
rect 15470 21972 15476 22024
rect 15528 22012 15534 22024
rect 15746 22012 15752 22024
rect 15528 21984 15573 22012
rect 15707 21984 15752 22012
rect 15528 21972 15534 21984
rect 15746 21972 15752 21984
rect 15804 21972 15810 22024
rect 16022 22012 16028 22024
rect 15983 21984 16028 22012
rect 16022 21972 16028 21984
rect 16080 21972 16086 22024
rect 16114 21972 16120 22024
rect 16172 22012 16178 22024
rect 16301 22015 16359 22021
rect 16301 22012 16313 22015
rect 16172 21984 16313 22012
rect 16172 21972 16178 21984
rect 16301 21981 16313 21984
rect 16347 21981 16359 22015
rect 16301 21975 16359 21981
rect 15396 21916 15884 21944
rect 15105 21907 15163 21913
rect 13357 21879 13415 21885
rect 13044 21848 13089 21876
rect 13044 21836 13050 21848
rect 13357 21845 13369 21879
rect 13403 21845 13415 21879
rect 13357 21839 13415 21845
rect 13814 21836 13820 21888
rect 13872 21876 13878 21888
rect 13909 21879 13967 21885
rect 13909 21876 13921 21879
rect 13872 21848 13921 21876
rect 13872 21836 13878 21848
rect 13909 21845 13921 21848
rect 13955 21845 13967 21879
rect 14734 21876 14740 21888
rect 14695 21848 14740 21876
rect 13909 21839 13967 21845
rect 14734 21836 14740 21848
rect 14792 21836 14798 21888
rect 15194 21836 15200 21888
rect 15252 21876 15258 21888
rect 15289 21879 15347 21885
rect 15289 21876 15301 21879
rect 15252 21848 15301 21876
rect 15252 21836 15258 21848
rect 15289 21845 15301 21848
rect 15335 21845 15347 21879
rect 15289 21839 15347 21845
rect 15378 21836 15384 21888
rect 15436 21876 15442 21888
rect 15856 21885 15884 21916
rect 15930 21904 15936 21956
rect 15988 21944 15994 21956
rect 16592 21944 16620 22052
rect 16684 22012 16712 22120
rect 17310 22108 17316 22160
rect 17368 22148 17374 22160
rect 17368 22120 17724 22148
rect 17368 22108 17374 22120
rect 16942 22080 16948 22092
rect 16903 22052 16948 22080
rect 16942 22040 16948 22052
rect 17000 22040 17006 22092
rect 17696 22089 17724 22120
rect 19150 22108 19156 22160
rect 19208 22148 19214 22160
rect 19208 22120 20668 22148
rect 19208 22108 19214 22120
rect 20640 22089 20668 22120
rect 17681 22083 17739 22089
rect 17681 22049 17693 22083
rect 17727 22080 17739 22083
rect 20625 22083 20683 22089
rect 17727 22052 17761 22080
rect 17880 22052 19012 22080
rect 17727 22049 17739 22052
rect 17681 22043 17739 22049
rect 17880 22012 17908 22052
rect 16684 21984 17908 22012
rect 17954 21972 17960 22024
rect 18012 22012 18018 22024
rect 18693 22015 18751 22021
rect 18012 21984 18552 22012
rect 18012 21972 18018 21984
rect 17037 21947 17095 21953
rect 17037 21944 17049 21947
rect 15988 21916 16528 21944
rect 16592 21916 17049 21944
rect 15988 21904 15994 21916
rect 15565 21879 15623 21885
rect 15565 21876 15577 21879
rect 15436 21848 15577 21876
rect 15436 21836 15442 21848
rect 15565 21845 15577 21848
rect 15611 21845 15623 21879
rect 15565 21839 15623 21845
rect 15841 21879 15899 21885
rect 15841 21845 15853 21879
rect 15887 21845 15899 21879
rect 16114 21876 16120 21888
rect 16075 21848 16120 21876
rect 15841 21839 15899 21845
rect 16114 21836 16120 21848
rect 16172 21836 16178 21888
rect 16298 21836 16304 21888
rect 16356 21876 16362 21888
rect 16393 21879 16451 21885
rect 16393 21876 16405 21879
rect 16356 21848 16405 21876
rect 16356 21836 16362 21848
rect 16393 21845 16405 21848
rect 16439 21845 16451 21879
rect 16500 21876 16528 21916
rect 17037 21913 17049 21916
rect 17083 21944 17095 21947
rect 17586 21944 17592 21956
rect 17083 21916 17592 21944
rect 17083 21913 17095 21916
rect 17037 21907 17095 21913
rect 17586 21904 17592 21916
rect 17644 21904 17650 21956
rect 17865 21947 17923 21953
rect 17865 21913 17877 21947
rect 17911 21944 17923 21947
rect 18138 21944 18144 21956
rect 17911 21916 18144 21944
rect 17911 21913 17923 21916
rect 17865 21907 17923 21913
rect 18138 21904 18144 21916
rect 18196 21904 18202 21956
rect 17126 21876 17132 21888
rect 16500 21848 17132 21876
rect 16393 21839 16451 21845
rect 17126 21836 17132 21848
rect 17184 21836 17190 21888
rect 17494 21876 17500 21888
rect 17455 21848 17500 21876
rect 17494 21836 17500 21848
rect 17552 21836 17558 21888
rect 17957 21879 18015 21885
rect 17957 21845 17969 21879
rect 18003 21876 18015 21879
rect 18230 21876 18236 21888
rect 18003 21848 18236 21876
rect 18003 21845 18015 21848
rect 17957 21839 18015 21845
rect 18230 21836 18236 21848
rect 18288 21836 18294 21888
rect 18322 21836 18328 21888
rect 18380 21876 18386 21888
rect 18524 21885 18552 21984
rect 18693 21981 18705 22015
rect 18739 22012 18751 22015
rect 18874 22012 18880 22024
rect 18739 21984 18880 22012
rect 18739 21981 18751 21984
rect 18693 21975 18751 21981
rect 18874 21972 18880 21984
rect 18932 21972 18938 22024
rect 18984 22021 19012 22052
rect 20625 22049 20637 22083
rect 20671 22080 20683 22083
rect 24118 22080 24124 22092
rect 20671 22052 20705 22080
rect 20824 22052 24124 22080
rect 20671 22049 20683 22052
rect 20625 22043 20683 22049
rect 18969 22015 19027 22021
rect 18969 21981 18981 22015
rect 19015 21981 19027 22015
rect 19334 22012 19340 22024
rect 19295 21984 19340 22012
rect 18969 21975 19027 21981
rect 19334 21972 19340 21984
rect 19392 21972 19398 22024
rect 19702 22012 19708 22024
rect 19663 21984 19708 22012
rect 19702 21972 19708 21984
rect 19760 21972 19766 22024
rect 20162 22012 20168 22024
rect 20123 21984 20168 22012
rect 20162 21972 20168 21984
rect 20220 21972 20226 22024
rect 20824 21944 20852 22052
rect 24118 22040 24124 22052
rect 24176 22040 24182 22092
rect 20901 22015 20959 22021
rect 20901 21981 20913 22015
rect 20947 22012 20959 22015
rect 20990 22012 20996 22024
rect 20947 21984 20996 22012
rect 20947 21981 20959 21984
rect 20901 21975 20959 21981
rect 20990 21972 20996 21984
rect 21048 21972 21054 22024
rect 21082 21972 21088 22024
rect 21140 22012 21146 22024
rect 21361 22015 21419 22021
rect 21361 22012 21373 22015
rect 21140 21984 21373 22012
rect 21140 21972 21146 21984
rect 21361 21981 21373 21984
rect 21407 21981 21419 22015
rect 21361 21975 21419 21981
rect 21450 21972 21456 22024
rect 21508 22012 21514 22024
rect 21818 22012 21824 22024
rect 21508 21984 21680 22012
rect 21779 21984 21824 22012
rect 21508 21972 21514 21984
rect 21652 21944 21680 21984
rect 21818 21972 21824 21984
rect 21876 21972 21882 22024
rect 22281 22015 22339 22021
rect 22281 22012 22293 22015
rect 22066 21984 22293 22012
rect 22066 21944 22094 21984
rect 22281 21981 22293 21984
rect 22327 21981 22339 22015
rect 22281 21975 22339 21981
rect 22462 21972 22468 22024
rect 22520 22012 22526 22024
rect 22833 22015 22891 22021
rect 22833 22012 22845 22015
rect 22520 21984 22845 22012
rect 22520 21972 22526 21984
rect 22833 21981 22845 21984
rect 22879 21981 22891 22015
rect 22833 21975 22891 21981
rect 19536 21916 20852 21944
rect 20916 21916 21588 21944
rect 21652 21916 22094 21944
rect 22741 21947 22799 21953
rect 18509 21879 18567 21885
rect 18380 21848 18425 21876
rect 18380 21836 18386 21848
rect 18509 21845 18521 21879
rect 18555 21845 18567 21879
rect 18509 21839 18567 21845
rect 18690 21836 18696 21888
rect 18748 21876 18754 21888
rect 19536 21885 19564 21916
rect 20916 21888 20944 21916
rect 18785 21879 18843 21885
rect 18785 21876 18797 21879
rect 18748 21848 18797 21876
rect 18748 21836 18754 21848
rect 18785 21845 18797 21848
rect 18831 21845 18843 21879
rect 18785 21839 18843 21845
rect 19521 21879 19579 21885
rect 19521 21845 19533 21879
rect 19567 21845 19579 21879
rect 19521 21839 19579 21845
rect 19610 21836 19616 21888
rect 19668 21876 19674 21888
rect 19889 21879 19947 21885
rect 19889 21876 19901 21879
rect 19668 21848 19901 21876
rect 19668 21836 19674 21848
rect 19889 21845 19901 21848
rect 19935 21845 19947 21879
rect 19889 21839 19947 21845
rect 20254 21836 20260 21888
rect 20312 21876 20318 21888
rect 20349 21879 20407 21885
rect 20349 21876 20361 21879
rect 20312 21848 20361 21876
rect 20312 21836 20318 21848
rect 20349 21845 20361 21848
rect 20395 21845 20407 21879
rect 20806 21876 20812 21888
rect 20767 21848 20812 21876
rect 20349 21839 20407 21845
rect 20806 21836 20812 21848
rect 20864 21836 20870 21888
rect 20898 21836 20904 21888
rect 20956 21836 20962 21888
rect 21266 21876 21272 21888
rect 21227 21848 21272 21876
rect 21266 21836 21272 21848
rect 21324 21836 21330 21888
rect 21560 21885 21588 21916
rect 22741 21913 22753 21947
rect 22787 21944 22799 21947
rect 23198 21944 23204 21956
rect 22787 21916 23204 21944
rect 22787 21913 22799 21916
rect 22741 21907 22799 21913
rect 23198 21904 23204 21916
rect 23256 21904 23262 21956
rect 21545 21879 21603 21885
rect 21545 21845 21557 21879
rect 21591 21845 21603 21879
rect 21545 21839 21603 21845
rect 21634 21836 21640 21888
rect 21692 21876 21698 21888
rect 22005 21879 22063 21885
rect 22005 21876 22017 21879
rect 21692 21848 22017 21876
rect 21692 21836 21698 21848
rect 22005 21845 22017 21848
rect 22051 21845 22063 21879
rect 22005 21839 22063 21845
rect 22186 21836 22192 21888
rect 22244 21876 22250 21888
rect 22465 21879 22523 21885
rect 22465 21876 22477 21879
rect 22244 21848 22477 21876
rect 22244 21836 22250 21848
rect 22465 21845 22477 21848
rect 22511 21845 22523 21879
rect 22465 21839 22523 21845
rect 22830 21836 22836 21888
rect 22888 21876 22894 21888
rect 23017 21879 23075 21885
rect 23017 21876 23029 21879
rect 22888 21848 23029 21876
rect 22888 21836 22894 21848
rect 23017 21845 23029 21848
rect 23063 21845 23075 21879
rect 23017 21839 23075 21845
rect 1104 21786 23460 21808
rect 1104 21734 6548 21786
rect 6600 21734 6612 21786
rect 6664 21734 6676 21786
rect 6728 21734 6740 21786
rect 6792 21734 6804 21786
rect 6856 21734 12146 21786
rect 12198 21734 12210 21786
rect 12262 21734 12274 21786
rect 12326 21734 12338 21786
rect 12390 21734 12402 21786
rect 12454 21734 17744 21786
rect 17796 21734 17808 21786
rect 17860 21734 17872 21786
rect 17924 21734 17936 21786
rect 17988 21734 18000 21786
rect 18052 21734 23460 21786
rect 1104 21712 23460 21734
rect 290 21632 296 21684
rect 348 21672 354 21684
rect 1489 21675 1547 21681
rect 1489 21672 1501 21675
rect 348 21644 1501 21672
rect 348 21632 354 21644
rect 1489 21641 1501 21644
rect 1535 21641 1547 21675
rect 2406 21672 2412 21684
rect 2367 21644 2412 21672
rect 1489 21635 1547 21641
rect 2406 21632 2412 21644
rect 2464 21632 2470 21684
rect 2958 21672 2964 21684
rect 2919 21644 2964 21672
rect 2958 21632 2964 21644
rect 3016 21632 3022 21684
rect 3234 21672 3240 21684
rect 3195 21644 3240 21672
rect 3234 21632 3240 21644
rect 3292 21632 3298 21684
rect 3694 21672 3700 21684
rect 3655 21644 3700 21672
rect 3694 21632 3700 21644
rect 3752 21632 3758 21684
rect 4982 21672 4988 21684
rect 4943 21644 4988 21672
rect 4982 21632 4988 21644
rect 5040 21632 5046 21684
rect 5626 21632 5632 21684
rect 5684 21672 5690 21684
rect 6454 21672 6460 21684
rect 5684 21644 6460 21672
rect 5684 21632 5690 21644
rect 6454 21632 6460 21644
rect 6512 21632 6518 21684
rect 7745 21675 7803 21681
rect 7745 21641 7757 21675
rect 7791 21672 7803 21675
rect 7834 21672 7840 21684
rect 7791 21644 7840 21672
rect 7791 21641 7803 21644
rect 7745 21635 7803 21641
rect 7834 21632 7840 21644
rect 7892 21632 7898 21684
rect 8297 21675 8355 21681
rect 8297 21641 8309 21675
rect 8343 21672 8355 21675
rect 8478 21672 8484 21684
rect 8343 21644 8484 21672
rect 8343 21641 8355 21644
rect 8297 21635 8355 21641
rect 8478 21632 8484 21644
rect 8536 21632 8542 21684
rect 9490 21632 9496 21684
rect 9548 21672 9554 21684
rect 10321 21675 10379 21681
rect 10321 21672 10333 21675
rect 9548 21644 10333 21672
rect 9548 21632 9554 21644
rect 10321 21641 10333 21644
rect 10367 21641 10379 21675
rect 10321 21635 10379 21641
rect 10965 21675 11023 21681
rect 10965 21641 10977 21675
rect 11011 21672 11023 21675
rect 11514 21672 11520 21684
rect 11011 21644 11520 21672
rect 11011 21641 11023 21644
rect 10965 21635 11023 21641
rect 11514 21632 11520 21644
rect 11572 21632 11578 21684
rect 11701 21675 11759 21681
rect 11701 21641 11713 21675
rect 11747 21672 11759 21675
rect 12526 21672 12532 21684
rect 11747 21644 12434 21672
rect 12487 21644 12532 21672
rect 11747 21641 11759 21644
rect 11701 21635 11759 21641
rect 4246 21604 4252 21616
rect 2332 21576 4252 21604
rect 2332 21545 2360 21576
rect 4246 21564 4252 21576
rect 4304 21564 4310 21616
rect 4433 21607 4491 21613
rect 4433 21573 4445 21607
rect 4479 21604 4491 21607
rect 5442 21604 5448 21616
rect 4479 21576 5448 21604
rect 4479 21573 4491 21576
rect 4433 21567 4491 21573
rect 5442 21564 5448 21576
rect 5500 21564 5506 21616
rect 5905 21607 5963 21613
rect 5905 21573 5917 21607
rect 5951 21604 5963 21607
rect 6362 21604 6368 21616
rect 5951 21576 6368 21604
rect 5951 21573 5963 21576
rect 5905 21567 5963 21573
rect 6362 21564 6368 21576
rect 6420 21564 6426 21616
rect 7558 21604 7564 21616
rect 6656 21576 7564 21604
rect 1673 21539 1731 21545
rect 1673 21505 1685 21539
rect 1719 21505 1731 21539
rect 1673 21499 1731 21505
rect 2041 21539 2099 21545
rect 2041 21505 2053 21539
rect 2087 21536 2099 21539
rect 2317 21539 2375 21545
rect 2087 21508 2268 21536
rect 2087 21505 2099 21508
rect 2041 21499 2099 21505
rect 1688 21468 1716 21499
rect 1688 21440 2176 21468
rect 934 21360 940 21412
rect 992 21400 998 21412
rect 2148 21409 2176 21440
rect 1857 21403 1915 21409
rect 1857 21400 1869 21403
rect 992 21372 1869 21400
rect 992 21360 998 21372
rect 1857 21369 1869 21372
rect 1903 21369 1915 21403
rect 1857 21363 1915 21369
rect 2133 21403 2191 21409
rect 2133 21369 2145 21403
rect 2179 21369 2191 21403
rect 2240 21400 2268 21508
rect 2317 21505 2329 21539
rect 2363 21505 2375 21539
rect 2317 21499 2375 21505
rect 2593 21539 2651 21545
rect 2593 21505 2605 21539
rect 2639 21536 2651 21539
rect 2774 21536 2780 21548
rect 2639 21508 2780 21536
rect 2639 21505 2651 21508
rect 2593 21499 2651 21505
rect 2774 21496 2780 21508
rect 2832 21496 2838 21548
rect 2869 21539 2927 21545
rect 2869 21505 2881 21539
rect 2915 21536 2927 21539
rect 2958 21536 2964 21548
rect 2915 21508 2964 21536
rect 2915 21505 2927 21508
rect 2869 21499 2927 21505
rect 2958 21496 2964 21508
rect 3016 21496 3022 21548
rect 3142 21536 3148 21548
rect 3103 21508 3148 21536
rect 3142 21496 3148 21508
rect 3200 21496 3206 21548
rect 3418 21536 3424 21548
rect 3379 21508 3424 21536
rect 3418 21496 3424 21508
rect 3476 21496 3482 21548
rect 3513 21539 3571 21545
rect 3513 21505 3525 21539
rect 3559 21536 3571 21539
rect 3602 21536 3608 21548
rect 3559 21508 3608 21536
rect 3559 21505 3571 21508
rect 3513 21499 3571 21505
rect 3602 21496 3608 21508
rect 3660 21496 3666 21548
rect 3970 21536 3976 21548
rect 3931 21508 3976 21536
rect 3970 21496 3976 21508
rect 4028 21496 4034 21548
rect 4893 21539 4951 21545
rect 4893 21505 4905 21539
rect 4939 21505 4951 21539
rect 5166 21536 5172 21548
rect 5127 21508 5172 21536
rect 4893 21499 4951 21505
rect 3234 21428 3240 21480
rect 3292 21468 3298 21480
rect 3789 21471 3847 21477
rect 3789 21468 3801 21471
rect 3292 21440 3801 21468
rect 3292 21428 3298 21440
rect 3789 21437 3801 21440
rect 3835 21437 3847 21471
rect 3789 21431 3847 21437
rect 4249 21471 4307 21477
rect 4249 21437 4261 21471
rect 4295 21468 4307 21471
rect 4798 21468 4804 21480
rect 4295 21440 4804 21468
rect 4295 21437 4307 21440
rect 4249 21431 4307 21437
rect 4798 21428 4804 21440
rect 4856 21428 4862 21480
rect 4908 21468 4936 21499
rect 5166 21496 5172 21508
rect 5224 21496 5230 21548
rect 5535 21540 5593 21545
rect 5535 21539 5672 21540
rect 5535 21505 5547 21539
rect 5581 21536 5672 21539
rect 5718 21536 5724 21548
rect 5581 21512 5724 21536
rect 5581 21505 5593 21512
rect 5644 21508 5724 21512
rect 5535 21499 5593 21505
rect 5718 21496 5724 21508
rect 5776 21496 5782 21548
rect 6656 21545 6684 21576
rect 7558 21564 7564 21576
rect 7616 21564 7622 21616
rect 8757 21607 8815 21613
rect 8757 21573 8769 21607
rect 8803 21604 8815 21607
rect 10597 21607 10655 21613
rect 10597 21604 10609 21607
rect 8803 21576 10609 21604
rect 8803 21573 8815 21576
rect 8757 21567 8815 21573
rect 10597 21573 10609 21576
rect 10643 21573 10655 21607
rect 10597 21567 10655 21573
rect 11333 21607 11391 21613
rect 11333 21573 11345 21607
rect 11379 21604 11391 21607
rect 11882 21604 11888 21616
rect 11379 21576 11888 21604
rect 11379 21573 11391 21576
rect 11333 21567 11391 21573
rect 11882 21564 11888 21576
rect 11940 21564 11946 21616
rect 12406 21604 12434 21644
rect 12526 21632 12532 21644
rect 12584 21632 12590 21684
rect 13081 21675 13139 21681
rect 13081 21641 13093 21675
rect 13127 21672 13139 21675
rect 13354 21672 13360 21684
rect 13127 21644 13360 21672
rect 13127 21641 13139 21644
rect 13081 21635 13139 21641
rect 13354 21632 13360 21644
rect 13412 21632 13418 21684
rect 13449 21675 13507 21681
rect 13449 21641 13461 21675
rect 13495 21672 13507 21675
rect 13722 21672 13728 21684
rect 13495 21644 13728 21672
rect 13495 21641 13507 21644
rect 13449 21635 13507 21641
rect 13722 21632 13728 21644
rect 13780 21632 13786 21684
rect 15286 21672 15292 21684
rect 13924 21644 15292 21672
rect 13924 21613 13952 21644
rect 15286 21632 15292 21644
rect 15344 21632 15350 21684
rect 15466 21675 15524 21681
rect 15466 21641 15478 21675
rect 15512 21672 15524 21675
rect 15654 21672 15660 21684
rect 15512 21644 15660 21672
rect 15512 21641 15524 21644
rect 15466 21635 15524 21641
rect 15654 21632 15660 21644
rect 15712 21632 15718 21684
rect 15930 21632 15936 21684
rect 15988 21672 15994 21684
rect 15988 21644 16252 21672
rect 15988 21632 15994 21644
rect 12989 21607 13047 21613
rect 12989 21604 13001 21607
rect 12406 21576 13001 21604
rect 12989 21573 13001 21576
rect 13035 21573 13047 21607
rect 12989 21567 13047 21573
rect 13909 21607 13967 21613
rect 13909 21573 13921 21607
rect 13955 21573 13967 21607
rect 13909 21567 13967 21573
rect 16025 21607 16083 21613
rect 16025 21573 16037 21607
rect 16071 21604 16083 21607
rect 16114 21604 16120 21616
rect 16071 21576 16120 21604
rect 16071 21573 16083 21576
rect 16025 21567 16083 21573
rect 16114 21564 16120 21576
rect 16172 21564 16178 21616
rect 16224 21613 16252 21644
rect 16942 21632 16948 21684
rect 17000 21672 17006 21684
rect 17497 21675 17555 21681
rect 17497 21672 17509 21675
rect 17000 21644 17509 21672
rect 17000 21632 17006 21644
rect 17497 21641 17509 21644
rect 17543 21641 17555 21675
rect 17497 21635 17555 21641
rect 17586 21632 17592 21684
rect 17644 21672 17650 21684
rect 18874 21672 18880 21684
rect 17644 21644 17816 21672
rect 18835 21644 18880 21672
rect 17644 21632 17650 21644
rect 16209 21607 16267 21613
rect 16209 21573 16221 21607
rect 16255 21573 16267 21607
rect 16209 21567 16267 21573
rect 16393 21607 16451 21613
rect 16393 21573 16405 21607
rect 16439 21604 16451 21607
rect 16439 21576 17724 21604
rect 16439 21573 16451 21576
rect 16393 21567 16451 21573
rect 6641 21539 6699 21545
rect 6641 21505 6653 21539
rect 6687 21505 6699 21539
rect 6641 21499 6699 21505
rect 7009 21539 7067 21545
rect 7009 21505 7021 21539
rect 7055 21536 7067 21539
rect 9490 21536 9496 21548
rect 7055 21508 7972 21536
rect 7055 21505 7067 21508
rect 7009 21499 7067 21505
rect 7650 21468 7656 21480
rect 4908 21440 7656 21468
rect 7650 21428 7656 21440
rect 7708 21428 7714 21480
rect 7834 21468 7840 21480
rect 7795 21440 7840 21468
rect 7834 21428 7840 21440
rect 7892 21428 7898 21480
rect 2685 21403 2743 21409
rect 2685 21400 2697 21403
rect 2240 21372 2697 21400
rect 2133 21363 2191 21369
rect 2685 21369 2697 21372
rect 2731 21369 2743 21403
rect 5353 21403 5411 21409
rect 5353 21400 5365 21403
rect 2685 21363 2743 21369
rect 3804 21372 5365 21400
rect 1394 21292 1400 21344
rect 1452 21332 1458 21344
rect 3804 21332 3832 21372
rect 5353 21369 5365 21372
rect 5399 21369 5411 21403
rect 5353 21363 5411 21369
rect 6086 21360 6092 21412
rect 6144 21400 6150 21412
rect 6825 21403 6883 21409
rect 6825 21400 6837 21403
rect 6144 21372 6837 21400
rect 6144 21360 6150 21372
rect 6825 21369 6837 21372
rect 6871 21369 6883 21403
rect 7944 21400 7972 21508
rect 8680 21508 9496 21536
rect 8021 21471 8079 21477
rect 8021 21437 8033 21471
rect 8067 21468 8079 21471
rect 8680 21468 8708 21508
rect 9490 21496 9496 21508
rect 9548 21496 9554 21548
rect 9585 21539 9643 21545
rect 9585 21505 9597 21539
rect 9631 21536 9643 21539
rect 10045 21539 10103 21545
rect 10045 21536 10057 21539
rect 9631 21508 10057 21536
rect 9631 21505 9643 21508
rect 9585 21499 9643 21505
rect 10045 21505 10057 21508
rect 10091 21505 10103 21539
rect 10045 21499 10103 21505
rect 10962 21496 10968 21548
rect 11020 21536 11026 21548
rect 11149 21539 11207 21545
rect 11149 21536 11161 21539
rect 11020 21508 11161 21536
rect 11020 21496 11026 21508
rect 11149 21505 11161 21508
rect 11195 21505 11207 21539
rect 11514 21536 11520 21548
rect 11475 21508 11520 21536
rect 11149 21499 11207 21505
rect 11514 21496 11520 21508
rect 11572 21496 11578 21548
rect 11790 21496 11796 21548
rect 11848 21536 11854 21548
rect 12069 21539 12127 21545
rect 12069 21536 12081 21539
rect 11848 21508 12081 21536
rect 11848 21496 11854 21508
rect 12069 21505 12081 21508
rect 12115 21505 12127 21539
rect 12069 21499 12127 21505
rect 12161 21539 12219 21545
rect 12161 21505 12173 21539
rect 12207 21536 12219 21539
rect 15102 21536 15108 21548
rect 12207 21508 12940 21536
rect 12207 21505 12219 21508
rect 12161 21499 12219 21505
rect 8846 21468 8852 21480
rect 8067 21440 8708 21468
rect 8807 21440 8852 21468
rect 8067 21437 8079 21440
rect 8021 21431 8079 21437
rect 8846 21428 8852 21440
rect 8904 21428 8910 21480
rect 9030 21468 9036 21480
rect 8991 21440 9036 21468
rect 9030 21428 9036 21440
rect 9088 21428 9094 21480
rect 9214 21428 9220 21480
rect 9272 21468 9278 21480
rect 9677 21471 9735 21477
rect 9677 21468 9689 21471
rect 9272 21440 9689 21468
rect 9272 21428 9278 21440
rect 9677 21437 9689 21440
rect 9723 21437 9735 21471
rect 9858 21468 9864 21480
rect 9819 21440 9864 21468
rect 9677 21431 9735 21437
rect 9858 21428 9864 21440
rect 9916 21428 9922 21480
rect 10318 21428 10324 21480
rect 10376 21468 10382 21480
rect 10376 21440 11284 21468
rect 10376 21428 10382 21440
rect 11146 21400 11152 21412
rect 7944 21372 11152 21400
rect 6825 21363 6883 21369
rect 11146 21360 11152 21372
rect 11204 21360 11210 21412
rect 11256 21400 11284 21440
rect 11698 21428 11704 21480
rect 11756 21468 11762 21480
rect 11885 21471 11943 21477
rect 11885 21468 11897 21471
rect 11756 21440 11897 21468
rect 11756 21428 11762 21440
rect 11885 21437 11897 21440
rect 11931 21437 11943 21471
rect 11885 21431 11943 21437
rect 12710 21428 12716 21480
rect 12768 21468 12774 21480
rect 12805 21471 12863 21477
rect 12805 21468 12817 21471
rect 12768 21440 12817 21468
rect 12768 21428 12774 21440
rect 12805 21437 12817 21440
rect 12851 21437 12863 21471
rect 12912 21468 12940 21508
rect 13280 21508 15108 21536
rect 13170 21468 13176 21480
rect 12912 21440 13176 21468
rect 12805 21431 12863 21437
rect 13170 21428 13176 21440
rect 13228 21428 13234 21480
rect 13280 21400 13308 21508
rect 15102 21496 15108 21508
rect 15160 21496 15166 21548
rect 15197 21539 15255 21545
rect 15197 21505 15209 21539
rect 15243 21536 15255 21539
rect 17313 21539 17371 21545
rect 15243 21508 16160 21536
rect 15243 21505 15255 21508
rect 15197 21499 15255 21505
rect 16132 21480 16160 21508
rect 17313 21505 17325 21539
rect 17359 21536 17371 21539
rect 17402 21536 17408 21548
rect 17359 21508 17408 21536
rect 17359 21505 17371 21508
rect 17313 21499 17371 21505
rect 17402 21496 17408 21508
rect 17460 21496 17466 21548
rect 17696 21545 17724 21576
rect 17681 21539 17739 21545
rect 17681 21505 17693 21539
rect 17727 21505 17739 21539
rect 17788 21536 17816 21644
rect 18874 21632 18880 21644
rect 18932 21632 18938 21684
rect 19153 21675 19211 21681
rect 19153 21641 19165 21675
rect 19199 21641 19211 21675
rect 19153 21635 19211 21641
rect 18230 21564 18236 21616
rect 18288 21604 18294 21616
rect 19168 21604 19196 21635
rect 19334 21632 19340 21684
rect 19392 21672 19398 21684
rect 19521 21675 19579 21681
rect 19521 21672 19533 21675
rect 19392 21644 19533 21672
rect 19392 21632 19398 21644
rect 19521 21641 19533 21644
rect 19567 21641 19579 21675
rect 20530 21672 20536 21684
rect 20491 21644 20536 21672
rect 19521 21635 19579 21641
rect 20530 21632 20536 21644
rect 20588 21632 20594 21684
rect 20622 21632 20628 21684
rect 20680 21672 20686 21684
rect 21358 21672 21364 21684
rect 20680 21644 21364 21672
rect 20680 21632 20686 21644
rect 21358 21632 21364 21644
rect 21416 21632 21422 21684
rect 21453 21675 21511 21681
rect 21453 21641 21465 21675
rect 21499 21672 21511 21675
rect 22281 21675 22339 21681
rect 22281 21672 22293 21675
rect 21499 21644 22293 21672
rect 21499 21641 21511 21644
rect 21453 21635 21511 21641
rect 22281 21641 22293 21644
rect 22327 21641 22339 21675
rect 22281 21635 22339 21641
rect 18288 21576 19196 21604
rect 19981 21607 20039 21613
rect 18288 21564 18294 21576
rect 19981 21573 19993 21607
rect 20027 21604 20039 21607
rect 21818 21604 21824 21616
rect 20027 21576 21824 21604
rect 20027 21573 20039 21576
rect 19981 21567 20039 21573
rect 21818 21564 21824 21576
rect 21876 21564 21882 21616
rect 22066 21576 22876 21604
rect 19058 21536 19064 21548
rect 17788 21508 18920 21536
rect 19019 21508 19064 21536
rect 17681 21499 17739 21505
rect 14366 21468 14372 21480
rect 11256 21372 13308 21400
rect 13372 21440 14372 21468
rect 1452 21304 3832 21332
rect 1452 21292 1458 21304
rect 4522 21292 4528 21344
rect 4580 21332 4586 21344
rect 4709 21335 4767 21341
rect 4709 21332 4721 21335
rect 4580 21304 4721 21332
rect 4580 21292 4586 21304
rect 4709 21301 4721 21304
rect 4755 21301 4767 21335
rect 4709 21295 4767 21301
rect 5718 21292 5724 21344
rect 5776 21332 5782 21344
rect 5813 21335 5871 21341
rect 5813 21332 5825 21335
rect 5776 21304 5825 21332
rect 5776 21292 5782 21304
rect 5813 21301 5825 21304
rect 5859 21301 5871 21335
rect 5813 21295 5871 21301
rect 6270 21292 6276 21344
rect 6328 21332 6334 21344
rect 6457 21335 6515 21341
rect 6457 21332 6469 21335
rect 6328 21304 6469 21332
rect 6328 21292 6334 21304
rect 6457 21301 6469 21304
rect 6503 21301 6515 21335
rect 7374 21332 7380 21344
rect 7335 21304 7380 21332
rect 6457 21295 6515 21301
rect 7374 21292 7380 21304
rect 7432 21292 7438 21344
rect 8386 21332 8392 21344
rect 8347 21304 8392 21332
rect 8386 21292 8392 21304
rect 8444 21292 8450 21344
rect 8478 21292 8484 21344
rect 8536 21332 8542 21344
rect 8938 21332 8944 21344
rect 8536 21304 8944 21332
rect 8536 21292 8542 21304
rect 8938 21292 8944 21304
rect 8996 21332 9002 21344
rect 9217 21335 9275 21341
rect 9217 21332 9229 21335
rect 8996 21304 9229 21332
rect 8996 21292 9002 21304
rect 9217 21301 9229 21304
rect 9263 21301 9275 21335
rect 9217 21295 9275 21301
rect 10502 21292 10508 21344
rect 10560 21332 10566 21344
rect 13372 21332 13400 21440
rect 14366 21428 14372 21440
rect 14424 21428 14430 21480
rect 15010 21468 15016 21480
rect 14568 21440 15016 21468
rect 13630 21360 13636 21412
rect 13688 21400 13694 21412
rect 13725 21403 13783 21409
rect 13725 21400 13737 21403
rect 13688 21372 13737 21400
rect 13688 21360 13694 21372
rect 13725 21369 13737 21372
rect 13771 21369 13783 21403
rect 14182 21400 14188 21412
rect 13725 21363 13783 21369
rect 13924 21372 14188 21400
rect 10560 21304 13400 21332
rect 13541 21335 13599 21341
rect 10560 21292 10566 21304
rect 13541 21301 13553 21335
rect 13587 21332 13599 21335
rect 13924 21332 13952 21372
rect 14182 21360 14188 21372
rect 14240 21400 14246 21412
rect 14568 21400 14596 21440
rect 15010 21428 15016 21440
rect 15068 21428 15074 21480
rect 15286 21428 15292 21480
rect 15344 21468 15350 21480
rect 15427 21471 15485 21477
rect 15427 21468 15439 21471
rect 15344 21440 15439 21468
rect 15344 21428 15350 21440
rect 15427 21437 15439 21440
rect 15473 21437 15485 21471
rect 15427 21431 15485 21437
rect 15933 21471 15991 21477
rect 15933 21437 15945 21471
rect 15979 21437 15991 21471
rect 15933 21431 15991 21437
rect 14240 21372 14596 21400
rect 14240 21360 14246 21372
rect 13587 21304 13952 21332
rect 13587 21301 13599 21304
rect 13541 21295 13599 21301
rect 13998 21292 14004 21344
rect 14056 21332 14062 21344
rect 14093 21335 14151 21341
rect 14093 21332 14105 21335
rect 14056 21304 14105 21332
rect 14056 21292 14062 21304
rect 14093 21301 14105 21304
rect 14139 21301 14151 21335
rect 14093 21295 14151 21301
rect 15194 21292 15200 21344
rect 15252 21332 15258 21344
rect 15948 21332 15976 21431
rect 16114 21428 16120 21480
rect 16172 21428 16178 21480
rect 16758 21468 16764 21480
rect 16719 21440 16764 21468
rect 16758 21428 16764 21440
rect 16816 21428 16822 21480
rect 17957 21471 18015 21477
rect 17957 21468 17969 21471
rect 17696 21440 17969 21468
rect 16776 21400 16804 21428
rect 17402 21400 17408 21412
rect 16776 21372 17408 21400
rect 17402 21360 17408 21372
rect 17460 21400 17466 21412
rect 17696 21400 17724 21440
rect 17957 21437 17969 21440
rect 18003 21437 18015 21471
rect 17957 21431 18015 21437
rect 18233 21471 18291 21477
rect 18233 21437 18245 21471
rect 18279 21468 18291 21471
rect 18892 21468 18920 21508
rect 19058 21496 19064 21508
rect 19116 21496 19122 21548
rect 19337 21539 19395 21545
rect 19337 21505 19349 21539
rect 19383 21505 19395 21539
rect 19886 21536 19892 21548
rect 19847 21508 19892 21536
rect 19337 21499 19395 21505
rect 19352 21468 19380 21499
rect 19886 21496 19892 21508
rect 19944 21496 19950 21548
rect 20346 21536 20352 21548
rect 20307 21508 20352 21536
rect 20346 21496 20352 21508
rect 20404 21496 20410 21548
rect 21082 21536 21088 21548
rect 21043 21508 21088 21536
rect 21082 21496 21088 21508
rect 21140 21496 21146 21548
rect 22066 21536 22094 21576
rect 21284 21508 22094 21536
rect 18279 21440 18828 21468
rect 18892 21440 19380 21468
rect 18279 21437 18291 21440
rect 18233 21431 18291 21437
rect 17460 21372 17724 21400
rect 18800 21400 18828 21440
rect 19518 21428 19524 21480
rect 19576 21468 19582 21480
rect 20073 21471 20131 21477
rect 20073 21468 20085 21471
rect 19576 21440 20085 21468
rect 19576 21428 19582 21440
rect 20073 21437 20085 21440
rect 20119 21437 20131 21471
rect 20073 21431 20131 21437
rect 20162 21428 20168 21480
rect 20220 21468 20226 21480
rect 20809 21471 20867 21477
rect 20809 21468 20821 21471
rect 20220 21440 20821 21468
rect 20220 21428 20226 21440
rect 20809 21437 20821 21440
rect 20855 21437 20867 21471
rect 20809 21431 20867 21437
rect 20993 21471 21051 21477
rect 20993 21437 21005 21471
rect 21039 21468 21051 21471
rect 21174 21468 21180 21480
rect 21039 21440 21180 21468
rect 21039 21437 21051 21440
rect 20993 21431 21051 21437
rect 21174 21428 21180 21440
rect 21232 21428 21238 21480
rect 19702 21400 19708 21412
rect 18800 21372 19708 21400
rect 17460 21360 17466 21372
rect 19702 21360 19708 21372
rect 19760 21360 19766 21412
rect 19794 21360 19800 21412
rect 19852 21400 19858 21412
rect 21284 21400 21312 21508
rect 22186 21496 22192 21548
rect 22244 21536 22250 21548
rect 22848 21545 22876 21576
rect 22833 21539 22891 21545
rect 22244 21508 22289 21536
rect 22244 21496 22250 21508
rect 22833 21505 22845 21539
rect 22879 21505 22891 21539
rect 22833 21499 22891 21505
rect 21726 21428 21732 21480
rect 21784 21468 21790 21480
rect 22373 21471 22431 21477
rect 21784 21440 22094 21468
rect 21784 21428 21790 21440
rect 19852 21372 21312 21400
rect 21637 21403 21695 21409
rect 19852 21360 19858 21372
rect 21637 21369 21649 21403
rect 21683 21400 21695 21403
rect 22066 21400 22094 21440
rect 22373 21437 22385 21471
rect 22419 21437 22431 21471
rect 22373 21431 22431 21437
rect 22388 21400 22416 21431
rect 21683 21372 21956 21400
rect 22066 21372 22416 21400
rect 21683 21369 21695 21372
rect 21637 21363 21695 21369
rect 15252 21304 15976 21332
rect 15252 21292 15258 21304
rect 16022 21292 16028 21344
rect 16080 21332 16086 21344
rect 17773 21335 17831 21341
rect 17773 21332 17785 21335
rect 16080 21304 17785 21332
rect 16080 21292 16086 21304
rect 17773 21301 17785 21304
rect 17819 21301 17831 21335
rect 17773 21295 17831 21301
rect 17862 21292 17868 21344
rect 17920 21332 17926 21344
rect 20622 21332 20628 21344
rect 17920 21304 20628 21332
rect 17920 21292 17926 21304
rect 20622 21292 20628 21304
rect 20680 21292 20686 21344
rect 21358 21292 21364 21344
rect 21416 21332 21422 21344
rect 21821 21335 21879 21341
rect 21821 21332 21833 21335
rect 21416 21304 21833 21332
rect 21416 21292 21422 21304
rect 21821 21301 21833 21304
rect 21867 21301 21879 21335
rect 21928 21332 21956 21372
rect 22094 21332 22100 21344
rect 21928 21304 22100 21332
rect 21821 21295 21879 21301
rect 22094 21292 22100 21304
rect 22152 21332 22158 21344
rect 22649 21335 22707 21341
rect 22649 21332 22661 21335
rect 22152 21304 22661 21332
rect 22152 21292 22158 21304
rect 22649 21301 22661 21304
rect 22695 21301 22707 21335
rect 23014 21332 23020 21344
rect 22975 21304 23020 21332
rect 22649 21295 22707 21301
rect 23014 21292 23020 21304
rect 23072 21292 23078 21344
rect 1104 21242 23460 21264
rect 1104 21190 3749 21242
rect 3801 21190 3813 21242
rect 3865 21190 3877 21242
rect 3929 21190 3941 21242
rect 3993 21190 4005 21242
rect 4057 21190 9347 21242
rect 9399 21190 9411 21242
rect 9463 21190 9475 21242
rect 9527 21190 9539 21242
rect 9591 21190 9603 21242
rect 9655 21190 14945 21242
rect 14997 21190 15009 21242
rect 15061 21190 15073 21242
rect 15125 21190 15137 21242
rect 15189 21190 15201 21242
rect 15253 21190 20543 21242
rect 20595 21190 20607 21242
rect 20659 21190 20671 21242
rect 20723 21190 20735 21242
rect 20787 21190 20799 21242
rect 20851 21190 23460 21242
rect 1104 21168 23460 21190
rect 3973 21131 4031 21137
rect 3973 21097 3985 21131
rect 4019 21128 4031 21131
rect 4062 21128 4068 21140
rect 4019 21100 4068 21128
rect 4019 21097 4031 21100
rect 3973 21091 4031 21097
rect 4062 21088 4068 21100
rect 4120 21088 4126 21140
rect 4338 21128 4344 21140
rect 4299 21100 4344 21128
rect 4338 21088 4344 21100
rect 4396 21088 4402 21140
rect 5920 21100 7788 21128
rect 2774 21020 2780 21072
rect 2832 21060 2838 21072
rect 2832 21032 2877 21060
rect 2832 21020 2838 21032
rect 2958 21020 2964 21072
rect 3016 21060 3022 21072
rect 5920 21060 5948 21100
rect 3016 21032 5948 21060
rect 7760 21060 7788 21100
rect 7834 21088 7840 21140
rect 7892 21128 7898 21140
rect 8021 21131 8079 21137
rect 8021 21128 8033 21131
rect 7892 21100 8033 21128
rect 7892 21088 7898 21100
rect 8021 21097 8033 21100
rect 8067 21097 8079 21131
rect 9766 21128 9772 21140
rect 9727 21100 9772 21128
rect 8021 21091 8079 21097
rect 9766 21088 9772 21100
rect 9824 21088 9830 21140
rect 9953 21131 10011 21137
rect 9953 21097 9965 21131
rect 9999 21128 10011 21131
rect 10226 21128 10232 21140
rect 9999 21100 10232 21128
rect 9999 21097 10011 21100
rect 9953 21091 10011 21097
rect 10226 21088 10232 21100
rect 10284 21088 10290 21140
rect 12805 21131 12863 21137
rect 11900 21100 12756 21128
rect 8478 21060 8484 21072
rect 7760 21032 8484 21060
rect 3016 21020 3022 21032
rect 8478 21020 8484 21032
rect 8536 21020 8542 21072
rect 8662 21020 8668 21072
rect 8720 21060 8726 21072
rect 9858 21060 9864 21072
rect 8720 21032 9864 21060
rect 8720 21020 8726 21032
rect 9858 21020 9864 21032
rect 9916 21020 9922 21072
rect 4801 20995 4859 21001
rect 4801 20961 4813 20995
rect 4847 20992 4859 20995
rect 5442 20992 5448 21004
rect 4847 20964 5448 20992
rect 4847 20961 4859 20964
rect 4801 20955 4859 20961
rect 5442 20952 5448 20964
rect 5500 20952 5506 21004
rect 7282 20992 7288 21004
rect 7243 20964 7288 20992
rect 7282 20952 7288 20964
rect 7340 20952 7346 21004
rect 8294 20992 8300 21004
rect 7760 20964 8300 20992
rect 3418 20884 3424 20936
rect 3476 20924 3482 20936
rect 3605 20927 3663 20933
rect 3605 20924 3617 20927
rect 3476 20896 3617 20924
rect 3476 20884 3482 20896
rect 3605 20893 3617 20896
rect 3651 20924 3663 20927
rect 3694 20924 3700 20936
rect 3651 20896 3700 20924
rect 3651 20893 3663 20896
rect 3605 20887 3663 20893
rect 3694 20884 3700 20896
rect 3752 20884 3758 20936
rect 4157 20927 4215 20933
rect 4157 20893 4169 20927
rect 4203 20924 4215 20927
rect 4338 20924 4344 20936
rect 4203 20896 4344 20924
rect 4203 20893 4215 20896
rect 4157 20887 4215 20893
rect 4338 20884 4344 20896
rect 4396 20884 4402 20936
rect 6178 20884 6184 20936
rect 6236 20924 6242 20936
rect 6825 20927 6883 20933
rect 6825 20924 6837 20927
rect 6236 20896 6837 20924
rect 6236 20884 6242 20896
rect 6825 20893 6837 20896
rect 6871 20893 6883 20927
rect 7760 20924 7788 20964
rect 8294 20952 8300 20964
rect 8352 20952 8358 21004
rect 8570 20992 8576 21004
rect 8531 20964 8576 20992
rect 8570 20952 8576 20964
rect 8628 20952 8634 21004
rect 9125 20995 9183 21001
rect 9125 20961 9137 20995
rect 9171 20961 9183 20995
rect 9125 20955 9183 20961
rect 10045 20995 10103 21001
rect 10045 20961 10057 20995
rect 10091 20992 10103 20995
rect 10318 20992 10324 21004
rect 10091 20964 10324 20992
rect 10091 20961 10103 20964
rect 10045 20955 10103 20961
rect 6825 20887 6883 20893
rect 7024 20896 7788 20924
rect 3142 20816 3148 20868
rect 3200 20856 3206 20868
rect 3329 20859 3387 20865
rect 3329 20856 3341 20859
rect 3200 20828 3341 20856
rect 3200 20816 3206 20828
rect 3329 20825 3341 20828
rect 3375 20856 3387 20859
rect 3375 20828 6408 20856
rect 3375 20825 3387 20828
rect 3329 20819 3387 20825
rect 3602 20748 3608 20800
rect 3660 20788 3666 20800
rect 3878 20788 3884 20800
rect 3660 20760 3884 20788
rect 3660 20748 3666 20760
rect 3878 20748 3884 20760
rect 3936 20748 3942 20800
rect 4338 20748 4344 20800
rect 4396 20788 4402 20800
rect 4893 20791 4951 20797
rect 4893 20788 4905 20791
rect 4396 20760 4905 20788
rect 4396 20748 4402 20760
rect 4893 20757 4905 20760
rect 4939 20757 4951 20791
rect 4893 20751 4951 20757
rect 4982 20748 4988 20800
rect 5040 20788 5046 20800
rect 5350 20788 5356 20800
rect 5040 20760 5085 20788
rect 5311 20760 5356 20788
rect 5040 20748 5046 20760
rect 5350 20748 5356 20760
rect 5408 20748 5414 20800
rect 5442 20748 5448 20800
rect 5500 20788 5506 20800
rect 6380 20788 6408 20828
rect 6454 20816 6460 20868
rect 6512 20856 6518 20868
rect 6558 20859 6616 20865
rect 6558 20856 6570 20859
rect 6512 20828 6570 20856
rect 6512 20816 6518 20828
rect 6558 20825 6570 20828
rect 6604 20825 6616 20859
rect 6558 20819 6616 20825
rect 7024 20788 7052 20896
rect 7834 20884 7840 20936
rect 7892 20924 7898 20936
rect 9140 20924 9168 20955
rect 10318 20952 10324 20964
rect 10376 20952 10382 21004
rect 10508 20995 10566 21001
rect 10508 20961 10520 20995
rect 10554 20992 10566 20995
rect 10594 20992 10600 21004
rect 10554 20964 10600 20992
rect 10554 20961 10566 20964
rect 10508 20955 10566 20961
rect 10594 20952 10600 20964
rect 10652 20952 10658 21004
rect 10781 20927 10839 20933
rect 10781 20924 10793 20927
rect 7892 20896 9168 20924
rect 10152 20896 10793 20924
rect 7892 20884 7898 20896
rect 7101 20859 7159 20865
rect 7101 20825 7113 20859
rect 7147 20856 7159 20859
rect 7561 20859 7619 20865
rect 7561 20856 7573 20859
rect 7147 20828 7573 20856
rect 7147 20825 7159 20828
rect 7101 20819 7159 20825
rect 7561 20825 7573 20828
rect 7607 20825 7619 20859
rect 8938 20856 8944 20868
rect 7561 20819 7619 20825
rect 8496 20828 8944 20856
rect 8496 20800 8524 20828
rect 8938 20816 8944 20828
rect 8996 20816 9002 20868
rect 9309 20859 9367 20865
rect 9309 20825 9321 20859
rect 9355 20856 9367 20859
rect 9950 20856 9956 20868
rect 9355 20828 9956 20856
rect 9355 20825 9367 20828
rect 9309 20819 9367 20825
rect 9950 20816 9956 20828
rect 10008 20856 10014 20868
rect 10152 20856 10180 20896
rect 10781 20893 10793 20896
rect 10827 20893 10839 20927
rect 10781 20887 10839 20893
rect 10008 20828 10180 20856
rect 10008 20816 10014 20828
rect 7466 20788 7472 20800
rect 5500 20760 5545 20788
rect 6380 20760 7052 20788
rect 7427 20760 7472 20788
rect 5500 20748 5506 20760
rect 7466 20748 7472 20760
rect 7524 20748 7530 20800
rect 7926 20788 7932 20800
rect 7887 20760 7932 20788
rect 7926 20748 7932 20760
rect 7984 20748 7990 20800
rect 8294 20748 8300 20800
rect 8352 20788 8358 20800
rect 8389 20791 8447 20797
rect 8389 20788 8401 20791
rect 8352 20760 8401 20788
rect 8352 20748 8358 20760
rect 8389 20757 8401 20760
rect 8435 20757 8447 20791
rect 8389 20751 8447 20757
rect 8478 20748 8484 20800
rect 8536 20788 8542 20800
rect 8536 20760 8581 20788
rect 8536 20748 8542 20760
rect 8754 20748 8760 20800
rect 8812 20788 8818 20800
rect 9401 20791 9459 20797
rect 9401 20788 9413 20791
rect 8812 20760 9413 20788
rect 8812 20748 8818 20760
rect 9401 20757 9413 20760
rect 9447 20757 9459 20791
rect 9401 20751 9459 20757
rect 9766 20748 9772 20800
rect 9824 20788 9830 20800
rect 10502 20788 10508 20800
rect 10560 20797 10566 20800
rect 9824 20760 10508 20788
rect 9824 20748 9830 20760
rect 10502 20748 10508 20760
rect 10560 20788 10569 20797
rect 10560 20760 10605 20788
rect 10560 20751 10569 20760
rect 10560 20748 10566 20751
rect 10686 20748 10692 20800
rect 10744 20788 10750 20800
rect 11900 20797 11928 21100
rect 12066 21020 12072 21072
rect 12124 21060 12130 21072
rect 12124 21032 12388 21060
rect 12124 21020 12130 21032
rect 12360 21001 12388 21032
rect 12253 20995 12311 21001
rect 12253 20961 12265 20995
rect 12299 20961 12311 20995
rect 12253 20955 12311 20961
rect 12345 20995 12403 21001
rect 12345 20961 12357 20995
rect 12391 20961 12403 20995
rect 12728 20992 12756 21100
rect 12805 21097 12817 21131
rect 12851 21128 12863 21131
rect 13538 21128 13544 21140
rect 12851 21100 13544 21128
rect 12851 21097 12863 21100
rect 12805 21091 12863 21097
rect 13538 21088 13544 21100
rect 13596 21088 13602 21140
rect 13722 21128 13728 21140
rect 13683 21100 13728 21128
rect 13722 21088 13728 21100
rect 13780 21088 13786 21140
rect 14461 21131 14519 21137
rect 14461 21097 14473 21131
rect 14507 21128 14519 21131
rect 14826 21128 14832 21140
rect 14507 21100 14832 21128
rect 14507 21097 14519 21100
rect 14461 21091 14519 21097
rect 14826 21088 14832 21100
rect 14884 21088 14890 21140
rect 14918 21088 14924 21140
rect 14976 21128 14982 21140
rect 15470 21128 15476 21140
rect 14976 21100 15476 21128
rect 14976 21088 14982 21100
rect 15470 21088 15476 21100
rect 15528 21088 15534 21140
rect 15746 21088 15752 21140
rect 15804 21128 15810 21140
rect 17037 21131 17095 21137
rect 17037 21128 17049 21131
rect 15804 21100 17049 21128
rect 15804 21088 15810 21100
rect 17037 21097 17049 21100
rect 17083 21097 17095 21131
rect 18049 21131 18107 21137
rect 17037 21091 17095 21097
rect 17144 21100 17448 21128
rect 12894 21020 12900 21072
rect 12952 21060 12958 21072
rect 14093 21063 14151 21069
rect 14093 21060 14105 21063
rect 12952 21032 14105 21060
rect 12952 21020 12958 21032
rect 14093 21029 14105 21032
rect 14139 21029 14151 21063
rect 14093 21023 14151 21029
rect 16942 21020 16948 21072
rect 17000 21060 17006 21072
rect 17144 21060 17172 21100
rect 17000 21032 17172 21060
rect 17000 21020 17006 21032
rect 17218 21020 17224 21072
rect 17276 21060 17282 21072
rect 17420 21060 17448 21100
rect 18049 21097 18061 21131
rect 18095 21128 18107 21131
rect 18138 21128 18144 21140
rect 18095 21100 18144 21128
rect 18095 21097 18107 21100
rect 18049 21091 18107 21097
rect 18138 21088 18144 21100
rect 18196 21088 18202 21140
rect 18598 21128 18604 21140
rect 18559 21100 18604 21128
rect 18598 21088 18604 21100
rect 18656 21088 18662 21140
rect 18966 21088 18972 21140
rect 19024 21128 19030 21140
rect 20073 21131 20131 21137
rect 20073 21128 20085 21131
rect 19024 21100 20085 21128
rect 19024 21088 19030 21100
rect 20073 21097 20085 21100
rect 20119 21097 20131 21131
rect 20073 21091 20131 21097
rect 20438 21088 20444 21140
rect 20496 21128 20502 21140
rect 22646 21128 22652 21140
rect 20496 21100 22094 21128
rect 22607 21100 22652 21128
rect 20496 21088 20502 21100
rect 17276 21032 17321 21060
rect 17420 21032 18092 21060
rect 17276 21020 17282 21032
rect 13541 20995 13599 21001
rect 12728 20964 13492 20992
rect 12345 20955 12403 20961
rect 12268 20924 12296 20955
rect 12802 20924 12808 20936
rect 12268 20896 12808 20924
rect 12802 20884 12808 20896
rect 12860 20884 12866 20936
rect 12066 20816 12072 20868
rect 12124 20856 12130 20868
rect 13265 20859 13323 20865
rect 13265 20856 13277 20859
rect 12124 20828 13277 20856
rect 12124 20816 12130 20828
rect 13265 20825 13277 20828
rect 13311 20825 13323 20859
rect 13464 20856 13492 20964
rect 13541 20961 13553 20995
rect 13587 20992 13599 20995
rect 13630 20992 13636 21004
rect 13587 20964 13636 20992
rect 13587 20961 13599 20964
rect 13541 20955 13599 20961
rect 13630 20952 13636 20964
rect 13688 20952 13694 21004
rect 14553 20995 14611 21001
rect 14553 20961 14565 20995
rect 14599 20992 14611 20995
rect 14918 20992 14924 21004
rect 14599 20964 14924 20992
rect 14599 20961 14611 20964
rect 14553 20955 14611 20961
rect 14918 20952 14924 20964
rect 14976 20952 14982 21004
rect 15059 20995 15117 21001
rect 15059 20961 15071 20995
rect 15105 20992 15117 20995
rect 16298 20992 16304 21004
rect 15105 20964 16304 20992
rect 15105 20961 15117 20964
rect 15059 20955 15117 20961
rect 16298 20952 16304 20964
rect 16356 20952 16362 21004
rect 16850 20952 16856 21004
rect 16908 20992 16914 21004
rect 17586 20992 17592 21004
rect 16908 20964 17592 20992
rect 16908 20952 16914 20964
rect 17586 20952 17592 20964
rect 17644 20952 17650 21004
rect 17862 20952 17868 21004
rect 17920 20992 17926 21004
rect 18064 20992 18092 21032
rect 18322 21020 18328 21072
rect 18380 21060 18386 21072
rect 22066 21060 22094 21100
rect 22646 21088 22652 21100
rect 22704 21088 22710 21140
rect 23198 21060 23204 21072
rect 18380 21032 19564 21060
rect 22066 21032 23204 21060
rect 18380 21020 18386 21032
rect 19536 21001 19564 21032
rect 23198 21020 23204 21032
rect 23256 21020 23262 21072
rect 19337 20995 19395 21001
rect 19337 20992 19349 20995
rect 17920 20964 17965 20992
rect 18064 20964 19349 20992
rect 17920 20952 17926 20964
rect 19337 20961 19349 20964
rect 19383 20961 19395 20995
rect 19337 20955 19395 20961
rect 19521 20995 19579 21001
rect 19521 20961 19533 20995
rect 19567 20961 19579 20995
rect 20904 20995 20962 21001
rect 20904 20992 20916 20995
rect 19521 20955 19579 20961
rect 20088 20964 20916 20992
rect 13906 20924 13912 20936
rect 13867 20896 13912 20924
rect 13906 20884 13912 20896
rect 13964 20884 13970 20936
rect 14274 20924 14280 20936
rect 14235 20896 14280 20924
rect 14274 20884 14280 20896
rect 14332 20884 14338 20936
rect 15289 20927 15347 20933
rect 15289 20924 15301 20927
rect 14660 20896 15301 20924
rect 14660 20856 14688 20896
rect 15289 20893 15301 20896
rect 15335 20924 15347 20927
rect 15378 20924 15384 20936
rect 15335 20896 15384 20924
rect 15335 20893 15347 20896
rect 15289 20887 15347 20893
rect 15378 20884 15384 20896
rect 15436 20884 15442 20936
rect 17494 20884 17500 20936
rect 17552 20924 17558 20936
rect 18233 20927 18291 20933
rect 18233 20924 18245 20927
rect 17552 20920 17632 20924
rect 17788 20920 18245 20924
rect 17552 20896 18245 20920
rect 17552 20884 17558 20896
rect 17604 20892 17816 20896
rect 18233 20893 18245 20896
rect 18279 20893 18291 20927
rect 18506 20924 18512 20936
rect 18467 20896 18512 20924
rect 18233 20887 18291 20893
rect 18506 20884 18512 20896
rect 18564 20884 18570 20936
rect 18598 20884 18604 20936
rect 18656 20924 18662 20936
rect 18785 20927 18843 20933
rect 18785 20924 18797 20927
rect 18656 20896 18797 20924
rect 18656 20884 18662 20896
rect 18785 20893 18797 20896
rect 18831 20893 18843 20927
rect 18785 20887 18843 20893
rect 18874 20884 18880 20936
rect 18932 20924 18938 20936
rect 20088 20924 20116 20964
rect 20904 20961 20916 20964
rect 20950 20992 20962 20995
rect 21082 20992 21088 21004
rect 20950 20964 21088 20992
rect 20950 20961 20962 20964
rect 20904 20955 20962 20961
rect 21082 20952 21088 20964
rect 21140 20952 21146 21004
rect 20254 20924 20260 20936
rect 18932 20896 20116 20924
rect 20215 20896 20260 20924
rect 18932 20884 18938 20896
rect 20254 20884 20260 20896
rect 20312 20884 20318 20936
rect 20441 20927 20499 20933
rect 20441 20893 20453 20927
rect 20487 20924 20499 20927
rect 20990 20924 20996 20936
rect 20487 20896 20996 20924
rect 20487 20893 20499 20896
rect 20441 20887 20499 20893
rect 13464 20828 14688 20856
rect 13265 20819 13323 20825
rect 16114 20816 16120 20868
rect 16172 20856 16178 20868
rect 19061 20859 19119 20865
rect 16172 20828 18368 20856
rect 16172 20816 16178 20828
rect 11885 20791 11943 20797
rect 11885 20788 11897 20791
rect 10744 20760 11897 20788
rect 10744 20748 10750 20760
rect 11885 20757 11897 20760
rect 11931 20757 11943 20791
rect 11885 20751 11943 20757
rect 12437 20791 12495 20797
rect 12437 20757 12449 20791
rect 12483 20788 12495 20791
rect 12526 20788 12532 20800
rect 12483 20760 12532 20788
rect 12483 20757 12495 20760
rect 12437 20751 12495 20757
rect 12526 20748 12532 20760
rect 12584 20748 12590 20800
rect 12894 20748 12900 20800
rect 12952 20788 12958 20800
rect 13357 20791 13415 20797
rect 12952 20760 12997 20788
rect 12952 20748 12958 20760
rect 13357 20757 13369 20791
rect 13403 20788 13415 20791
rect 13446 20788 13452 20800
rect 13403 20760 13452 20788
rect 13403 20757 13415 20760
rect 13357 20751 13415 20757
rect 13446 20748 13452 20760
rect 13504 20748 13510 20800
rect 14826 20748 14832 20800
rect 14884 20788 14890 20800
rect 15019 20791 15077 20797
rect 15019 20788 15031 20791
rect 14884 20760 15031 20788
rect 14884 20748 14890 20760
rect 15019 20757 15031 20760
rect 15065 20757 15077 20791
rect 15019 20751 15077 20757
rect 15378 20748 15384 20800
rect 15436 20788 15442 20800
rect 16022 20788 16028 20800
rect 15436 20760 16028 20788
rect 15436 20748 15442 20760
rect 16022 20748 16028 20760
rect 16080 20748 16086 20800
rect 16206 20748 16212 20800
rect 16264 20788 16270 20800
rect 16393 20791 16451 20797
rect 16393 20788 16405 20791
rect 16264 20760 16405 20788
rect 16264 20748 16270 20760
rect 16393 20757 16405 20760
rect 16439 20757 16451 20791
rect 16393 20751 16451 20757
rect 16482 20748 16488 20800
rect 16540 20788 16546 20800
rect 16758 20788 16764 20800
rect 16540 20760 16585 20788
rect 16719 20760 16764 20788
rect 16540 20748 16546 20760
rect 16758 20748 16764 20760
rect 16816 20748 16822 20800
rect 17494 20748 17500 20800
rect 17552 20788 17558 20800
rect 17589 20791 17647 20797
rect 17589 20788 17601 20791
rect 17552 20760 17601 20788
rect 17552 20748 17558 20760
rect 17589 20757 17601 20760
rect 17635 20757 17647 20791
rect 17589 20751 17647 20757
rect 17678 20748 17684 20800
rect 17736 20788 17742 20800
rect 18340 20797 18368 20828
rect 19061 20825 19073 20859
rect 19107 20856 19119 20859
rect 19613 20859 19671 20865
rect 19613 20856 19625 20859
rect 19107 20828 19625 20856
rect 19107 20825 19119 20828
rect 19061 20819 19119 20825
rect 19613 20825 19625 20828
rect 19659 20825 19671 20859
rect 19613 20819 19671 20825
rect 19702 20816 19708 20868
rect 19760 20856 19766 20868
rect 20456 20856 20484 20887
rect 20990 20884 20996 20896
rect 21048 20884 21054 20936
rect 21177 20927 21235 20933
rect 21177 20893 21189 20927
rect 21223 20924 21235 20927
rect 22278 20924 22284 20936
rect 21223 20896 22284 20924
rect 21223 20893 21235 20896
rect 21177 20887 21235 20893
rect 22278 20884 22284 20896
rect 22336 20884 22342 20936
rect 22465 20927 22523 20933
rect 22465 20893 22477 20927
rect 22511 20893 22523 20927
rect 22465 20887 22523 20893
rect 19760 20828 20484 20856
rect 22480 20856 22508 20887
rect 22554 20884 22560 20936
rect 22612 20924 22618 20936
rect 22833 20927 22891 20933
rect 22833 20924 22845 20927
rect 22612 20896 22845 20924
rect 22612 20884 22618 20896
rect 22833 20893 22845 20896
rect 22879 20893 22891 20927
rect 22833 20887 22891 20893
rect 23106 20856 23112 20868
rect 22480 20828 23112 20856
rect 19760 20816 19766 20828
rect 23106 20816 23112 20828
rect 23164 20816 23170 20868
rect 18325 20791 18383 20797
rect 17736 20760 17781 20788
rect 17736 20748 17742 20760
rect 18325 20757 18337 20791
rect 18371 20757 18383 20791
rect 18325 20751 18383 20757
rect 19981 20791 20039 20797
rect 19981 20757 19993 20791
rect 20027 20788 20039 20791
rect 20714 20788 20720 20800
rect 20027 20760 20720 20788
rect 20027 20757 20039 20760
rect 19981 20751 20039 20757
rect 20714 20748 20720 20760
rect 20772 20748 20778 20800
rect 20806 20748 20812 20800
rect 20864 20788 20870 20800
rect 20907 20791 20965 20797
rect 20907 20788 20919 20791
rect 20864 20760 20919 20788
rect 20864 20748 20870 20760
rect 20907 20757 20919 20760
rect 20953 20788 20965 20791
rect 21542 20788 21548 20800
rect 20953 20760 21548 20788
rect 20953 20757 20965 20760
rect 20907 20751 20965 20757
rect 21542 20748 21548 20760
rect 21600 20748 21606 20800
rect 21634 20748 21640 20800
rect 21692 20788 21698 20800
rect 22281 20791 22339 20797
rect 22281 20788 22293 20791
rect 21692 20760 22293 20788
rect 21692 20748 21698 20760
rect 22281 20757 22293 20760
rect 22327 20757 22339 20791
rect 23014 20788 23020 20800
rect 22975 20760 23020 20788
rect 22281 20751 22339 20757
rect 23014 20748 23020 20760
rect 23072 20748 23078 20800
rect 1104 20698 23460 20720
rect 1104 20646 6548 20698
rect 6600 20646 6612 20698
rect 6664 20646 6676 20698
rect 6728 20646 6740 20698
rect 6792 20646 6804 20698
rect 6856 20646 12146 20698
rect 12198 20646 12210 20698
rect 12262 20646 12274 20698
rect 12326 20646 12338 20698
rect 12390 20646 12402 20698
rect 12454 20646 17744 20698
rect 17796 20646 17808 20698
rect 17860 20646 17872 20698
rect 17924 20646 17936 20698
rect 17988 20646 18000 20698
rect 18052 20646 23460 20698
rect 1104 20624 23460 20646
rect 4709 20587 4767 20593
rect 4709 20553 4721 20587
rect 4755 20584 4767 20587
rect 4982 20584 4988 20596
rect 4755 20556 4988 20584
rect 4755 20553 4767 20556
rect 4709 20547 4767 20553
rect 4982 20544 4988 20556
rect 5040 20544 5046 20596
rect 5350 20544 5356 20596
rect 5408 20584 5414 20596
rect 7377 20587 7435 20593
rect 5408 20556 7328 20584
rect 5408 20544 5414 20556
rect 6365 20519 6423 20525
rect 6365 20516 6377 20519
rect 4448 20488 6377 20516
rect 4448 20457 4476 20488
rect 6365 20485 6377 20488
rect 6411 20485 6423 20519
rect 6365 20479 6423 20485
rect 6549 20519 6607 20525
rect 6549 20485 6561 20519
rect 6595 20516 6607 20519
rect 7190 20516 7196 20528
rect 6595 20488 7196 20516
rect 6595 20485 6607 20488
rect 6549 20479 6607 20485
rect 7190 20476 7196 20488
rect 7248 20476 7254 20528
rect 4433 20451 4491 20457
rect 4433 20417 4445 20451
rect 4479 20417 4491 20451
rect 4433 20411 4491 20417
rect 4706 20408 4712 20460
rect 4764 20448 4770 20460
rect 5914 20451 5972 20457
rect 5914 20448 5926 20451
rect 4764 20420 5926 20448
rect 4764 20408 4770 20420
rect 5914 20417 5926 20420
rect 5960 20417 5972 20451
rect 5914 20411 5972 20417
rect 6733 20451 6791 20457
rect 6733 20417 6745 20451
rect 6779 20448 6791 20451
rect 7098 20448 7104 20460
rect 6779 20420 7104 20448
rect 6779 20417 6791 20420
rect 6733 20411 6791 20417
rect 7098 20408 7104 20420
rect 7156 20408 7162 20460
rect 6178 20380 6184 20392
rect 6139 20352 6184 20380
rect 6178 20340 6184 20352
rect 6236 20340 6242 20392
rect 7300 20380 7328 20556
rect 7377 20553 7389 20587
rect 7423 20584 7435 20587
rect 7466 20584 7472 20596
rect 7423 20556 7472 20584
rect 7423 20553 7435 20556
rect 7377 20547 7435 20553
rect 7466 20544 7472 20556
rect 7524 20544 7530 20596
rect 8478 20584 8484 20596
rect 7760 20556 8484 20584
rect 7760 20460 7788 20556
rect 8478 20544 8484 20556
rect 8536 20544 8542 20596
rect 8671 20587 8729 20593
rect 8671 20553 8683 20587
rect 8717 20584 8729 20587
rect 9766 20584 9772 20596
rect 8717 20556 9772 20584
rect 8717 20553 8729 20556
rect 8671 20547 8729 20553
rect 9766 20544 9772 20556
rect 9824 20544 9830 20596
rect 9950 20544 9956 20596
rect 10008 20584 10014 20596
rect 10045 20587 10103 20593
rect 10045 20584 10057 20587
rect 10008 20556 10057 20584
rect 10008 20544 10014 20556
rect 10045 20553 10057 20556
rect 10091 20553 10103 20587
rect 10686 20584 10692 20596
rect 10647 20556 10692 20584
rect 10045 20547 10103 20553
rect 10686 20544 10692 20556
rect 10744 20544 10750 20596
rect 11054 20544 11060 20596
rect 11112 20584 11118 20596
rect 11149 20587 11207 20593
rect 11149 20584 11161 20587
rect 11112 20556 11161 20584
rect 11112 20544 11118 20556
rect 11149 20553 11161 20556
rect 11195 20553 11207 20587
rect 11149 20547 11207 20553
rect 11977 20587 12035 20593
rect 11977 20553 11989 20587
rect 12023 20584 12035 20587
rect 12526 20584 12532 20596
rect 12023 20556 12532 20584
rect 12023 20553 12035 20556
rect 11977 20547 12035 20553
rect 12526 20544 12532 20556
rect 12584 20544 12590 20596
rect 13633 20587 13691 20593
rect 13633 20553 13645 20587
rect 13679 20553 13691 20587
rect 13633 20547 13691 20553
rect 13725 20587 13783 20593
rect 13725 20553 13737 20587
rect 13771 20584 13783 20587
rect 13906 20584 13912 20596
rect 13771 20556 13912 20584
rect 13771 20553 13783 20556
rect 13725 20547 13783 20553
rect 12894 20516 12900 20528
rect 11532 20488 12900 20516
rect 7742 20448 7748 20460
rect 7703 20420 7748 20448
rect 7742 20408 7748 20420
rect 7800 20408 7806 20460
rect 7926 20408 7932 20460
rect 7984 20448 7990 20460
rect 8938 20448 8944 20460
rect 7984 20420 8524 20448
rect 8899 20420 8944 20448
rect 7984 20408 7990 20420
rect 7837 20383 7895 20389
rect 7837 20380 7849 20383
rect 7300 20352 7849 20380
rect 7837 20349 7849 20352
rect 7883 20349 7895 20383
rect 8018 20380 8024 20392
rect 7979 20352 8024 20380
rect 7837 20343 7895 20349
rect 1578 20272 1584 20324
rect 1636 20312 1642 20324
rect 4614 20312 4620 20324
rect 1636 20284 4620 20312
rect 1636 20272 1642 20284
rect 4614 20272 4620 20284
rect 4672 20272 4678 20324
rect 2130 20204 2136 20256
rect 2188 20244 2194 20256
rect 4249 20247 4307 20253
rect 4249 20244 4261 20247
rect 2188 20216 4261 20244
rect 2188 20204 2194 20216
rect 4249 20213 4261 20216
rect 4295 20213 4307 20247
rect 4798 20244 4804 20256
rect 4759 20216 4804 20244
rect 4249 20207 4307 20213
rect 4798 20204 4804 20216
rect 4856 20204 4862 20256
rect 6822 20204 6828 20256
rect 6880 20244 6886 20256
rect 6917 20247 6975 20253
rect 6917 20244 6929 20247
rect 6880 20216 6929 20244
rect 6880 20204 6886 20216
rect 6917 20213 6929 20216
rect 6963 20244 6975 20247
rect 7101 20247 7159 20253
rect 7101 20244 7113 20247
rect 6963 20216 7113 20244
rect 6963 20213 6975 20216
rect 6917 20207 6975 20213
rect 7101 20213 7113 20216
rect 7147 20213 7159 20247
rect 7852 20244 7880 20343
rect 8018 20340 8024 20352
rect 8076 20340 8082 20392
rect 8205 20383 8263 20389
rect 8205 20349 8217 20383
rect 8251 20380 8263 20383
rect 8386 20380 8392 20392
rect 8251 20352 8392 20380
rect 8251 20349 8263 20352
rect 8205 20343 8263 20349
rect 8386 20340 8392 20352
rect 8444 20340 8450 20392
rect 8496 20380 8524 20420
rect 8938 20408 8944 20420
rect 8996 20408 9002 20460
rect 10594 20448 10600 20460
rect 10555 20420 10600 20448
rect 10594 20408 10600 20420
rect 10652 20408 10658 20460
rect 11532 20457 11560 20488
rect 12894 20476 12900 20488
rect 12952 20476 12958 20528
rect 13648 20516 13676 20547
rect 13906 20544 13912 20556
rect 13964 20544 13970 20596
rect 14185 20587 14243 20593
rect 14185 20553 14197 20587
rect 14231 20584 14243 20587
rect 14642 20584 14648 20596
rect 14231 20556 14648 20584
rect 14231 20553 14243 20556
rect 14185 20547 14243 20553
rect 14642 20544 14648 20556
rect 14700 20544 14706 20596
rect 14737 20587 14795 20593
rect 14737 20553 14749 20587
rect 14783 20584 14795 20587
rect 15286 20584 15292 20596
rect 14783 20556 15292 20584
rect 14783 20553 14795 20556
rect 14737 20547 14795 20553
rect 15286 20544 15292 20556
rect 15344 20544 15350 20596
rect 15565 20587 15623 20593
rect 15565 20553 15577 20587
rect 15611 20584 15623 20587
rect 15654 20584 15660 20596
rect 15611 20556 15660 20584
rect 15611 20553 15623 20556
rect 15565 20547 15623 20553
rect 15654 20544 15660 20556
rect 15712 20544 15718 20596
rect 15933 20587 15991 20593
rect 15933 20553 15945 20587
rect 15979 20584 15991 20587
rect 16758 20584 16764 20596
rect 15979 20556 16764 20584
rect 15979 20553 15991 20556
rect 15933 20547 15991 20553
rect 16758 20544 16764 20556
rect 16816 20544 16822 20596
rect 17494 20544 17500 20596
rect 17552 20584 17558 20596
rect 17589 20587 17647 20593
rect 17589 20584 17601 20587
rect 17552 20556 17601 20584
rect 17552 20544 17558 20556
rect 17589 20553 17601 20556
rect 17635 20553 17647 20587
rect 17589 20547 17647 20553
rect 18138 20544 18144 20596
rect 18196 20584 18202 20596
rect 18331 20587 18389 20593
rect 18331 20584 18343 20587
rect 18196 20556 18343 20584
rect 18196 20544 18202 20556
rect 18331 20553 18343 20556
rect 18377 20553 18389 20587
rect 18331 20547 18389 20553
rect 19886 20544 19892 20596
rect 19944 20584 19950 20596
rect 19981 20587 20039 20593
rect 19981 20584 19993 20587
rect 19944 20556 19993 20584
rect 19944 20544 19950 20556
rect 19981 20553 19993 20556
rect 20027 20553 20039 20587
rect 19981 20547 20039 20553
rect 20625 20587 20683 20593
rect 20625 20553 20637 20587
rect 20671 20584 20683 20587
rect 20714 20584 20720 20596
rect 20671 20556 20720 20584
rect 20671 20553 20683 20556
rect 20625 20547 20683 20553
rect 20714 20544 20720 20556
rect 20772 20544 20778 20596
rect 20898 20544 20904 20596
rect 20956 20584 20962 20596
rect 21085 20587 21143 20593
rect 21085 20584 21097 20587
rect 20956 20556 21097 20584
rect 20956 20544 20962 20556
rect 21085 20553 21097 20556
rect 21131 20553 21143 20587
rect 21085 20547 21143 20553
rect 21269 20587 21327 20593
rect 21269 20553 21281 20587
rect 21315 20584 21327 20587
rect 22002 20584 22008 20596
rect 21315 20556 22008 20584
rect 21315 20553 21327 20556
rect 21269 20547 21327 20553
rect 22002 20544 22008 20556
rect 22060 20544 22066 20596
rect 14274 20516 14280 20528
rect 13648 20488 14280 20516
rect 14274 20476 14280 20488
rect 14332 20476 14338 20528
rect 16206 20476 16212 20528
rect 16264 20516 16270 20528
rect 20732 20516 20760 20544
rect 22189 20519 22247 20525
rect 22189 20516 22201 20519
rect 16264 20488 17448 20516
rect 20732 20488 22201 20516
rect 16264 20476 16270 20488
rect 11517 20451 11575 20457
rect 11517 20417 11529 20451
rect 11563 20417 11575 20451
rect 11790 20448 11796 20460
rect 11751 20420 11796 20448
rect 11517 20411 11575 20417
rect 11790 20408 11796 20420
rect 11848 20408 11854 20460
rect 12434 20408 12440 20460
rect 12492 20448 12498 20460
rect 12492 20420 12537 20448
rect 12492 20408 12498 20420
rect 13078 20408 13084 20460
rect 13136 20448 13142 20460
rect 13265 20451 13323 20457
rect 13265 20448 13277 20451
rect 13136 20420 13277 20448
rect 13136 20408 13142 20420
rect 13265 20417 13277 20420
rect 13311 20417 13323 20451
rect 13265 20411 13323 20417
rect 14093 20451 14151 20457
rect 14093 20417 14105 20451
rect 14139 20448 14151 20451
rect 14366 20448 14372 20460
rect 14139 20420 14372 20448
rect 14139 20417 14151 20420
rect 14093 20411 14151 20417
rect 14366 20408 14372 20420
rect 14424 20408 14430 20460
rect 15105 20451 15163 20457
rect 15105 20417 15117 20451
rect 15151 20448 15163 20451
rect 15838 20448 15844 20460
rect 15151 20420 15844 20448
rect 15151 20417 15163 20420
rect 15105 20411 15163 20417
rect 15838 20408 15844 20420
rect 15896 20408 15902 20460
rect 16025 20451 16083 20457
rect 16025 20417 16037 20451
rect 16071 20448 16083 20451
rect 16071 20420 16528 20448
rect 16071 20417 16083 20420
rect 16025 20411 16083 20417
rect 8668 20385 8726 20391
rect 8668 20382 8680 20385
rect 8588 20380 8680 20382
rect 8496 20354 8680 20380
rect 8496 20352 8616 20354
rect 8668 20351 8680 20354
rect 8714 20351 8726 20385
rect 8668 20345 8726 20351
rect 10778 20340 10784 20392
rect 10836 20380 10842 20392
rect 10836 20352 10881 20380
rect 10836 20340 10842 20352
rect 12250 20340 12256 20392
rect 12308 20380 12314 20392
rect 12529 20383 12587 20389
rect 12529 20380 12541 20383
rect 12308 20352 12541 20380
rect 12308 20340 12314 20352
rect 12529 20349 12541 20352
rect 12575 20349 12587 20383
rect 12529 20343 12587 20349
rect 12713 20383 12771 20389
rect 12713 20349 12725 20383
rect 12759 20380 12771 20383
rect 12989 20383 13047 20389
rect 12989 20380 13001 20383
rect 12759 20352 13001 20380
rect 12759 20349 12771 20352
rect 12713 20343 12771 20349
rect 12989 20349 13001 20352
rect 13035 20349 13047 20383
rect 13170 20380 13176 20392
rect 13131 20352 13176 20380
rect 12989 20343 13047 20349
rect 11701 20315 11759 20321
rect 11701 20281 11713 20315
rect 11747 20312 11759 20315
rect 13004 20312 13032 20343
rect 13170 20340 13176 20352
rect 13228 20340 13234 20392
rect 14277 20383 14335 20389
rect 14277 20349 14289 20383
rect 14323 20349 14335 20383
rect 15194 20380 15200 20392
rect 15155 20352 15200 20380
rect 14277 20343 14335 20349
rect 13630 20312 13636 20324
rect 11747 20284 12434 20312
rect 13004 20284 13636 20312
rect 11747 20281 11759 20284
rect 11701 20275 11759 20281
rect 8754 20244 8760 20256
rect 7852 20216 8760 20244
rect 7101 20207 7159 20213
rect 8754 20204 8760 20216
rect 8812 20204 8818 20256
rect 8846 20204 8852 20256
rect 8904 20244 8910 20256
rect 10229 20247 10287 20253
rect 10229 20244 10241 20247
rect 8904 20216 10241 20244
rect 8904 20204 8910 20216
rect 10229 20213 10241 20216
rect 10275 20213 10287 20247
rect 10229 20207 10287 20213
rect 11514 20204 11520 20256
rect 11572 20244 11578 20256
rect 12069 20247 12127 20253
rect 12069 20244 12081 20247
rect 11572 20216 12081 20244
rect 11572 20204 11578 20216
rect 12069 20213 12081 20216
rect 12115 20213 12127 20247
rect 12406 20244 12434 20284
rect 13630 20272 13636 20284
rect 13688 20312 13694 20324
rect 14292 20312 14320 20343
rect 15194 20340 15200 20352
rect 15252 20340 15258 20392
rect 15289 20383 15347 20389
rect 15289 20349 15301 20383
rect 15335 20349 15347 20383
rect 15289 20343 15347 20349
rect 15304 20312 15332 20343
rect 15378 20340 15384 20392
rect 15436 20380 15442 20392
rect 16117 20383 16175 20389
rect 16117 20380 16129 20383
rect 15436 20352 16129 20380
rect 15436 20340 15442 20352
rect 16117 20349 16129 20352
rect 16163 20349 16175 20383
rect 16500 20380 16528 20420
rect 16574 20408 16580 20460
rect 16632 20448 16638 20460
rect 17037 20451 17095 20457
rect 17037 20448 17049 20451
rect 16632 20420 17049 20448
rect 16632 20408 16638 20420
rect 17037 20417 17049 20420
rect 17083 20417 17095 20451
rect 17420 20448 17448 20488
rect 22189 20485 22201 20488
rect 22235 20485 22247 20519
rect 22189 20479 22247 20485
rect 18601 20451 18659 20457
rect 18601 20448 18613 20451
rect 17420 20420 18613 20448
rect 17037 20411 17095 20417
rect 18601 20417 18613 20420
rect 18647 20417 18659 20451
rect 18601 20411 18659 20417
rect 19978 20408 19984 20460
rect 20036 20448 20042 20460
rect 20073 20451 20131 20457
rect 20073 20448 20085 20451
rect 20036 20420 20085 20448
rect 20036 20408 20042 20420
rect 20073 20417 20085 20420
rect 20119 20417 20131 20451
rect 20073 20411 20131 20417
rect 20717 20451 20775 20457
rect 20717 20417 20729 20451
rect 20763 20417 20775 20451
rect 21358 20448 21364 20460
rect 21319 20420 21364 20448
rect 20717 20411 20775 20417
rect 16666 20380 16672 20392
rect 16500 20352 16672 20380
rect 16117 20343 16175 20349
rect 16666 20340 16672 20352
rect 16724 20340 16730 20392
rect 16850 20340 16856 20392
rect 16908 20380 16914 20392
rect 17129 20383 17187 20389
rect 17129 20380 17141 20383
rect 16908 20352 17141 20380
rect 16908 20340 16914 20352
rect 17129 20349 17141 20352
rect 17175 20349 17187 20383
rect 17129 20343 17187 20349
rect 17218 20340 17224 20392
rect 17276 20380 17282 20392
rect 17276 20352 17321 20380
rect 17276 20340 17282 20352
rect 17402 20340 17408 20392
rect 17460 20380 17466 20392
rect 17865 20383 17923 20389
rect 17865 20380 17877 20383
rect 17460 20352 17877 20380
rect 17460 20340 17466 20352
rect 17865 20349 17877 20352
rect 17911 20349 17923 20383
rect 17865 20343 17923 20349
rect 18322 20340 18328 20392
rect 18380 20380 18386 20392
rect 18380 20352 18425 20380
rect 18380 20340 18386 20352
rect 18506 20340 18512 20392
rect 18564 20380 18570 20392
rect 20441 20383 20499 20389
rect 20441 20380 20453 20383
rect 18564 20352 20453 20380
rect 18564 20340 18570 20352
rect 20441 20349 20453 20352
rect 20487 20349 20499 20383
rect 20441 20343 20499 20349
rect 13688 20284 14320 20312
rect 14384 20284 15332 20312
rect 13688 20272 13694 20284
rect 12986 20244 12992 20256
rect 12406 20216 12992 20244
rect 12069 20207 12127 20213
rect 12986 20204 12992 20216
rect 13044 20204 13050 20256
rect 13906 20204 13912 20256
rect 13964 20244 13970 20256
rect 14384 20244 14412 20284
rect 16298 20272 16304 20324
rect 16356 20312 16362 20324
rect 20732 20312 20760 20411
rect 21358 20408 21364 20420
rect 21416 20408 21422 20460
rect 22830 20448 22836 20460
rect 22791 20420 22836 20448
rect 22830 20408 22836 20420
rect 22888 20408 22894 20460
rect 22278 20380 22284 20392
rect 22239 20352 22284 20380
rect 22278 20340 22284 20352
rect 22336 20340 22342 20392
rect 22465 20383 22523 20389
rect 22465 20349 22477 20383
rect 22511 20380 22523 20383
rect 22554 20380 22560 20392
rect 22511 20352 22560 20380
rect 22511 20349 22523 20352
rect 22465 20343 22523 20349
rect 22554 20340 22560 20352
rect 22612 20340 22618 20392
rect 21450 20312 21456 20324
rect 16356 20284 16712 20312
rect 16356 20272 16362 20284
rect 13964 20216 14412 20244
rect 13964 20204 13970 20216
rect 14458 20204 14464 20256
rect 14516 20244 14522 20256
rect 14553 20247 14611 20253
rect 14553 20244 14565 20247
rect 14516 20216 14565 20244
rect 14516 20204 14522 20216
rect 14553 20213 14565 20216
rect 14599 20213 14611 20247
rect 16390 20244 16396 20256
rect 16351 20216 16396 20244
rect 14553 20207 14611 20213
rect 16390 20204 16396 20216
rect 16448 20204 16454 20256
rect 16684 20253 16712 20284
rect 19720 20284 21456 20312
rect 16669 20247 16727 20253
rect 16669 20213 16681 20247
rect 16715 20213 16727 20247
rect 16669 20207 16727 20213
rect 18138 20204 18144 20256
rect 18196 20244 18202 20256
rect 19720 20253 19748 20284
rect 21450 20272 21456 20284
rect 21508 20272 21514 20324
rect 21545 20315 21603 20321
rect 21545 20281 21557 20315
rect 21591 20312 21603 20315
rect 23474 20312 23480 20324
rect 21591 20284 23480 20312
rect 21591 20281 21603 20284
rect 21545 20275 21603 20281
rect 23474 20272 23480 20284
rect 23532 20272 23538 20324
rect 19705 20247 19763 20253
rect 19705 20244 19717 20247
rect 18196 20216 19717 20244
rect 18196 20204 18202 20216
rect 19705 20213 19717 20216
rect 19751 20213 19763 20247
rect 19705 20207 19763 20213
rect 20257 20247 20315 20253
rect 20257 20213 20269 20247
rect 20303 20244 20315 20247
rect 21082 20244 21088 20256
rect 20303 20216 21088 20244
rect 20303 20213 20315 20216
rect 20257 20207 20315 20213
rect 21082 20204 21088 20216
rect 21140 20204 21146 20256
rect 21818 20244 21824 20256
rect 21779 20216 21824 20244
rect 21818 20204 21824 20216
rect 21876 20204 21882 20256
rect 22646 20244 22652 20256
rect 22607 20216 22652 20244
rect 22646 20204 22652 20216
rect 22704 20204 22710 20256
rect 23014 20244 23020 20256
rect 22975 20216 23020 20244
rect 23014 20204 23020 20216
rect 23072 20204 23078 20256
rect 1104 20154 23460 20176
rect 1104 20102 3749 20154
rect 3801 20102 3813 20154
rect 3865 20102 3877 20154
rect 3929 20102 3941 20154
rect 3993 20102 4005 20154
rect 4057 20102 9347 20154
rect 9399 20102 9411 20154
rect 9463 20102 9475 20154
rect 9527 20102 9539 20154
rect 9591 20102 9603 20154
rect 9655 20102 14945 20154
rect 14997 20102 15009 20154
rect 15061 20102 15073 20154
rect 15125 20102 15137 20154
rect 15189 20102 15201 20154
rect 15253 20102 20543 20154
rect 20595 20102 20607 20154
rect 20659 20102 20671 20154
rect 20723 20102 20735 20154
rect 20787 20102 20799 20154
rect 20851 20102 23460 20154
rect 1104 20080 23460 20102
rect 3237 20043 3295 20049
rect 3237 20009 3249 20043
rect 3283 20040 3295 20043
rect 3283 20012 9168 20040
rect 3283 20009 3295 20012
rect 3237 20003 3295 20009
rect 3142 19932 3148 19984
rect 3200 19972 3206 19984
rect 4065 19975 4123 19981
rect 4065 19972 4077 19975
rect 3200 19944 4077 19972
rect 3200 19932 3206 19944
rect 4065 19941 4077 19944
rect 4111 19941 4123 19975
rect 4065 19935 4123 19941
rect 8386 19932 8392 19984
rect 8444 19972 8450 19984
rect 9140 19972 9168 20012
rect 9214 20000 9220 20052
rect 9272 20040 9278 20052
rect 9861 20043 9919 20049
rect 9861 20040 9873 20043
rect 9272 20012 9873 20040
rect 9272 20000 9278 20012
rect 9861 20009 9873 20012
rect 9907 20009 9919 20043
rect 10870 20040 10876 20052
rect 10831 20012 10876 20040
rect 9861 20003 9919 20009
rect 10870 20000 10876 20012
rect 10928 20000 10934 20052
rect 11057 20043 11115 20049
rect 11057 20009 11069 20043
rect 11103 20040 11115 20043
rect 11146 20040 11152 20052
rect 11103 20012 11152 20040
rect 11103 20009 11115 20012
rect 11057 20003 11115 20009
rect 11146 20000 11152 20012
rect 11204 20000 11210 20052
rect 12250 20040 12256 20052
rect 12211 20012 12256 20040
rect 12250 20000 12256 20012
rect 12308 20000 12314 20052
rect 13998 20040 14004 20052
rect 13188 20012 14004 20040
rect 10594 19972 10600 19984
rect 8444 19944 8616 19972
rect 9140 19944 10600 19972
rect 8444 19932 8450 19944
rect 2222 19796 2228 19848
rect 2280 19836 2286 19848
rect 3053 19839 3111 19845
rect 3053 19836 3065 19839
rect 2280 19808 3065 19836
rect 2280 19796 2286 19808
rect 3053 19805 3065 19808
rect 3099 19805 3111 19839
rect 3510 19836 3516 19848
rect 3471 19808 3516 19836
rect 3053 19799 3111 19805
rect 3510 19796 3516 19808
rect 3568 19796 3574 19848
rect 5445 19839 5503 19845
rect 5445 19805 5457 19839
rect 5491 19836 5503 19839
rect 6178 19836 6184 19848
rect 5491 19808 6184 19836
rect 5491 19805 5503 19808
rect 5445 19799 5503 19805
rect 6178 19796 6184 19808
rect 6236 19836 6242 19848
rect 6822 19836 6828 19848
rect 6236 19808 6828 19836
rect 6236 19796 6242 19808
rect 6822 19796 6828 19808
rect 6880 19836 6886 19848
rect 6917 19839 6975 19845
rect 6917 19836 6929 19839
rect 6880 19808 6929 19836
rect 6880 19796 6886 19808
rect 6917 19805 6929 19808
rect 6963 19805 6975 19839
rect 6917 19799 6975 19805
rect 7190 19796 7196 19848
rect 7248 19836 7254 19848
rect 8122 19839 8180 19845
rect 8122 19836 8134 19839
rect 7248 19808 8134 19836
rect 7248 19796 7254 19808
rect 8122 19805 8134 19808
rect 8168 19805 8180 19839
rect 8122 19799 8180 19805
rect 8389 19839 8447 19845
rect 8389 19805 8401 19839
rect 8435 19805 8447 19839
rect 8389 19799 8447 19805
rect 2746 19740 3372 19768
rect 2498 19660 2504 19712
rect 2556 19700 2562 19712
rect 2746 19700 2774 19740
rect 3344 19709 3372 19740
rect 5166 19728 5172 19780
rect 5224 19777 5230 19780
rect 5224 19768 5236 19777
rect 5224 19740 5580 19768
rect 5224 19731 5236 19740
rect 5224 19728 5230 19731
rect 2556 19672 2774 19700
rect 3329 19703 3387 19709
rect 2556 19660 2562 19672
rect 3329 19669 3341 19703
rect 3375 19669 3387 19703
rect 3970 19700 3976 19712
rect 3931 19672 3976 19700
rect 3329 19663 3387 19669
rect 3970 19660 3976 19672
rect 4028 19660 4034 19712
rect 5552 19709 5580 19740
rect 5902 19728 5908 19780
rect 5960 19768 5966 19780
rect 6672 19771 6730 19777
rect 6672 19768 6684 19771
rect 5960 19740 6684 19768
rect 5960 19728 5966 19740
rect 6672 19737 6684 19740
rect 6718 19768 6730 19771
rect 7282 19768 7288 19780
rect 6718 19740 7288 19768
rect 6718 19737 6730 19740
rect 6672 19731 6730 19737
rect 7282 19728 7288 19740
rect 7340 19728 7346 19780
rect 5537 19703 5595 19709
rect 5537 19669 5549 19703
rect 5583 19669 5595 19703
rect 5537 19663 5595 19669
rect 5626 19660 5632 19712
rect 5684 19700 5690 19712
rect 6454 19700 6460 19712
rect 5684 19672 6460 19700
rect 5684 19660 5690 19672
rect 6454 19660 6460 19672
rect 6512 19700 6518 19712
rect 7009 19703 7067 19709
rect 7009 19700 7021 19703
rect 6512 19672 7021 19700
rect 6512 19660 6518 19672
rect 7009 19669 7021 19672
rect 7055 19669 7067 19703
rect 7009 19663 7067 19669
rect 8294 19660 8300 19712
rect 8352 19700 8358 19712
rect 8404 19700 8432 19799
rect 8481 19703 8539 19709
rect 8481 19700 8493 19703
rect 8352 19672 8493 19700
rect 8352 19660 8358 19672
rect 8481 19669 8493 19672
rect 8527 19669 8539 19703
rect 8588 19700 8616 19944
rect 10594 19932 10600 19944
rect 10652 19932 10658 19984
rect 10689 19975 10747 19981
rect 10689 19941 10701 19975
rect 10735 19972 10747 19975
rect 11238 19972 11244 19984
rect 10735 19944 11244 19972
rect 10735 19941 10747 19944
rect 10689 19935 10747 19941
rect 11238 19932 11244 19944
rect 11296 19932 11302 19984
rect 11974 19972 11980 19984
rect 11935 19944 11980 19972
rect 11974 19932 11980 19944
rect 12032 19932 12038 19984
rect 12158 19972 12164 19984
rect 12119 19944 12164 19972
rect 12158 19932 12164 19944
rect 12216 19932 12222 19984
rect 9214 19904 9220 19916
rect 9175 19876 9220 19904
rect 9214 19864 9220 19876
rect 9272 19864 9278 19916
rect 11609 19907 11667 19913
rect 11609 19873 11621 19907
rect 11655 19904 11667 19907
rect 12618 19904 12624 19916
rect 11655 19876 12624 19904
rect 11655 19873 11667 19876
rect 11609 19867 11667 19873
rect 12618 19864 12624 19876
rect 12676 19864 12682 19916
rect 12894 19904 12900 19916
rect 12855 19876 12900 19904
rect 12894 19864 12900 19876
rect 12952 19864 12958 19916
rect 8846 19796 8852 19848
rect 8904 19836 8910 19848
rect 9401 19839 9459 19845
rect 9401 19836 9413 19839
rect 8904 19808 9413 19836
rect 8904 19796 8910 19808
rect 9401 19805 9413 19808
rect 9447 19836 9459 19839
rect 13188 19836 13216 20012
rect 13998 20000 14004 20012
rect 14056 20000 14062 20052
rect 14366 20040 14372 20052
rect 14327 20012 14372 20040
rect 14366 20000 14372 20012
rect 14424 20000 14430 20052
rect 15197 20043 15255 20049
rect 15197 20009 15209 20043
rect 15243 20040 15255 20043
rect 15286 20040 15292 20052
rect 15243 20012 15292 20040
rect 15243 20009 15255 20012
rect 15197 20003 15255 20009
rect 15286 20000 15292 20012
rect 15344 20000 15350 20052
rect 16850 20040 16856 20052
rect 16811 20012 16856 20040
rect 16850 20000 16856 20012
rect 16908 20000 16914 20052
rect 17586 20000 17592 20052
rect 17644 20040 17650 20052
rect 17681 20043 17739 20049
rect 17681 20040 17693 20043
rect 17644 20012 17693 20040
rect 17644 20000 17650 20012
rect 17681 20009 17693 20012
rect 17727 20009 17739 20043
rect 18782 20040 18788 20052
rect 18743 20012 18788 20040
rect 17681 20003 17739 20009
rect 18782 20000 18788 20012
rect 18840 20000 18846 20052
rect 20438 20040 20444 20052
rect 18892 20012 20444 20040
rect 13449 19975 13507 19981
rect 13449 19941 13461 19975
rect 13495 19972 13507 19975
rect 13722 19972 13728 19984
rect 13495 19944 13728 19972
rect 13495 19941 13507 19944
rect 13449 19935 13507 19941
rect 13722 19932 13728 19944
rect 13780 19932 13786 19984
rect 14090 19972 14096 19984
rect 13924 19944 14096 19972
rect 13924 19913 13952 19944
rect 14090 19932 14096 19944
rect 14148 19932 14154 19984
rect 14277 19975 14335 19981
rect 14277 19941 14289 19975
rect 14323 19972 14335 19975
rect 14550 19972 14556 19984
rect 14323 19944 14556 19972
rect 14323 19941 14335 19944
rect 14277 19935 14335 19941
rect 14550 19932 14556 19944
rect 14608 19932 14614 19984
rect 15470 19932 15476 19984
rect 15528 19972 15534 19984
rect 15528 19944 18276 19972
rect 15528 19932 15534 19944
rect 13909 19907 13967 19913
rect 13909 19873 13921 19907
rect 13955 19873 13967 19907
rect 13909 19867 13967 19873
rect 14921 19907 14979 19913
rect 14921 19873 14933 19907
rect 14967 19873 14979 19907
rect 14921 19867 14979 19873
rect 9447 19808 13216 19836
rect 13265 19839 13323 19845
rect 9447 19805 9459 19808
rect 9401 19799 9459 19805
rect 13265 19805 13277 19839
rect 13311 19836 13323 19839
rect 13354 19836 13360 19848
rect 13311 19808 13360 19836
rect 13311 19805 13323 19808
rect 13265 19799 13323 19805
rect 13354 19796 13360 19808
rect 13412 19796 13418 19848
rect 13538 19796 13544 19848
rect 13596 19836 13602 19848
rect 14093 19839 14151 19845
rect 13596 19808 14044 19836
rect 13596 19796 13602 19808
rect 9490 19768 9496 19780
rect 9451 19740 9496 19768
rect 9490 19728 9496 19740
rect 9548 19728 9554 19780
rect 11422 19768 11428 19780
rect 11383 19740 11428 19768
rect 11422 19728 11428 19740
rect 11480 19728 11486 19780
rect 14016 19768 14044 19808
rect 14093 19805 14105 19839
rect 14139 19836 14151 19839
rect 14458 19836 14464 19848
rect 14139 19808 14464 19836
rect 14139 19805 14151 19808
rect 14093 19799 14151 19805
rect 14458 19796 14464 19808
rect 14516 19796 14522 19848
rect 14550 19796 14556 19848
rect 14608 19836 14614 19848
rect 14936 19836 14964 19867
rect 15286 19864 15292 19916
rect 15344 19904 15350 19916
rect 15749 19907 15807 19913
rect 15749 19904 15761 19907
rect 15344 19876 15761 19904
rect 15344 19864 15350 19876
rect 15749 19873 15761 19876
rect 15795 19873 15807 19907
rect 16114 19904 16120 19916
rect 16075 19876 16120 19904
rect 15749 19867 15807 19873
rect 16114 19864 16120 19876
rect 16172 19864 16178 19916
rect 17494 19904 17500 19916
rect 16316 19876 17356 19904
rect 17455 19876 17500 19904
rect 14608 19808 14964 19836
rect 15565 19839 15623 19845
rect 14608 19796 14614 19808
rect 15565 19805 15577 19839
rect 15611 19836 15623 19839
rect 16316 19836 16344 19876
rect 15611 19808 16344 19836
rect 16393 19839 16451 19845
rect 15611 19805 15623 19808
rect 15565 19799 15623 19805
rect 16393 19805 16405 19839
rect 16439 19836 16451 19839
rect 16482 19836 16488 19848
rect 16439 19808 16488 19836
rect 16439 19805 16451 19808
rect 16393 19799 16451 19805
rect 16482 19796 16488 19808
rect 16540 19796 16546 19848
rect 17221 19839 17279 19845
rect 17221 19836 17233 19839
rect 16583 19808 17233 19836
rect 16301 19771 16359 19777
rect 16301 19768 16313 19771
rect 14016 19740 16313 19768
rect 16301 19737 16313 19740
rect 16347 19737 16359 19771
rect 16301 19731 16359 19737
rect 9858 19700 9864 19712
rect 8588 19672 9864 19700
rect 8481 19663 8539 19669
rect 9858 19660 9864 19672
rect 9916 19700 9922 19712
rect 10318 19700 10324 19712
rect 9916 19672 10324 19700
rect 9916 19660 9922 19672
rect 10318 19660 10324 19672
rect 10376 19660 10382 19712
rect 11146 19700 11152 19712
rect 11107 19672 11152 19700
rect 11146 19660 11152 19672
rect 11204 19660 11210 19712
rect 11514 19660 11520 19712
rect 11572 19700 11578 19712
rect 11701 19703 11759 19709
rect 11701 19700 11713 19703
rect 11572 19672 11713 19700
rect 11572 19660 11578 19672
rect 11701 19669 11713 19672
rect 11747 19700 11759 19703
rect 11882 19700 11888 19712
rect 11747 19672 11888 19700
rect 11747 19669 11759 19672
rect 11701 19663 11759 19669
rect 11882 19660 11888 19672
rect 11940 19660 11946 19712
rect 12618 19700 12624 19712
rect 12579 19672 12624 19700
rect 12618 19660 12624 19672
rect 12676 19660 12682 19712
rect 12710 19660 12716 19712
rect 12768 19700 12774 19712
rect 13081 19703 13139 19709
rect 12768 19672 12813 19700
rect 12768 19660 12774 19672
rect 13081 19669 13093 19703
rect 13127 19700 13139 19703
rect 13630 19700 13636 19712
rect 13127 19672 13636 19700
rect 13127 19669 13139 19672
rect 13081 19663 13139 19669
rect 13630 19660 13636 19672
rect 13688 19660 13694 19712
rect 14734 19700 14740 19712
rect 14695 19672 14740 19700
rect 14734 19660 14740 19672
rect 14792 19660 14798 19712
rect 14826 19660 14832 19712
rect 14884 19700 14890 19712
rect 14884 19672 14929 19700
rect 14884 19660 14890 19672
rect 15654 19660 15660 19712
rect 15712 19700 15718 19712
rect 15712 19672 15757 19700
rect 15712 19660 15718 19672
rect 16022 19660 16028 19712
rect 16080 19700 16086 19712
rect 16583 19700 16611 19808
rect 17221 19805 17233 19808
rect 17267 19805 17279 19839
rect 17328 19836 17356 19876
rect 17494 19864 17500 19876
rect 17552 19864 17558 19916
rect 18138 19904 18144 19916
rect 18099 19876 18144 19904
rect 18138 19864 18144 19876
rect 18196 19864 18202 19916
rect 18248 19913 18276 19944
rect 18233 19907 18291 19913
rect 18233 19873 18245 19907
rect 18279 19873 18291 19907
rect 18233 19867 18291 19873
rect 18046 19836 18052 19848
rect 17328 19808 17908 19836
rect 18007 19808 18052 19836
rect 17221 19799 17279 19805
rect 17034 19768 17040 19780
rect 16776 19740 17040 19768
rect 16776 19709 16804 19740
rect 17034 19728 17040 19740
rect 17092 19768 17098 19780
rect 17313 19771 17371 19777
rect 17313 19768 17325 19771
rect 17092 19740 17325 19768
rect 17092 19728 17098 19740
rect 17313 19737 17325 19740
rect 17359 19737 17371 19771
rect 17880 19768 17908 19808
rect 18046 19796 18052 19808
rect 18104 19836 18110 19848
rect 18322 19836 18328 19848
rect 18104 19808 18328 19836
rect 18104 19796 18110 19808
rect 18322 19796 18328 19808
rect 18380 19796 18386 19848
rect 18414 19796 18420 19848
rect 18472 19836 18478 19848
rect 18892 19845 18920 20012
rect 20438 20000 20444 20012
rect 20496 20000 20502 20052
rect 20530 20000 20536 20052
rect 20588 20040 20594 20052
rect 20809 20043 20867 20049
rect 20809 20040 20821 20043
rect 20588 20012 20821 20040
rect 20588 20000 20594 20012
rect 20809 20009 20821 20012
rect 20855 20040 20867 20043
rect 22002 20040 22008 20052
rect 20855 20012 22008 20040
rect 20855 20009 20867 20012
rect 20809 20003 20867 20009
rect 22002 20000 22008 20012
rect 22060 20000 22066 20052
rect 22278 20000 22284 20052
rect 22336 20040 22342 20052
rect 22741 20043 22799 20049
rect 22741 20040 22753 20043
rect 22336 20012 22753 20040
rect 22336 20000 22342 20012
rect 22741 20009 22753 20012
rect 22787 20009 22799 20043
rect 22741 20003 22799 20009
rect 21266 19864 21272 19916
rect 21324 19904 21330 19916
rect 21364 19907 21422 19913
rect 21364 19904 21376 19907
rect 21324 19876 21376 19904
rect 21324 19864 21330 19876
rect 21364 19873 21376 19876
rect 21410 19873 21422 19907
rect 21364 19867 21422 19873
rect 21450 19864 21456 19916
rect 21508 19904 21514 19916
rect 21637 19907 21695 19913
rect 21637 19904 21649 19907
rect 21508 19876 21649 19904
rect 21508 19864 21514 19876
rect 21637 19873 21649 19876
rect 21683 19873 21695 19907
rect 21637 19867 21695 19873
rect 18601 19839 18659 19845
rect 18601 19836 18613 19839
rect 18472 19808 18613 19836
rect 18472 19796 18478 19808
rect 18601 19805 18613 19808
rect 18647 19805 18659 19839
rect 18601 19799 18659 19805
rect 18877 19839 18935 19845
rect 18877 19805 18889 19839
rect 18923 19805 18935 19839
rect 19242 19836 19248 19848
rect 19155 19808 19248 19836
rect 18877 19799 18935 19805
rect 19242 19796 19248 19808
rect 19300 19836 19306 19848
rect 20530 19836 20536 19848
rect 19300 19808 20536 19836
rect 19300 19796 19306 19808
rect 20530 19796 20536 19808
rect 20588 19796 20594 19848
rect 20898 19836 20904 19848
rect 20859 19808 20904 19836
rect 20898 19796 20904 19808
rect 20956 19796 20962 19848
rect 21726 19836 21732 19848
rect 21008 19808 21732 19836
rect 18690 19768 18696 19780
rect 17880 19740 18696 19768
rect 17313 19731 17371 19737
rect 18690 19728 18696 19740
rect 18748 19728 18754 19780
rect 19512 19771 19570 19777
rect 19512 19737 19524 19771
rect 19558 19768 19570 19771
rect 20162 19768 20168 19780
rect 19558 19740 20168 19768
rect 19558 19737 19570 19740
rect 19512 19731 19570 19737
rect 16080 19672 16611 19700
rect 16761 19703 16819 19709
rect 16080 19660 16086 19672
rect 16761 19669 16773 19703
rect 16807 19669 16819 19703
rect 16761 19663 16819 19669
rect 19061 19703 19119 19709
rect 19061 19669 19073 19703
rect 19107 19700 19119 19703
rect 19150 19700 19156 19712
rect 19107 19672 19156 19700
rect 19107 19669 19119 19672
rect 19061 19663 19119 19669
rect 19150 19660 19156 19672
rect 19208 19660 19214 19712
rect 19426 19660 19432 19712
rect 19484 19700 19490 19712
rect 19527 19700 19555 19731
rect 20162 19728 20168 19740
rect 20220 19728 20226 19780
rect 19484 19672 19555 19700
rect 20625 19703 20683 19709
rect 19484 19660 19490 19672
rect 20625 19669 20637 19703
rect 20671 19700 20683 19703
rect 20714 19700 20720 19712
rect 20671 19672 20720 19700
rect 20671 19669 20683 19672
rect 20625 19663 20683 19669
rect 20714 19660 20720 19672
rect 20772 19700 20778 19712
rect 21008 19700 21036 19808
rect 21726 19796 21732 19808
rect 21784 19796 21790 19848
rect 22833 19839 22891 19845
rect 22833 19805 22845 19839
rect 22879 19836 22891 19839
rect 22922 19836 22928 19848
rect 22879 19808 22928 19836
rect 22879 19805 22891 19808
rect 22833 19799 22891 19805
rect 22922 19796 22928 19808
rect 22980 19796 22986 19848
rect 20772 19672 21036 19700
rect 21367 19703 21425 19709
rect 20772 19660 20778 19672
rect 21367 19669 21379 19703
rect 21413 19700 21425 19703
rect 21542 19700 21548 19712
rect 21413 19672 21548 19700
rect 21413 19669 21425 19672
rect 21367 19663 21425 19669
rect 21542 19660 21548 19672
rect 21600 19660 21606 19712
rect 23014 19700 23020 19712
rect 22975 19672 23020 19700
rect 23014 19660 23020 19672
rect 23072 19660 23078 19712
rect 1104 19610 23460 19632
rect 1104 19558 6548 19610
rect 6600 19558 6612 19610
rect 6664 19558 6676 19610
rect 6728 19558 6740 19610
rect 6792 19558 6804 19610
rect 6856 19558 12146 19610
rect 12198 19558 12210 19610
rect 12262 19558 12274 19610
rect 12326 19558 12338 19610
rect 12390 19558 12402 19610
rect 12454 19558 17744 19610
rect 17796 19558 17808 19610
rect 17860 19558 17872 19610
rect 17924 19558 17936 19610
rect 17988 19558 18000 19610
rect 18052 19558 23460 19610
rect 1104 19536 23460 19558
rect 2406 19456 2412 19508
rect 2464 19496 2470 19508
rect 2869 19499 2927 19505
rect 2869 19496 2881 19499
rect 2464 19468 2881 19496
rect 2464 19456 2470 19468
rect 2869 19465 2881 19468
rect 2915 19465 2927 19499
rect 2869 19459 2927 19465
rect 3970 19456 3976 19508
rect 4028 19496 4034 19508
rect 4065 19499 4123 19505
rect 4065 19496 4077 19499
rect 4028 19468 4077 19496
rect 4028 19456 4034 19468
rect 4065 19465 4077 19468
rect 4111 19465 4123 19499
rect 4430 19496 4436 19508
rect 4391 19468 4436 19496
rect 4065 19459 4123 19465
rect 4430 19456 4436 19468
rect 4488 19456 4494 19508
rect 4706 19496 4712 19508
rect 4619 19468 4712 19496
rect 4706 19456 4712 19468
rect 4764 19456 4770 19508
rect 7742 19496 7748 19508
rect 7703 19468 7748 19496
rect 7742 19456 7748 19468
rect 7800 19456 7806 19508
rect 8570 19456 8576 19508
rect 8628 19496 8634 19508
rect 10870 19496 10876 19508
rect 8628 19468 10876 19496
rect 8628 19456 8634 19468
rect 2133 19431 2191 19437
rect 2133 19397 2145 19431
rect 2179 19428 2191 19431
rect 2590 19428 2596 19440
rect 2179 19400 2596 19428
rect 2179 19397 2191 19400
rect 2133 19391 2191 19397
rect 2590 19388 2596 19400
rect 2648 19388 2654 19440
rect 3237 19431 3295 19437
rect 3237 19397 3249 19431
rect 3283 19428 3295 19431
rect 3418 19428 3424 19440
rect 3283 19400 3424 19428
rect 3283 19397 3295 19400
rect 3237 19391 3295 19397
rect 3418 19388 3424 19400
rect 3476 19388 3482 19440
rect 4724 19428 4752 19456
rect 4448 19400 4752 19428
rect 4448 19372 4476 19400
rect 2038 19320 2044 19372
rect 2096 19360 2102 19372
rect 2225 19363 2283 19369
rect 2225 19360 2237 19363
rect 2096 19332 2237 19360
rect 2096 19320 2102 19332
rect 2225 19329 2237 19332
rect 2271 19329 2283 19363
rect 2682 19360 2688 19372
rect 2225 19323 2283 19329
rect 2608 19332 2688 19360
rect 1949 19295 2007 19301
rect 1949 19261 1961 19295
rect 1995 19261 2007 19295
rect 1949 19255 2007 19261
rect 1964 19168 1992 19255
rect 2608 19233 2636 19332
rect 2682 19320 2688 19332
rect 2740 19320 2746 19372
rect 3326 19320 3332 19372
rect 3384 19360 3390 19372
rect 3384 19332 3429 19360
rect 3896 19332 4108 19360
rect 3384 19320 3390 19332
rect 2774 19252 2780 19304
rect 2832 19292 2838 19304
rect 3234 19292 3240 19304
rect 2832 19264 3240 19292
rect 2832 19252 2838 19264
rect 3234 19252 3240 19264
rect 3292 19292 3298 19304
rect 3896 19301 3924 19332
rect 3421 19295 3479 19301
rect 3421 19292 3433 19295
rect 3292 19264 3433 19292
rect 3292 19252 3298 19264
rect 3421 19261 3433 19264
rect 3467 19261 3479 19295
rect 3421 19255 3479 19261
rect 3881 19295 3939 19301
rect 3881 19261 3893 19295
rect 3927 19261 3939 19295
rect 3881 19255 3939 19261
rect 3973 19295 4031 19301
rect 3973 19261 3985 19295
rect 4019 19261 4031 19295
rect 4080 19292 4108 19332
rect 4430 19320 4436 19372
rect 4488 19320 4494 19372
rect 5534 19320 5540 19372
rect 5592 19360 5598 19372
rect 5822 19363 5880 19369
rect 5822 19360 5834 19363
rect 5592 19332 5834 19360
rect 5592 19320 5598 19332
rect 5822 19329 5834 19332
rect 5868 19329 5880 19363
rect 8846 19360 8852 19372
rect 8807 19332 8852 19360
rect 5822 19323 5880 19329
rect 8846 19320 8852 19332
rect 8904 19320 8910 19372
rect 9262 19363 9320 19369
rect 9262 19329 9274 19363
rect 9308 19360 9320 19363
rect 9766 19360 9772 19372
rect 9308 19332 9772 19360
rect 9308 19329 9320 19332
rect 9262 19323 9320 19329
rect 9766 19320 9772 19332
rect 9824 19320 9830 19372
rect 9858 19320 9864 19372
rect 9916 19320 9922 19372
rect 10805 19369 10833 19468
rect 10870 19456 10876 19468
rect 10928 19456 10934 19508
rect 11517 19499 11575 19505
rect 11517 19465 11529 19499
rect 11563 19496 11575 19499
rect 11606 19496 11612 19508
rect 11563 19468 11612 19496
rect 11563 19465 11575 19468
rect 11517 19459 11575 19465
rect 11606 19456 11612 19468
rect 11664 19496 11670 19508
rect 13449 19499 13507 19505
rect 13449 19496 13461 19499
rect 11664 19468 13461 19496
rect 11664 19456 11670 19468
rect 13449 19465 13461 19468
rect 13495 19465 13507 19499
rect 13449 19459 13507 19465
rect 14369 19499 14427 19505
rect 14369 19465 14381 19499
rect 14415 19496 14427 19499
rect 14734 19496 14740 19508
rect 14415 19468 14740 19496
rect 14415 19465 14427 19468
rect 14369 19459 14427 19465
rect 14734 19456 14740 19468
rect 14792 19456 14798 19508
rect 15838 19496 15844 19508
rect 15799 19468 15844 19496
rect 15838 19456 15844 19468
rect 15896 19456 15902 19508
rect 16209 19499 16267 19505
rect 16209 19465 16221 19499
rect 16255 19496 16267 19499
rect 16390 19496 16396 19508
rect 16255 19468 16396 19496
rect 16255 19465 16267 19468
rect 16209 19459 16267 19465
rect 12894 19388 12900 19440
rect 12952 19428 12958 19440
rect 12952 19400 13584 19428
rect 12952 19388 12958 19400
rect 10790 19363 10848 19369
rect 10790 19329 10802 19363
rect 10836 19329 10848 19363
rect 10790 19323 10848 19329
rect 12641 19363 12699 19369
rect 12641 19329 12653 19363
rect 12687 19360 12699 19363
rect 12986 19360 12992 19372
rect 12687 19332 12992 19360
rect 12687 19329 12699 19332
rect 12641 19323 12699 19329
rect 12986 19320 12992 19332
rect 13044 19320 13050 19372
rect 13262 19320 13268 19372
rect 13320 19360 13326 19372
rect 13357 19363 13415 19369
rect 13357 19360 13369 19363
rect 13320 19332 13369 19360
rect 13320 19320 13326 19332
rect 13357 19329 13369 19332
rect 13403 19329 13415 19363
rect 13357 19323 13415 19329
rect 5074 19292 5080 19304
rect 4080 19264 5080 19292
rect 3973 19255 4031 19261
rect 2593 19227 2651 19233
rect 2593 19193 2605 19227
rect 2639 19193 2651 19227
rect 2593 19187 2651 19193
rect 3602 19184 3608 19236
rect 3660 19224 3666 19236
rect 3988 19224 4016 19255
rect 5074 19252 5080 19264
rect 5132 19252 5138 19304
rect 6089 19295 6147 19301
rect 6089 19261 6101 19295
rect 6135 19292 6147 19295
rect 6135 19264 6224 19292
rect 6135 19261 6147 19264
rect 6089 19255 6147 19261
rect 3660 19196 4016 19224
rect 3660 19184 3666 19196
rect 6196 19168 6224 19264
rect 8110 19252 8116 19304
rect 8168 19292 8174 19304
rect 9079 19295 9137 19301
rect 9079 19292 9091 19295
rect 8168 19264 9091 19292
rect 8168 19252 8174 19264
rect 9079 19261 9091 19264
rect 9125 19261 9137 19295
rect 9079 19255 9137 19261
rect 9585 19295 9643 19301
rect 9585 19261 9597 19295
rect 9631 19292 9643 19295
rect 9876 19292 9904 19320
rect 13556 19304 13584 19400
rect 14826 19388 14832 19440
rect 14884 19428 14890 19440
rect 15482 19431 15540 19437
rect 15482 19428 15494 19431
rect 14884 19400 15494 19428
rect 14884 19388 14890 19400
rect 15482 19397 15494 19400
rect 15528 19397 15540 19431
rect 15482 19391 15540 19397
rect 14001 19363 14059 19369
rect 14001 19329 14013 19363
rect 14047 19360 14059 19363
rect 14550 19360 14556 19372
rect 14047 19332 14556 19360
rect 14047 19329 14059 19332
rect 14001 19323 14059 19329
rect 14550 19320 14556 19332
rect 14608 19320 14614 19372
rect 15746 19360 15752 19372
rect 15659 19332 15752 19360
rect 15746 19320 15752 19332
rect 15804 19360 15810 19372
rect 16224 19360 16252 19459
rect 16390 19456 16396 19468
rect 16448 19456 16454 19508
rect 16485 19499 16543 19505
rect 16485 19465 16497 19499
rect 16531 19496 16543 19499
rect 16574 19496 16580 19508
rect 16531 19468 16580 19496
rect 16531 19465 16543 19468
rect 16485 19459 16543 19465
rect 16574 19456 16580 19468
rect 16632 19456 16638 19508
rect 16666 19456 16672 19508
rect 16724 19496 16730 19508
rect 17034 19496 17040 19508
rect 16724 19468 16769 19496
rect 16995 19468 17040 19496
rect 16724 19456 16730 19468
rect 17034 19456 17040 19468
rect 17092 19456 17098 19508
rect 17497 19499 17555 19505
rect 17497 19465 17509 19499
rect 17543 19496 17555 19499
rect 18138 19496 18144 19508
rect 17543 19468 18144 19496
rect 17543 19465 17555 19468
rect 17497 19459 17555 19465
rect 18138 19456 18144 19468
rect 18196 19496 18202 19508
rect 18506 19496 18512 19508
rect 18196 19468 18512 19496
rect 18196 19456 18202 19468
rect 18506 19456 18512 19468
rect 18564 19456 18570 19508
rect 19334 19456 19340 19508
rect 19392 19496 19398 19508
rect 20625 19499 20683 19505
rect 20625 19496 20637 19499
rect 19392 19468 20637 19496
rect 19392 19456 19398 19468
rect 20625 19465 20637 19468
rect 20671 19465 20683 19499
rect 20625 19459 20683 19465
rect 21177 19499 21235 19505
rect 21177 19465 21189 19499
rect 21223 19496 21235 19499
rect 21821 19499 21879 19505
rect 21821 19496 21833 19499
rect 21223 19468 21833 19496
rect 21223 19465 21235 19468
rect 21177 19459 21235 19465
rect 21821 19465 21833 19468
rect 21867 19465 21879 19499
rect 21821 19459 21879 19465
rect 16298 19388 16304 19440
rect 16356 19428 16362 19440
rect 17129 19431 17187 19437
rect 17129 19428 17141 19431
rect 16356 19400 17141 19428
rect 16356 19388 16362 19400
rect 17129 19397 17141 19400
rect 17175 19397 17187 19431
rect 17129 19391 17187 19397
rect 18632 19431 18690 19437
rect 18632 19397 18644 19431
rect 18678 19428 18690 19431
rect 20714 19428 20720 19440
rect 18678 19400 20720 19428
rect 18678 19397 18690 19400
rect 18632 19391 18690 19397
rect 20714 19388 20720 19400
rect 20772 19388 20778 19440
rect 21082 19388 21088 19440
rect 21140 19428 21146 19440
rect 21140 19400 22876 19428
rect 21140 19388 21146 19400
rect 15804 19332 16252 19360
rect 15804 19320 15810 19332
rect 17402 19320 17408 19372
rect 17460 19360 17466 19372
rect 19058 19360 19064 19372
rect 17460 19332 19064 19360
rect 17460 19320 17466 19332
rect 19058 19320 19064 19332
rect 19116 19320 19122 19372
rect 20070 19360 20076 19372
rect 20128 19369 20134 19372
rect 20040 19332 20076 19360
rect 20070 19320 20076 19332
rect 20128 19323 20140 19369
rect 20530 19360 20536 19372
rect 20364 19332 20536 19360
rect 20128 19320 20134 19323
rect 9631 19264 9904 19292
rect 11057 19295 11115 19301
rect 9631 19261 9643 19264
rect 9585 19255 9643 19261
rect 11057 19261 11069 19295
rect 11103 19292 11115 19295
rect 11103 19264 11192 19292
rect 11103 19261 11115 19264
rect 11057 19255 11115 19261
rect 9674 19224 9680 19236
rect 9635 19196 9680 19224
rect 9674 19184 9680 19196
rect 9732 19184 9738 19236
rect 11164 19168 11192 19264
rect 12894 19252 12900 19304
rect 12952 19292 12958 19304
rect 13538 19292 13544 19304
rect 12952 19264 13400 19292
rect 13499 19264 13544 19292
rect 12952 19252 12958 19264
rect 13372 19224 13400 19264
rect 13538 19252 13544 19264
rect 13596 19292 13602 19304
rect 13817 19295 13875 19301
rect 13817 19292 13829 19295
rect 13596 19264 13829 19292
rect 13596 19252 13602 19264
rect 13817 19261 13829 19264
rect 13863 19261 13875 19295
rect 13817 19255 13875 19261
rect 17221 19295 17279 19301
rect 17221 19261 17233 19295
rect 17267 19261 17279 19295
rect 17221 19255 17279 19261
rect 18877 19295 18935 19301
rect 18877 19261 18889 19295
rect 18923 19292 18935 19295
rect 19242 19292 19248 19304
rect 18923 19264 19248 19292
rect 18923 19261 18935 19264
rect 18877 19255 18935 19261
rect 13372 19196 13676 19224
rect 13648 19168 13676 19196
rect 1946 19156 1952 19168
rect 1859 19128 1952 19156
rect 1946 19116 1952 19128
rect 2004 19156 2010 19168
rect 6086 19156 6092 19168
rect 2004 19128 6092 19156
rect 2004 19116 2010 19128
rect 6086 19116 6092 19128
rect 6144 19116 6150 19168
rect 6178 19116 6184 19168
rect 6236 19156 6242 19168
rect 6365 19159 6423 19165
rect 6365 19156 6377 19159
rect 6236 19128 6377 19156
rect 6236 19116 6242 19128
rect 6365 19125 6377 19128
rect 6411 19156 6423 19159
rect 6549 19159 6607 19165
rect 6549 19156 6561 19159
rect 6411 19128 6561 19156
rect 6411 19125 6423 19128
rect 6365 19119 6423 19125
rect 6549 19125 6561 19128
rect 6595 19156 6607 19159
rect 6733 19159 6791 19165
rect 6733 19156 6745 19159
rect 6595 19128 6745 19156
rect 6595 19125 6607 19128
rect 6549 19119 6607 19125
rect 6733 19125 6745 19128
rect 6779 19156 6791 19159
rect 7009 19159 7067 19165
rect 7009 19156 7021 19159
rect 6779 19128 7021 19156
rect 6779 19125 6791 19128
rect 6733 19119 6791 19125
rect 7009 19125 7021 19128
rect 7055 19156 7067 19159
rect 7377 19159 7435 19165
rect 7377 19156 7389 19159
rect 7055 19128 7389 19156
rect 7055 19125 7067 19128
rect 7009 19119 7067 19125
rect 7377 19125 7389 19128
rect 7423 19125 7435 19159
rect 11146 19156 11152 19168
rect 11107 19128 11152 19156
rect 7377 19119 7435 19125
rect 11146 19116 11152 19128
rect 11204 19116 11210 19168
rect 12989 19159 13047 19165
rect 12989 19125 13001 19159
rect 13035 19156 13047 19159
rect 13078 19156 13084 19168
rect 13035 19128 13084 19156
rect 13035 19125 13047 19128
rect 12989 19119 13047 19125
rect 13078 19116 13084 19128
rect 13136 19116 13142 19168
rect 13630 19116 13636 19168
rect 13688 19156 13694 19168
rect 14274 19156 14280 19168
rect 13688 19128 14280 19156
rect 13688 19116 13694 19128
rect 14274 19116 14280 19128
rect 14332 19116 14338 19168
rect 14366 19116 14372 19168
rect 14424 19156 14430 19168
rect 17236 19156 17264 19255
rect 19242 19252 19248 19264
rect 19300 19252 19306 19304
rect 20364 19301 20392 19332
rect 20530 19320 20536 19332
rect 20588 19320 20594 19372
rect 20809 19363 20867 19369
rect 20809 19329 20821 19363
rect 20855 19360 20867 19363
rect 20898 19360 20904 19372
rect 20855 19332 20904 19360
rect 20855 19329 20867 19332
rect 20809 19323 20867 19329
rect 20898 19320 20904 19332
rect 20956 19320 20962 19372
rect 21269 19363 21327 19369
rect 21269 19329 21281 19363
rect 21315 19360 21327 19363
rect 22094 19360 22100 19372
rect 21315 19332 22100 19360
rect 21315 19329 21327 19332
rect 21269 19323 21327 19329
rect 22094 19320 22100 19332
rect 22152 19320 22158 19372
rect 22189 19363 22247 19369
rect 22189 19329 22201 19363
rect 22235 19360 22247 19363
rect 22370 19360 22376 19372
rect 22235 19332 22376 19360
rect 22235 19329 22247 19332
rect 22189 19323 22247 19329
rect 22370 19320 22376 19332
rect 22428 19320 22434 19372
rect 22848 19369 22876 19400
rect 22833 19363 22891 19369
rect 22833 19329 22845 19363
rect 22879 19329 22891 19363
rect 22833 19323 22891 19329
rect 20349 19295 20407 19301
rect 20349 19261 20361 19295
rect 20395 19292 20407 19295
rect 21085 19295 21143 19301
rect 20395 19264 20429 19292
rect 20395 19261 20407 19264
rect 20349 19255 20407 19261
rect 21085 19261 21097 19295
rect 21131 19292 21143 19295
rect 21726 19292 21732 19304
rect 21131 19264 21732 19292
rect 21131 19261 21143 19264
rect 21085 19255 21143 19261
rect 21726 19252 21732 19264
rect 21784 19252 21790 19304
rect 21910 19252 21916 19304
rect 21968 19292 21974 19304
rect 22281 19295 22339 19301
rect 22281 19292 22293 19295
rect 21968 19264 22293 19292
rect 21968 19252 21974 19264
rect 22281 19261 22293 19264
rect 22327 19261 22339 19295
rect 22462 19292 22468 19304
rect 22423 19264 22468 19292
rect 22281 19255 22339 19261
rect 22462 19252 22468 19264
rect 22520 19252 22526 19304
rect 21100 19196 21956 19224
rect 14424 19128 17264 19156
rect 14424 19116 14430 19128
rect 18506 19116 18512 19168
rect 18564 19156 18570 19168
rect 18969 19159 19027 19165
rect 18969 19156 18981 19159
rect 18564 19128 18981 19156
rect 18564 19116 18570 19128
rect 18969 19125 18981 19128
rect 19015 19156 19027 19159
rect 21100 19156 21128 19196
rect 19015 19128 21128 19156
rect 19015 19125 19027 19128
rect 18969 19119 19027 19125
rect 21174 19116 21180 19168
rect 21232 19156 21238 19168
rect 21637 19159 21695 19165
rect 21637 19156 21649 19159
rect 21232 19128 21649 19156
rect 21232 19116 21238 19128
rect 21637 19125 21649 19128
rect 21683 19125 21695 19159
rect 21928 19156 21956 19196
rect 22002 19184 22008 19236
rect 22060 19224 22066 19236
rect 22830 19224 22836 19236
rect 22060 19196 22836 19224
rect 22060 19184 22066 19196
rect 22830 19184 22836 19196
rect 22888 19184 22894 19236
rect 22278 19156 22284 19168
rect 21928 19128 22284 19156
rect 21637 19119 21695 19125
rect 22278 19116 22284 19128
rect 22336 19116 22342 19168
rect 22738 19156 22744 19168
rect 22699 19128 22744 19156
rect 22738 19116 22744 19128
rect 22796 19116 22802 19168
rect 23014 19156 23020 19168
rect 22975 19128 23020 19156
rect 23014 19116 23020 19128
rect 23072 19116 23078 19168
rect 1104 19066 23460 19088
rect 1104 19014 3749 19066
rect 3801 19014 3813 19066
rect 3865 19014 3877 19066
rect 3929 19014 3941 19066
rect 3993 19014 4005 19066
rect 4057 19014 9347 19066
rect 9399 19014 9411 19066
rect 9463 19014 9475 19066
rect 9527 19014 9539 19066
rect 9591 19014 9603 19066
rect 9655 19014 14945 19066
rect 14997 19014 15009 19066
rect 15061 19014 15073 19066
rect 15125 19014 15137 19066
rect 15189 19014 15201 19066
rect 15253 19014 20543 19066
rect 20595 19014 20607 19066
rect 20659 19014 20671 19066
rect 20723 19014 20735 19066
rect 20787 19014 20799 19066
rect 20851 19014 23460 19066
rect 1104 18992 23460 19014
rect 3510 18912 3516 18964
rect 3568 18952 3574 18964
rect 3973 18955 4031 18961
rect 3973 18952 3985 18955
rect 3568 18924 3985 18952
rect 3568 18912 3574 18924
rect 3973 18921 3985 18924
rect 4019 18921 4031 18955
rect 5626 18952 5632 18964
rect 3973 18915 4031 18921
rect 4816 18924 5632 18952
rect 3605 18887 3663 18893
rect 3605 18853 3617 18887
rect 3651 18884 3663 18887
rect 4338 18884 4344 18896
rect 3651 18856 4344 18884
rect 3651 18853 3663 18856
rect 3605 18847 3663 18853
rect 4338 18844 4344 18856
rect 4396 18844 4402 18896
rect 1946 18776 1952 18828
rect 2004 18816 2010 18828
rect 2041 18819 2099 18825
rect 2041 18816 2053 18819
rect 2004 18788 2053 18816
rect 2004 18776 2010 18788
rect 2041 18785 2053 18788
rect 2087 18785 2099 18819
rect 2041 18779 2099 18785
rect 3053 18819 3111 18825
rect 3053 18785 3065 18819
rect 3099 18816 3111 18819
rect 4816 18816 4844 18924
rect 5626 18912 5632 18924
rect 5684 18912 5690 18964
rect 5902 18952 5908 18964
rect 5863 18924 5908 18952
rect 5902 18912 5908 18924
rect 5960 18912 5966 18964
rect 7377 18955 7435 18961
rect 7377 18921 7389 18955
rect 7423 18952 7435 18955
rect 8018 18952 8024 18964
rect 7423 18924 8024 18952
rect 7423 18921 7435 18924
rect 7377 18915 7435 18921
rect 3099 18788 4844 18816
rect 3099 18785 3111 18788
rect 3053 18779 3111 18785
rect 4246 18708 4252 18760
rect 4304 18748 4310 18760
rect 4798 18748 4804 18760
rect 4304 18720 4804 18748
rect 4304 18708 4310 18720
rect 4798 18708 4804 18720
rect 4856 18748 4862 18760
rect 5546 18751 5604 18757
rect 5546 18748 5558 18751
rect 4856 18720 5558 18748
rect 4856 18708 4862 18720
rect 5546 18717 5558 18720
rect 5592 18717 5604 18751
rect 5546 18711 5604 18717
rect 5813 18751 5871 18757
rect 5813 18717 5825 18751
rect 5859 18748 5871 18751
rect 6178 18748 6184 18760
rect 5859 18720 6184 18748
rect 5859 18717 5871 18720
rect 5813 18711 5871 18717
rect 6178 18708 6184 18720
rect 6236 18748 6242 18760
rect 7285 18751 7343 18757
rect 7285 18748 7297 18751
rect 6236 18720 7297 18748
rect 6236 18708 6242 18720
rect 7285 18717 7297 18720
rect 7331 18717 7343 18751
rect 7285 18711 7343 18717
rect 1946 18640 1952 18692
rect 2004 18680 2010 18692
rect 3145 18683 3203 18689
rect 3145 18680 3157 18683
rect 2004 18652 3157 18680
rect 2004 18640 2010 18652
rect 3145 18649 3157 18652
rect 3191 18649 3203 18683
rect 4154 18680 4160 18692
rect 4115 18652 4160 18680
rect 3145 18643 3203 18649
rect 4154 18640 4160 18652
rect 4212 18640 4218 18692
rect 4341 18683 4399 18689
rect 4341 18649 4353 18683
rect 4387 18680 4399 18683
rect 6914 18680 6920 18692
rect 4387 18652 6920 18680
rect 4387 18649 4399 18652
rect 4341 18643 4399 18649
rect 6914 18640 6920 18652
rect 6972 18640 6978 18692
rect 7040 18683 7098 18689
rect 7040 18649 7052 18683
rect 7086 18680 7098 18683
rect 7392 18680 7420 18915
rect 8018 18912 8024 18924
rect 8076 18912 8082 18964
rect 10870 18912 10876 18964
rect 10928 18952 10934 18964
rect 11057 18955 11115 18961
rect 11057 18952 11069 18955
rect 10928 18924 11069 18952
rect 10928 18912 10934 18924
rect 11057 18921 11069 18924
rect 11103 18921 11115 18955
rect 12986 18952 12992 18964
rect 12947 18924 12992 18952
rect 11057 18915 11115 18921
rect 12986 18912 12992 18924
rect 13044 18952 13050 18964
rect 13630 18952 13636 18964
rect 13044 18924 13636 18952
rect 13044 18912 13050 18924
rect 13630 18912 13636 18924
rect 13688 18912 13694 18964
rect 15286 18952 15292 18964
rect 13740 18924 15292 18952
rect 13078 18844 13084 18896
rect 13136 18884 13142 18896
rect 13740 18884 13768 18924
rect 15286 18912 15292 18924
rect 15344 18912 15350 18964
rect 15749 18955 15807 18961
rect 15749 18921 15761 18955
rect 15795 18952 15807 18955
rect 15838 18952 15844 18964
rect 15795 18924 15844 18952
rect 15795 18921 15807 18924
rect 15749 18915 15807 18921
rect 15838 18912 15844 18924
rect 15896 18952 15902 18964
rect 17310 18952 17316 18964
rect 15896 18924 17316 18952
rect 15896 18912 15902 18924
rect 17310 18912 17316 18924
rect 17368 18912 17374 18964
rect 19061 18955 19119 18961
rect 19061 18921 19073 18955
rect 19107 18952 19119 18955
rect 22002 18952 22008 18964
rect 19107 18924 22008 18952
rect 19107 18921 19119 18924
rect 19061 18915 19119 18921
rect 22002 18912 22008 18924
rect 22060 18912 22066 18964
rect 22094 18912 22100 18964
rect 22152 18952 22158 18964
rect 22373 18955 22431 18961
rect 22373 18952 22385 18955
rect 22152 18924 22385 18952
rect 22152 18912 22158 18924
rect 22373 18921 22385 18924
rect 22419 18921 22431 18955
rect 22373 18915 22431 18921
rect 13136 18856 13768 18884
rect 18693 18887 18751 18893
rect 13136 18844 13142 18856
rect 18693 18853 18705 18887
rect 18739 18884 18751 18887
rect 19426 18884 19432 18896
rect 18739 18856 19432 18884
rect 18739 18853 18751 18856
rect 18693 18847 18751 18853
rect 19426 18844 19432 18856
rect 19484 18844 19490 18896
rect 20806 18844 20812 18896
rect 20864 18884 20870 18896
rect 20901 18887 20959 18893
rect 20901 18884 20913 18887
rect 20864 18856 20913 18884
rect 20864 18844 20870 18856
rect 20901 18853 20913 18856
rect 20947 18853 20959 18887
rect 20901 18847 20959 18853
rect 9030 18816 9036 18828
rect 8680 18788 9036 18816
rect 8501 18751 8559 18757
rect 8501 18717 8513 18751
rect 8547 18748 8559 18751
rect 8680 18748 8708 18788
rect 9030 18776 9036 18788
rect 9088 18776 9094 18828
rect 13814 18776 13820 18828
rect 13872 18816 13878 18828
rect 13909 18819 13967 18825
rect 13909 18816 13921 18819
rect 13872 18788 13921 18816
rect 13872 18776 13878 18788
rect 13909 18785 13921 18788
rect 13955 18785 13967 18819
rect 13909 18779 13967 18785
rect 15746 18776 15752 18828
rect 15804 18816 15810 18828
rect 15841 18819 15899 18825
rect 15841 18816 15853 18819
rect 15804 18788 15853 18816
rect 15804 18776 15810 18788
rect 15841 18785 15853 18788
rect 15887 18785 15899 18819
rect 15841 18779 15899 18785
rect 8547 18720 8708 18748
rect 8757 18751 8815 18757
rect 8547 18717 8559 18720
rect 8501 18711 8559 18717
rect 8757 18717 8769 18751
rect 8803 18748 8815 18751
rect 9582 18748 9588 18760
rect 8803 18720 9588 18748
rect 8803 18717 8815 18720
rect 8757 18711 8815 18717
rect 7086 18652 7420 18680
rect 7086 18649 7098 18652
rect 7040 18643 7098 18649
rect 1670 18572 1676 18624
rect 1728 18612 1734 18624
rect 2225 18615 2283 18621
rect 2225 18612 2237 18615
rect 1728 18584 2237 18612
rect 1728 18572 1734 18584
rect 2225 18581 2237 18584
rect 2271 18581 2283 18615
rect 2225 18575 2283 18581
rect 2314 18572 2320 18624
rect 2372 18612 2378 18624
rect 2682 18612 2688 18624
rect 2372 18584 2417 18612
rect 2643 18584 2688 18612
rect 2372 18572 2378 18584
rect 2682 18572 2688 18584
rect 2740 18572 2746 18624
rect 3234 18612 3240 18624
rect 3195 18584 3240 18612
rect 3234 18572 3240 18584
rect 3292 18572 3298 18624
rect 4430 18612 4436 18624
rect 4391 18584 4436 18612
rect 4430 18572 4436 18584
rect 4488 18572 4494 18624
rect 5350 18572 5356 18624
rect 5408 18612 5414 18624
rect 8110 18612 8116 18624
rect 5408 18584 8116 18612
rect 5408 18572 5414 18584
rect 8110 18572 8116 18584
rect 8168 18572 8174 18624
rect 8294 18572 8300 18624
rect 8352 18612 8358 18624
rect 8772 18612 8800 18711
rect 9582 18708 9588 18720
rect 9640 18748 9646 18760
rect 9677 18751 9735 18757
rect 9677 18748 9689 18751
rect 9640 18720 9689 18748
rect 9640 18708 9646 18720
rect 9677 18717 9689 18720
rect 9723 18748 9735 18751
rect 11146 18748 11152 18760
rect 9723 18720 11152 18748
rect 9723 18717 9735 18720
rect 9677 18711 9735 18717
rect 11146 18708 11152 18720
rect 11204 18748 11210 18760
rect 11425 18751 11483 18757
rect 11425 18748 11437 18751
rect 11204 18720 11437 18748
rect 11204 18708 11210 18720
rect 11425 18717 11437 18720
rect 11471 18748 11483 18751
rect 11609 18751 11667 18757
rect 11609 18748 11621 18751
rect 11471 18720 11621 18748
rect 11471 18717 11483 18720
rect 11425 18711 11483 18717
rect 11609 18717 11621 18720
rect 11655 18748 11667 18751
rect 12894 18748 12900 18760
rect 11655 18720 12900 18748
rect 11655 18717 11667 18720
rect 11609 18711 11667 18717
rect 12894 18708 12900 18720
rect 12952 18708 12958 18760
rect 13446 18708 13452 18760
rect 13504 18748 13510 18760
rect 13633 18751 13691 18757
rect 13633 18748 13645 18751
rect 13504 18720 13645 18748
rect 13504 18708 13510 18720
rect 13633 18717 13645 18720
rect 13679 18748 13691 18751
rect 14185 18751 14243 18757
rect 13679 18720 13860 18748
rect 13679 18717 13691 18720
rect 13633 18711 13691 18717
rect 8846 18640 8852 18692
rect 8904 18680 8910 18692
rect 9922 18683 9980 18689
rect 9922 18680 9934 18683
rect 8904 18652 9934 18680
rect 8904 18640 8910 18652
rect 9922 18649 9934 18652
rect 9968 18649 9980 18683
rect 9922 18643 9980 18649
rect 11876 18683 11934 18689
rect 11876 18649 11888 18683
rect 11922 18680 11934 18683
rect 13722 18680 13728 18692
rect 11922 18652 13728 18680
rect 11922 18649 11934 18652
rect 11876 18643 11934 18649
rect 13722 18640 13728 18652
rect 13780 18640 13786 18692
rect 8941 18615 8999 18621
rect 8941 18612 8953 18615
rect 8352 18584 8953 18612
rect 8352 18572 8358 18584
rect 8941 18581 8953 18584
rect 8987 18581 8999 18615
rect 13832 18612 13860 18720
rect 14185 18717 14197 18751
rect 14231 18748 14243 18751
rect 14274 18748 14280 18760
rect 14231 18720 14280 18748
rect 14231 18717 14243 18720
rect 14185 18711 14243 18717
rect 14274 18708 14280 18720
rect 14332 18748 14338 18760
rect 14369 18751 14427 18757
rect 14369 18748 14381 18751
rect 14332 18720 14381 18748
rect 14332 18708 14338 18720
rect 14369 18717 14381 18720
rect 14415 18748 14427 18751
rect 15856 18748 15884 18779
rect 22462 18776 22468 18828
rect 22520 18816 22526 18828
rect 22646 18816 22652 18828
rect 22520 18788 22652 18816
rect 22520 18776 22526 18788
rect 22646 18776 22652 18788
rect 22704 18816 22710 18828
rect 22925 18819 22983 18825
rect 22925 18816 22937 18819
rect 22704 18788 22937 18816
rect 22704 18776 22710 18788
rect 22925 18785 22937 18788
rect 22971 18785 22983 18819
rect 22925 18779 22983 18785
rect 17313 18751 17371 18757
rect 17313 18748 17325 18751
rect 14415 18720 17325 18748
rect 14415 18717 14427 18720
rect 14369 18711 14427 18717
rect 17313 18717 17325 18720
rect 17359 18717 17371 18751
rect 18874 18748 18880 18760
rect 18835 18720 18880 18748
rect 17313 18711 17371 18717
rect 18874 18708 18880 18720
rect 18932 18708 18938 18760
rect 19242 18708 19248 18760
rect 19300 18748 19306 18760
rect 19337 18751 19395 18757
rect 19337 18748 19349 18751
rect 19300 18720 19349 18748
rect 19300 18708 19306 18720
rect 19337 18717 19349 18720
rect 19383 18748 19395 18751
rect 20714 18748 20720 18760
rect 19383 18720 20720 18748
rect 19383 18717 19395 18720
rect 19337 18711 19395 18717
rect 20714 18708 20720 18720
rect 20772 18748 20778 18760
rect 20809 18751 20867 18757
rect 20809 18748 20821 18751
rect 20772 18720 20821 18748
rect 20772 18708 20778 18720
rect 20809 18717 20821 18720
rect 20855 18748 20867 18751
rect 22281 18751 22339 18757
rect 22281 18748 22293 18751
rect 20855 18720 22293 18748
rect 20855 18717 20867 18720
rect 20809 18711 20867 18717
rect 22281 18717 22293 18720
rect 22327 18717 22339 18751
rect 22281 18711 22339 18717
rect 22370 18708 22376 18760
rect 22428 18748 22434 18760
rect 22833 18751 22891 18757
rect 22833 18748 22845 18751
rect 22428 18720 22845 18748
rect 22428 18708 22434 18720
rect 22833 18717 22845 18720
rect 22879 18717 22891 18751
rect 22833 18711 22891 18717
rect 14636 18683 14694 18689
rect 14636 18649 14648 18683
rect 14682 18680 14694 18683
rect 15930 18680 15936 18692
rect 14682 18652 15936 18680
rect 14682 18649 14694 18652
rect 14636 18643 14694 18649
rect 15930 18640 15936 18652
rect 15988 18640 15994 18692
rect 16108 18683 16166 18689
rect 16108 18649 16120 18683
rect 16154 18680 16166 18683
rect 16942 18680 16948 18692
rect 16154 18652 16948 18680
rect 16154 18649 16166 18652
rect 16108 18643 16166 18649
rect 16942 18640 16948 18652
rect 17000 18640 17006 18692
rect 17586 18689 17592 18692
rect 17580 18680 17592 18689
rect 17547 18652 17592 18680
rect 17580 18643 17592 18652
rect 17586 18640 17592 18643
rect 17644 18640 17650 18692
rect 19794 18680 19800 18692
rect 17696 18652 19800 18680
rect 14550 18612 14556 18624
rect 13832 18584 14556 18612
rect 8941 18575 8999 18581
rect 14550 18572 14556 18584
rect 14608 18572 14614 18624
rect 17218 18612 17224 18624
rect 17179 18584 17224 18612
rect 17218 18572 17224 18584
rect 17276 18572 17282 18624
rect 17402 18572 17408 18624
rect 17460 18612 17466 18624
rect 17696 18612 17724 18652
rect 19794 18640 19800 18652
rect 19852 18640 19858 18692
rect 20438 18640 20444 18692
rect 20496 18680 20502 18692
rect 20542 18683 20600 18689
rect 20542 18680 20554 18683
rect 20496 18652 20554 18680
rect 20496 18640 20502 18652
rect 20542 18649 20554 18652
rect 20588 18649 20600 18683
rect 20542 18643 20600 18649
rect 21910 18640 21916 18692
rect 21968 18680 21974 18692
rect 22025 18683 22083 18689
rect 22025 18680 22037 18683
rect 21968 18652 22037 18680
rect 21968 18640 21974 18652
rect 22025 18649 22037 18652
rect 22071 18649 22083 18683
rect 22025 18643 22083 18649
rect 17460 18584 17724 18612
rect 19429 18615 19487 18621
rect 17460 18572 17466 18584
rect 19429 18581 19441 18615
rect 19475 18612 19487 18615
rect 19702 18612 19708 18624
rect 19475 18584 19708 18612
rect 19475 18581 19487 18584
rect 19429 18575 19487 18581
rect 19702 18572 19708 18584
rect 19760 18572 19766 18624
rect 22462 18572 22468 18624
rect 22520 18612 22526 18624
rect 22741 18615 22799 18621
rect 22741 18612 22753 18615
rect 22520 18584 22753 18612
rect 22520 18572 22526 18584
rect 22741 18581 22753 18584
rect 22787 18581 22799 18615
rect 22741 18575 22799 18581
rect 1104 18522 23460 18544
rect 1104 18470 6548 18522
rect 6600 18470 6612 18522
rect 6664 18470 6676 18522
rect 6728 18470 6740 18522
rect 6792 18470 6804 18522
rect 6856 18470 12146 18522
rect 12198 18470 12210 18522
rect 12262 18470 12274 18522
rect 12326 18470 12338 18522
rect 12390 18470 12402 18522
rect 12454 18470 17744 18522
rect 17796 18470 17808 18522
rect 17860 18470 17872 18522
rect 17924 18470 17936 18522
rect 17988 18470 18000 18522
rect 18052 18470 23460 18522
rect 1104 18448 23460 18470
rect 2041 18411 2099 18417
rect 2041 18377 2053 18411
rect 2087 18377 2099 18411
rect 2041 18371 2099 18377
rect 2133 18411 2191 18417
rect 2133 18377 2145 18411
rect 2179 18408 2191 18411
rect 2314 18408 2320 18420
rect 2179 18380 2320 18408
rect 2179 18377 2191 18380
rect 2133 18371 2191 18377
rect 2056 18340 2084 18371
rect 2314 18368 2320 18380
rect 2372 18368 2378 18420
rect 5350 18408 5356 18420
rect 2746 18380 5356 18408
rect 2746 18340 2774 18380
rect 5350 18368 5356 18380
rect 5408 18368 5414 18420
rect 5442 18368 5448 18420
rect 5500 18408 5506 18420
rect 5500 18380 6316 18408
rect 5500 18368 5506 18380
rect 6288 18340 6316 18380
rect 7834 18368 7840 18420
rect 7892 18408 7898 18420
rect 8113 18411 8171 18417
rect 8113 18408 8125 18411
rect 7892 18380 8125 18408
rect 7892 18368 7898 18380
rect 8113 18377 8125 18380
rect 8159 18377 8171 18411
rect 8113 18371 8171 18377
rect 9582 18368 9588 18420
rect 9640 18408 9646 18420
rect 9677 18411 9735 18417
rect 9677 18408 9689 18411
rect 9640 18380 9689 18408
rect 9640 18368 9646 18380
rect 9677 18377 9689 18380
rect 9723 18377 9735 18411
rect 9677 18371 9735 18377
rect 6978 18343 7036 18349
rect 6978 18340 6990 18343
rect 2056 18312 2774 18340
rect 4816 18312 6224 18340
rect 6288 18312 6990 18340
rect 1854 18272 1860 18284
rect 1815 18244 1860 18272
rect 1854 18232 1860 18244
rect 1912 18232 1918 18284
rect 2317 18275 2375 18281
rect 2317 18241 2329 18275
rect 2363 18272 2375 18275
rect 2406 18272 2412 18284
rect 2363 18244 2412 18272
rect 2363 18241 2375 18244
rect 2317 18235 2375 18241
rect 2406 18232 2412 18244
rect 2464 18232 2470 18284
rect 3237 18275 3295 18281
rect 3237 18241 3249 18275
rect 3283 18272 3295 18275
rect 4062 18272 4068 18284
rect 3283 18244 4068 18272
rect 3283 18241 3295 18244
rect 3237 18235 3295 18241
rect 4062 18232 4068 18244
rect 4120 18232 4126 18284
rect 4154 18232 4160 18284
rect 4212 18272 4218 18284
rect 4453 18275 4511 18281
rect 4453 18272 4465 18275
rect 4212 18244 4465 18272
rect 4212 18232 4218 18244
rect 4453 18241 4465 18244
rect 4499 18272 4511 18275
rect 4614 18272 4620 18284
rect 4499 18244 4620 18272
rect 4499 18241 4511 18244
rect 4453 18235 4511 18241
rect 4614 18232 4620 18244
rect 4672 18232 4678 18284
rect 4816 18281 4844 18312
rect 4709 18275 4767 18281
rect 4709 18241 4721 18275
rect 4755 18272 4767 18275
rect 4801 18275 4859 18281
rect 4801 18272 4813 18275
rect 4755 18244 4813 18272
rect 4755 18241 4767 18244
rect 4709 18235 4767 18241
rect 4801 18241 4813 18244
rect 4847 18241 4859 18275
rect 5057 18275 5115 18281
rect 5057 18272 5069 18275
rect 4801 18235 4859 18241
rect 4908 18244 5069 18272
rect 2961 18207 3019 18213
rect 2961 18173 2973 18207
rect 3007 18204 3019 18207
rect 3510 18204 3516 18216
rect 3007 18176 3516 18204
rect 3007 18173 3019 18176
rect 2961 18167 3019 18173
rect 3510 18164 3516 18176
rect 3568 18164 3574 18216
rect 4908 18204 4936 18244
rect 5057 18241 5069 18244
rect 5103 18241 5115 18275
rect 5057 18235 5115 18241
rect 6196 18216 6224 18312
rect 6978 18309 6990 18312
rect 7024 18309 7036 18343
rect 8450 18343 8508 18349
rect 8450 18340 8462 18343
rect 6978 18303 7036 18309
rect 7760 18312 8462 18340
rect 4724 18176 4936 18204
rect 2958 18028 2964 18080
rect 3016 18068 3022 18080
rect 3329 18071 3387 18077
rect 3329 18068 3341 18071
rect 3016 18040 3341 18068
rect 3016 18028 3022 18040
rect 3329 18037 3341 18040
rect 3375 18068 3387 18071
rect 4724 18068 4752 18176
rect 6178 18164 6184 18216
rect 6236 18204 6242 18216
rect 6365 18207 6423 18213
rect 6365 18204 6377 18207
rect 6236 18176 6377 18204
rect 6236 18164 6242 18176
rect 6365 18173 6377 18176
rect 6411 18204 6423 18207
rect 6549 18207 6607 18213
rect 6549 18204 6561 18207
rect 6411 18176 6561 18204
rect 6411 18173 6423 18176
rect 6365 18167 6423 18173
rect 6549 18173 6561 18176
rect 6595 18204 6607 18207
rect 6733 18207 6791 18213
rect 6733 18204 6745 18207
rect 6595 18176 6745 18204
rect 6595 18173 6607 18176
rect 6549 18167 6607 18173
rect 6733 18173 6745 18176
rect 6779 18173 6791 18207
rect 6733 18167 6791 18173
rect 3375 18040 4752 18068
rect 3375 18037 3387 18040
rect 3329 18031 3387 18037
rect 5074 18028 5080 18080
rect 5132 18068 5138 18080
rect 6181 18071 6239 18077
rect 6181 18068 6193 18071
rect 5132 18040 6193 18068
rect 5132 18028 5138 18040
rect 6181 18037 6193 18040
rect 6227 18068 6239 18071
rect 7760 18068 7788 18312
rect 8450 18309 8462 18312
rect 8496 18309 8508 18343
rect 8450 18303 8508 18309
rect 8205 18275 8263 18281
rect 8205 18241 8217 18275
rect 8251 18272 8263 18275
rect 8294 18272 8300 18284
rect 8251 18244 8300 18272
rect 8251 18241 8263 18244
rect 8205 18235 8263 18241
rect 8294 18232 8300 18244
rect 8352 18232 8358 18284
rect 9692 18272 9720 18371
rect 9766 18368 9772 18420
rect 9824 18368 9830 18420
rect 11333 18411 11391 18417
rect 11333 18377 11345 18411
rect 11379 18408 11391 18411
rect 11379 18380 12434 18408
rect 11379 18377 11391 18380
rect 11333 18371 11391 18377
rect 9784 18340 9812 18368
rect 10198 18343 10256 18349
rect 10198 18340 10210 18343
rect 9784 18312 10210 18340
rect 10198 18309 10210 18312
rect 10244 18309 10256 18343
rect 12406 18340 12434 18380
rect 14274 18368 14280 18420
rect 14332 18368 14338 18420
rect 14642 18368 14648 18420
rect 14700 18408 14706 18420
rect 15565 18411 15623 18417
rect 15565 18408 15577 18411
rect 14700 18380 15577 18408
rect 14700 18368 14706 18380
rect 15565 18377 15577 18380
rect 15611 18377 15623 18411
rect 15565 18371 15623 18377
rect 15746 18368 15752 18420
rect 15804 18408 15810 18420
rect 16393 18411 16451 18417
rect 16393 18408 16405 18411
rect 15804 18380 16405 18408
rect 15804 18368 15810 18380
rect 16393 18377 16405 18380
rect 16439 18377 16451 18411
rect 16393 18371 16451 18377
rect 12744 18343 12802 18349
rect 12744 18340 12756 18343
rect 12406 18312 12756 18340
rect 10198 18303 10256 18309
rect 12744 18309 12756 18312
rect 12790 18340 12802 18343
rect 13078 18340 13084 18352
rect 12790 18312 13084 18340
rect 12790 18309 12802 18312
rect 12744 18303 12802 18309
rect 13078 18300 13084 18312
rect 13136 18300 13142 18352
rect 13630 18340 13636 18352
rect 13591 18312 13636 18340
rect 13630 18300 13636 18312
rect 13688 18300 13694 18352
rect 9953 18275 10011 18281
rect 9953 18272 9965 18275
rect 9692 18244 9965 18272
rect 9953 18241 9965 18244
rect 9999 18241 10011 18275
rect 9953 18235 10011 18241
rect 12989 18275 13047 18281
rect 12989 18241 13001 18275
rect 13035 18272 13047 18275
rect 13173 18275 13231 18281
rect 13173 18272 13185 18275
rect 13035 18244 13185 18272
rect 13035 18241 13047 18244
rect 12989 18235 13047 18241
rect 13173 18241 13185 18244
rect 13219 18272 13231 18275
rect 14093 18275 14151 18281
rect 14093 18272 14105 18275
rect 13219 18244 14105 18272
rect 13219 18241 13231 18244
rect 13173 18235 13231 18241
rect 14093 18241 14105 18244
rect 14139 18272 14151 18275
rect 14292 18272 14320 18368
rect 14360 18343 14418 18349
rect 14360 18309 14372 18343
rect 14406 18340 14418 18343
rect 14734 18340 14740 18352
rect 14406 18312 14740 18340
rect 14406 18309 14418 18312
rect 14360 18303 14418 18309
rect 14734 18300 14740 18312
rect 14792 18300 14798 18352
rect 15120 18312 16160 18340
rect 14139 18244 14320 18272
rect 14139 18241 14151 18244
rect 14093 18235 14151 18241
rect 14642 18232 14648 18284
rect 14700 18272 14706 18284
rect 15120 18272 15148 18312
rect 14700 18244 15148 18272
rect 14700 18232 14706 18244
rect 15286 18232 15292 18284
rect 15344 18272 15350 18284
rect 15933 18275 15991 18281
rect 15933 18272 15945 18275
rect 15344 18244 15945 18272
rect 15344 18232 15350 18244
rect 15933 18241 15945 18244
rect 15979 18241 15991 18275
rect 15933 18235 15991 18241
rect 13722 18204 13728 18216
rect 13683 18176 13728 18204
rect 13722 18164 13728 18176
rect 13780 18164 13786 18216
rect 13814 18164 13820 18216
rect 13872 18204 13878 18216
rect 16132 18213 16160 18312
rect 16408 18272 16436 18371
rect 17586 18368 17592 18420
rect 17644 18408 17650 18420
rect 18049 18411 18107 18417
rect 18049 18408 18061 18411
rect 17644 18380 18061 18408
rect 17644 18368 17650 18380
rect 18049 18377 18061 18380
rect 18095 18408 18107 18411
rect 19426 18408 19432 18420
rect 18095 18380 19432 18408
rect 18095 18377 18107 18380
rect 18049 18371 18107 18377
rect 19426 18368 19432 18380
rect 19484 18368 19490 18420
rect 19521 18411 19579 18417
rect 19521 18377 19533 18411
rect 19567 18408 19579 18411
rect 19610 18408 19616 18420
rect 19567 18380 19616 18408
rect 19567 18377 19579 18380
rect 19521 18371 19579 18377
rect 19610 18368 19616 18380
rect 19668 18408 19674 18420
rect 20622 18408 20628 18420
rect 19668 18380 20628 18408
rect 19668 18368 19674 18380
rect 20622 18368 20628 18380
rect 20680 18368 20686 18420
rect 21361 18411 21419 18417
rect 21361 18377 21373 18411
rect 21407 18377 21419 18411
rect 21361 18371 21419 18377
rect 21637 18411 21695 18417
rect 21637 18377 21649 18411
rect 21683 18408 21695 18411
rect 22281 18411 22339 18417
rect 22281 18408 22293 18411
rect 21683 18380 22293 18408
rect 21683 18377 21695 18380
rect 21637 18371 21695 18377
rect 22281 18377 22293 18380
rect 22327 18377 22339 18411
rect 22738 18408 22744 18420
rect 22699 18380 22744 18408
rect 22281 18371 22339 18377
rect 18408 18343 18466 18349
rect 16684 18312 18184 18340
rect 16684 18281 16712 18312
rect 16669 18275 16727 18281
rect 16669 18272 16681 18275
rect 16408 18244 16681 18272
rect 16669 18241 16681 18244
rect 16715 18241 16727 18275
rect 16669 18235 16727 18241
rect 16936 18275 16994 18281
rect 16936 18241 16948 18275
rect 16982 18272 16994 18275
rect 17218 18272 17224 18284
rect 16982 18244 17224 18272
rect 16982 18241 16994 18244
rect 16936 18235 16994 18241
rect 17218 18232 17224 18244
rect 17276 18272 17282 18284
rect 18156 18281 18184 18312
rect 18408 18309 18420 18343
rect 18454 18340 18466 18343
rect 18506 18340 18512 18352
rect 18454 18312 18512 18340
rect 18454 18309 18466 18312
rect 18408 18303 18466 18309
rect 18506 18300 18512 18312
rect 18564 18300 18570 18352
rect 18966 18300 18972 18352
rect 19024 18340 19030 18352
rect 20254 18340 20260 18352
rect 19024 18312 20260 18340
rect 19024 18300 19030 18312
rect 20254 18300 20260 18312
rect 20312 18300 20318 18352
rect 21266 18340 21272 18352
rect 20364 18312 21272 18340
rect 18141 18275 18199 18281
rect 17276 18244 18092 18272
rect 17276 18232 17282 18244
rect 16025 18207 16083 18213
rect 13872 18176 13917 18204
rect 13872 18164 13878 18176
rect 16025 18173 16037 18207
rect 16071 18173 16083 18207
rect 16025 18167 16083 18173
rect 16117 18207 16175 18213
rect 16117 18173 16129 18207
rect 16163 18173 16175 18207
rect 18064 18204 18092 18244
rect 18141 18241 18153 18275
rect 18187 18241 18199 18275
rect 18141 18235 18199 18241
rect 19242 18232 19248 18284
rect 19300 18272 19306 18284
rect 19613 18275 19671 18281
rect 19613 18272 19625 18275
rect 19300 18244 19625 18272
rect 19300 18232 19306 18244
rect 19613 18241 19625 18244
rect 19659 18241 19671 18275
rect 19613 18235 19671 18241
rect 19702 18232 19708 18284
rect 19760 18272 19766 18284
rect 19880 18275 19938 18281
rect 19880 18272 19892 18275
rect 19760 18244 19892 18272
rect 19760 18232 19766 18244
rect 19880 18241 19892 18244
rect 19926 18272 19938 18275
rect 20364 18272 20392 18312
rect 21266 18300 21272 18312
rect 21324 18300 21330 18352
rect 21376 18340 21404 18371
rect 22738 18368 22744 18380
rect 22796 18368 22802 18420
rect 23014 18408 23020 18420
rect 22975 18380 23020 18408
rect 23014 18368 23020 18380
rect 23072 18368 23078 18420
rect 22189 18343 22247 18349
rect 22189 18340 22201 18343
rect 21376 18312 22201 18340
rect 22189 18309 22201 18312
rect 22235 18309 22247 18343
rect 22189 18303 22247 18309
rect 21174 18272 21180 18284
rect 19926 18244 20392 18272
rect 21135 18244 21180 18272
rect 19926 18241 19938 18244
rect 19880 18235 19938 18241
rect 21174 18232 21180 18244
rect 21232 18232 21238 18284
rect 21450 18272 21456 18284
rect 21411 18244 21456 18272
rect 21450 18232 21456 18244
rect 21508 18232 21514 18284
rect 22830 18272 22836 18284
rect 22791 18244 22836 18272
rect 22830 18232 22836 18244
rect 22888 18232 22894 18284
rect 22186 18204 22192 18216
rect 18064 18176 18184 18204
rect 16117 18167 16175 18173
rect 13170 18096 13176 18148
rect 13228 18136 13234 18148
rect 13265 18139 13323 18145
rect 13265 18136 13277 18139
rect 13228 18108 13277 18136
rect 13228 18096 13234 18108
rect 13265 18105 13277 18108
rect 13311 18105 13323 18139
rect 13265 18099 13323 18105
rect 13630 18096 13636 18148
rect 13688 18136 13694 18148
rect 16040 18136 16068 18167
rect 13688 18108 14044 18136
rect 13688 18096 13694 18108
rect 6227 18040 7788 18068
rect 6227 18037 6239 18040
rect 6181 18031 6239 18037
rect 8570 18028 8576 18080
rect 8628 18068 8634 18080
rect 9214 18068 9220 18080
rect 8628 18040 9220 18068
rect 8628 18028 8634 18040
rect 9214 18028 9220 18040
rect 9272 18068 9278 18080
rect 9585 18071 9643 18077
rect 9585 18068 9597 18071
rect 9272 18040 9597 18068
rect 9272 18028 9278 18040
rect 9585 18037 9597 18040
rect 9631 18037 9643 18071
rect 9585 18031 9643 18037
rect 9674 18028 9680 18080
rect 9732 18068 9738 18080
rect 11609 18071 11667 18077
rect 11609 18068 11621 18071
rect 9732 18040 11621 18068
rect 9732 18028 9738 18040
rect 11609 18037 11621 18040
rect 11655 18068 11667 18071
rect 13906 18068 13912 18080
rect 11655 18040 13912 18068
rect 11655 18037 11667 18040
rect 11609 18031 11667 18037
rect 13906 18028 13912 18040
rect 13964 18028 13970 18080
rect 14016 18068 14044 18108
rect 15028 18108 16068 18136
rect 14274 18068 14280 18080
rect 14016 18040 14280 18068
rect 14274 18028 14280 18040
rect 14332 18028 14338 18080
rect 14366 18028 14372 18080
rect 14424 18068 14430 18080
rect 15028 18068 15056 18108
rect 14424 18040 15056 18068
rect 15473 18071 15531 18077
rect 14424 18028 14430 18040
rect 15473 18037 15485 18071
rect 15519 18068 15531 18071
rect 15930 18068 15936 18080
rect 15519 18040 15936 18068
rect 15519 18037 15531 18040
rect 15473 18031 15531 18037
rect 15930 18028 15936 18040
rect 15988 18028 15994 18080
rect 18156 18068 18184 18176
rect 20640 18176 22192 18204
rect 19076 18108 19656 18136
rect 19076 18068 19104 18108
rect 18156 18040 19104 18068
rect 19628 18068 19656 18108
rect 20640 18068 20668 18176
rect 22186 18164 22192 18176
rect 22244 18164 22250 18216
rect 22370 18204 22376 18216
rect 22331 18176 22376 18204
rect 22370 18164 22376 18176
rect 22428 18164 22434 18216
rect 20714 18096 20720 18148
rect 20772 18136 20778 18148
rect 22462 18136 22468 18148
rect 20772 18108 22468 18136
rect 20772 18096 20778 18108
rect 22462 18096 22468 18108
rect 22520 18096 22526 18148
rect 20990 18068 20996 18080
rect 19628 18040 20668 18068
rect 20951 18040 20996 18068
rect 20990 18028 20996 18040
rect 21048 18028 21054 18080
rect 21821 18071 21879 18077
rect 21821 18037 21833 18071
rect 21867 18068 21879 18071
rect 22094 18068 22100 18080
rect 21867 18040 22100 18068
rect 21867 18037 21879 18040
rect 21821 18031 21879 18037
rect 22094 18028 22100 18040
rect 22152 18028 22158 18080
rect 22186 18028 22192 18080
rect 22244 18068 22250 18080
rect 22554 18068 22560 18080
rect 22244 18040 22560 18068
rect 22244 18028 22250 18040
rect 22554 18028 22560 18040
rect 22612 18028 22618 18080
rect 1104 17978 23460 18000
rect 1104 17926 3749 17978
rect 3801 17926 3813 17978
rect 3865 17926 3877 17978
rect 3929 17926 3941 17978
rect 3993 17926 4005 17978
rect 4057 17926 9347 17978
rect 9399 17926 9411 17978
rect 9463 17926 9475 17978
rect 9527 17926 9539 17978
rect 9591 17926 9603 17978
rect 9655 17926 14945 17978
rect 14997 17926 15009 17978
rect 15061 17926 15073 17978
rect 15125 17926 15137 17978
rect 15189 17926 15201 17978
rect 15253 17926 20543 17978
rect 20595 17926 20607 17978
rect 20659 17926 20671 17978
rect 20723 17926 20735 17978
rect 20787 17926 20799 17978
rect 20851 17926 23460 17978
rect 1104 17904 23460 17926
rect 1946 17864 1952 17876
rect 1907 17836 1952 17864
rect 1946 17824 1952 17836
rect 2004 17824 2010 17876
rect 2869 17867 2927 17873
rect 2869 17833 2881 17867
rect 2915 17864 2927 17867
rect 3326 17864 3332 17876
rect 2915 17836 3332 17864
rect 2915 17833 2927 17836
rect 2869 17827 2927 17833
rect 3326 17824 3332 17836
rect 3384 17824 3390 17876
rect 3418 17824 3424 17876
rect 3476 17864 3482 17876
rect 3789 17867 3847 17873
rect 3789 17864 3801 17867
rect 3476 17836 3801 17864
rect 3476 17824 3482 17836
rect 3789 17833 3801 17836
rect 3835 17833 3847 17867
rect 5534 17864 5540 17876
rect 3789 17827 3847 17833
rect 3896 17836 5540 17864
rect 3896 17796 3924 17836
rect 5534 17824 5540 17836
rect 5592 17824 5598 17876
rect 7190 17824 7196 17876
rect 7248 17864 7254 17876
rect 7469 17867 7527 17873
rect 7469 17864 7481 17867
rect 7248 17836 7481 17864
rect 7248 17824 7254 17836
rect 7469 17833 7481 17836
rect 7515 17833 7527 17867
rect 7469 17827 7527 17833
rect 9030 17824 9036 17876
rect 9088 17864 9094 17876
rect 9493 17867 9551 17873
rect 9493 17864 9505 17867
rect 9088 17836 9505 17864
rect 9088 17824 9094 17836
rect 9493 17833 9505 17836
rect 9539 17833 9551 17867
rect 10962 17864 10968 17876
rect 10923 17836 10968 17864
rect 9493 17827 9551 17833
rect 10962 17824 10968 17836
rect 11020 17824 11026 17876
rect 12526 17824 12532 17876
rect 12584 17864 12590 17876
rect 12713 17867 12771 17873
rect 12713 17864 12725 17867
rect 12584 17836 12725 17864
rect 12584 17824 12590 17836
rect 12713 17833 12725 17836
rect 12759 17833 12771 17867
rect 13906 17864 13912 17876
rect 13867 17836 13912 17864
rect 12713 17827 12771 17833
rect 13906 17824 13912 17836
rect 13964 17824 13970 17876
rect 15194 17864 15200 17876
rect 14108 17836 15200 17864
rect 3344 17768 3924 17796
rect 2130 17688 2136 17740
rect 2188 17728 2194 17740
rect 3344 17737 3372 17768
rect 4154 17756 4160 17808
rect 4212 17796 4218 17808
rect 13725 17799 13783 17805
rect 4212 17768 4476 17796
rect 4212 17756 4218 17768
rect 2593 17731 2651 17737
rect 2593 17728 2605 17731
rect 2188 17700 2605 17728
rect 2188 17688 2194 17700
rect 2593 17697 2605 17700
rect 2639 17697 2651 17731
rect 2593 17691 2651 17697
rect 3329 17731 3387 17737
rect 3329 17697 3341 17731
rect 3375 17697 3387 17731
rect 3510 17728 3516 17740
rect 3471 17700 3516 17728
rect 3329 17691 3387 17697
rect 3510 17688 3516 17700
rect 3568 17688 3574 17740
rect 4246 17728 4252 17740
rect 4207 17700 4252 17728
rect 4246 17688 4252 17700
rect 4304 17688 4310 17740
rect 4448 17737 4476 17768
rect 13725 17765 13737 17799
rect 13771 17796 13783 17799
rect 14108 17796 14136 17836
rect 15194 17824 15200 17836
rect 15252 17824 15258 17876
rect 15470 17864 15476 17876
rect 15431 17836 15476 17864
rect 15470 17824 15476 17836
rect 15528 17824 15534 17876
rect 15746 17864 15752 17876
rect 15580 17836 15752 17864
rect 13771 17768 14136 17796
rect 13771 17765 13783 17768
rect 13725 17759 13783 17765
rect 4433 17731 4491 17737
rect 4433 17697 4445 17731
rect 4479 17728 4491 17731
rect 4522 17728 4528 17740
rect 4479 17700 4528 17728
rect 4479 17697 4491 17700
rect 4433 17691 4491 17697
rect 4522 17688 4528 17700
rect 4580 17688 4586 17740
rect 13357 17731 13415 17737
rect 13357 17697 13369 17731
rect 13403 17728 13415 17731
rect 13446 17728 13452 17740
rect 13403 17700 13452 17728
rect 13403 17697 13415 17700
rect 13357 17691 13415 17697
rect 13446 17688 13452 17700
rect 13504 17688 13510 17740
rect 15580 17737 15608 17836
rect 15746 17824 15752 17836
rect 15804 17824 15810 17876
rect 16942 17864 16948 17876
rect 16903 17836 16948 17864
rect 16942 17824 16948 17836
rect 17000 17824 17006 17876
rect 17034 17824 17040 17876
rect 17092 17864 17098 17876
rect 20346 17864 20352 17876
rect 17092 17836 20352 17864
rect 17092 17824 17098 17836
rect 20346 17824 20352 17836
rect 20404 17824 20410 17876
rect 20438 17824 20444 17876
rect 20496 17864 20502 17876
rect 20625 17867 20683 17873
rect 20625 17864 20637 17867
rect 20496 17836 20637 17864
rect 20496 17824 20502 17836
rect 20625 17833 20637 17836
rect 20671 17864 20683 17867
rect 21082 17864 21088 17876
rect 20671 17836 21088 17864
rect 20671 17833 20683 17836
rect 20625 17827 20683 17833
rect 21082 17824 21088 17836
rect 21140 17824 21146 17876
rect 21726 17824 21732 17876
rect 21784 17864 21790 17876
rect 21784 17836 22968 17864
rect 21784 17824 21790 17836
rect 19058 17796 19064 17808
rect 19019 17768 19064 17796
rect 19058 17756 19064 17768
rect 19116 17756 19122 17808
rect 21453 17799 21511 17805
rect 21453 17765 21465 17799
rect 21499 17796 21511 17799
rect 21499 17768 22876 17796
rect 21499 17765 21511 17768
rect 21453 17759 21511 17765
rect 15565 17731 15623 17737
rect 15565 17697 15577 17731
rect 15611 17697 15623 17731
rect 15565 17691 15623 17697
rect 1765 17663 1823 17669
rect 1765 17629 1777 17663
rect 1811 17660 1823 17663
rect 1811 17632 2084 17660
rect 1811 17629 1823 17632
rect 1765 17623 1823 17629
rect 2056 17533 2084 17632
rect 2222 17620 2228 17672
rect 2280 17660 2286 17672
rect 2409 17663 2467 17669
rect 2409 17660 2421 17663
rect 2280 17632 2421 17660
rect 2280 17620 2286 17632
rect 2409 17629 2421 17632
rect 2455 17629 2467 17663
rect 2409 17623 2467 17629
rect 3237 17663 3295 17669
rect 3237 17629 3249 17663
rect 3283 17660 3295 17663
rect 4338 17660 4344 17672
rect 3283 17632 4344 17660
rect 3283 17629 3295 17632
rect 3237 17623 3295 17629
rect 4338 17620 4344 17632
rect 4396 17620 4402 17672
rect 4617 17663 4675 17669
rect 4617 17629 4629 17663
rect 4663 17660 4675 17663
rect 6089 17663 6147 17669
rect 6089 17660 6101 17663
rect 4663 17632 6101 17660
rect 4663 17629 4675 17632
rect 4617 17623 4675 17629
rect 6089 17629 6101 17632
rect 6135 17660 6147 17663
rect 6178 17660 6184 17672
rect 6135 17632 6184 17660
rect 6135 17629 6147 17632
rect 6089 17623 6147 17629
rect 6178 17620 6184 17632
rect 6236 17620 6242 17672
rect 10617 17663 10675 17669
rect 10617 17629 10629 17663
rect 10663 17660 10675 17663
rect 10778 17660 10784 17672
rect 10663 17632 10784 17660
rect 10663 17629 10675 17632
rect 10617 17623 10675 17629
rect 10778 17620 10784 17632
rect 10836 17620 10842 17672
rect 10873 17663 10931 17669
rect 10873 17629 10885 17663
rect 10919 17660 10931 17663
rect 12345 17663 12403 17669
rect 12345 17660 12357 17663
rect 10919 17632 12357 17660
rect 10919 17629 10931 17632
rect 10873 17623 10931 17629
rect 12345 17629 12357 17632
rect 12391 17660 12403 17663
rect 14093 17663 14151 17669
rect 12391 17632 12480 17660
rect 12391 17629 12403 17632
rect 12345 17623 12403 17629
rect 3142 17552 3148 17604
rect 3200 17592 3206 17604
rect 6362 17601 6368 17604
rect 4862 17595 4920 17601
rect 4862 17592 4874 17595
rect 3200 17564 4874 17592
rect 3200 17552 3206 17564
rect 4862 17561 4874 17564
rect 4908 17561 4920 17595
rect 4862 17555 4920 17561
rect 5920 17564 6316 17592
rect 2041 17527 2099 17533
rect 2041 17493 2053 17527
rect 2087 17493 2099 17527
rect 2041 17487 2099 17493
rect 2501 17527 2559 17533
rect 2501 17493 2513 17527
rect 2547 17524 2559 17527
rect 2682 17524 2688 17536
rect 2547 17496 2688 17524
rect 2547 17493 2559 17496
rect 2501 17487 2559 17493
rect 2682 17484 2688 17496
rect 2740 17484 2746 17536
rect 4157 17527 4215 17533
rect 4157 17493 4169 17527
rect 4203 17524 4215 17527
rect 4430 17524 4436 17536
rect 4203 17496 4436 17524
rect 4203 17493 4215 17496
rect 4157 17487 4215 17493
rect 4430 17484 4436 17496
rect 4488 17524 4494 17536
rect 5920 17524 5948 17564
rect 4488 17496 5948 17524
rect 4488 17484 4494 17496
rect 5994 17484 6000 17536
rect 6052 17524 6058 17536
rect 6288 17524 6316 17564
rect 6356 17555 6368 17601
rect 6420 17592 6426 17604
rect 12078 17595 12136 17601
rect 12078 17592 12090 17595
rect 6420 17564 6456 17592
rect 6932 17564 12090 17592
rect 6362 17552 6368 17555
rect 6420 17552 6426 17564
rect 6932 17524 6960 17564
rect 12078 17561 12090 17564
rect 12124 17561 12136 17595
rect 12452 17592 12480 17632
rect 14093 17629 14105 17663
rect 14139 17660 14151 17663
rect 14182 17660 14188 17672
rect 14139 17632 14188 17660
rect 14139 17629 14151 17632
rect 14093 17623 14151 17629
rect 14182 17620 14188 17632
rect 14240 17660 14246 17672
rect 15580 17660 15608 17691
rect 18414 17688 18420 17740
rect 18472 17728 18478 17740
rect 19242 17728 19248 17740
rect 18472 17700 19248 17728
rect 18472 17688 18478 17700
rect 19242 17688 19248 17700
rect 19300 17688 19306 17740
rect 20901 17731 20959 17737
rect 20901 17697 20913 17731
rect 20947 17728 20959 17731
rect 21542 17728 21548 17740
rect 20947 17700 21548 17728
rect 20947 17697 20959 17700
rect 20901 17691 20959 17697
rect 21542 17688 21548 17700
rect 21600 17728 21606 17740
rect 21637 17731 21695 17737
rect 21637 17728 21649 17731
rect 21600 17700 21649 17728
rect 21600 17688 21606 17700
rect 21637 17697 21649 17700
rect 21683 17728 21695 17731
rect 22646 17728 22652 17740
rect 21683 17700 22652 17728
rect 21683 17697 21695 17700
rect 21637 17691 21695 17697
rect 22646 17688 22652 17700
rect 22704 17688 22710 17740
rect 22848 17737 22876 17768
rect 22940 17740 22968 17836
rect 22833 17731 22891 17737
rect 22833 17697 22845 17731
rect 22879 17697 22891 17731
rect 22833 17691 22891 17697
rect 22922 17688 22928 17740
rect 22980 17728 22986 17740
rect 22980 17700 23073 17728
rect 22980 17688 22986 17700
rect 15838 17669 15844 17672
rect 15832 17660 15844 17669
rect 14240 17632 15608 17660
rect 15799 17632 15844 17660
rect 14240 17620 14246 17632
rect 15832 17623 15844 17632
rect 15838 17620 15844 17623
rect 15896 17620 15902 17672
rect 18138 17620 18144 17672
rect 18196 17669 18202 17672
rect 18196 17660 18208 17669
rect 18601 17663 18659 17669
rect 18196 17632 18241 17660
rect 18196 17623 18208 17632
rect 18601 17629 18613 17663
rect 18647 17629 18659 17663
rect 18874 17660 18880 17672
rect 18835 17632 18880 17660
rect 18601 17623 18659 17629
rect 18196 17620 18202 17623
rect 12452 17564 12572 17592
rect 12078 17555 12136 17561
rect 12544 17536 12572 17564
rect 13998 17552 14004 17604
rect 14056 17592 14062 17604
rect 14360 17595 14418 17601
rect 14360 17592 14372 17595
rect 14056 17564 14372 17592
rect 14056 17552 14062 17564
rect 14360 17561 14372 17564
rect 14406 17592 14418 17595
rect 15378 17592 15384 17604
rect 14406 17564 15384 17592
rect 14406 17561 14418 17564
rect 14360 17555 14418 17561
rect 15378 17552 15384 17564
rect 15436 17552 15442 17604
rect 16022 17552 16028 17604
rect 16080 17592 16086 17604
rect 18506 17592 18512 17604
rect 16080 17564 18512 17592
rect 16080 17552 16086 17564
rect 18506 17552 18512 17564
rect 18564 17552 18570 17604
rect 18616 17592 18644 17623
rect 18874 17620 18880 17632
rect 18932 17620 18938 17672
rect 20990 17620 20996 17672
rect 21048 17620 21054 17672
rect 21082 17620 21088 17672
rect 21140 17660 21146 17672
rect 21140 17632 21185 17660
rect 21140 17620 21146 17632
rect 21266 17620 21272 17672
rect 21324 17660 21330 17672
rect 21821 17663 21879 17669
rect 21821 17660 21833 17663
rect 21324 17632 21833 17660
rect 21324 17620 21330 17632
rect 21821 17629 21833 17632
rect 21867 17629 21879 17663
rect 21821 17623 21879 17629
rect 19334 17592 19340 17604
rect 18616 17564 19340 17592
rect 19334 17552 19340 17564
rect 19392 17552 19398 17604
rect 19512 17595 19570 17601
rect 19512 17561 19524 17595
rect 19558 17592 19570 17595
rect 19794 17592 19800 17604
rect 19558 17564 19800 17592
rect 19558 17561 19570 17564
rect 19512 17555 19570 17561
rect 19794 17552 19800 17564
rect 19852 17592 19858 17604
rect 21008 17592 21036 17620
rect 21913 17595 21971 17601
rect 21913 17592 21925 17595
rect 19852 17564 20852 17592
rect 21008 17564 21925 17592
rect 19852 17552 19858 17564
rect 6052 17496 6097 17524
rect 6288 17496 6960 17524
rect 7653 17527 7711 17533
rect 6052 17484 6058 17496
rect 7653 17493 7665 17527
rect 7699 17524 7711 17527
rect 8205 17527 8263 17533
rect 8205 17524 8217 17527
rect 7699 17496 8217 17524
rect 7699 17493 7711 17496
rect 7653 17487 7711 17493
rect 8205 17493 8217 17496
rect 8251 17524 8263 17527
rect 8294 17524 8300 17536
rect 8251 17496 8300 17524
rect 8251 17493 8263 17496
rect 8205 17487 8263 17493
rect 8294 17484 8300 17496
rect 8352 17524 8358 17536
rect 8478 17524 8484 17536
rect 8352 17496 8484 17524
rect 8352 17484 8358 17496
rect 8478 17484 8484 17496
rect 8536 17484 8542 17536
rect 12526 17524 12532 17536
rect 12487 17496 12532 17524
rect 12526 17484 12532 17496
rect 12584 17484 12590 17536
rect 13078 17524 13084 17536
rect 13039 17496 13084 17524
rect 13078 17484 13084 17496
rect 13136 17484 13142 17536
rect 13173 17527 13231 17533
rect 13173 17493 13185 17527
rect 13219 17524 13231 17527
rect 13354 17524 13360 17536
rect 13219 17496 13360 17524
rect 13219 17493 13231 17496
rect 13173 17487 13231 17493
rect 13354 17484 13360 17496
rect 13412 17484 13418 17536
rect 14274 17484 14280 17536
rect 14332 17524 14338 17536
rect 14642 17524 14648 17536
rect 14332 17496 14648 17524
rect 14332 17484 14338 17496
rect 14642 17484 14648 17496
rect 14700 17484 14706 17536
rect 15194 17484 15200 17536
rect 15252 17524 15258 17536
rect 15562 17524 15568 17536
rect 15252 17496 15568 17524
rect 15252 17484 15258 17496
rect 15562 17484 15568 17496
rect 15620 17484 15626 17536
rect 17037 17527 17095 17533
rect 17037 17493 17049 17527
rect 17083 17524 17095 17527
rect 17218 17524 17224 17536
rect 17083 17496 17224 17524
rect 17083 17493 17095 17496
rect 17037 17487 17095 17493
rect 17218 17484 17224 17496
rect 17276 17484 17282 17536
rect 18785 17527 18843 17533
rect 18785 17493 18797 17527
rect 18831 17524 18843 17527
rect 20714 17524 20720 17536
rect 18831 17496 20720 17524
rect 18831 17493 18843 17496
rect 18785 17487 18843 17493
rect 20714 17484 20720 17496
rect 20772 17484 20778 17536
rect 20824 17524 20852 17564
rect 21913 17561 21925 17564
rect 21959 17561 21971 17595
rect 22741 17595 22799 17601
rect 22741 17592 22753 17595
rect 21913 17555 21971 17561
rect 22296 17564 22753 17592
rect 22296 17533 22324 17564
rect 22741 17561 22753 17564
rect 22787 17561 22799 17595
rect 22741 17555 22799 17561
rect 20993 17527 21051 17533
rect 20993 17524 21005 17527
rect 20824 17496 21005 17524
rect 20993 17493 21005 17496
rect 21039 17493 21051 17527
rect 20993 17487 21051 17493
rect 22281 17527 22339 17533
rect 22281 17493 22293 17527
rect 22327 17493 22339 17527
rect 22281 17487 22339 17493
rect 22373 17527 22431 17533
rect 22373 17493 22385 17527
rect 22419 17524 22431 17527
rect 22646 17524 22652 17536
rect 22419 17496 22652 17524
rect 22419 17493 22431 17496
rect 22373 17487 22431 17493
rect 22646 17484 22652 17496
rect 22704 17484 22710 17536
rect 1104 17434 23460 17456
rect 1104 17382 6548 17434
rect 6600 17382 6612 17434
rect 6664 17382 6676 17434
rect 6728 17382 6740 17434
rect 6792 17382 6804 17434
rect 6856 17382 12146 17434
rect 12198 17382 12210 17434
rect 12262 17382 12274 17434
rect 12326 17382 12338 17434
rect 12390 17382 12402 17434
rect 12454 17382 17744 17434
rect 17796 17382 17808 17434
rect 17860 17382 17872 17434
rect 17924 17382 17936 17434
rect 17988 17382 18000 17434
rect 18052 17382 23460 17434
rect 1104 17360 23460 17382
rect 1854 17280 1860 17332
rect 1912 17320 1918 17332
rect 2130 17320 2136 17332
rect 1912 17292 2136 17320
rect 1912 17280 1918 17292
rect 2130 17280 2136 17292
rect 2188 17320 2194 17332
rect 2225 17323 2283 17329
rect 2225 17320 2237 17323
rect 2188 17292 2237 17320
rect 2188 17280 2194 17292
rect 2225 17289 2237 17292
rect 2271 17289 2283 17323
rect 2225 17283 2283 17289
rect 2590 17280 2596 17332
rect 2648 17320 2654 17332
rect 2685 17323 2743 17329
rect 2685 17320 2697 17323
rect 2648 17292 2697 17320
rect 2648 17280 2654 17292
rect 2685 17289 2697 17292
rect 2731 17289 2743 17323
rect 2685 17283 2743 17289
rect 3145 17323 3203 17329
rect 3145 17289 3157 17323
rect 3191 17320 3203 17323
rect 3234 17320 3240 17332
rect 3191 17292 3240 17320
rect 3191 17289 3203 17292
rect 3145 17283 3203 17289
rect 3234 17280 3240 17292
rect 3292 17280 3298 17332
rect 3605 17323 3663 17329
rect 3605 17289 3617 17323
rect 3651 17320 3663 17323
rect 5166 17320 5172 17332
rect 3651 17292 5172 17320
rect 3651 17289 3663 17292
rect 3605 17283 3663 17289
rect 5166 17280 5172 17292
rect 5224 17280 5230 17332
rect 8389 17323 8447 17329
rect 8389 17289 8401 17323
rect 8435 17320 8447 17323
rect 8846 17320 8852 17332
rect 8435 17292 8852 17320
rect 8435 17289 8447 17292
rect 8389 17283 8447 17289
rect 8846 17280 8852 17292
rect 8904 17280 8910 17332
rect 9861 17323 9919 17329
rect 9861 17289 9873 17323
rect 9907 17320 9919 17323
rect 10778 17320 10784 17332
rect 9907 17292 10784 17320
rect 9907 17289 9919 17292
rect 9861 17283 9919 17289
rect 10778 17280 10784 17292
rect 10836 17280 10842 17332
rect 12066 17280 12072 17332
rect 12124 17320 12130 17332
rect 12345 17323 12403 17329
rect 12345 17320 12357 17323
rect 12124 17292 12357 17320
rect 12124 17280 12130 17292
rect 12345 17289 12357 17292
rect 12391 17289 12403 17323
rect 12345 17283 12403 17289
rect 12526 17280 12532 17332
rect 12584 17320 12590 17332
rect 14182 17320 14188 17332
rect 12584 17292 14188 17320
rect 12584 17280 12590 17292
rect 4522 17212 4528 17264
rect 4580 17252 4586 17264
rect 6270 17252 6276 17264
rect 4580 17224 6276 17252
rect 4580 17212 4586 17224
rect 6270 17212 6276 17224
rect 6328 17212 6334 17264
rect 7276 17255 7334 17261
rect 7276 17221 7288 17255
rect 7322 17252 7334 17255
rect 8570 17252 8576 17264
rect 7322 17224 8576 17252
rect 7322 17221 7334 17224
rect 7276 17215 7334 17221
rect 8570 17212 8576 17224
rect 8628 17212 8634 17264
rect 8754 17261 8760 17264
rect 8748 17252 8760 17261
rect 8667 17224 8760 17252
rect 8748 17215 8760 17224
rect 8812 17252 8818 17264
rect 9122 17252 9128 17264
rect 8812 17224 9128 17252
rect 8754 17212 8760 17215
rect 8812 17212 8818 17224
rect 9122 17212 9128 17224
rect 9180 17212 9186 17264
rect 10220 17255 10278 17261
rect 10220 17221 10232 17255
rect 10266 17252 10278 17255
rect 10962 17252 10968 17264
rect 10266 17224 10968 17252
rect 10266 17221 10278 17224
rect 10220 17215 10278 17221
rect 10962 17212 10968 17224
rect 11020 17212 11026 17264
rect 11330 17212 11336 17264
rect 11388 17252 11394 17264
rect 11977 17255 12035 17261
rect 11977 17252 11989 17255
rect 11388 17224 11989 17252
rect 11388 17212 11394 17224
rect 11977 17221 11989 17224
rect 12023 17221 12035 17255
rect 11977 17215 12035 17221
rect 2866 17184 2872 17196
rect 2827 17156 2872 17184
rect 2866 17144 2872 17156
rect 2924 17144 2930 17196
rect 2961 17187 3019 17193
rect 2961 17153 2973 17187
rect 3007 17153 3019 17187
rect 2961 17147 3019 17153
rect 1854 17076 1860 17128
rect 1912 17116 1918 17128
rect 2317 17119 2375 17125
rect 2317 17116 2329 17119
rect 1912 17088 2329 17116
rect 1912 17076 1918 17088
rect 2317 17085 2329 17088
rect 2363 17085 2375 17119
rect 2498 17116 2504 17128
rect 2459 17088 2504 17116
rect 2317 17079 2375 17085
rect 2498 17076 2504 17088
rect 2556 17076 2562 17128
rect 2590 17076 2596 17128
rect 2648 17116 2654 17128
rect 2976 17116 3004 17147
rect 3142 17144 3148 17196
rect 3200 17184 3206 17196
rect 3697 17187 3755 17193
rect 3697 17184 3709 17187
rect 3200 17156 3709 17184
rect 3200 17144 3206 17156
rect 3697 17153 3709 17156
rect 3743 17153 3755 17187
rect 3697 17147 3755 17153
rect 4338 17144 4344 17196
rect 4396 17184 4402 17196
rect 5914 17187 5972 17193
rect 5914 17184 5926 17187
rect 4396 17156 5926 17184
rect 4396 17144 4402 17156
rect 5914 17153 5926 17156
rect 5960 17153 5972 17187
rect 5914 17147 5972 17153
rect 10502 17144 10508 17196
rect 10560 17184 10566 17196
rect 12636 17193 12664 17292
rect 14182 17280 14188 17292
rect 14240 17280 14246 17332
rect 14553 17323 14611 17329
rect 14553 17289 14565 17323
rect 14599 17320 14611 17323
rect 16022 17320 16028 17332
rect 14599 17292 16028 17320
rect 14599 17289 14611 17292
rect 14553 17283 14611 17289
rect 16022 17280 16028 17292
rect 16080 17280 16086 17332
rect 17126 17320 17132 17332
rect 16132 17292 17132 17320
rect 12888 17255 12946 17261
rect 12888 17221 12900 17255
rect 12934 17252 12946 17255
rect 13170 17252 13176 17264
rect 12934 17224 13176 17252
rect 12934 17221 12946 17224
rect 12888 17215 12946 17221
rect 13170 17212 13176 17224
rect 13228 17252 13234 17264
rect 13630 17252 13636 17264
rect 13228 17224 13636 17252
rect 13228 17212 13234 17224
rect 13630 17212 13636 17224
rect 13688 17212 13694 17264
rect 15780 17255 15838 17261
rect 15780 17221 15792 17255
rect 15826 17252 15838 17255
rect 16132 17252 16160 17292
rect 17126 17280 17132 17292
rect 17184 17280 17190 17332
rect 17310 17320 17316 17332
rect 17271 17292 17316 17320
rect 17310 17280 17316 17292
rect 17368 17280 17374 17332
rect 17402 17280 17408 17332
rect 17460 17320 17466 17332
rect 17589 17323 17647 17329
rect 17589 17320 17601 17323
rect 17460 17292 17601 17320
rect 17460 17280 17466 17292
rect 17589 17289 17601 17292
rect 17635 17289 17647 17323
rect 17589 17283 17647 17289
rect 17954 17280 17960 17332
rect 18012 17320 18018 17332
rect 18506 17320 18512 17332
rect 18012 17292 18512 17320
rect 18012 17280 18018 17292
rect 18506 17280 18512 17292
rect 18564 17280 18570 17332
rect 19429 17323 19487 17329
rect 19429 17289 19441 17323
rect 19475 17320 19487 17323
rect 21177 17323 21235 17329
rect 21177 17320 21189 17323
rect 19475 17292 21189 17320
rect 19475 17289 19487 17292
rect 19429 17283 19487 17289
rect 21177 17289 21189 17292
rect 21223 17289 21235 17323
rect 22370 17320 22376 17332
rect 21177 17283 21235 17289
rect 21928 17292 22376 17320
rect 15826 17224 16160 17252
rect 16209 17255 16267 17261
rect 15826 17221 15838 17224
rect 15780 17215 15838 17221
rect 16209 17221 16221 17255
rect 16255 17252 16267 17255
rect 16393 17255 16451 17261
rect 16393 17252 16405 17255
rect 16255 17224 16405 17252
rect 16255 17221 16267 17224
rect 16209 17215 16267 17221
rect 16393 17221 16405 17224
rect 16439 17252 16451 17255
rect 18414 17252 18420 17264
rect 16439 17224 18420 17252
rect 16439 17221 16451 17224
rect 16393 17215 16451 17221
rect 11885 17187 11943 17193
rect 11885 17184 11897 17187
rect 10560 17156 11897 17184
rect 10560 17144 10566 17156
rect 11885 17153 11897 17156
rect 11931 17153 11943 17187
rect 11885 17147 11943 17153
rect 12621 17187 12679 17193
rect 12621 17153 12633 17187
rect 12667 17153 12679 17187
rect 12621 17147 12679 17153
rect 16025 17187 16083 17193
rect 16025 17153 16037 17187
rect 16071 17184 16083 17187
rect 16224 17184 16252 17215
rect 16071 17156 16252 17184
rect 16853 17187 16911 17193
rect 16071 17153 16083 17156
rect 16025 17147 16083 17153
rect 16853 17153 16865 17187
rect 16899 17153 16911 17187
rect 16853 17147 16911 17153
rect 3510 17116 3516 17128
rect 2648 17088 3004 17116
rect 3471 17088 3516 17116
rect 2648 17076 2654 17088
rect 3510 17076 3516 17088
rect 3568 17076 3574 17128
rect 6181 17119 6239 17125
rect 6181 17085 6193 17119
rect 6227 17116 6239 17119
rect 7009 17119 7067 17125
rect 7009 17116 7021 17119
rect 6227 17088 7021 17116
rect 6227 17085 6239 17088
rect 6181 17079 6239 17085
rect 7009 17085 7021 17088
rect 7055 17085 7067 17119
rect 8478 17116 8484 17128
rect 8439 17088 8484 17116
rect 7009 17079 7067 17085
rect 2774 17008 2780 17060
rect 2832 17048 2838 17060
rect 4430 17048 4436 17060
rect 2832 17020 4436 17048
rect 2832 17008 2838 17020
rect 4430 17008 4436 17020
rect 4488 17008 4494 17060
rect 4709 17051 4767 17057
rect 4709 17017 4721 17051
rect 4755 17048 4767 17051
rect 4755 17020 5304 17048
rect 4755 17017 4767 17020
rect 4709 17011 4767 17017
rect 1762 16940 1768 16992
rect 1820 16980 1826 16992
rect 1857 16983 1915 16989
rect 1857 16980 1869 16983
rect 1820 16952 1869 16980
rect 1820 16940 1826 16952
rect 1857 16949 1869 16952
rect 1903 16949 1915 16983
rect 1857 16943 1915 16949
rect 4065 16983 4123 16989
rect 4065 16949 4077 16983
rect 4111 16980 4123 16983
rect 4246 16980 4252 16992
rect 4111 16952 4252 16980
rect 4111 16949 4123 16952
rect 4065 16943 4123 16949
rect 4246 16940 4252 16952
rect 4304 16940 4310 16992
rect 4801 16983 4859 16989
rect 4801 16949 4813 16983
rect 4847 16980 4859 16983
rect 5166 16980 5172 16992
rect 4847 16952 5172 16980
rect 4847 16949 4859 16952
rect 4801 16943 4859 16949
rect 5166 16940 5172 16952
rect 5224 16940 5230 16992
rect 5276 16980 5304 17020
rect 6196 16992 6224 17079
rect 8478 17076 8484 17088
rect 8536 17076 8542 17128
rect 9766 17076 9772 17128
rect 9824 17116 9830 17128
rect 9953 17119 10011 17125
rect 9953 17116 9965 17119
rect 9824 17088 9965 17116
rect 9824 17076 9830 17088
rect 9953 17085 9965 17088
rect 9999 17085 10011 17119
rect 11790 17116 11796 17128
rect 11751 17088 11796 17116
rect 9953 17079 10011 17085
rect 11790 17076 11796 17088
rect 11848 17076 11854 17128
rect 11333 17051 11391 17057
rect 11333 17017 11345 17051
rect 11379 17048 11391 17051
rect 11379 17020 12434 17048
rect 11379 17017 11391 17020
rect 11333 17011 11391 17017
rect 6178 16980 6184 16992
rect 5276 16952 6184 16980
rect 6178 16940 6184 16952
rect 6236 16980 6242 16992
rect 6365 16983 6423 16989
rect 6365 16980 6377 16983
rect 6236 16952 6377 16980
rect 6236 16940 6242 16952
rect 6365 16949 6377 16952
rect 6411 16949 6423 16983
rect 12406 16980 12434 17020
rect 13722 17008 13728 17060
rect 13780 17048 13786 17060
rect 14645 17051 14703 17057
rect 14645 17048 14657 17051
rect 13780 17020 14657 17048
rect 13780 17008 13786 17020
rect 14645 17017 14657 17020
rect 14691 17017 14703 17051
rect 16868 17048 16896 17147
rect 16942 17144 16948 17196
rect 17000 17184 17006 17196
rect 17129 17187 17187 17193
rect 17129 17184 17141 17187
rect 17000 17156 17141 17184
rect 17000 17144 17006 17156
rect 17129 17153 17141 17156
rect 17175 17153 17187 17187
rect 17129 17147 17187 17153
rect 17405 17187 17463 17193
rect 17405 17153 17417 17187
rect 17451 17184 17463 17187
rect 17586 17184 17592 17196
rect 17451 17156 17592 17184
rect 17451 17153 17463 17156
rect 17405 17147 17463 17153
rect 17586 17144 17592 17156
rect 17644 17144 17650 17196
rect 17681 17187 17739 17193
rect 17681 17153 17693 17187
rect 17727 17184 17739 17187
rect 17862 17184 17868 17196
rect 17727 17156 17868 17184
rect 17727 17153 17739 17156
rect 17681 17147 17739 17153
rect 17862 17144 17868 17156
rect 17920 17144 17926 17196
rect 17972 17193 18000 17224
rect 18414 17212 18420 17224
rect 18472 17212 18478 17264
rect 17957 17187 18015 17193
rect 17957 17153 17969 17187
rect 18003 17153 18015 17187
rect 17957 17147 18015 17153
rect 18224 17187 18282 17193
rect 18224 17153 18236 17187
rect 18270 17184 18282 17187
rect 19444 17184 19472 17283
rect 20564 17255 20622 17261
rect 20564 17221 20576 17255
rect 20610 17252 20622 17255
rect 20990 17252 20996 17264
rect 20610 17224 20996 17252
rect 20610 17221 20622 17224
rect 20564 17215 20622 17221
rect 20990 17212 20996 17224
rect 21048 17212 21054 17264
rect 18270 17156 19472 17184
rect 18270 17153 18282 17156
rect 18224 17147 18282 17153
rect 20714 17144 20720 17196
rect 20772 17184 20778 17196
rect 20772 17156 21220 17184
rect 20772 17144 20778 17156
rect 20809 17119 20867 17125
rect 20809 17085 20821 17119
rect 20855 17116 20867 17119
rect 20898 17116 20904 17128
rect 20855 17088 20904 17116
rect 20855 17085 20867 17088
rect 20809 17079 20867 17085
rect 20898 17076 20904 17088
rect 20956 17076 20962 17128
rect 21082 17116 21088 17128
rect 21043 17088 21088 17116
rect 21082 17076 21088 17088
rect 21140 17076 21146 17128
rect 21192 17116 21220 17156
rect 21266 17144 21272 17196
rect 21324 17184 21330 17196
rect 21324 17156 21369 17184
rect 21324 17144 21330 17156
rect 21928 17125 21956 17292
rect 22370 17280 22376 17292
rect 22428 17280 22434 17332
rect 22741 17323 22799 17329
rect 22741 17289 22753 17323
rect 22787 17320 22799 17323
rect 22922 17320 22928 17332
rect 22787 17292 22928 17320
rect 22787 17289 22799 17292
rect 22741 17283 22799 17289
rect 22922 17280 22928 17292
rect 22980 17280 22986 17332
rect 22186 17184 22192 17196
rect 22147 17156 22192 17184
rect 22186 17144 22192 17156
rect 22244 17144 22250 17196
rect 22833 17187 22891 17193
rect 22833 17184 22845 17187
rect 22480 17156 22845 17184
rect 21913 17119 21971 17125
rect 21913 17116 21925 17119
rect 21192 17088 21925 17116
rect 21913 17085 21925 17088
rect 21959 17085 21971 17119
rect 21913 17079 21971 17085
rect 22097 17119 22155 17125
rect 22097 17085 22109 17119
rect 22143 17116 22155 17119
rect 22370 17116 22376 17128
rect 22143 17088 22376 17116
rect 22143 17085 22155 17088
rect 22097 17079 22155 17085
rect 22370 17076 22376 17088
rect 22428 17076 22434 17128
rect 17402 17048 17408 17060
rect 16868 17020 17408 17048
rect 14645 17011 14703 17017
rect 17402 17008 17408 17020
rect 17460 17008 17466 17060
rect 22480 17048 22508 17156
rect 22833 17153 22845 17156
rect 22879 17153 22891 17187
rect 22833 17147 22891 17153
rect 22738 17076 22744 17128
rect 22796 17116 22802 17128
rect 23017 17119 23075 17125
rect 23017 17116 23029 17119
rect 22796 17088 23029 17116
rect 22796 17076 22802 17088
rect 23017 17085 23029 17088
rect 23063 17085 23075 17119
rect 23017 17079 23075 17085
rect 19260 17020 19932 17048
rect 12802 16980 12808 16992
rect 12406 16952 12808 16980
rect 6365 16943 6423 16949
rect 12802 16940 12808 16952
rect 12860 16940 12866 16992
rect 13998 16980 14004 16992
rect 13959 16952 14004 16980
rect 13998 16940 14004 16952
rect 14056 16940 14062 16992
rect 16758 16980 16764 16992
rect 16719 16952 16764 16980
rect 16758 16940 16764 16952
rect 16816 16940 16822 16992
rect 17034 16980 17040 16992
rect 16995 16952 17040 16980
rect 17034 16940 17040 16952
rect 17092 16940 17098 16992
rect 17865 16983 17923 16989
rect 17865 16949 17877 16983
rect 17911 16980 17923 16983
rect 19260 16980 19288 17020
rect 17911 16952 19288 16980
rect 17911 16949 17923 16952
rect 17865 16943 17923 16949
rect 19334 16940 19340 16992
rect 19392 16980 19398 16992
rect 19904 16980 19932 17020
rect 20824 17020 22508 17048
rect 20824 16980 20852 17020
rect 21634 16980 21640 16992
rect 19392 16952 19437 16980
rect 19904 16952 20852 16980
rect 21595 16952 21640 16980
rect 19392 16940 19398 16952
rect 21634 16940 21640 16952
rect 21692 16940 21698 16992
rect 22554 16980 22560 16992
rect 22515 16952 22560 16980
rect 22554 16940 22560 16952
rect 22612 16940 22618 16992
rect 1104 16890 23460 16912
rect 1104 16838 3749 16890
rect 3801 16838 3813 16890
rect 3865 16838 3877 16890
rect 3929 16838 3941 16890
rect 3993 16838 4005 16890
rect 4057 16838 9347 16890
rect 9399 16838 9411 16890
rect 9463 16838 9475 16890
rect 9527 16838 9539 16890
rect 9591 16838 9603 16890
rect 9655 16838 14945 16890
rect 14997 16838 15009 16890
rect 15061 16838 15073 16890
rect 15125 16838 15137 16890
rect 15189 16838 15201 16890
rect 15253 16838 20543 16890
rect 20595 16838 20607 16890
rect 20659 16838 20671 16890
rect 20723 16838 20735 16890
rect 20787 16838 20799 16890
rect 20851 16838 23460 16890
rect 1104 16816 23460 16838
rect 2866 16736 2872 16788
rect 2924 16776 2930 16788
rect 3789 16779 3847 16785
rect 3789 16776 3801 16779
rect 2924 16748 3801 16776
rect 2924 16736 2930 16748
rect 3789 16745 3801 16748
rect 3835 16745 3847 16779
rect 3789 16739 3847 16745
rect 4982 16736 4988 16788
rect 5040 16776 5046 16788
rect 5718 16776 5724 16788
rect 5040 16748 5724 16776
rect 5040 16736 5046 16748
rect 5718 16736 5724 16748
rect 5776 16736 5782 16788
rect 8754 16776 8760 16788
rect 8715 16748 8760 16776
rect 8754 16736 8760 16748
rect 8812 16736 8818 16788
rect 16669 16779 16727 16785
rect 16669 16745 16681 16779
rect 16715 16776 16727 16779
rect 17126 16776 17132 16788
rect 16715 16748 17132 16776
rect 16715 16745 16727 16748
rect 16669 16739 16727 16745
rect 17126 16736 17132 16748
rect 17184 16736 17190 16788
rect 18233 16779 18291 16785
rect 18233 16745 18245 16779
rect 18279 16776 18291 16779
rect 18414 16776 18420 16788
rect 18279 16748 18420 16776
rect 18279 16745 18291 16748
rect 18233 16739 18291 16745
rect 1946 16668 1952 16720
rect 2004 16708 2010 16720
rect 2004 16680 3188 16708
rect 2004 16668 2010 16680
rect 2685 16643 2743 16649
rect 2685 16609 2697 16643
rect 2731 16640 2743 16643
rect 2774 16640 2780 16652
rect 2731 16612 2780 16640
rect 2731 16609 2743 16612
rect 2685 16603 2743 16609
rect 2774 16600 2780 16612
rect 2832 16600 2838 16652
rect 2958 16640 2964 16652
rect 2919 16612 2964 16640
rect 2958 16600 2964 16612
rect 3016 16600 3022 16652
rect 3160 16649 3188 16680
rect 3970 16668 3976 16720
rect 4028 16708 4034 16720
rect 4617 16711 4675 16717
rect 4617 16708 4629 16711
rect 4028 16680 4629 16708
rect 4028 16668 4034 16680
rect 4617 16677 4629 16680
rect 4663 16677 4675 16711
rect 4617 16671 4675 16677
rect 3145 16643 3203 16649
rect 3145 16609 3157 16643
rect 3191 16609 3203 16643
rect 4246 16640 4252 16652
rect 4207 16612 4252 16640
rect 3145 16603 3203 16609
rect 4246 16600 4252 16612
rect 4304 16600 4310 16652
rect 4430 16640 4436 16652
rect 4391 16612 4436 16640
rect 4430 16600 4436 16612
rect 4488 16600 4494 16652
rect 5445 16643 5503 16649
rect 5445 16609 5457 16643
rect 5491 16640 5503 16643
rect 5491 16612 5580 16640
rect 5491 16609 5503 16612
rect 5445 16603 5503 16609
rect 2314 16532 2320 16584
rect 2372 16572 2378 16584
rect 3237 16575 3295 16581
rect 3237 16572 3249 16575
rect 2372 16544 3249 16572
rect 2372 16532 2378 16544
rect 3237 16541 3249 16544
rect 3283 16541 3295 16575
rect 3237 16535 3295 16541
rect 3510 16532 3516 16584
rect 3568 16572 3574 16584
rect 4801 16575 4859 16581
rect 4801 16572 4813 16575
rect 3568 16544 4813 16572
rect 3568 16532 3574 16544
rect 4801 16541 4813 16544
rect 4847 16541 4859 16575
rect 5552 16572 5580 16612
rect 8478 16600 8484 16652
rect 8536 16600 8542 16652
rect 11609 16643 11667 16649
rect 11609 16609 11621 16643
rect 11655 16640 11667 16643
rect 11790 16640 11796 16652
rect 11655 16612 11796 16640
rect 11655 16609 11667 16612
rect 11609 16603 11667 16609
rect 11790 16600 11796 16612
rect 11848 16640 11854 16652
rect 13538 16640 13544 16652
rect 11848 16612 13544 16640
rect 11848 16600 11854 16612
rect 13538 16600 13544 16612
rect 13596 16600 13602 16652
rect 18049 16643 18107 16649
rect 18049 16609 18061 16643
rect 18095 16640 18107 16643
rect 18248 16640 18276 16739
rect 18414 16736 18420 16748
rect 18472 16736 18478 16788
rect 19334 16736 19340 16788
rect 19392 16776 19398 16788
rect 21266 16776 21272 16788
rect 19392 16748 21272 16776
rect 19392 16736 19398 16748
rect 21266 16736 21272 16748
rect 21324 16736 21330 16788
rect 22186 16736 22192 16788
rect 22244 16776 22250 16788
rect 22465 16779 22523 16785
rect 22465 16776 22477 16779
rect 22244 16748 22477 16776
rect 22244 16736 22250 16748
rect 22465 16745 22477 16748
rect 22511 16745 22523 16779
rect 22738 16776 22744 16788
rect 22699 16748 22744 16776
rect 22465 16739 22523 16745
rect 22738 16736 22744 16748
rect 22796 16736 22802 16788
rect 20898 16708 20904 16720
rect 20640 16680 20904 16708
rect 19426 16640 19432 16652
rect 18095 16612 18276 16640
rect 18708 16612 19432 16640
rect 18095 16609 18107 16612
rect 18049 16603 18107 16609
rect 7377 16575 7435 16581
rect 7377 16572 7389 16575
rect 5552 16544 6224 16572
rect 4801 16535 4859 16541
rect 6196 16516 6224 16544
rect 6932 16544 7389 16572
rect 2409 16507 2467 16513
rect 2409 16473 2421 16507
rect 2455 16504 2467 16507
rect 3694 16504 3700 16516
rect 2455 16476 3700 16504
rect 2455 16473 2467 16476
rect 2409 16467 2467 16473
rect 3694 16464 3700 16476
rect 3752 16464 3758 16516
rect 5534 16464 5540 16516
rect 5592 16504 5598 16516
rect 5690 16507 5748 16513
rect 5690 16504 5702 16507
rect 5592 16476 5702 16504
rect 5592 16464 5598 16476
rect 5690 16473 5702 16476
rect 5736 16504 5748 16507
rect 5994 16504 6000 16516
rect 5736 16476 6000 16504
rect 5736 16473 5748 16476
rect 5690 16467 5748 16473
rect 5994 16464 6000 16476
rect 6052 16464 6058 16516
rect 6178 16464 6184 16516
rect 6236 16504 6242 16516
rect 6932 16513 6960 16544
rect 7377 16541 7389 16544
rect 7423 16572 7435 16575
rect 8496 16572 8524 16600
rect 8941 16575 8999 16581
rect 8941 16572 8953 16575
rect 7423 16544 8953 16572
rect 7423 16541 7435 16544
rect 7377 16535 7435 16541
rect 8941 16541 8953 16544
rect 8987 16572 8999 16575
rect 9585 16575 9643 16581
rect 9585 16572 9597 16575
rect 8987 16544 9597 16572
rect 8987 16541 8999 16544
rect 8941 16535 8999 16541
rect 9585 16541 9597 16544
rect 9631 16572 9643 16575
rect 9766 16572 9772 16584
rect 9631 16544 9772 16572
rect 9631 16541 9643 16544
rect 9585 16535 9643 16541
rect 9766 16532 9772 16544
rect 9824 16572 9830 16584
rect 11333 16575 11391 16581
rect 11333 16572 11345 16575
rect 9824 16544 11345 16572
rect 9824 16532 9830 16544
rect 11333 16541 11345 16544
rect 11379 16572 11391 16575
rect 12253 16575 12311 16581
rect 12253 16572 12265 16575
rect 11379 16544 12265 16572
rect 11379 16541 11391 16544
rect 11333 16535 11391 16541
rect 12253 16541 12265 16544
rect 12299 16572 12311 16575
rect 13725 16575 13783 16581
rect 13725 16572 13737 16575
rect 12299 16544 13737 16572
rect 12299 16541 12311 16544
rect 12253 16535 12311 16541
rect 13725 16541 13737 16544
rect 13771 16572 13783 16575
rect 14737 16575 14795 16581
rect 14737 16572 14749 16575
rect 13771 16544 14749 16572
rect 13771 16541 13783 16544
rect 13725 16535 13783 16541
rect 14737 16541 14749 16544
rect 14783 16541 14795 16575
rect 14737 16535 14795 16541
rect 15004 16575 15062 16581
rect 15004 16541 15016 16575
rect 15050 16572 15062 16575
rect 15470 16572 15476 16584
rect 15050 16544 15476 16572
rect 15050 16541 15062 16544
rect 15004 16535 15062 16541
rect 15470 16532 15476 16544
rect 15528 16532 15534 16584
rect 17494 16532 17500 16584
rect 17552 16572 17558 16584
rect 17782 16575 17840 16581
rect 17782 16572 17794 16575
rect 17552 16544 17794 16572
rect 17552 16532 17558 16544
rect 17782 16541 17794 16544
rect 17828 16541 17840 16575
rect 17782 16535 17840 16541
rect 18138 16532 18144 16584
rect 18196 16572 18202 16584
rect 18601 16575 18659 16581
rect 18601 16572 18613 16575
rect 18196 16544 18613 16572
rect 18196 16532 18202 16544
rect 18601 16541 18613 16544
rect 18647 16572 18659 16575
rect 18708 16572 18736 16612
rect 19426 16600 19432 16612
rect 19484 16600 19490 16652
rect 20640 16649 20668 16680
rect 20898 16668 20904 16680
rect 20956 16708 20962 16720
rect 21818 16708 21824 16720
rect 20956 16680 21824 16708
rect 20956 16668 20962 16680
rect 21818 16668 21824 16680
rect 21876 16708 21882 16720
rect 22756 16708 22784 16736
rect 21876 16680 22784 16708
rect 21876 16668 21882 16680
rect 20625 16643 20683 16649
rect 20625 16609 20637 16643
rect 20671 16609 20683 16643
rect 20625 16603 20683 16609
rect 20717 16643 20775 16649
rect 20717 16609 20729 16643
rect 20763 16640 20775 16643
rect 21082 16640 21088 16652
rect 20763 16612 21088 16640
rect 20763 16609 20775 16612
rect 20717 16603 20775 16609
rect 18877 16575 18935 16581
rect 18877 16572 18889 16575
rect 18647 16544 18736 16572
rect 18800 16544 18889 16572
rect 18647 16541 18659 16544
rect 18601 16535 18659 16541
rect 6917 16507 6975 16513
rect 6917 16504 6929 16507
rect 6236 16476 6929 16504
rect 6236 16464 6242 16476
rect 6917 16473 6929 16476
rect 6963 16473 6975 16507
rect 6917 16467 6975 16473
rect 7644 16507 7702 16513
rect 7644 16473 7656 16507
rect 7690 16504 7702 16507
rect 7834 16504 7840 16516
rect 7690 16476 7840 16504
rect 7690 16473 7702 16476
rect 7644 16467 7702 16473
rect 7834 16464 7840 16476
rect 7892 16464 7898 16516
rect 11054 16464 11060 16516
rect 11112 16513 11118 16516
rect 11112 16504 11124 16513
rect 16666 16504 16672 16516
rect 11112 16476 11157 16504
rect 16132 16476 16672 16504
rect 11112 16467 11124 16476
rect 11112 16464 11118 16467
rect 1486 16396 1492 16448
rect 1544 16436 1550 16448
rect 2041 16439 2099 16445
rect 2041 16436 2053 16439
rect 1544 16408 2053 16436
rect 1544 16396 1550 16408
rect 2041 16405 2053 16408
rect 2087 16405 2099 16439
rect 2041 16399 2099 16405
rect 2501 16439 2559 16445
rect 2501 16405 2513 16439
rect 2547 16436 2559 16439
rect 2866 16436 2872 16448
rect 2547 16408 2872 16436
rect 2547 16405 2559 16408
rect 2501 16399 2559 16405
rect 2866 16396 2872 16408
rect 2924 16396 2930 16448
rect 3602 16436 3608 16448
rect 3563 16408 3608 16436
rect 3602 16396 3608 16408
rect 3660 16396 3666 16448
rect 4154 16436 4160 16448
rect 4115 16408 4160 16436
rect 4154 16396 4160 16408
rect 4212 16396 4218 16448
rect 6270 16396 6276 16448
rect 6328 16436 6334 16448
rect 6825 16439 6883 16445
rect 6825 16436 6837 16439
rect 6328 16408 6837 16436
rect 6328 16396 6334 16408
rect 6825 16405 6837 16408
rect 6871 16405 6883 16439
rect 6825 16399 6883 16405
rect 9953 16439 10011 16445
rect 9953 16405 9965 16439
rect 9999 16436 10011 16439
rect 11238 16436 11244 16448
rect 9999 16408 11244 16436
rect 9999 16405 10011 16408
rect 9953 16399 10011 16405
rect 11238 16396 11244 16408
rect 11296 16436 11302 16448
rect 11701 16439 11759 16445
rect 11701 16436 11713 16439
rect 11296 16408 11713 16436
rect 11296 16396 11302 16408
rect 11701 16405 11713 16408
rect 11747 16405 11759 16439
rect 11701 16399 11759 16405
rect 11790 16396 11796 16448
rect 11848 16436 11854 16448
rect 12161 16439 12219 16445
rect 11848 16408 11893 16436
rect 11848 16396 11854 16408
rect 12161 16405 12173 16439
rect 12207 16436 12219 16439
rect 12986 16436 12992 16448
rect 12207 16408 12992 16436
rect 12207 16405 12219 16408
rect 12161 16399 12219 16405
rect 12986 16396 12992 16408
rect 13044 16396 13050 16448
rect 16132 16445 16160 16476
rect 16666 16464 16672 16476
rect 16724 16464 16730 16516
rect 16117 16439 16175 16445
rect 16117 16405 16129 16439
rect 16163 16405 16175 16439
rect 16298 16436 16304 16448
rect 16259 16408 16304 16436
rect 16117 16399 16175 16405
rect 16298 16396 16304 16408
rect 16356 16436 16362 16448
rect 16485 16439 16543 16445
rect 16485 16436 16497 16439
rect 16356 16408 16497 16436
rect 16356 16396 16362 16408
rect 16485 16405 16497 16408
rect 16531 16405 16543 16439
rect 16485 16399 16543 16405
rect 18509 16439 18567 16445
rect 18509 16405 18521 16439
rect 18555 16436 18567 16439
rect 18598 16436 18604 16448
rect 18555 16408 18604 16436
rect 18555 16405 18567 16408
rect 18509 16399 18567 16405
rect 18598 16396 18604 16408
rect 18656 16396 18662 16448
rect 18800 16445 18828 16544
rect 18877 16541 18889 16544
rect 18923 16541 18935 16575
rect 20732 16572 20760 16603
rect 21082 16600 21088 16612
rect 21140 16600 21146 16652
rect 21634 16600 21640 16652
rect 21692 16640 21698 16652
rect 22097 16643 22155 16649
rect 22097 16640 22109 16643
rect 21692 16612 22109 16640
rect 21692 16600 21698 16612
rect 22097 16609 22109 16612
rect 22143 16609 22155 16643
rect 22097 16603 22155 16609
rect 22189 16643 22247 16649
rect 22189 16609 22201 16643
rect 22235 16609 22247 16643
rect 22189 16603 22247 16609
rect 18877 16535 18935 16541
rect 19076 16544 20760 16572
rect 19076 16445 19104 16544
rect 20898 16532 20904 16584
rect 20956 16572 20962 16584
rect 20993 16575 21051 16581
rect 20993 16572 21005 16575
rect 20956 16544 21005 16572
rect 20956 16532 20962 16544
rect 20993 16541 21005 16544
rect 21039 16541 21051 16575
rect 20993 16535 21051 16541
rect 21726 16532 21732 16584
rect 21784 16572 21790 16584
rect 22204 16572 22232 16603
rect 22646 16572 22652 16584
rect 21784 16544 22232 16572
rect 22607 16544 22652 16572
rect 21784 16532 21790 16544
rect 22646 16532 22652 16544
rect 22704 16532 22710 16584
rect 23109 16575 23167 16581
rect 23109 16541 23121 16575
rect 23155 16572 23167 16575
rect 23198 16572 23204 16584
rect 23155 16544 23204 16572
rect 23155 16541 23167 16544
rect 23109 16535 23167 16541
rect 20346 16504 20352 16516
rect 20404 16513 20410 16516
rect 20316 16476 20352 16504
rect 20346 16464 20352 16476
rect 20404 16467 20416 16513
rect 20404 16464 20410 16467
rect 20530 16464 20536 16516
rect 20588 16504 20594 16516
rect 23124 16504 23152 16535
rect 23198 16532 23204 16544
rect 23256 16532 23262 16584
rect 20588 16476 23152 16504
rect 20588 16464 20594 16476
rect 18785 16439 18843 16445
rect 18785 16405 18797 16439
rect 18831 16405 18843 16439
rect 18785 16399 18843 16405
rect 19061 16439 19119 16445
rect 19061 16405 19073 16439
rect 19107 16405 19119 16439
rect 19061 16399 19119 16405
rect 19245 16439 19303 16445
rect 19245 16405 19257 16439
rect 19291 16436 19303 16439
rect 19886 16436 19892 16448
rect 19291 16408 19892 16436
rect 19291 16405 19303 16408
rect 19245 16399 19303 16405
rect 19886 16396 19892 16408
rect 19944 16396 19950 16448
rect 21450 16396 21456 16448
rect 21508 16436 21514 16448
rect 21637 16439 21695 16445
rect 21637 16436 21649 16439
rect 21508 16408 21649 16436
rect 21508 16396 21514 16408
rect 21637 16405 21649 16408
rect 21683 16405 21695 16439
rect 22002 16436 22008 16448
rect 21963 16408 22008 16436
rect 21637 16399 21695 16405
rect 22002 16396 22008 16408
rect 22060 16396 22066 16448
rect 22925 16439 22983 16445
rect 22925 16405 22937 16439
rect 22971 16436 22983 16439
rect 23014 16436 23020 16448
rect 22971 16408 23020 16436
rect 22971 16405 22983 16408
rect 22925 16399 22983 16405
rect 23014 16396 23020 16408
rect 23072 16396 23078 16448
rect 1104 16346 23460 16368
rect 1104 16294 6548 16346
rect 6600 16294 6612 16346
rect 6664 16294 6676 16346
rect 6728 16294 6740 16346
rect 6792 16294 6804 16346
rect 6856 16294 12146 16346
rect 12198 16294 12210 16346
rect 12262 16294 12274 16346
rect 12326 16294 12338 16346
rect 12390 16294 12402 16346
rect 12454 16294 17744 16346
rect 17796 16294 17808 16346
rect 17860 16294 17872 16346
rect 17924 16294 17936 16346
rect 17988 16294 18000 16346
rect 18052 16294 23460 16346
rect 1104 16272 23460 16294
rect 1670 16232 1676 16244
rect 1631 16204 1676 16232
rect 1670 16192 1676 16204
rect 1728 16192 1734 16244
rect 1946 16232 1952 16244
rect 1907 16204 1952 16232
rect 1946 16192 1952 16204
rect 2004 16192 2010 16244
rect 2406 16232 2412 16244
rect 2367 16204 2412 16232
rect 2406 16192 2412 16204
rect 2464 16192 2470 16244
rect 2866 16232 2872 16244
rect 2827 16204 2872 16232
rect 2866 16192 2872 16204
rect 2924 16192 2930 16244
rect 3510 16232 3516 16244
rect 3160 16204 3516 16232
rect 3160 16164 3188 16204
rect 3510 16192 3516 16204
rect 3568 16192 3574 16244
rect 3694 16232 3700 16244
rect 3655 16204 3700 16232
rect 3694 16192 3700 16204
rect 3752 16192 3758 16244
rect 4157 16235 4215 16241
rect 4157 16201 4169 16235
rect 4203 16232 4215 16235
rect 4798 16232 4804 16244
rect 4203 16204 4804 16232
rect 4203 16201 4215 16204
rect 4157 16195 4215 16201
rect 4798 16192 4804 16204
rect 4856 16192 4862 16244
rect 9582 16232 9588 16244
rect 9508 16204 9588 16232
rect 2240 16136 3188 16164
rect 3237 16167 3295 16173
rect 1486 16096 1492 16108
rect 1447 16068 1492 16096
rect 1486 16056 1492 16068
rect 1544 16056 1550 16108
rect 1762 16096 1768 16108
rect 1723 16068 1768 16096
rect 1762 16056 1768 16068
rect 1820 16056 1826 16108
rect 2240 16037 2268 16136
rect 3237 16133 3249 16167
rect 3283 16164 3295 16167
rect 5718 16164 5724 16176
rect 3283 16136 5724 16164
rect 3283 16133 3295 16136
rect 3237 16127 3295 16133
rect 5718 16124 5724 16136
rect 5776 16164 5782 16176
rect 9508 16173 9536 16204
rect 9582 16192 9588 16204
rect 9640 16192 9646 16244
rect 9858 16232 9864 16244
rect 9771 16204 9864 16232
rect 9858 16192 9864 16204
rect 9916 16232 9922 16244
rect 11790 16232 11796 16244
rect 9916 16204 11796 16232
rect 9916 16192 9922 16204
rect 11790 16192 11796 16204
rect 11848 16192 11854 16244
rect 14001 16235 14059 16241
rect 14001 16201 14013 16235
rect 14047 16232 14059 16235
rect 14826 16232 14832 16244
rect 14047 16204 14832 16232
rect 14047 16201 14059 16204
rect 14001 16195 14059 16201
rect 14826 16192 14832 16204
rect 14884 16192 14890 16244
rect 15657 16235 15715 16241
rect 15657 16201 15669 16235
rect 15703 16232 15715 16235
rect 15841 16235 15899 16241
rect 15841 16232 15853 16235
rect 15703 16204 15853 16232
rect 15703 16201 15715 16204
rect 15657 16195 15715 16201
rect 15841 16201 15853 16204
rect 15887 16232 15899 16235
rect 16209 16235 16267 16241
rect 16209 16232 16221 16235
rect 15887 16204 16221 16232
rect 15887 16201 15899 16204
rect 15841 16195 15899 16201
rect 16209 16201 16221 16204
rect 16255 16232 16267 16235
rect 16298 16232 16304 16244
rect 16255 16204 16304 16232
rect 16255 16201 16267 16204
rect 16209 16195 16267 16201
rect 5914 16167 5972 16173
rect 5914 16164 5926 16167
rect 5776 16136 5926 16164
rect 5776 16124 5782 16136
rect 5914 16133 5926 16136
rect 5960 16133 5972 16167
rect 5914 16127 5972 16133
rect 9502 16167 9560 16173
rect 9502 16133 9514 16167
rect 9548 16133 9560 16167
rect 11517 16167 11575 16173
rect 11517 16164 11529 16167
rect 9502 16127 9560 16133
rect 9784 16136 11529 16164
rect 9784 16108 9812 16136
rect 4065 16099 4123 16105
rect 4065 16065 4077 16099
rect 4111 16096 4123 16099
rect 4338 16096 4344 16108
rect 4111 16068 4344 16096
rect 4111 16065 4123 16068
rect 4065 16059 4123 16065
rect 4338 16056 4344 16068
rect 4396 16056 4402 16108
rect 9766 16096 9772 16108
rect 9727 16068 9772 16096
rect 9766 16056 9772 16068
rect 9824 16056 9830 16108
rect 10985 16099 11043 16105
rect 10985 16065 10997 16099
rect 11031 16096 11043 16099
rect 11146 16096 11152 16108
rect 11031 16068 11152 16096
rect 11031 16065 11043 16068
rect 10985 16059 11043 16065
rect 11146 16056 11152 16068
rect 11204 16056 11210 16108
rect 11256 16105 11284 16136
rect 11517 16133 11529 16136
rect 11563 16133 11575 16167
rect 13909 16167 13967 16173
rect 13909 16164 13921 16167
rect 11517 16127 11575 16133
rect 12268 16136 13921 16164
rect 11241 16099 11299 16105
rect 11241 16065 11253 16099
rect 11287 16065 11299 16099
rect 11532 16096 11560 16127
rect 11974 16096 11980 16108
rect 11532 16068 11980 16096
rect 11241 16059 11299 16065
rect 11974 16056 11980 16068
rect 12032 16096 12038 16108
rect 12268 16105 12296 16136
rect 13909 16133 13921 16136
rect 13955 16164 13967 16167
rect 13955 16136 15424 16164
rect 13955 16133 13967 16136
rect 13909 16127 13967 16133
rect 12253 16099 12311 16105
rect 12253 16096 12265 16099
rect 12032 16068 12265 16096
rect 12032 16056 12038 16068
rect 12253 16065 12265 16068
rect 12299 16065 12311 16099
rect 12253 16059 12311 16065
rect 12520 16099 12578 16105
rect 12520 16065 12532 16099
rect 12566 16096 12578 16099
rect 12802 16096 12808 16108
rect 12566 16068 12808 16096
rect 12566 16065 12578 16068
rect 12520 16059 12578 16065
rect 12802 16056 12808 16068
rect 12860 16056 12866 16108
rect 15125 16099 15183 16105
rect 15125 16065 15137 16099
rect 15171 16096 15183 16099
rect 15286 16096 15292 16108
rect 15171 16068 15292 16096
rect 15171 16065 15183 16068
rect 15125 16059 15183 16065
rect 15286 16056 15292 16068
rect 15344 16056 15350 16108
rect 15396 16105 15424 16136
rect 15381 16099 15439 16105
rect 15381 16065 15393 16099
rect 15427 16096 15439 16099
rect 15672 16096 15700 16195
rect 16298 16192 16304 16204
rect 16356 16232 16362 16244
rect 16853 16235 16911 16241
rect 16853 16232 16865 16235
rect 16356 16204 16865 16232
rect 16356 16192 16362 16204
rect 16853 16201 16865 16204
rect 16899 16232 16911 16235
rect 17037 16235 17095 16241
rect 17037 16232 17049 16235
rect 16899 16204 17049 16232
rect 16899 16201 16911 16204
rect 16853 16195 16911 16201
rect 17037 16201 17049 16204
rect 17083 16232 17095 16235
rect 17221 16235 17279 16241
rect 17221 16232 17233 16235
rect 17083 16204 17233 16232
rect 17083 16201 17095 16204
rect 17037 16195 17095 16201
rect 17221 16201 17233 16204
rect 17267 16232 17279 16235
rect 17497 16235 17555 16241
rect 17497 16232 17509 16235
rect 17267 16204 17509 16232
rect 17267 16201 17279 16204
rect 17221 16195 17279 16201
rect 17497 16201 17509 16204
rect 17543 16232 17555 16235
rect 17681 16235 17739 16241
rect 17681 16232 17693 16235
rect 17543 16204 17693 16232
rect 17543 16201 17555 16204
rect 17497 16195 17555 16201
rect 17681 16201 17693 16204
rect 17727 16232 17739 16235
rect 18233 16235 18291 16241
rect 18233 16232 18245 16235
rect 17727 16204 18245 16232
rect 17727 16201 17739 16204
rect 17681 16195 17739 16201
rect 18233 16201 18245 16204
rect 18279 16232 18291 16235
rect 18414 16232 18420 16244
rect 18279 16204 18420 16232
rect 18279 16201 18291 16204
rect 18233 16195 18291 16201
rect 18414 16192 18420 16204
rect 18472 16232 18478 16244
rect 18598 16232 18604 16244
rect 18472 16204 18604 16232
rect 18472 16192 18478 16204
rect 18598 16192 18604 16204
rect 18656 16192 18662 16244
rect 20530 16232 20536 16244
rect 19168 16204 20536 16232
rect 17865 16167 17923 16173
rect 17865 16133 17877 16167
rect 17911 16164 17923 16167
rect 18138 16164 18144 16176
rect 17911 16136 18144 16164
rect 17911 16133 17923 16136
rect 17865 16127 17923 16133
rect 18138 16124 18144 16136
rect 18196 16124 18202 16176
rect 15427 16068 15700 16096
rect 16485 16099 16543 16105
rect 15427 16065 15439 16068
rect 15381 16059 15439 16065
rect 16485 16065 16497 16099
rect 16531 16096 16543 16099
rect 19168 16096 19196 16204
rect 20530 16192 20536 16204
rect 20588 16192 20594 16244
rect 21177 16235 21235 16241
rect 21177 16201 21189 16235
rect 21223 16232 21235 16235
rect 21910 16232 21916 16244
rect 21223 16204 21916 16232
rect 21223 16201 21235 16204
rect 21177 16195 21235 16201
rect 21910 16192 21916 16204
rect 21968 16192 21974 16244
rect 22557 16235 22615 16241
rect 22557 16201 22569 16235
rect 22603 16201 22615 16235
rect 22557 16195 22615 16201
rect 20162 16164 20168 16176
rect 19812 16136 20168 16164
rect 16531 16068 19196 16096
rect 19449 16099 19507 16105
rect 16531 16065 16543 16068
rect 16485 16059 16543 16065
rect 19449 16065 19461 16099
rect 19495 16096 19507 16099
rect 19610 16096 19616 16108
rect 19495 16068 19616 16096
rect 19495 16065 19507 16068
rect 19449 16059 19507 16065
rect 19610 16056 19616 16068
rect 19668 16056 19674 16108
rect 19812 16105 19840 16136
rect 20162 16124 20168 16136
rect 20220 16124 20226 16176
rect 21542 16164 21548 16176
rect 21503 16136 21548 16164
rect 21542 16124 21548 16136
rect 21600 16124 21606 16176
rect 19705 16099 19763 16105
rect 19705 16065 19717 16099
rect 19751 16096 19763 16099
rect 19797 16099 19855 16105
rect 19797 16096 19809 16099
rect 19751 16068 19809 16096
rect 19751 16065 19763 16068
rect 19705 16059 19763 16065
rect 19797 16065 19809 16068
rect 19843 16065 19855 16099
rect 19797 16059 19855 16065
rect 19886 16056 19892 16108
rect 19944 16096 19950 16108
rect 20053 16099 20111 16105
rect 20053 16096 20065 16099
rect 19944 16068 20065 16096
rect 19944 16056 19950 16068
rect 20053 16065 20065 16068
rect 20099 16065 20111 16099
rect 20053 16059 20111 16065
rect 20898 16056 20904 16108
rect 20956 16096 20962 16108
rect 21361 16099 21419 16105
rect 21361 16096 21373 16099
rect 20956 16068 21373 16096
rect 20956 16056 20962 16068
rect 21361 16065 21373 16068
rect 21407 16065 21419 16099
rect 21361 16059 21419 16065
rect 21450 16056 21456 16108
rect 21508 16096 21514 16108
rect 22097 16099 22155 16105
rect 22097 16096 22109 16099
rect 21508 16068 22109 16096
rect 21508 16056 21514 16068
rect 22097 16065 22109 16068
rect 22143 16065 22155 16099
rect 22097 16059 22155 16065
rect 22189 16099 22247 16105
rect 22189 16065 22201 16099
rect 22235 16065 22247 16099
rect 22572 16096 22600 16195
rect 22833 16099 22891 16105
rect 22833 16096 22845 16099
rect 22572 16068 22845 16096
rect 22189 16059 22247 16065
rect 22833 16065 22845 16068
rect 22879 16065 22891 16099
rect 23106 16096 23112 16108
rect 23067 16068 23112 16096
rect 22833 16059 22891 16065
rect 2225 16031 2283 16037
rect 2225 15997 2237 16031
rect 2271 15997 2283 16031
rect 2225 15991 2283 15997
rect 2317 16031 2375 16037
rect 2317 15997 2329 16031
rect 2363 15997 2375 16031
rect 3326 16028 3332 16040
rect 3287 16000 3332 16028
rect 2317 15991 2375 15997
rect 2332 15892 2360 15991
rect 3326 15988 3332 16000
rect 3384 15988 3390 16040
rect 3510 15988 3516 16040
rect 3568 16028 3574 16040
rect 3970 16028 3976 16040
rect 3568 16000 3976 16028
rect 3568 15988 3574 16000
rect 3970 15988 3976 16000
rect 4028 16028 4034 16040
rect 4249 16031 4307 16037
rect 4249 16028 4261 16031
rect 4028 16000 4261 16028
rect 4028 15988 4034 16000
rect 4249 15997 4261 16000
rect 4295 15997 4307 16031
rect 4249 15991 4307 15997
rect 6181 16031 6239 16037
rect 6181 15997 6193 16031
rect 6227 15997 6239 16031
rect 6181 15991 6239 15997
rect 18049 16031 18107 16037
rect 18049 15997 18061 16031
rect 18095 16028 18107 16031
rect 18506 16028 18512 16040
rect 18095 16000 18512 16028
rect 18095 15997 18107 16000
rect 18049 15991 18107 15997
rect 2777 15963 2835 15969
rect 2777 15929 2789 15963
rect 2823 15960 2835 15963
rect 4154 15960 4160 15972
rect 2823 15932 4160 15960
rect 2823 15929 2835 15932
rect 2777 15923 2835 15929
rect 4154 15920 4160 15932
rect 4212 15920 4218 15972
rect 6196 15904 6224 15991
rect 18506 15988 18512 16000
rect 18564 15988 18570 16040
rect 21726 15988 21732 16040
rect 21784 16028 21790 16040
rect 21913 16031 21971 16037
rect 21913 16028 21925 16031
rect 21784 16000 21925 16028
rect 21784 15988 21790 16000
rect 21913 15997 21925 16000
rect 21959 15997 21971 16031
rect 21913 15991 21971 15997
rect 21266 15920 21272 15972
rect 21324 15960 21330 15972
rect 22204 15960 22232 16059
rect 23106 16056 23112 16068
rect 23164 16056 23170 16108
rect 21324 15932 22232 15960
rect 21324 15920 21330 15932
rect 22370 15920 22376 15972
rect 22428 15960 22434 15972
rect 22649 15963 22707 15969
rect 22649 15960 22661 15963
rect 22428 15932 22661 15960
rect 22428 15920 22434 15932
rect 22649 15929 22661 15932
rect 22695 15929 22707 15963
rect 22649 15923 22707 15929
rect 5534 15892 5540 15904
rect 2332 15864 5540 15892
rect 5534 15852 5540 15864
rect 5592 15852 5598 15904
rect 6178 15852 6184 15904
rect 6236 15892 6242 15904
rect 6365 15895 6423 15901
rect 6365 15892 6377 15895
rect 6236 15864 6377 15892
rect 6236 15852 6242 15864
rect 6365 15861 6377 15864
rect 6411 15861 6423 15895
rect 8386 15892 8392 15904
rect 8347 15864 8392 15892
rect 6365 15855 6423 15861
rect 8386 15852 8392 15864
rect 8444 15852 8450 15904
rect 13633 15895 13691 15901
rect 13633 15861 13645 15895
rect 13679 15892 13691 15895
rect 14274 15892 14280 15904
rect 13679 15864 14280 15892
rect 13679 15861 13691 15864
rect 13633 15855 13691 15861
rect 14274 15852 14280 15864
rect 14332 15892 14338 15904
rect 16114 15892 16120 15904
rect 14332 15864 16120 15892
rect 14332 15852 14338 15864
rect 16114 15852 16120 15864
rect 16172 15852 16178 15904
rect 18325 15895 18383 15901
rect 18325 15861 18337 15895
rect 18371 15892 18383 15895
rect 18414 15892 18420 15904
rect 18371 15864 18420 15892
rect 18371 15861 18383 15864
rect 18325 15855 18383 15861
rect 18414 15852 18420 15864
rect 18472 15892 18478 15904
rect 21082 15892 21088 15904
rect 18472 15864 21088 15892
rect 18472 15852 18478 15864
rect 21082 15852 21088 15864
rect 21140 15852 21146 15904
rect 22922 15892 22928 15904
rect 22883 15864 22928 15892
rect 22922 15852 22928 15864
rect 22980 15852 22986 15904
rect 1104 15802 23460 15824
rect 1104 15750 3749 15802
rect 3801 15750 3813 15802
rect 3865 15750 3877 15802
rect 3929 15750 3941 15802
rect 3993 15750 4005 15802
rect 4057 15750 9347 15802
rect 9399 15750 9411 15802
rect 9463 15750 9475 15802
rect 9527 15750 9539 15802
rect 9591 15750 9603 15802
rect 9655 15750 14945 15802
rect 14997 15750 15009 15802
rect 15061 15750 15073 15802
rect 15125 15750 15137 15802
rect 15189 15750 15201 15802
rect 15253 15750 20543 15802
rect 20595 15750 20607 15802
rect 20659 15750 20671 15802
rect 20723 15750 20735 15802
rect 20787 15750 20799 15802
rect 20851 15750 23460 15802
rect 1104 15728 23460 15750
rect 1949 15691 2007 15697
rect 1949 15657 1961 15691
rect 1995 15688 2007 15691
rect 2038 15688 2044 15700
rect 1995 15660 2044 15688
rect 1995 15657 2007 15660
rect 1949 15651 2007 15657
rect 2038 15648 2044 15660
rect 2096 15648 2102 15700
rect 4249 15691 4307 15697
rect 4249 15657 4261 15691
rect 4295 15688 4307 15691
rect 4338 15688 4344 15700
rect 4295 15660 4344 15688
rect 4295 15657 4307 15660
rect 4249 15651 4307 15657
rect 4338 15648 4344 15660
rect 4396 15648 4402 15700
rect 10413 15691 10471 15697
rect 4724 15660 5672 15688
rect 4724 15620 4752 15660
rect 4172 15592 4752 15620
rect 5644 15620 5672 15660
rect 10413 15657 10425 15691
rect 10459 15688 10471 15691
rect 10502 15688 10508 15700
rect 10459 15660 10508 15688
rect 10459 15657 10471 15660
rect 10413 15651 10471 15657
rect 10502 15648 10508 15660
rect 10560 15648 10566 15700
rect 11974 15688 11980 15700
rect 11935 15660 11980 15688
rect 11974 15648 11980 15660
rect 12032 15688 12038 15700
rect 12161 15691 12219 15697
rect 12161 15688 12173 15691
rect 12032 15660 12173 15688
rect 12032 15648 12038 15660
rect 12161 15657 12173 15660
rect 12207 15657 12219 15691
rect 12161 15651 12219 15657
rect 15286 15648 15292 15700
rect 15344 15688 15350 15700
rect 15473 15691 15531 15697
rect 15473 15688 15485 15691
rect 15344 15660 15485 15688
rect 15344 15648 15350 15660
rect 15473 15657 15485 15660
rect 15519 15657 15531 15691
rect 15473 15651 15531 15657
rect 17037 15691 17095 15697
rect 17037 15657 17049 15691
rect 17083 15688 17095 15691
rect 18230 15688 18236 15700
rect 17083 15660 18236 15688
rect 17083 15657 17095 15660
rect 17037 15651 17095 15657
rect 18230 15648 18236 15660
rect 18288 15648 18294 15700
rect 18598 15688 18604 15700
rect 18559 15660 18604 15688
rect 18598 15648 18604 15660
rect 18656 15648 18662 15700
rect 20162 15688 20168 15700
rect 19260 15660 20168 15688
rect 5810 15620 5816 15632
rect 5644 15592 5816 15620
rect 2682 15552 2688 15564
rect 2643 15524 2688 15552
rect 2682 15512 2688 15524
rect 2740 15512 2746 15564
rect 3513 15555 3571 15561
rect 3513 15521 3525 15555
rect 3559 15552 3571 15555
rect 4062 15552 4068 15564
rect 3559 15524 4068 15552
rect 3559 15521 3571 15524
rect 3513 15515 3571 15521
rect 4062 15512 4068 15524
rect 4120 15512 4126 15564
rect 1670 15484 1676 15496
rect 1631 15456 1676 15484
rect 1670 15444 1676 15456
rect 1728 15444 1734 15496
rect 1765 15487 1823 15493
rect 1765 15453 1777 15487
rect 1811 15484 1823 15487
rect 3234 15484 3240 15496
rect 1811 15456 2084 15484
rect 3195 15456 3240 15484
rect 1811 15453 1823 15456
rect 1765 15447 1823 15453
rect 1486 15348 1492 15360
rect 1447 15320 1492 15348
rect 1486 15308 1492 15320
rect 1544 15308 1550 15360
rect 2056 15357 2084 15456
rect 3234 15444 3240 15456
rect 3292 15444 3298 15496
rect 4172 15493 4200 15592
rect 5810 15580 5816 15592
rect 5868 15580 5874 15632
rect 11885 15555 11943 15561
rect 11885 15521 11897 15555
rect 11931 15552 11943 15555
rect 11992 15552 12020 15648
rect 17129 15623 17187 15629
rect 17129 15589 17141 15623
rect 17175 15620 17187 15623
rect 17494 15620 17500 15632
rect 17175 15592 17500 15620
rect 17175 15589 17187 15592
rect 17129 15583 17187 15589
rect 17494 15580 17500 15592
rect 17552 15580 17558 15632
rect 12529 15555 12587 15561
rect 12529 15552 12541 15555
rect 11931 15524 12541 15552
rect 11931 15521 11943 15524
rect 11885 15515 11943 15521
rect 12529 15521 12541 15524
rect 12575 15521 12587 15555
rect 12529 15515 12587 15521
rect 18509 15555 18567 15561
rect 18509 15521 18521 15555
rect 18555 15552 18567 15555
rect 18616 15552 18644 15648
rect 19260 15561 19288 15660
rect 20162 15648 20168 15660
rect 20220 15648 20226 15700
rect 20346 15648 20352 15700
rect 20404 15688 20410 15700
rect 20625 15691 20683 15697
rect 20625 15688 20637 15691
rect 20404 15660 20637 15688
rect 20404 15648 20410 15660
rect 20625 15657 20637 15660
rect 20671 15688 20683 15691
rect 21453 15691 21511 15697
rect 20671 15660 21036 15688
rect 20671 15657 20683 15660
rect 20625 15651 20683 15657
rect 19245 15555 19303 15561
rect 19245 15552 19257 15555
rect 18555 15524 19257 15552
rect 18555 15521 18567 15524
rect 18509 15515 18567 15521
rect 19245 15521 19257 15524
rect 19291 15521 19303 15555
rect 20806 15552 20812 15564
rect 20767 15524 20812 15552
rect 19245 15515 19303 15521
rect 4157 15487 4215 15493
rect 4157 15453 4169 15487
rect 4203 15453 4215 15487
rect 4157 15447 4215 15453
rect 4798 15444 4804 15496
rect 4856 15484 4862 15496
rect 5362 15487 5420 15493
rect 5362 15484 5374 15487
rect 4856 15456 5374 15484
rect 4856 15444 4862 15456
rect 5362 15453 5374 15456
rect 5408 15453 5420 15487
rect 5362 15447 5420 15453
rect 5629 15487 5687 15493
rect 5629 15453 5641 15487
rect 5675 15484 5687 15487
rect 7101 15487 7159 15493
rect 7101 15484 7113 15487
rect 5675 15456 7113 15484
rect 5675 15453 5687 15456
rect 5629 15447 5687 15453
rect 6196 15428 6224 15456
rect 7101 15453 7113 15456
rect 7147 15484 7159 15487
rect 7285 15487 7343 15493
rect 7285 15484 7297 15487
rect 7147 15456 7297 15484
rect 7147 15453 7159 15456
rect 7101 15447 7159 15453
rect 7285 15453 7297 15456
rect 7331 15484 7343 15487
rect 9033 15487 9091 15493
rect 9033 15484 9045 15487
rect 7331 15456 9045 15484
rect 7331 15453 7343 15456
rect 7285 15447 7343 15453
rect 9033 15453 9045 15456
rect 9079 15453 9091 15487
rect 9033 15447 9091 15453
rect 9300 15487 9358 15493
rect 9300 15453 9312 15487
rect 9346 15484 9358 15487
rect 9858 15484 9864 15496
rect 9346 15456 9864 15484
rect 9346 15453 9358 15456
rect 9300 15447 9358 15453
rect 9858 15444 9864 15456
rect 9916 15444 9922 15496
rect 11606 15484 11612 15496
rect 11664 15493 11670 15496
rect 11576 15456 11612 15484
rect 11606 15444 11612 15456
rect 11664 15447 11676 15493
rect 12544 15484 12572 15515
rect 20806 15512 20812 15524
rect 20864 15512 20870 15564
rect 21008 15561 21036 15660
rect 21453 15657 21465 15691
rect 21499 15688 21511 15691
rect 22002 15688 22008 15700
rect 21499 15660 22008 15688
rect 21499 15657 21511 15660
rect 21453 15651 21511 15657
rect 22002 15648 22008 15660
rect 22060 15648 22066 15700
rect 21082 15580 21088 15632
rect 21140 15580 21146 15632
rect 22741 15623 22799 15629
rect 21836 15592 22692 15620
rect 20993 15555 21051 15561
rect 20993 15521 21005 15555
rect 21039 15521 21051 15555
rect 21100 15552 21128 15580
rect 21100 15524 21772 15552
rect 20993 15515 21051 15521
rect 14093 15487 14151 15493
rect 14093 15484 14105 15487
rect 12544 15456 14105 15484
rect 14093 15453 14105 15456
rect 14139 15484 14151 15487
rect 15657 15487 15715 15493
rect 15657 15484 15669 15487
rect 14139 15456 15669 15484
rect 14139 15453 14151 15456
rect 14093 15447 14151 15453
rect 11664 15444 11670 15447
rect 14568 15428 14596 15456
rect 15657 15453 15669 15456
rect 15703 15453 15715 15487
rect 15657 15447 15715 15453
rect 15924 15487 15982 15493
rect 15924 15453 15936 15487
rect 15970 15484 15982 15487
rect 18414 15484 18420 15496
rect 15970 15456 18420 15484
rect 15970 15453 15982 15456
rect 15924 15447 15982 15453
rect 18414 15444 18420 15456
rect 18472 15444 18478 15496
rect 18874 15484 18880 15496
rect 18787 15456 18880 15484
rect 18874 15444 18880 15456
rect 18932 15484 18938 15496
rect 19150 15484 19156 15496
rect 18932 15456 19156 15484
rect 18932 15444 18938 15456
rect 19150 15444 19156 15456
rect 19208 15444 19214 15496
rect 19334 15444 19340 15496
rect 19392 15484 19398 15496
rect 19501 15487 19559 15493
rect 19501 15484 19513 15487
rect 19392 15456 19513 15484
rect 19392 15444 19398 15456
rect 19501 15453 19513 15456
rect 19547 15453 19559 15487
rect 19501 15447 19559 15453
rect 19886 15444 19892 15496
rect 19944 15484 19950 15496
rect 21085 15487 21143 15493
rect 21085 15484 21097 15487
rect 19944 15456 21097 15484
rect 19944 15444 19950 15456
rect 21085 15453 21097 15456
rect 21131 15453 21143 15487
rect 21542 15484 21548 15496
rect 21503 15456 21548 15484
rect 21085 15447 21143 15453
rect 21542 15444 21548 15456
rect 21600 15444 21606 15496
rect 21744 15493 21772 15524
rect 21729 15487 21787 15493
rect 21729 15453 21741 15487
rect 21775 15453 21787 15487
rect 21729 15447 21787 15453
rect 2501 15419 2559 15425
rect 2501 15385 2513 15419
rect 2547 15416 2559 15419
rect 2774 15416 2780 15428
rect 2547 15388 2780 15416
rect 2547 15385 2559 15388
rect 2501 15379 2559 15385
rect 2774 15376 2780 15388
rect 2832 15376 2838 15428
rect 3329 15419 3387 15425
rect 3329 15385 3341 15419
rect 3375 15416 3387 15419
rect 3375 15388 6132 15416
rect 3375 15385 3387 15388
rect 3329 15379 3387 15385
rect 2041 15351 2099 15357
rect 2041 15317 2053 15351
rect 2087 15317 2099 15351
rect 2406 15348 2412 15360
rect 2367 15320 2412 15348
rect 2041 15311 2099 15317
rect 2406 15308 2412 15320
rect 2464 15308 2470 15360
rect 2866 15348 2872 15360
rect 2827 15320 2872 15348
rect 2866 15308 2872 15320
rect 2924 15308 2930 15360
rect 3602 15308 3608 15360
rect 3660 15348 3666 15360
rect 3973 15351 4031 15357
rect 3973 15348 3985 15351
rect 3660 15320 3985 15348
rect 3660 15308 3666 15320
rect 3973 15317 3985 15320
rect 4019 15317 4031 15351
rect 5718 15348 5724 15360
rect 5679 15320 5724 15348
rect 3973 15311 4031 15317
rect 5718 15308 5724 15320
rect 5776 15308 5782 15360
rect 6104 15348 6132 15388
rect 6178 15376 6184 15428
rect 6236 15376 6242 15428
rect 6454 15376 6460 15428
rect 6512 15416 6518 15428
rect 6834 15419 6892 15425
rect 6834 15416 6846 15419
rect 6512 15388 6846 15416
rect 6512 15376 6518 15388
rect 6834 15385 6846 15388
rect 6880 15385 6892 15419
rect 7530 15419 7588 15425
rect 7530 15416 7542 15419
rect 6834 15379 6892 15385
rect 6932 15388 7542 15416
rect 6932 15348 6960 15388
rect 7530 15385 7542 15388
rect 7576 15416 7588 15419
rect 8386 15416 8392 15428
rect 7576 15388 8392 15416
rect 7576 15385 7588 15388
rect 7530 15379 7588 15385
rect 8386 15376 8392 15388
rect 8444 15376 8450 15428
rect 12526 15376 12532 15428
rect 12584 15416 12590 15428
rect 12796 15419 12854 15425
rect 12796 15416 12808 15419
rect 12584 15388 12808 15416
rect 12584 15376 12590 15388
rect 12796 15385 12808 15388
rect 12842 15416 12854 15419
rect 13078 15416 13084 15428
rect 12842 15388 13084 15416
rect 12842 15385 12854 15388
rect 12796 15379 12854 15385
rect 13078 15376 13084 15388
rect 13136 15376 13142 15428
rect 14366 15425 14372 15428
rect 14360 15416 14372 15425
rect 13924 15388 14372 15416
rect 8662 15348 8668 15360
rect 6104 15320 6960 15348
rect 8623 15320 8668 15348
rect 8662 15308 8668 15320
rect 8720 15308 8726 15360
rect 10505 15351 10563 15357
rect 10505 15317 10517 15351
rect 10551 15348 10563 15351
rect 11054 15348 11060 15360
rect 10551 15320 11060 15348
rect 10551 15317 10563 15320
rect 10505 15311 10563 15317
rect 11054 15308 11060 15320
rect 11112 15348 11118 15360
rect 13262 15348 13268 15360
rect 11112 15320 13268 15348
rect 11112 15308 11118 15320
rect 13262 15308 13268 15320
rect 13320 15308 13326 15360
rect 13924 15357 13952 15388
rect 14360 15379 14372 15388
rect 14366 15376 14372 15379
rect 14424 15376 14430 15428
rect 14550 15376 14556 15428
rect 14608 15376 14614 15428
rect 16666 15376 16672 15428
rect 16724 15416 16730 15428
rect 18242 15419 18300 15425
rect 18242 15416 18254 15419
rect 16724 15388 18254 15416
rect 16724 15376 16730 15388
rect 18242 15385 18254 15388
rect 18288 15385 18300 15419
rect 18242 15379 18300 15385
rect 19978 15376 19984 15428
rect 20036 15416 20042 15428
rect 21836 15416 21864 15592
rect 22189 15555 22247 15561
rect 22189 15521 22201 15555
rect 22235 15552 22247 15555
rect 22462 15552 22468 15564
rect 22235 15524 22468 15552
rect 22235 15521 22247 15524
rect 22189 15515 22247 15521
rect 22462 15512 22468 15524
rect 22520 15512 22526 15564
rect 22664 15552 22692 15592
rect 22741 15589 22753 15623
rect 22787 15620 22799 15623
rect 23290 15620 23296 15632
rect 22787 15592 23296 15620
rect 22787 15589 22799 15592
rect 22741 15583 22799 15589
rect 23290 15580 23296 15592
rect 23348 15580 23354 15632
rect 23658 15552 23664 15564
rect 22664 15524 23664 15552
rect 23658 15512 23664 15524
rect 23716 15512 23722 15564
rect 21913 15487 21971 15493
rect 21913 15453 21925 15487
rect 21959 15484 21971 15487
rect 23017 15487 23075 15493
rect 23017 15484 23029 15487
rect 21959 15456 23029 15484
rect 21959 15453 21971 15456
rect 21913 15447 21971 15453
rect 23017 15453 23029 15456
rect 23063 15453 23075 15487
rect 23017 15447 23075 15453
rect 20036 15388 21864 15416
rect 20036 15376 20042 15388
rect 13909 15351 13967 15357
rect 13909 15317 13921 15351
rect 13955 15317 13967 15351
rect 13909 15311 13967 15317
rect 19061 15351 19119 15357
rect 19061 15317 19073 15351
rect 19107 15348 19119 15351
rect 21634 15348 21640 15360
rect 19107 15320 21640 15348
rect 19107 15317 19119 15320
rect 19061 15311 19119 15317
rect 21634 15308 21640 15320
rect 21692 15308 21698 15360
rect 22278 15348 22284 15360
rect 22239 15320 22284 15348
rect 22278 15308 22284 15320
rect 22336 15308 22342 15360
rect 22370 15308 22376 15360
rect 22428 15348 22434 15360
rect 22428 15320 22473 15348
rect 22428 15308 22434 15320
rect 22646 15308 22652 15360
rect 22704 15348 22710 15360
rect 22833 15351 22891 15357
rect 22833 15348 22845 15351
rect 22704 15320 22845 15348
rect 22704 15308 22710 15320
rect 22833 15317 22845 15320
rect 22879 15317 22891 15351
rect 22833 15311 22891 15317
rect 1104 15258 23460 15280
rect 1104 15206 6548 15258
rect 6600 15206 6612 15258
rect 6664 15206 6676 15258
rect 6728 15206 6740 15258
rect 6792 15206 6804 15258
rect 6856 15206 12146 15258
rect 12198 15206 12210 15258
rect 12262 15206 12274 15258
rect 12326 15206 12338 15258
rect 12390 15206 12402 15258
rect 12454 15206 17744 15258
rect 17796 15206 17808 15258
rect 17860 15206 17872 15258
rect 17924 15206 17936 15258
rect 17988 15206 18000 15258
rect 18052 15206 23460 15258
rect 1104 15184 23460 15206
rect 1949 15147 2007 15153
rect 1949 15113 1961 15147
rect 1995 15144 2007 15147
rect 2314 15144 2320 15156
rect 1995 15116 2320 15144
rect 1995 15113 2007 15116
rect 1949 15107 2007 15113
rect 2314 15104 2320 15116
rect 2372 15104 2378 15156
rect 2774 15104 2780 15156
rect 2832 15144 2838 15156
rect 2869 15147 2927 15153
rect 2869 15144 2881 15147
rect 2832 15116 2881 15144
rect 2832 15104 2838 15116
rect 2869 15113 2881 15116
rect 2915 15113 2927 15147
rect 2869 15107 2927 15113
rect 3326 15104 3332 15156
rect 3384 15144 3390 15156
rect 4801 15147 4859 15153
rect 4801 15144 4813 15147
rect 3384 15116 4813 15144
rect 3384 15104 3390 15116
rect 4801 15113 4813 15116
rect 4847 15144 4859 15147
rect 6454 15144 6460 15156
rect 4847 15116 6460 15144
rect 4847 15113 4859 15116
rect 4801 15107 4859 15113
rect 6454 15104 6460 15116
rect 6512 15104 6518 15156
rect 11330 15144 11336 15156
rect 11291 15116 11336 15144
rect 11330 15104 11336 15116
rect 11388 15144 11394 15156
rect 11606 15144 11612 15156
rect 11388 15116 11612 15144
rect 11388 15104 11394 15116
rect 11606 15104 11612 15116
rect 11664 15104 11670 15156
rect 13170 15144 13176 15156
rect 13131 15116 13176 15144
rect 13170 15104 13176 15116
rect 13228 15104 13234 15156
rect 16025 15147 16083 15153
rect 16025 15113 16037 15147
rect 16071 15144 16083 15147
rect 18233 15147 18291 15153
rect 16071 15116 16896 15144
rect 16071 15113 16083 15116
rect 16025 15107 16083 15113
rect 3237 15079 3295 15085
rect 3237 15045 3249 15079
rect 3283 15076 3295 15079
rect 3283 15048 6408 15076
rect 3283 15045 3295 15048
rect 3237 15039 3295 15045
rect 1762 15008 1768 15020
rect 1723 14980 1768 15008
rect 1762 14968 1768 14980
rect 1820 14968 1826 15020
rect 2409 15011 2467 15017
rect 2409 14977 2421 15011
rect 2455 15008 2467 15011
rect 2590 15008 2596 15020
rect 2455 14980 2596 15008
rect 2455 14977 2467 14980
rect 2409 14971 2467 14977
rect 2590 14968 2596 14980
rect 2648 14968 2654 15020
rect 4249 15011 4307 15017
rect 4249 14977 4261 15011
rect 4295 15008 4307 15011
rect 4706 15008 4712 15020
rect 4295 14980 4712 15008
rect 4295 14977 4307 14980
rect 4249 14971 4307 14977
rect 4706 14968 4712 14980
rect 4764 14968 4770 15020
rect 5914 15011 5972 15017
rect 5914 15008 5926 15011
rect 5175 14980 5926 15008
rect 1578 14900 1584 14952
rect 1636 14940 1642 14952
rect 2133 14943 2191 14949
rect 2133 14940 2145 14943
rect 1636 14912 2145 14940
rect 1636 14900 1642 14912
rect 2133 14909 2145 14912
rect 2179 14909 2191 14943
rect 2314 14940 2320 14952
rect 2275 14912 2320 14940
rect 2133 14903 2191 14909
rect 2148 14804 2176 14903
rect 2314 14900 2320 14912
rect 2372 14900 2378 14952
rect 3329 14943 3387 14949
rect 3329 14909 3341 14943
rect 3375 14909 3387 14943
rect 3510 14940 3516 14952
rect 3471 14912 3516 14940
rect 3329 14903 3387 14909
rect 2682 14832 2688 14884
rect 2740 14872 2746 14884
rect 2777 14875 2835 14881
rect 2777 14872 2789 14875
rect 2740 14844 2789 14872
rect 2740 14832 2746 14844
rect 2777 14841 2789 14844
rect 2823 14841 2835 14875
rect 2777 14835 2835 14841
rect 3142 14804 3148 14816
rect 2148 14776 3148 14804
rect 3142 14764 3148 14776
rect 3200 14764 3206 14816
rect 3344 14804 3372 14903
rect 3510 14900 3516 14912
rect 3568 14900 3574 14952
rect 4522 14940 4528 14952
rect 4483 14912 4528 14940
rect 4522 14900 4528 14912
rect 4580 14900 4586 14952
rect 3418 14832 3424 14884
rect 3476 14872 3482 14884
rect 5175 14872 5203 14980
rect 5914 14977 5926 14980
rect 5960 15008 5972 15011
rect 6270 15008 6276 15020
rect 5960 14980 6276 15008
rect 5960 14977 5972 14980
rect 5914 14971 5972 14977
rect 6270 14968 6276 14980
rect 6328 14968 6334 15020
rect 6380 15008 6408 15048
rect 8662 15036 8668 15088
rect 8720 15085 8726 15088
rect 8720 15079 8784 15085
rect 8720 15045 8738 15079
rect 8772 15045 8784 15079
rect 8720 15039 8784 15045
rect 10220 15079 10278 15085
rect 10220 15045 10232 15079
rect 10266 15076 10278 15079
rect 10502 15076 10508 15088
rect 10266 15048 10508 15076
rect 10266 15045 10278 15048
rect 10220 15039 10278 15045
rect 8720 15036 8726 15039
rect 10502 15036 10508 15048
rect 10560 15036 10566 15088
rect 14274 15036 14280 15088
rect 14332 15085 14338 15088
rect 14332 15076 14344 15085
rect 16117 15079 16175 15085
rect 16117 15076 16129 15079
rect 14332 15048 14377 15076
rect 14660 15048 16129 15076
rect 14332 15039 14344 15048
rect 14332 15036 14338 15039
rect 6454 15008 6460 15020
rect 6380 14980 6460 15008
rect 6454 14968 6460 14980
rect 6512 14968 6518 15020
rect 14550 15008 14556 15020
rect 14511 14980 14556 15008
rect 14550 14968 14556 14980
rect 14608 15008 14614 15020
rect 14660 15017 14688 15048
rect 16117 15045 16129 15048
rect 16163 15076 16175 15079
rect 16301 15079 16359 15085
rect 16301 15076 16313 15079
rect 16163 15048 16313 15076
rect 16163 15045 16175 15048
rect 16117 15039 16175 15045
rect 16301 15045 16313 15048
rect 16347 15045 16359 15079
rect 16868 15076 16896 15116
rect 18233 15113 18245 15147
rect 18279 15144 18291 15147
rect 18414 15144 18420 15156
rect 18279 15116 18420 15144
rect 18279 15113 18291 15116
rect 18233 15107 18291 15113
rect 18414 15104 18420 15116
rect 18472 15144 18478 15156
rect 18598 15144 18604 15156
rect 18472 15116 18604 15144
rect 18472 15104 18478 15116
rect 18598 15104 18604 15116
rect 18656 15104 18662 15156
rect 19794 15144 19800 15156
rect 19755 15116 19800 15144
rect 19794 15104 19800 15116
rect 19852 15104 19858 15156
rect 20625 15147 20683 15153
rect 20625 15113 20637 15147
rect 20671 15144 20683 15147
rect 21266 15144 21272 15156
rect 20671 15116 21272 15144
rect 20671 15113 20683 15116
rect 20625 15107 20683 15113
rect 21266 15104 21272 15116
rect 21324 15104 21330 15156
rect 21450 15144 21456 15156
rect 21411 15116 21456 15144
rect 21450 15104 21456 15116
rect 21508 15104 21514 15156
rect 21637 15147 21695 15153
rect 21637 15113 21649 15147
rect 21683 15144 21695 15147
rect 21726 15144 21732 15156
rect 21683 15116 21732 15144
rect 21683 15113 21695 15116
rect 21637 15107 21695 15113
rect 21726 15104 21732 15116
rect 21784 15104 21790 15156
rect 21818 15104 21824 15156
rect 21876 15144 21882 15156
rect 22097 15147 22155 15153
rect 22097 15144 22109 15147
rect 21876 15116 22109 15144
rect 21876 15104 21882 15116
rect 22097 15113 22109 15116
rect 22143 15113 22155 15147
rect 22097 15107 22155 15113
rect 16936 15079 16994 15085
rect 16936 15076 16948 15079
rect 16868 15048 16948 15076
rect 16301 15039 16359 15045
rect 16936 15045 16948 15048
rect 16982 15076 16994 15079
rect 20165 15079 20223 15085
rect 20165 15076 20177 15079
rect 16982 15048 20177 15076
rect 16982 15045 16994 15048
rect 16936 15039 16994 15045
rect 20165 15045 20177 15048
rect 20211 15045 20223 15079
rect 20165 15039 20223 15045
rect 22833 15079 22891 15085
rect 22833 15045 22845 15079
rect 22879 15076 22891 15079
rect 22922 15076 22928 15088
rect 22879 15048 22928 15076
rect 22879 15045 22891 15048
rect 22833 15039 22891 15045
rect 14645 15011 14703 15017
rect 14645 15008 14657 15011
rect 14608 14980 14657 15008
rect 14608 14968 14614 14980
rect 14645 14977 14657 14980
rect 14691 14977 14703 15011
rect 14645 14971 14703 14977
rect 14912 15011 14970 15017
rect 14912 14977 14924 15011
rect 14958 15008 14970 15011
rect 16316 15008 16344 15039
rect 22922 15036 22928 15048
rect 22980 15036 22986 15088
rect 16669 15011 16727 15017
rect 16669 15008 16681 15011
rect 14958 14980 16252 15008
rect 16316 14980 16681 15008
rect 14958 14977 14970 14980
rect 14912 14971 14970 14977
rect 6181 14943 6239 14949
rect 6181 14909 6193 14943
rect 6227 14909 6239 14943
rect 8481 14943 8539 14949
rect 8481 14940 8493 14943
rect 6181 14903 6239 14909
rect 8312 14912 8493 14940
rect 3476 14844 5203 14872
rect 3476 14832 3482 14844
rect 6196 14816 6224 14903
rect 5994 14804 6000 14816
rect 3344 14776 6000 14804
rect 5994 14764 6000 14776
rect 6052 14764 6058 14816
rect 6178 14764 6184 14816
rect 6236 14804 6242 14816
rect 8312 14813 8340 14912
rect 8481 14909 8493 14912
rect 8527 14909 8539 14943
rect 8481 14903 8539 14909
rect 9858 14900 9864 14952
rect 9916 14940 9922 14952
rect 9953 14943 10011 14949
rect 9953 14940 9965 14943
rect 9916 14912 9965 14940
rect 9916 14900 9922 14912
rect 9953 14909 9965 14912
rect 9999 14909 10011 14943
rect 16224 14940 16252 14980
rect 16669 14977 16681 14980
rect 16715 14977 16727 15011
rect 18414 15008 18420 15020
rect 18375 14980 18420 15008
rect 16669 14971 16727 14977
rect 18414 14968 18420 14980
rect 18472 14968 18478 15020
rect 18684 15011 18742 15017
rect 18684 15008 18696 15011
rect 18524 14980 18696 15008
rect 16574 14940 16580 14952
rect 16224 14912 16580 14940
rect 9953 14903 10011 14909
rect 16574 14900 16580 14912
rect 16632 14900 16638 14952
rect 18524 14940 18552 14980
rect 18684 14977 18696 14980
rect 18730 15008 18742 15011
rect 20257 15011 20315 15017
rect 20257 15008 20269 15011
rect 18730 14980 20269 15008
rect 18730 14977 18742 14980
rect 18684 14971 18742 14977
rect 20257 14977 20269 14980
rect 20303 14977 20315 15011
rect 21082 15008 21088 15020
rect 21043 14980 21088 15008
rect 20257 14971 20315 14977
rect 21082 14968 21088 14980
rect 21140 14968 21146 15020
rect 21450 14968 21456 15020
rect 21508 15008 21514 15020
rect 22189 15011 22247 15017
rect 22189 15008 22201 15011
rect 21508 14980 22201 15008
rect 21508 14968 21514 14980
rect 22189 14977 22201 14980
rect 22235 14977 22247 15011
rect 22189 14971 22247 14977
rect 18064 14912 18552 14940
rect 20073 14943 20131 14949
rect 10962 14832 10968 14884
rect 11020 14872 11026 14884
rect 18064 14881 18092 14912
rect 20073 14909 20085 14943
rect 20119 14940 20131 14943
rect 20806 14940 20812 14952
rect 20119 14912 20812 14940
rect 20119 14909 20131 14912
rect 20073 14903 20131 14909
rect 20806 14900 20812 14912
rect 20864 14900 20870 14952
rect 20990 14940 20996 14952
rect 20951 14912 20996 14940
rect 20990 14900 20996 14912
rect 21048 14900 21054 14952
rect 22005 14943 22063 14949
rect 22005 14909 22017 14943
rect 22051 14940 22063 14943
rect 22462 14940 22468 14952
rect 22051 14912 22468 14940
rect 22051 14909 22063 14912
rect 22005 14903 22063 14909
rect 22462 14900 22468 14912
rect 22520 14940 22526 14952
rect 22649 14943 22707 14949
rect 22649 14940 22661 14943
rect 22520 14912 22661 14940
rect 22520 14900 22526 14912
rect 22649 14909 22661 14912
rect 22695 14909 22707 14943
rect 22649 14903 22707 14909
rect 11517 14875 11575 14881
rect 11517 14872 11529 14875
rect 11020 14844 11529 14872
rect 11020 14832 11026 14844
rect 11517 14841 11529 14844
rect 11563 14841 11575 14875
rect 11517 14835 11575 14841
rect 18049 14875 18107 14881
rect 18049 14841 18061 14875
rect 18095 14841 18107 14875
rect 18049 14835 18107 14841
rect 22557 14875 22615 14881
rect 22557 14841 22569 14875
rect 22603 14872 22615 14875
rect 23382 14872 23388 14884
rect 22603 14844 23388 14872
rect 22603 14841 22615 14844
rect 22557 14835 22615 14841
rect 23382 14832 23388 14844
rect 23440 14832 23446 14884
rect 6365 14807 6423 14813
rect 6365 14804 6377 14807
rect 6236 14776 6377 14804
rect 6236 14764 6242 14776
rect 6365 14773 6377 14776
rect 6411 14804 6423 14807
rect 6549 14807 6607 14813
rect 6549 14804 6561 14807
rect 6411 14776 6561 14804
rect 6411 14773 6423 14776
rect 6365 14767 6423 14773
rect 6549 14773 6561 14776
rect 6595 14804 6607 14807
rect 7193 14807 7251 14813
rect 7193 14804 7205 14807
rect 6595 14776 7205 14804
rect 6595 14773 6607 14776
rect 6549 14767 6607 14773
rect 7193 14773 7205 14776
rect 7239 14804 7251 14807
rect 8297 14807 8355 14813
rect 8297 14804 8309 14807
rect 7239 14776 8309 14804
rect 7239 14773 7251 14776
rect 7193 14767 7251 14773
rect 8297 14773 8309 14776
rect 8343 14773 8355 14807
rect 8297 14767 8355 14773
rect 9766 14764 9772 14816
rect 9824 14804 9830 14816
rect 9861 14807 9919 14813
rect 9861 14804 9873 14807
rect 9824 14776 9873 14804
rect 9824 14764 9830 14776
rect 9861 14773 9873 14776
rect 9907 14773 9919 14807
rect 9861 14767 9919 14773
rect 18138 14764 18144 14816
rect 18196 14804 18202 14816
rect 21726 14804 21732 14816
rect 18196 14776 21732 14804
rect 18196 14764 18202 14776
rect 21726 14764 21732 14776
rect 21784 14764 21790 14816
rect 23106 14804 23112 14816
rect 23067 14776 23112 14804
rect 23106 14764 23112 14776
rect 23164 14764 23170 14816
rect 1104 14714 23460 14736
rect 1104 14662 3749 14714
rect 3801 14662 3813 14714
rect 3865 14662 3877 14714
rect 3929 14662 3941 14714
rect 3993 14662 4005 14714
rect 4057 14662 9347 14714
rect 9399 14662 9411 14714
rect 9463 14662 9475 14714
rect 9527 14662 9539 14714
rect 9591 14662 9603 14714
rect 9655 14662 14945 14714
rect 14997 14662 15009 14714
rect 15061 14662 15073 14714
rect 15125 14662 15137 14714
rect 15189 14662 15201 14714
rect 15253 14662 20543 14714
rect 20595 14662 20607 14714
rect 20659 14662 20671 14714
rect 20723 14662 20735 14714
rect 20787 14662 20799 14714
rect 20851 14662 23460 14714
rect 1104 14640 23460 14662
rect 1673 14603 1731 14609
rect 1673 14569 1685 14603
rect 1719 14600 1731 14603
rect 2314 14600 2320 14612
rect 1719 14572 2320 14600
rect 1719 14569 1731 14572
rect 1673 14563 1731 14569
rect 2314 14560 2320 14572
rect 2372 14560 2378 14612
rect 2406 14560 2412 14612
rect 2464 14600 2470 14612
rect 2869 14603 2927 14609
rect 2869 14600 2881 14603
rect 2464 14572 2881 14600
rect 2464 14560 2470 14572
rect 2869 14569 2881 14572
rect 2915 14569 2927 14603
rect 8478 14600 8484 14612
rect 2869 14563 2927 14569
rect 4172 14572 8484 14600
rect 1949 14535 2007 14541
rect 1949 14501 1961 14535
rect 1995 14532 2007 14535
rect 2958 14532 2964 14544
rect 1995 14504 2964 14532
rect 1995 14501 2007 14504
rect 1949 14495 2007 14501
rect 2958 14492 2964 14504
rect 3016 14492 3022 14544
rect 3418 14532 3424 14544
rect 3252 14504 3424 14532
rect 1394 14424 1400 14476
rect 1452 14464 1458 14476
rect 2593 14467 2651 14473
rect 2593 14464 2605 14467
rect 1452 14436 2605 14464
rect 1452 14424 1458 14436
rect 2593 14433 2605 14436
rect 2639 14464 2651 14467
rect 2682 14464 2688 14476
rect 2639 14436 2688 14464
rect 2639 14433 2651 14436
rect 2593 14427 2651 14433
rect 2682 14424 2688 14436
rect 2740 14424 2746 14476
rect 1489 14399 1547 14405
rect 1489 14365 1501 14399
rect 1535 14365 1547 14399
rect 1489 14359 1547 14365
rect 1765 14399 1823 14405
rect 1765 14365 1777 14399
rect 1811 14396 1823 14399
rect 2314 14396 2320 14408
rect 1811 14368 2320 14396
rect 1811 14365 1823 14368
rect 1765 14359 1823 14365
rect 1504 14328 1532 14359
rect 2314 14356 2320 14368
rect 2372 14356 2378 14408
rect 2501 14399 2559 14405
rect 2501 14365 2513 14399
rect 2547 14396 2559 14399
rect 2866 14396 2872 14408
rect 2547 14368 2872 14396
rect 2547 14365 2559 14368
rect 2501 14359 2559 14365
rect 2866 14356 2872 14368
rect 2924 14356 2930 14408
rect 3252 14405 3280 14504
rect 3418 14492 3424 14504
rect 3476 14492 3482 14544
rect 3510 14464 3516 14476
rect 3471 14436 3516 14464
rect 3510 14424 3516 14436
rect 3568 14424 3574 14476
rect 3237 14399 3295 14405
rect 3237 14365 3249 14399
rect 3283 14365 3295 14399
rect 3237 14359 3295 14365
rect 3329 14399 3387 14405
rect 3329 14365 3341 14399
rect 3375 14396 3387 14399
rect 4062 14396 4068 14408
rect 3375 14368 4068 14396
rect 3375 14365 3387 14368
rect 3329 14359 3387 14365
rect 4062 14356 4068 14368
rect 4120 14356 4126 14408
rect 4172 14337 4200 14572
rect 8478 14560 8484 14572
rect 8536 14560 8542 14612
rect 12253 14603 12311 14609
rect 12253 14569 12265 14603
rect 12299 14600 12311 14603
rect 12526 14600 12532 14612
rect 12299 14572 12532 14600
rect 12299 14569 12311 14572
rect 12253 14563 12311 14569
rect 12526 14560 12532 14572
rect 12584 14560 12590 14612
rect 15473 14603 15531 14609
rect 15473 14569 15485 14603
rect 15519 14600 15531 14603
rect 16574 14600 16580 14612
rect 15519 14572 16580 14600
rect 15519 14569 15531 14572
rect 15473 14563 15531 14569
rect 16574 14560 16580 14572
rect 16632 14560 16638 14612
rect 17129 14603 17187 14609
rect 17129 14569 17141 14603
rect 17175 14600 17187 14603
rect 18414 14600 18420 14612
rect 17175 14572 18420 14600
rect 17175 14569 17187 14572
rect 17129 14563 17187 14569
rect 4614 14492 4620 14544
rect 4672 14532 4678 14544
rect 4801 14535 4859 14541
rect 4801 14532 4813 14535
rect 4672 14504 4813 14532
rect 4672 14492 4678 14504
rect 4801 14501 4813 14504
rect 4847 14501 4859 14535
rect 6362 14532 6368 14544
rect 6323 14504 6368 14532
rect 4801 14495 4859 14501
rect 6362 14492 6368 14504
rect 6420 14492 6426 14544
rect 9125 14535 9183 14541
rect 9125 14532 9137 14535
rect 7944 14504 9137 14532
rect 4433 14467 4491 14473
rect 4433 14433 4445 14467
rect 4479 14464 4491 14467
rect 4706 14464 4712 14476
rect 4479 14436 4712 14464
rect 4479 14433 4491 14436
rect 4433 14427 4491 14433
rect 4706 14424 4712 14436
rect 4764 14424 4770 14476
rect 6178 14396 6184 14408
rect 6139 14368 6184 14396
rect 6178 14356 6184 14368
rect 6236 14396 6242 14408
rect 7745 14399 7803 14405
rect 7745 14396 7757 14399
rect 6236 14368 7757 14396
rect 6236 14356 6242 14368
rect 7745 14365 7757 14368
rect 7791 14396 7803 14399
rect 7837 14399 7895 14405
rect 7837 14396 7849 14399
rect 7791 14368 7849 14396
rect 7791 14365 7803 14368
rect 7745 14359 7803 14365
rect 7837 14365 7849 14368
rect 7883 14365 7895 14399
rect 7837 14359 7895 14365
rect 2409 14331 2467 14337
rect 1504 14300 2084 14328
rect 2056 14269 2084 14300
rect 2409 14297 2421 14331
rect 2455 14328 2467 14331
rect 4157 14331 4215 14337
rect 2455 14300 3832 14328
rect 2455 14297 2467 14300
rect 2409 14291 2467 14297
rect 3804 14269 3832 14300
rect 4157 14297 4169 14331
rect 4203 14297 4215 14331
rect 4157 14291 4215 14297
rect 4249 14331 4307 14337
rect 4249 14297 4261 14331
rect 4295 14328 4307 14331
rect 5810 14328 5816 14340
rect 4295 14300 5816 14328
rect 4295 14297 4307 14300
rect 4249 14291 4307 14297
rect 5810 14288 5816 14300
rect 5868 14288 5874 14340
rect 5902 14288 5908 14340
rect 5960 14337 5966 14340
rect 5960 14331 5994 14337
rect 5982 14328 5994 14331
rect 5982 14300 7420 14328
rect 5982 14297 5994 14300
rect 5960 14291 5994 14297
rect 5960 14288 5966 14291
rect 2041 14263 2099 14269
rect 2041 14229 2053 14263
rect 2087 14229 2099 14263
rect 2041 14223 2099 14229
rect 3789 14263 3847 14269
rect 3789 14229 3801 14263
rect 3835 14229 3847 14263
rect 3789 14223 3847 14229
rect 3878 14220 3884 14272
rect 3936 14260 3942 14272
rect 6362 14260 6368 14272
rect 3936 14232 6368 14260
rect 3936 14220 3942 14232
rect 6362 14220 6368 14232
rect 6420 14220 6426 14272
rect 7392 14260 7420 14300
rect 7466 14288 7472 14340
rect 7524 14337 7530 14340
rect 7524 14328 7536 14337
rect 7944 14328 7972 14504
rect 9125 14501 9137 14504
rect 9171 14501 9183 14535
rect 9125 14495 9183 14501
rect 16942 14424 16948 14476
rect 17000 14464 17006 14476
rect 17144 14464 17172 14563
rect 18414 14560 18420 14572
rect 18472 14600 18478 14612
rect 18785 14603 18843 14609
rect 18785 14600 18797 14603
rect 18472 14572 18797 14600
rect 18472 14560 18478 14572
rect 18785 14569 18797 14572
rect 18831 14600 18843 14603
rect 18969 14603 19027 14609
rect 18969 14600 18981 14603
rect 18831 14572 18981 14600
rect 18831 14569 18843 14572
rect 18785 14563 18843 14569
rect 18969 14569 18981 14572
rect 19015 14569 19027 14603
rect 18969 14563 19027 14569
rect 18693 14535 18751 14541
rect 18693 14501 18705 14535
rect 18739 14532 18751 14535
rect 18874 14532 18880 14544
rect 18739 14504 18880 14532
rect 18739 14501 18751 14504
rect 18693 14495 18751 14501
rect 18874 14492 18880 14504
rect 18932 14492 18938 14544
rect 17000 14436 17172 14464
rect 18984 14464 19012 14563
rect 19426 14560 19432 14612
rect 19484 14600 19490 14612
rect 21450 14600 21456 14612
rect 19484 14572 20208 14600
rect 21411 14572 21456 14600
rect 19484 14560 19490 14572
rect 20180 14532 20208 14572
rect 21450 14560 21456 14572
rect 21508 14560 21514 14612
rect 21542 14560 21548 14612
rect 21600 14600 21606 14612
rect 21910 14600 21916 14612
rect 21600 14572 21916 14600
rect 21600 14560 21606 14572
rect 21910 14560 21916 14572
rect 21968 14600 21974 14612
rect 22738 14600 22744 14612
rect 21968 14572 22744 14600
rect 21968 14560 21974 14572
rect 22738 14560 22744 14572
rect 22796 14600 22802 14612
rect 23017 14603 23075 14609
rect 23017 14600 23029 14603
rect 22796 14572 23029 14600
rect 22796 14560 22802 14572
rect 23017 14569 23029 14572
rect 23063 14569 23075 14603
rect 23017 14563 23075 14569
rect 23474 14532 23480 14544
rect 20180 14504 23480 14532
rect 23474 14492 23480 14504
rect 23532 14492 23538 14544
rect 19242 14464 19248 14476
rect 18984 14436 19248 14464
rect 17000 14424 17006 14436
rect 19242 14424 19248 14436
rect 19300 14424 19306 14476
rect 20806 14424 20812 14476
rect 20864 14464 20870 14476
rect 20901 14467 20959 14473
rect 20901 14464 20913 14467
rect 20864 14436 20913 14464
rect 20864 14424 20870 14436
rect 20901 14433 20913 14436
rect 20947 14464 20959 14467
rect 22373 14467 22431 14473
rect 22373 14464 22385 14467
rect 20947 14436 22385 14464
rect 20947 14433 20959 14436
rect 20901 14427 20959 14433
rect 22373 14433 22385 14436
rect 22419 14433 22431 14467
rect 22373 14427 22431 14433
rect 10505 14399 10563 14405
rect 10505 14365 10517 14399
rect 10551 14365 10563 14399
rect 10505 14359 10563 14365
rect 7524 14300 7972 14328
rect 7524 14291 7536 14300
rect 7524 14288 7530 14291
rect 9950 14288 9956 14340
rect 10008 14328 10014 14340
rect 10238 14331 10296 14337
rect 10238 14328 10250 14331
rect 10008 14300 10250 14328
rect 10008 14288 10014 14300
rect 10238 14297 10250 14300
rect 10284 14297 10296 14331
rect 10238 14291 10296 14297
rect 9674 14260 9680 14272
rect 7392 14232 9680 14260
rect 9674 14220 9680 14232
rect 9732 14220 9738 14272
rect 9858 14220 9864 14272
rect 9916 14260 9922 14272
rect 10520 14260 10548 14359
rect 13354 14356 13360 14408
rect 13412 14405 13418 14408
rect 13412 14396 13424 14405
rect 13538 14396 13544 14408
rect 13412 14368 13544 14396
rect 13412 14359 13424 14368
rect 13412 14356 13418 14359
rect 13538 14356 13544 14368
rect 13596 14356 13602 14408
rect 13633 14399 13691 14405
rect 13633 14365 13645 14399
rect 13679 14396 13691 14399
rect 13817 14399 13875 14405
rect 13817 14396 13829 14399
rect 13679 14368 13829 14396
rect 13679 14365 13691 14368
rect 13633 14359 13691 14365
rect 13817 14365 13829 14368
rect 13863 14396 13875 14399
rect 14090 14396 14096 14408
rect 13863 14368 14096 14396
rect 13863 14365 13875 14368
rect 13817 14359 13875 14365
rect 14090 14356 14096 14368
rect 14148 14356 14154 14408
rect 17218 14396 17224 14408
rect 14292 14368 17224 14396
rect 13262 14288 13268 14340
rect 13320 14328 13326 14340
rect 14292 14328 14320 14368
rect 17218 14356 17224 14368
rect 17276 14356 17282 14408
rect 19150 14356 19156 14408
rect 19208 14396 19214 14408
rect 19512 14399 19570 14405
rect 19512 14396 19524 14399
rect 19208 14368 19524 14396
rect 19208 14356 19214 14368
rect 19512 14365 19524 14368
rect 19558 14396 19570 14399
rect 20714 14396 20720 14408
rect 19558 14368 20720 14396
rect 19558 14365 19570 14368
rect 19512 14359 19570 14365
rect 20714 14356 20720 14368
rect 20772 14356 20778 14408
rect 21634 14396 21640 14408
rect 21595 14368 21640 14396
rect 21634 14356 21640 14368
rect 21692 14356 21698 14408
rect 21726 14356 21732 14408
rect 21784 14396 21790 14408
rect 21821 14399 21879 14405
rect 21821 14396 21833 14399
rect 21784 14368 21833 14396
rect 21784 14356 21790 14368
rect 21821 14365 21833 14368
rect 21867 14365 21879 14399
rect 21821 14359 21879 14365
rect 22097 14399 22155 14405
rect 22097 14365 22109 14399
rect 22143 14396 22155 14399
rect 22186 14396 22192 14408
rect 22143 14368 22192 14396
rect 22143 14365 22155 14368
rect 22097 14359 22155 14365
rect 22186 14356 22192 14368
rect 22244 14396 22250 14408
rect 22922 14396 22928 14408
rect 22244 14368 22928 14396
rect 22244 14356 22250 14368
rect 22922 14356 22928 14368
rect 22980 14356 22986 14408
rect 13320 14300 14320 14328
rect 14360 14331 14418 14337
rect 13320 14288 13326 14300
rect 14360 14297 14372 14331
rect 14406 14328 14418 14331
rect 14734 14328 14740 14340
rect 14406 14300 14740 14328
rect 14406 14297 14418 14300
rect 14360 14291 14418 14297
rect 14734 14288 14740 14300
rect 14792 14288 14798 14340
rect 16666 14288 16672 14340
rect 16724 14337 16730 14340
rect 16724 14328 16736 14337
rect 18325 14331 18383 14337
rect 16724 14300 16769 14328
rect 16724 14291 16736 14300
rect 18325 14297 18337 14331
rect 18371 14328 18383 14331
rect 19426 14328 19432 14340
rect 18371 14300 19432 14328
rect 18371 14297 18383 14300
rect 18325 14291 18383 14297
rect 16724 14288 16730 14291
rect 19426 14288 19432 14300
rect 19484 14288 19490 14340
rect 19610 14288 19616 14340
rect 19668 14328 19674 14340
rect 21085 14331 21143 14337
rect 21085 14328 21097 14331
rect 19668 14300 21097 14328
rect 19668 14288 19674 14300
rect 21085 14297 21097 14300
rect 21131 14297 21143 14331
rect 21085 14291 21143 14297
rect 10597 14263 10655 14269
rect 10597 14260 10609 14263
rect 9916 14232 10609 14260
rect 9916 14220 9922 14232
rect 10597 14229 10609 14232
rect 10643 14260 10655 14263
rect 10781 14263 10839 14269
rect 10781 14260 10793 14263
rect 10643 14232 10793 14260
rect 10643 14229 10655 14232
rect 10597 14223 10655 14229
rect 10781 14229 10793 14232
rect 10827 14260 10839 14263
rect 10962 14260 10968 14272
rect 10827 14232 10968 14260
rect 10827 14229 10839 14232
rect 10781 14223 10839 14229
rect 10962 14220 10968 14232
rect 11020 14260 11026 14272
rect 11425 14263 11483 14269
rect 11425 14260 11437 14263
rect 11020 14232 11437 14260
rect 11020 14220 11026 14232
rect 11425 14229 11437 14232
rect 11471 14229 11483 14263
rect 11425 14223 11483 14229
rect 15565 14263 15623 14269
rect 15565 14229 15577 14263
rect 15611 14260 15623 14263
rect 15746 14260 15752 14272
rect 15611 14232 15752 14260
rect 15611 14229 15623 14232
rect 15565 14223 15623 14229
rect 15746 14220 15752 14232
rect 15804 14220 15810 14272
rect 18509 14263 18567 14269
rect 18509 14229 18521 14263
rect 18555 14260 18567 14263
rect 20254 14260 20260 14272
rect 18555 14232 20260 14260
rect 18555 14229 18567 14232
rect 18509 14223 18567 14229
rect 20254 14220 20260 14232
rect 20312 14220 20318 14272
rect 20530 14220 20536 14272
rect 20588 14260 20594 14272
rect 20625 14263 20683 14269
rect 20625 14260 20637 14263
rect 20588 14232 20637 14260
rect 20588 14220 20594 14232
rect 20625 14229 20637 14232
rect 20671 14260 20683 14263
rect 20993 14263 21051 14269
rect 20993 14260 21005 14263
rect 20671 14232 21005 14260
rect 20671 14229 20683 14232
rect 20625 14223 20683 14229
rect 20993 14229 21005 14232
rect 21039 14229 21051 14263
rect 20993 14223 21051 14229
rect 21726 14220 21732 14272
rect 21784 14260 21790 14272
rect 22005 14263 22063 14269
rect 22005 14260 22017 14263
rect 21784 14232 22017 14260
rect 21784 14220 21790 14232
rect 22005 14229 22017 14232
rect 22051 14229 22063 14263
rect 22005 14223 22063 14229
rect 1104 14170 23460 14192
rect 1104 14118 6548 14170
rect 6600 14118 6612 14170
rect 6664 14118 6676 14170
rect 6728 14118 6740 14170
rect 6792 14118 6804 14170
rect 6856 14118 12146 14170
rect 12198 14118 12210 14170
rect 12262 14118 12274 14170
rect 12326 14118 12338 14170
rect 12390 14118 12402 14170
rect 12454 14118 17744 14170
rect 17796 14118 17808 14170
rect 17860 14118 17872 14170
rect 17924 14118 17936 14170
rect 17988 14118 18000 14170
rect 18052 14118 23460 14170
rect 1104 14096 23460 14118
rect 2314 14056 2320 14068
rect 2275 14028 2320 14056
rect 2314 14016 2320 14028
rect 2372 14016 2378 14068
rect 2685 14059 2743 14065
rect 2685 14025 2697 14059
rect 2731 14056 2743 14059
rect 3145 14059 3203 14065
rect 3145 14056 3157 14059
rect 2731 14028 3157 14056
rect 2731 14025 2743 14028
rect 2685 14019 2743 14025
rect 3145 14025 3157 14028
rect 3191 14025 3203 14059
rect 3145 14019 3203 14025
rect 3513 14059 3571 14065
rect 3513 14025 3525 14059
rect 3559 14056 3571 14059
rect 3878 14056 3884 14068
rect 3559 14028 3884 14056
rect 3559 14025 3571 14028
rect 3513 14019 3571 14025
rect 3878 14016 3884 14028
rect 3936 14016 3942 14068
rect 3973 14059 4031 14065
rect 3973 14025 3985 14059
rect 4019 14025 4031 14059
rect 3973 14019 4031 14025
rect 2777 13991 2835 13997
rect 2777 13957 2789 13991
rect 2823 13988 2835 13991
rect 3988 13988 4016 14019
rect 4154 14016 4160 14068
rect 4212 14056 4218 14068
rect 4801 14059 4859 14065
rect 4801 14056 4813 14059
rect 4212 14028 4813 14056
rect 4212 14016 4218 14028
rect 4801 14025 4813 14028
rect 4847 14056 4859 14059
rect 5166 14056 5172 14068
rect 4847 14028 5172 14056
rect 4847 14025 4859 14028
rect 4801 14019 4859 14025
rect 5166 14016 5172 14028
rect 5224 14016 5230 14068
rect 5810 14016 5816 14068
rect 5868 14056 5874 14068
rect 8478 14056 8484 14068
rect 5868 14028 8340 14056
rect 8439 14028 8484 14056
rect 5868 14016 5874 14028
rect 2823 13960 4016 13988
rect 4264 13960 6500 13988
rect 2823 13957 2835 13960
rect 2777 13951 2835 13957
rect 3605 13923 3663 13929
rect 3605 13889 3617 13923
rect 3651 13920 3663 13923
rect 4264 13920 4292 13960
rect 3651 13892 4292 13920
rect 4341 13923 4399 13929
rect 3651 13889 3663 13892
rect 3605 13883 3663 13889
rect 4341 13889 4353 13923
rect 4387 13920 4399 13923
rect 5626 13920 5632 13932
rect 4387 13892 5632 13920
rect 4387 13889 4399 13892
rect 4341 13883 4399 13889
rect 5626 13880 5632 13892
rect 5684 13880 5690 13932
rect 5925 13923 5983 13929
rect 5925 13889 5937 13923
rect 5971 13920 5983 13923
rect 6362 13920 6368 13932
rect 5971 13892 6368 13920
rect 5971 13889 5983 13892
rect 5925 13883 5983 13889
rect 6362 13880 6368 13892
rect 6420 13880 6426 13932
rect 6472 13920 6500 13960
rect 6546 13948 6552 14000
rect 6604 13988 6610 14000
rect 8312 13988 8340 14028
rect 8478 14016 8484 14028
rect 8536 14016 8542 14068
rect 9950 14056 9956 14068
rect 9863 14028 9956 14056
rect 9594 13991 9652 13997
rect 9594 13988 9606 13991
rect 6604 13960 8248 13988
rect 8312 13960 9606 13988
rect 6604 13948 6610 13960
rect 7466 13920 7472 13932
rect 6472 13892 7472 13920
rect 7466 13880 7472 13892
rect 7524 13880 7530 13932
rect 7834 13880 7840 13932
rect 7892 13929 7898 13932
rect 7892 13920 7904 13929
rect 8113 13923 8171 13929
rect 7892 13892 7937 13920
rect 7892 13883 7904 13892
rect 8113 13889 8125 13923
rect 8159 13889 8171 13923
rect 8220 13920 8248 13960
rect 9594 13957 9606 13960
rect 9640 13988 9652 13991
rect 9766 13988 9772 14000
rect 9640 13960 9772 13988
rect 9640 13957 9652 13960
rect 9594 13951 9652 13957
rect 9766 13948 9772 13960
rect 9824 13948 9830 14000
rect 9876 13920 9904 14028
rect 9950 14016 9956 14028
rect 10008 14016 10014 14068
rect 11238 14016 11244 14068
rect 11296 14056 11302 14068
rect 11517 14059 11575 14065
rect 11517 14056 11529 14059
rect 11296 14028 11529 14056
rect 11296 14016 11302 14028
rect 11517 14025 11529 14028
rect 11563 14025 11575 14059
rect 14734 14056 14740 14068
rect 14695 14028 14740 14056
rect 11517 14019 11575 14025
rect 14734 14016 14740 14028
rect 14792 14016 14798 14068
rect 16761 14059 16819 14065
rect 16761 14025 16773 14059
rect 16807 14056 16819 14059
rect 16942 14056 16948 14068
rect 16807 14028 16948 14056
rect 16807 14025 16819 14028
rect 16761 14019 16819 14025
rect 10962 13948 10968 14000
rect 11020 13988 11026 14000
rect 12652 13991 12710 13997
rect 11020 13960 11376 13988
rect 11020 13948 11026 13960
rect 11348 13929 11376 13960
rect 12652 13957 12664 13991
rect 12698 13988 12710 13991
rect 13262 13988 13268 14000
rect 12698 13960 13268 13988
rect 12698 13957 12710 13960
rect 12652 13951 12710 13957
rect 13262 13948 13268 13960
rect 13320 13948 13326 14000
rect 14090 13988 14096 14000
rect 13372 13960 14096 13988
rect 11066 13923 11124 13929
rect 11066 13920 11078 13923
rect 8220 13892 9904 13920
rect 10060 13892 11078 13920
rect 8113 13883 8171 13889
rect 7892 13880 7898 13883
rect 2682 13812 2688 13864
rect 2740 13852 2746 13864
rect 2869 13855 2927 13861
rect 2740 13812 2774 13852
rect 2869 13821 2881 13855
rect 2915 13821 2927 13855
rect 2869 13815 2927 13821
rect 3789 13855 3847 13861
rect 3789 13821 3801 13855
rect 3835 13821 3847 13855
rect 4430 13852 4436 13864
rect 4391 13824 4436 13852
rect 3789 13815 3847 13821
rect 2746 13784 2774 13812
rect 2884 13784 2912 13815
rect 2746 13756 2912 13784
rect 3804 13784 3832 13815
rect 4430 13812 4436 13824
rect 4488 13812 4494 13864
rect 4617 13855 4675 13861
rect 4617 13821 4629 13855
rect 4663 13852 4675 13855
rect 4706 13852 4712 13864
rect 4663 13824 4712 13852
rect 4663 13821 4675 13824
rect 4617 13815 4675 13821
rect 4632 13784 4660 13815
rect 4706 13812 4712 13824
rect 4764 13812 4770 13864
rect 6178 13852 6184 13864
rect 6139 13824 6184 13852
rect 6178 13812 6184 13824
rect 6236 13812 6242 13864
rect 6454 13812 6460 13864
rect 6512 13852 6518 13864
rect 8128 13852 8156 13883
rect 9858 13852 9864 13864
rect 6512 13824 6776 13852
rect 8128 13824 8248 13852
rect 9819 13824 9864 13852
rect 6512 13812 6518 13824
rect 6748 13793 6776 13824
rect 3804 13756 4660 13784
rect 6733 13787 6791 13793
rect 6733 13753 6745 13787
rect 6779 13753 6791 13787
rect 6733 13747 6791 13753
rect 6178 13676 6184 13728
rect 6236 13716 6242 13728
rect 8220 13725 8248 13824
rect 9858 13812 9864 13824
rect 9916 13812 9922 13864
rect 10060 13852 10088 13892
rect 11066 13889 11078 13892
rect 11112 13889 11124 13923
rect 11066 13883 11124 13889
rect 11333 13923 11391 13929
rect 11333 13889 11345 13923
rect 11379 13889 11391 13923
rect 11333 13883 11391 13889
rect 12897 13923 12955 13929
rect 12897 13889 12909 13923
rect 12943 13920 12955 13923
rect 13078 13920 13084 13932
rect 12943 13892 13084 13920
rect 12943 13889 12955 13892
rect 12897 13883 12955 13889
rect 13078 13880 13084 13892
rect 13136 13920 13142 13932
rect 13372 13929 13400 13960
rect 14090 13948 14096 13960
rect 14148 13988 14154 14000
rect 14921 13991 14979 13997
rect 14921 13988 14933 13991
rect 14148 13960 14933 13988
rect 14148 13948 14154 13960
rect 14921 13957 14933 13960
rect 14967 13988 14979 13991
rect 16776 13988 16804 14019
rect 16942 14016 16948 14028
rect 17000 14056 17006 14068
rect 17037 14059 17095 14065
rect 17037 14056 17049 14059
rect 17000 14028 17049 14056
rect 17000 14016 17006 14028
rect 17037 14025 17049 14028
rect 17083 14025 17095 14059
rect 17037 14019 17095 14025
rect 17773 14059 17831 14065
rect 17773 14025 17785 14059
rect 17819 14056 17831 14059
rect 18138 14056 18144 14068
rect 17819 14028 18144 14056
rect 17819 14025 17831 14028
rect 17773 14019 17831 14025
rect 18138 14016 18144 14028
rect 18196 14056 18202 14068
rect 18874 14056 18880 14068
rect 18196 14028 18880 14056
rect 18196 14016 18202 14028
rect 18874 14016 18880 14028
rect 18932 14016 18938 14068
rect 19242 14016 19248 14068
rect 19300 14056 19306 14068
rect 21542 14056 21548 14068
rect 19300 14028 21548 14056
rect 19300 14016 19306 14028
rect 19334 13988 19340 14000
rect 14967 13960 16804 13988
rect 18432 13960 19340 13988
rect 14967 13957 14979 13960
rect 14921 13951 14979 13957
rect 13357 13923 13415 13929
rect 13357 13920 13369 13923
rect 13136 13892 13369 13920
rect 13136 13880 13142 13892
rect 13357 13889 13369 13892
rect 13403 13889 13415 13923
rect 13357 13883 13415 13889
rect 13624 13923 13682 13929
rect 13624 13889 13636 13923
rect 13670 13920 13682 13923
rect 14182 13920 14188 13932
rect 13670 13892 14188 13920
rect 13670 13889 13682 13892
rect 13624 13883 13682 13889
rect 14182 13880 14188 13892
rect 14240 13880 14246 13932
rect 15120 13929 15148 13960
rect 15378 13929 15384 13932
rect 15105 13923 15163 13929
rect 15105 13889 15117 13923
rect 15151 13889 15163 13923
rect 15105 13883 15163 13889
rect 15372 13883 15384 13929
rect 15436 13920 15442 13932
rect 16666 13920 16672 13932
rect 15436 13892 15472 13920
rect 16500 13892 16672 13920
rect 15378 13880 15384 13883
rect 15436 13880 15442 13892
rect 9968 13824 10088 13852
rect 9968 13784 9996 13824
rect 16500 13793 16528 13892
rect 16666 13880 16672 13892
rect 16724 13920 16730 13932
rect 18432 13920 18460 13960
rect 19334 13948 19340 13960
rect 19392 13948 19398 14000
rect 16724 13892 18460 13920
rect 18897 13923 18955 13929
rect 16724 13880 16730 13892
rect 18897 13889 18909 13923
rect 18943 13920 18955 13923
rect 19153 13923 19211 13929
rect 18943 13892 19104 13920
rect 18943 13889 18955 13892
rect 18897 13883 18955 13889
rect 19076 13852 19104 13892
rect 19153 13889 19165 13923
rect 19199 13920 19211 13923
rect 19242 13920 19248 13932
rect 19199 13892 19248 13920
rect 19199 13889 19211 13892
rect 19153 13883 19211 13889
rect 19242 13880 19248 13892
rect 19300 13880 19306 13932
rect 20369 13923 20427 13929
rect 20369 13889 20381 13923
rect 20415 13920 20427 13923
rect 20530 13920 20536 13932
rect 20415 13892 20536 13920
rect 20415 13889 20427 13892
rect 20369 13883 20427 13889
rect 20530 13880 20536 13892
rect 20588 13880 20594 13932
rect 20640 13929 20668 14028
rect 21542 14016 21548 14028
rect 21600 14016 21606 14068
rect 22922 14056 22928 14068
rect 22883 14028 22928 14056
rect 22922 14016 22928 14028
rect 22980 14016 22986 14068
rect 20714 13948 20720 14000
rect 20772 13988 20778 14000
rect 21085 13991 21143 13997
rect 21085 13988 21097 13991
rect 20772 13960 21097 13988
rect 20772 13948 20778 13960
rect 21085 13957 21097 13960
rect 21131 13957 21143 13991
rect 21085 13951 21143 13957
rect 22097 13991 22155 13997
rect 22097 13957 22109 13991
rect 22143 13988 22155 13991
rect 22554 13988 22560 14000
rect 22143 13960 22560 13988
rect 22143 13957 22155 13960
rect 22097 13951 22155 13957
rect 22554 13948 22560 13960
rect 22612 13948 22618 14000
rect 20625 13923 20683 13929
rect 20625 13889 20637 13923
rect 20671 13889 20683 13923
rect 20625 13883 20683 13889
rect 21910 13880 21916 13932
rect 21968 13920 21974 13932
rect 22189 13923 22247 13929
rect 22189 13920 22201 13923
rect 21968 13892 22201 13920
rect 21968 13880 21974 13892
rect 22189 13889 22201 13892
rect 22235 13889 22247 13923
rect 22649 13923 22707 13929
rect 22649 13920 22661 13923
rect 22189 13883 22247 13889
rect 22572 13892 22661 13920
rect 19610 13852 19616 13864
rect 19076 13824 19616 13852
rect 19260 13793 19288 13824
rect 19610 13812 19616 13824
rect 19668 13812 19674 13864
rect 20806 13852 20812 13864
rect 20767 13824 20812 13852
rect 20806 13812 20812 13824
rect 20864 13812 20870 13864
rect 20990 13852 20996 13864
rect 20951 13824 20996 13852
rect 20990 13812 20996 13824
rect 21048 13812 21054 13864
rect 21818 13852 21824 13864
rect 21468 13824 21824 13852
rect 9876 13756 9996 13784
rect 16485 13787 16543 13793
rect 6365 13719 6423 13725
rect 6365 13716 6377 13719
rect 6236 13688 6377 13716
rect 6236 13676 6242 13688
rect 6365 13685 6377 13688
rect 6411 13716 6423 13719
rect 6549 13719 6607 13725
rect 6549 13716 6561 13719
rect 6411 13688 6561 13716
rect 6411 13685 6423 13688
rect 6365 13679 6423 13685
rect 6549 13685 6561 13688
rect 6595 13716 6607 13719
rect 8205 13719 8263 13725
rect 8205 13716 8217 13719
rect 6595 13688 8217 13716
rect 6595 13685 6607 13688
rect 6549 13679 6607 13685
rect 8205 13685 8217 13688
rect 8251 13685 8263 13719
rect 8205 13679 8263 13685
rect 8386 13676 8392 13728
rect 8444 13716 8450 13728
rect 9876 13716 9904 13756
rect 16485 13753 16497 13787
rect 16531 13753 16543 13787
rect 16485 13747 16543 13753
rect 19245 13787 19303 13793
rect 19245 13753 19257 13787
rect 19291 13753 19303 13787
rect 20824 13784 20852 13812
rect 21082 13784 21088 13796
rect 20824 13756 21088 13784
rect 19245 13747 19303 13753
rect 21082 13744 21088 13756
rect 21140 13744 21146 13796
rect 21468 13793 21496 13824
rect 21818 13812 21824 13824
rect 21876 13812 21882 13864
rect 22005 13855 22063 13861
rect 22005 13821 22017 13855
rect 22051 13821 22063 13855
rect 22005 13815 22063 13821
rect 21453 13787 21511 13793
rect 21453 13753 21465 13787
rect 21499 13753 21511 13787
rect 22020 13784 22048 13815
rect 22572 13793 22600 13892
rect 22649 13889 22661 13892
rect 22695 13889 22707 13923
rect 23106 13920 23112 13932
rect 23067 13892 23112 13920
rect 22649 13883 22707 13889
rect 23106 13880 23112 13892
rect 23164 13880 23170 13932
rect 22557 13787 22615 13793
rect 22020 13756 22094 13784
rect 21453 13747 21511 13753
rect 8444 13688 9904 13716
rect 8444 13676 8450 13688
rect 15746 13676 15752 13728
rect 15804 13716 15810 13728
rect 21266 13716 21272 13728
rect 15804 13688 21272 13716
rect 15804 13676 15810 13688
rect 21266 13676 21272 13688
rect 21324 13676 21330 13728
rect 21358 13676 21364 13728
rect 21416 13716 21422 13728
rect 21818 13716 21824 13728
rect 21416 13688 21824 13716
rect 21416 13676 21422 13688
rect 21818 13676 21824 13688
rect 21876 13676 21882 13728
rect 22066 13716 22094 13756
rect 22557 13753 22569 13787
rect 22603 13753 22615 13787
rect 22557 13747 22615 13753
rect 22646 13716 22652 13728
rect 22066 13688 22652 13716
rect 22646 13676 22652 13688
rect 22704 13676 22710 13728
rect 22830 13716 22836 13728
rect 22791 13688 22836 13716
rect 22830 13676 22836 13688
rect 22888 13676 22894 13728
rect 1104 13626 23460 13648
rect 1104 13574 3749 13626
rect 3801 13574 3813 13626
rect 3865 13574 3877 13626
rect 3929 13574 3941 13626
rect 3993 13574 4005 13626
rect 4057 13574 9347 13626
rect 9399 13574 9411 13626
rect 9463 13574 9475 13626
rect 9527 13574 9539 13626
rect 9591 13574 9603 13626
rect 9655 13574 14945 13626
rect 14997 13574 15009 13626
rect 15061 13574 15073 13626
rect 15125 13574 15137 13626
rect 15189 13574 15201 13626
rect 15253 13574 20543 13626
rect 20595 13574 20607 13626
rect 20659 13574 20671 13626
rect 20723 13574 20735 13626
rect 20787 13574 20799 13626
rect 20851 13574 23460 13626
rect 1104 13552 23460 13574
rect 1670 13472 1676 13524
rect 1728 13512 1734 13524
rect 1857 13515 1915 13521
rect 1857 13512 1869 13515
rect 1728 13484 1869 13512
rect 1728 13472 1734 13484
rect 1857 13481 1869 13484
rect 1903 13481 1915 13515
rect 1857 13475 1915 13481
rect 2222 13472 2228 13524
rect 2280 13512 2286 13524
rect 2593 13515 2651 13521
rect 2593 13512 2605 13515
rect 2280 13484 2605 13512
rect 2280 13472 2286 13484
rect 2593 13481 2605 13484
rect 2639 13481 2651 13515
rect 6270 13512 6276 13524
rect 6231 13484 6276 13512
rect 2593 13475 2651 13481
rect 6270 13472 6276 13484
rect 6328 13472 6334 13524
rect 7834 13512 7840 13524
rect 6380 13484 7840 13512
rect 3234 13404 3240 13456
rect 3292 13444 3298 13456
rect 4890 13444 4896 13456
rect 3292 13416 4896 13444
rect 3292 13404 3298 13416
rect 4890 13404 4896 13416
rect 4948 13404 4954 13456
rect 5994 13404 6000 13456
rect 6052 13444 6058 13456
rect 6380 13453 6408 13484
rect 7834 13472 7840 13484
rect 7892 13472 7898 13524
rect 9674 13472 9680 13524
rect 9732 13512 9738 13524
rect 10505 13515 10563 13521
rect 10505 13512 10517 13515
rect 9732 13484 10517 13512
rect 9732 13472 9738 13484
rect 10505 13481 10517 13484
rect 10551 13481 10563 13515
rect 10505 13475 10563 13481
rect 10962 13472 10968 13524
rect 11020 13512 11026 13524
rect 11977 13515 12035 13521
rect 11977 13512 11989 13515
rect 11020 13484 11989 13512
rect 11020 13472 11026 13484
rect 6365 13447 6423 13453
rect 6365 13444 6377 13447
rect 6052 13416 6377 13444
rect 6052 13404 6058 13416
rect 6365 13413 6377 13416
rect 6411 13413 6423 13447
rect 6365 13407 6423 13413
rect 3142 13376 3148 13388
rect 3103 13348 3148 13376
rect 3142 13336 3148 13348
rect 3200 13336 3206 13388
rect 11900 13385 11928 13484
rect 11977 13481 11989 13484
rect 12023 13512 12035 13515
rect 12161 13515 12219 13521
rect 12161 13512 12173 13515
rect 12023 13484 12173 13512
rect 12023 13481 12035 13484
rect 11977 13475 12035 13481
rect 12161 13481 12173 13484
rect 12207 13481 12219 13515
rect 12161 13475 12219 13481
rect 19150 13472 19156 13524
rect 19208 13512 19214 13524
rect 19245 13515 19303 13521
rect 19245 13512 19257 13515
rect 19208 13484 19257 13512
rect 19208 13472 19214 13484
rect 19245 13481 19257 13484
rect 19291 13481 19303 13515
rect 20898 13512 20904 13524
rect 19245 13475 19303 13481
rect 19352 13484 20904 13512
rect 14090 13444 14096 13456
rect 14051 13416 14096 13444
rect 14090 13404 14096 13416
rect 14148 13404 14154 13456
rect 18138 13404 18144 13456
rect 18196 13444 18202 13456
rect 18417 13447 18475 13453
rect 18417 13444 18429 13447
rect 18196 13416 18429 13444
rect 18196 13404 18202 13416
rect 18417 13413 18429 13416
rect 18463 13444 18475 13447
rect 19352 13444 19380 13484
rect 20898 13472 20904 13484
rect 20956 13472 20962 13524
rect 21542 13512 21548 13524
rect 21503 13484 21548 13512
rect 21542 13472 21548 13484
rect 21600 13472 21606 13524
rect 22278 13472 22284 13524
rect 22336 13512 22342 13524
rect 22465 13515 22523 13521
rect 22465 13512 22477 13515
rect 22336 13484 22477 13512
rect 22336 13472 22342 13484
rect 22465 13481 22477 13484
rect 22511 13481 22523 13515
rect 22465 13475 22523 13481
rect 22833 13515 22891 13521
rect 22833 13481 22845 13515
rect 22879 13512 22891 13515
rect 22922 13512 22928 13524
rect 22879 13484 22928 13512
rect 22879 13481 22891 13484
rect 22833 13475 22891 13481
rect 22922 13472 22928 13484
rect 22980 13472 22986 13524
rect 21560 13444 21588 13472
rect 22554 13444 22560 13456
rect 18463 13416 19380 13444
rect 20640 13416 21588 13444
rect 22480 13416 22560 13444
rect 18463 13413 18475 13416
rect 18417 13407 18475 13413
rect 11885 13379 11943 13385
rect 11885 13345 11897 13379
rect 11931 13345 11943 13379
rect 18598 13376 18604 13388
rect 18511 13348 18604 13376
rect 11885 13339 11943 13345
rect 18598 13336 18604 13348
rect 18656 13376 18662 13388
rect 18693 13379 18751 13385
rect 18693 13376 18705 13379
rect 18656 13348 18705 13376
rect 18656 13336 18662 13348
rect 18693 13345 18705 13348
rect 18739 13376 18751 13379
rect 19242 13376 19248 13388
rect 18739 13348 19248 13376
rect 18739 13345 18751 13348
rect 18693 13339 18751 13345
rect 19242 13336 19248 13348
rect 19300 13336 19306 13388
rect 20640 13385 20668 13416
rect 20625 13379 20683 13385
rect 20625 13345 20637 13379
rect 20671 13345 20683 13379
rect 20625 13339 20683 13345
rect 20901 13379 20959 13385
rect 20901 13345 20913 13379
rect 20947 13376 20959 13379
rect 21082 13376 21088 13388
rect 20947 13348 21088 13376
rect 20947 13345 20959 13348
rect 20901 13339 20959 13345
rect 21082 13336 21088 13348
rect 21140 13336 21146 13388
rect 21913 13379 21971 13385
rect 21913 13345 21925 13379
rect 21959 13376 21971 13379
rect 22186 13376 22192 13388
rect 21959 13348 22192 13376
rect 21959 13345 21971 13348
rect 21913 13339 21971 13345
rect 22186 13336 22192 13348
rect 22244 13336 22250 13388
rect 2041 13311 2099 13317
rect 2041 13277 2053 13311
rect 2087 13308 2099 13311
rect 2958 13308 2964 13320
rect 2087 13280 2176 13308
rect 2919 13280 2964 13308
rect 2087 13277 2099 13280
rect 2041 13271 2099 13277
rect 2148 13184 2176 13280
rect 2958 13268 2964 13280
rect 3016 13268 3022 13320
rect 4706 13308 4712 13320
rect 4667 13280 4712 13308
rect 4706 13268 4712 13280
rect 4764 13268 4770 13320
rect 5166 13317 5172 13320
rect 4893 13311 4951 13317
rect 4893 13277 4905 13311
rect 4939 13277 4951 13311
rect 4893 13271 4951 13277
rect 5160 13271 5172 13317
rect 5224 13308 5230 13320
rect 7745 13311 7803 13317
rect 5224 13280 5260 13308
rect 2682 13200 2688 13252
rect 2740 13240 2746 13252
rect 3418 13240 3424 13252
rect 2740 13212 3424 13240
rect 2740 13200 2746 13212
rect 3418 13200 3424 13212
rect 3476 13200 3482 13252
rect 2130 13172 2136 13184
rect 2091 13144 2136 13172
rect 2130 13132 2136 13144
rect 2188 13132 2194 13184
rect 3050 13132 3056 13184
rect 3108 13172 3114 13184
rect 4617 13175 4675 13181
rect 3108 13144 3153 13172
rect 3108 13132 3114 13144
rect 4617 13141 4629 13175
rect 4663 13172 4675 13175
rect 4798 13172 4804 13184
rect 4663 13144 4804 13172
rect 4663 13141 4675 13144
rect 4617 13135 4675 13141
rect 4798 13132 4804 13144
rect 4856 13132 4862 13184
rect 4908 13172 4936 13271
rect 5166 13268 5172 13271
rect 5224 13268 5230 13280
rect 7745 13277 7757 13311
rect 7791 13308 7803 13311
rect 8941 13311 8999 13317
rect 8941 13308 8953 13311
rect 7791 13280 8953 13308
rect 7791 13277 7803 13280
rect 7745 13271 7803 13277
rect 8941 13277 8953 13280
rect 8987 13277 8999 13311
rect 8941 13271 8999 13277
rect 15473 13311 15531 13317
rect 15473 13277 15485 13311
rect 15519 13308 15531 13311
rect 15565 13311 15623 13317
rect 15565 13308 15577 13311
rect 15519 13280 15577 13308
rect 15519 13277 15531 13280
rect 15473 13271 15531 13277
rect 15565 13277 15577 13280
rect 15611 13308 15623 13311
rect 17034 13308 17040 13320
rect 15611 13280 17040 13308
rect 15611 13277 15623 13280
rect 15565 13271 15623 13277
rect 6086 13200 6092 13252
rect 6144 13240 6150 13252
rect 7478 13243 7536 13249
rect 7478 13240 7490 13243
rect 6144 13212 7490 13240
rect 6144 13200 6150 13212
rect 7478 13209 7490 13212
rect 7524 13209 7536 13243
rect 7478 13203 7536 13209
rect 6178 13172 6184 13184
rect 4908 13144 6184 13172
rect 6178 13132 6184 13144
rect 6236 13172 6242 13184
rect 7760 13172 7788 13271
rect 17034 13268 17040 13280
rect 17092 13268 17098 13320
rect 18506 13268 18512 13320
rect 18564 13308 18570 13320
rect 18877 13311 18935 13317
rect 18877 13308 18889 13311
rect 18564 13280 18889 13308
rect 18564 13268 18570 13280
rect 18877 13277 18889 13280
rect 18923 13277 18935 13311
rect 18877 13271 18935 13277
rect 20369 13311 20427 13317
rect 20369 13277 20381 13311
rect 20415 13308 20427 13311
rect 20990 13308 20996 13320
rect 20415 13280 20996 13308
rect 20415 13277 20427 13280
rect 20369 13271 20427 13277
rect 20990 13268 20996 13280
rect 21048 13268 21054 13320
rect 21266 13268 21272 13320
rect 21324 13308 21330 13320
rect 22097 13311 22155 13317
rect 22097 13308 22109 13311
rect 21324 13280 22109 13308
rect 21324 13268 21330 13280
rect 22097 13277 22109 13280
rect 22143 13277 22155 13311
rect 22097 13271 22155 13277
rect 22480 13284 22508 13416
rect 22554 13404 22560 13416
rect 22612 13404 22618 13456
rect 22646 13336 22652 13388
rect 22704 13376 22710 13388
rect 22704 13348 23060 13376
rect 22704 13336 22710 13348
rect 23032 13317 23060 13348
rect 23017 13311 23075 13317
rect 22557 13287 22615 13293
rect 22557 13284 22569 13287
rect 22480 13256 22569 13284
rect 22557 13253 22569 13256
rect 22603 13253 22615 13287
rect 23017 13277 23029 13311
rect 23063 13277 23075 13311
rect 23017 13271 23075 13277
rect 8478 13200 8484 13252
rect 8536 13240 8542 13252
rect 9186 13243 9244 13249
rect 9186 13240 9198 13243
rect 8536 13212 9198 13240
rect 8536 13200 8542 13212
rect 9186 13209 9198 13212
rect 9232 13209 9244 13243
rect 9186 13203 9244 13209
rect 11514 13200 11520 13252
rect 11572 13240 11578 13252
rect 11618 13243 11676 13249
rect 11618 13240 11630 13243
rect 11572 13212 11630 13240
rect 11572 13200 11578 13212
rect 11618 13209 11630 13212
rect 11664 13209 11676 13243
rect 11618 13203 11676 13209
rect 15228 13243 15286 13249
rect 15228 13209 15240 13243
rect 15274 13240 15286 13243
rect 15654 13240 15660 13252
rect 15274 13212 15660 13240
rect 15274 13209 15286 13212
rect 15228 13203 15286 13209
rect 15654 13200 15660 13212
rect 15712 13200 15718 13252
rect 15832 13243 15890 13249
rect 15832 13209 15844 13243
rect 15878 13240 15890 13243
rect 16114 13240 16120 13252
rect 15878 13212 16120 13240
rect 15878 13209 15890 13212
rect 15832 13203 15890 13209
rect 16114 13200 16120 13212
rect 16172 13200 16178 13252
rect 17304 13243 17362 13249
rect 17304 13240 17316 13243
rect 16960 13212 17316 13240
rect 7837 13175 7895 13181
rect 7837 13172 7849 13175
rect 6236 13144 7849 13172
rect 6236 13132 6242 13144
rect 7837 13141 7849 13144
rect 7883 13141 7895 13175
rect 10318 13172 10324 13184
rect 10279 13144 10324 13172
rect 7837 13135 7895 13141
rect 10318 13132 10324 13144
rect 10376 13132 10382 13184
rect 16960 13181 16988 13212
rect 17304 13209 17316 13212
rect 17350 13240 17362 13243
rect 19610 13240 19616 13252
rect 17350 13212 19616 13240
rect 17350 13209 17362 13212
rect 17304 13203 17362 13209
rect 19610 13200 19616 13212
rect 19668 13200 19674 13252
rect 21085 13243 21143 13249
rect 21085 13240 21097 13243
rect 19720 13212 21097 13240
rect 16945 13175 17003 13181
rect 16945 13141 16957 13175
rect 16991 13141 17003 13175
rect 19058 13172 19064 13184
rect 19019 13144 19064 13172
rect 16945 13135 17003 13141
rect 19058 13132 19064 13144
rect 19116 13132 19122 13184
rect 19242 13132 19248 13184
rect 19300 13172 19306 13184
rect 19720 13172 19748 13212
rect 21085 13209 21097 13212
rect 21131 13209 21143 13243
rect 22186 13240 22192 13252
rect 21085 13203 21143 13209
rect 21468 13212 22192 13240
rect 19300 13144 19748 13172
rect 19300 13132 19306 13144
rect 20714 13132 20720 13184
rect 20772 13172 20778 13184
rect 21468 13181 21496 13212
rect 22186 13200 22192 13212
rect 22244 13200 22250 13252
rect 22557 13247 22615 13253
rect 20993 13175 21051 13181
rect 20993 13172 21005 13175
rect 20772 13144 21005 13172
rect 20772 13132 20778 13144
rect 20993 13141 21005 13144
rect 21039 13141 21051 13175
rect 20993 13135 21051 13141
rect 21453 13175 21511 13181
rect 21453 13141 21465 13175
rect 21499 13141 21511 13175
rect 22002 13172 22008 13184
rect 21963 13144 22008 13172
rect 21453 13135 21511 13141
rect 22002 13132 22008 13144
rect 22060 13132 22066 13184
rect 22646 13132 22652 13184
rect 22704 13172 22710 13184
rect 22741 13175 22799 13181
rect 22741 13172 22753 13175
rect 22704 13144 22753 13172
rect 22704 13132 22710 13144
rect 22741 13141 22753 13144
rect 22787 13141 22799 13175
rect 22741 13135 22799 13141
rect 1104 13082 23460 13104
rect 1104 13030 6548 13082
rect 6600 13030 6612 13082
rect 6664 13030 6676 13082
rect 6728 13030 6740 13082
rect 6792 13030 6804 13082
rect 6856 13030 12146 13082
rect 12198 13030 12210 13082
rect 12262 13030 12274 13082
rect 12326 13030 12338 13082
rect 12390 13030 12402 13082
rect 12454 13030 17744 13082
rect 17796 13030 17808 13082
rect 17860 13030 17872 13082
rect 17924 13030 17936 13082
rect 17988 13030 18000 13082
rect 18052 13030 23460 13082
rect 1104 13008 23460 13030
rect 2222 12928 2228 12980
rect 2280 12968 2286 12980
rect 2501 12971 2559 12977
rect 2501 12968 2513 12971
rect 2280 12940 2513 12968
rect 2280 12928 2286 12940
rect 2501 12937 2513 12940
rect 2547 12937 2559 12971
rect 2501 12931 2559 12937
rect 3789 12971 3847 12977
rect 3789 12937 3801 12971
rect 3835 12968 3847 12971
rect 4157 12971 4215 12977
rect 4157 12968 4169 12971
rect 3835 12940 4169 12968
rect 3835 12937 3847 12940
rect 3789 12931 3847 12937
rect 4157 12937 4169 12940
rect 4203 12937 4215 12971
rect 4157 12931 4215 12937
rect 6178 12928 6184 12980
rect 6236 12968 6242 12980
rect 6362 12968 6368 12980
rect 6236 12940 6368 12968
rect 6236 12928 6242 12940
rect 6362 12928 6368 12940
rect 6420 12928 6426 12980
rect 8386 12968 8392 12980
rect 8347 12940 8392 12968
rect 8386 12928 8392 12940
rect 8444 12928 8450 12980
rect 13078 12968 13084 12980
rect 13039 12940 13084 12968
rect 13078 12928 13084 12940
rect 13136 12928 13142 12980
rect 16206 12928 16212 12980
rect 16264 12968 16270 12980
rect 16301 12971 16359 12977
rect 16301 12968 16313 12971
rect 16264 12940 16313 12968
rect 16264 12928 16270 12940
rect 16301 12937 16313 12940
rect 16347 12968 16359 12971
rect 16485 12971 16543 12977
rect 16485 12968 16497 12971
rect 16347 12940 16497 12968
rect 16347 12937 16359 12940
rect 16301 12931 16359 12937
rect 16485 12937 16497 12940
rect 16531 12968 16543 12971
rect 17034 12968 17040 12980
rect 16531 12940 17040 12968
rect 16531 12937 16543 12940
rect 16485 12931 16543 12937
rect 17034 12928 17040 12940
rect 17092 12928 17098 12980
rect 18233 12971 18291 12977
rect 18233 12937 18245 12971
rect 18279 12968 18291 12971
rect 18598 12968 18604 12980
rect 18279 12940 18604 12968
rect 18279 12937 18291 12940
rect 18233 12931 18291 12937
rect 3602 12860 3608 12912
rect 3660 12900 3666 12912
rect 5169 12903 5227 12909
rect 5169 12900 5181 12903
rect 3660 12872 5181 12900
rect 3660 12860 3666 12872
rect 5169 12869 5181 12872
rect 5215 12869 5227 12903
rect 5169 12863 5227 12869
rect 6270 12860 6276 12912
rect 6328 12900 6334 12912
rect 7254 12903 7312 12909
rect 7254 12900 7266 12903
rect 6328 12872 7266 12900
rect 6328 12860 6334 12872
rect 7254 12869 7266 12872
rect 7300 12869 7312 12903
rect 7254 12863 7312 12869
rect 9858 12860 9864 12912
rect 9916 12900 9922 12912
rect 9916 12872 11376 12900
rect 9916 12860 9922 12872
rect 2866 12832 2872 12844
rect 2827 12804 2872 12832
rect 2866 12792 2872 12804
rect 2924 12792 2930 12844
rect 3697 12835 3755 12841
rect 3697 12801 3709 12835
rect 3743 12832 3755 12835
rect 4246 12832 4252 12844
rect 3743 12804 4252 12832
rect 3743 12801 3755 12804
rect 3697 12795 3755 12801
rect 4246 12792 4252 12804
rect 4304 12792 4310 12844
rect 4525 12835 4583 12841
rect 4525 12801 4537 12835
rect 4571 12801 4583 12835
rect 4525 12795 4583 12801
rect 4617 12835 4675 12841
rect 4617 12801 4629 12835
rect 4663 12832 4675 12835
rect 4663 12804 5120 12832
rect 4663 12801 4675 12804
rect 4617 12795 4675 12801
rect 2958 12764 2964 12776
rect 2919 12736 2964 12764
rect 2958 12724 2964 12736
rect 3016 12724 3022 12776
rect 3145 12767 3203 12773
rect 3145 12733 3157 12767
rect 3191 12764 3203 12767
rect 3234 12764 3240 12776
rect 3191 12736 3240 12764
rect 3191 12733 3203 12736
rect 3145 12727 3203 12733
rect 2682 12656 2688 12708
rect 2740 12696 2746 12708
rect 3160 12696 3188 12727
rect 3234 12724 3240 12736
rect 3292 12724 3298 12776
rect 3418 12724 3424 12776
rect 3476 12764 3482 12776
rect 3881 12767 3939 12773
rect 3881 12764 3893 12767
rect 3476 12736 3893 12764
rect 3476 12724 3482 12736
rect 3881 12733 3893 12736
rect 3927 12733 3939 12767
rect 4540 12764 4568 12795
rect 4798 12764 4804 12776
rect 3881 12727 3939 12733
rect 4448 12736 4568 12764
rect 4759 12736 4804 12764
rect 2740 12668 3188 12696
rect 2740 12656 2746 12668
rect 2774 12588 2780 12640
rect 2832 12628 2838 12640
rect 3329 12631 3387 12637
rect 3329 12628 3341 12631
rect 2832 12600 3341 12628
rect 2832 12588 2838 12600
rect 3329 12597 3341 12600
rect 3375 12597 3387 12631
rect 4448 12628 4476 12736
rect 4798 12724 4804 12736
rect 4856 12724 4862 12776
rect 5092 12764 5120 12804
rect 6362 12792 6368 12844
rect 6420 12832 6426 12844
rect 7009 12835 7067 12841
rect 7009 12832 7021 12835
rect 6420 12804 7021 12832
rect 6420 12792 6426 12804
rect 7009 12801 7021 12804
rect 7055 12801 7067 12835
rect 9594 12835 9652 12841
rect 9594 12832 9606 12835
rect 7009 12795 7067 12801
rect 7116 12804 9606 12832
rect 7116 12764 7144 12804
rect 9594 12801 9606 12804
rect 9640 12832 9652 12835
rect 10318 12832 10324 12844
rect 9640 12804 10324 12832
rect 9640 12801 9652 12804
rect 9594 12795 9652 12801
rect 10318 12792 10324 12804
rect 10376 12792 10382 12844
rect 11054 12832 11060 12844
rect 11112 12841 11118 12844
rect 11348 12841 11376 12872
rect 11112 12835 11135 12841
rect 10987 12804 11060 12832
rect 11054 12792 11060 12804
rect 11123 12832 11135 12835
rect 11333 12835 11391 12841
rect 11123 12804 11284 12832
rect 11123 12801 11135 12804
rect 11112 12795 11135 12801
rect 11112 12792 11118 12795
rect 9858 12764 9864 12776
rect 5092 12736 7144 12764
rect 9819 12736 9864 12764
rect 9858 12724 9864 12736
rect 9916 12724 9922 12776
rect 11256 12764 11284 12804
rect 11333 12801 11345 12835
rect 11379 12801 11391 12835
rect 11333 12795 11391 12801
rect 12733 12835 12791 12841
rect 12733 12801 12745 12835
rect 12779 12832 12791 12835
rect 12894 12832 12900 12844
rect 12779 12804 12900 12832
rect 12779 12801 12791 12804
rect 12733 12795 12791 12801
rect 12894 12792 12900 12804
rect 12952 12792 12958 12844
rect 12989 12835 13047 12841
rect 12989 12801 13001 12835
rect 13035 12832 13047 12835
rect 13096 12832 13124 12928
rect 16224 12900 16252 12928
rect 14752 12872 16252 12900
rect 17804 12903 17862 12909
rect 13265 12835 13323 12841
rect 13265 12832 13277 12835
rect 13035 12804 13277 12832
rect 13035 12801 13047 12804
rect 12989 12795 13047 12801
rect 13265 12801 13277 12804
rect 13311 12801 13323 12835
rect 13265 12795 13323 12801
rect 13532 12835 13590 12841
rect 13532 12801 13544 12835
rect 13578 12832 13590 12835
rect 13906 12832 13912 12844
rect 13578 12804 13912 12832
rect 13578 12801 13590 12804
rect 13532 12795 13590 12801
rect 13906 12792 13912 12804
rect 13964 12792 13970 12844
rect 14752 12841 14780 12872
rect 17804 12869 17816 12903
rect 17850 12900 17862 12903
rect 18138 12900 18144 12912
rect 17850 12872 18144 12900
rect 17850 12869 17862 12872
rect 17804 12863 17862 12869
rect 18138 12860 18144 12872
rect 18196 12860 18202 12912
rect 14737 12835 14795 12841
rect 14737 12801 14749 12835
rect 14783 12801 14795 12835
rect 15004 12835 15062 12841
rect 15004 12832 15016 12835
rect 14737 12795 14795 12801
rect 14844 12804 15016 12832
rect 14844 12764 14872 12804
rect 15004 12801 15016 12804
rect 15050 12832 15062 12835
rect 16574 12832 16580 12844
rect 15050 12804 16580 12832
rect 15050 12801 15062 12804
rect 15004 12795 15062 12801
rect 16574 12792 16580 12804
rect 16632 12792 16638 12844
rect 18049 12835 18107 12841
rect 18049 12801 18061 12835
rect 18095 12832 18107 12835
rect 18248 12832 18276 12931
rect 18598 12928 18604 12940
rect 18656 12928 18662 12980
rect 20990 12928 20996 12980
rect 21048 12968 21054 12980
rect 21177 12971 21235 12977
rect 21177 12968 21189 12971
rect 21048 12940 21189 12968
rect 21048 12928 21054 12940
rect 21177 12937 21189 12940
rect 21223 12937 21235 12971
rect 21177 12931 21235 12937
rect 22094 12928 22100 12980
rect 22152 12968 22158 12980
rect 22152 12940 22197 12968
rect 22152 12928 22158 12940
rect 22370 12928 22376 12980
rect 22428 12968 22434 12980
rect 22557 12971 22615 12977
rect 22557 12968 22569 12971
rect 22428 12940 22569 12968
rect 22428 12928 22434 12940
rect 22557 12937 22569 12940
rect 22603 12937 22615 12971
rect 23106 12968 23112 12980
rect 23067 12940 23112 12968
rect 22557 12931 22615 12937
rect 23106 12928 23112 12940
rect 23164 12928 23170 12980
rect 18616 12900 18644 12928
rect 19150 12900 19156 12912
rect 18616 12872 19156 12900
rect 19150 12860 19156 12872
rect 19208 12900 19214 12912
rect 19208 12872 19334 12900
rect 19208 12860 19214 12872
rect 18325 12835 18383 12841
rect 18325 12832 18337 12835
rect 18095 12804 18337 12832
rect 18095 12801 18107 12804
rect 18049 12795 18107 12801
rect 18325 12801 18337 12804
rect 18371 12832 18383 12835
rect 18414 12832 18420 12844
rect 18371 12804 18420 12832
rect 18371 12801 18383 12804
rect 18325 12795 18383 12801
rect 18414 12792 18420 12804
rect 18472 12792 18478 12844
rect 18592 12835 18650 12841
rect 18592 12801 18604 12835
rect 18638 12832 18650 12835
rect 18874 12832 18880 12844
rect 18638 12804 18880 12832
rect 18638 12801 18650 12804
rect 18592 12795 18650 12801
rect 18874 12792 18880 12804
rect 18932 12792 18938 12844
rect 19306 12832 19334 12872
rect 20254 12860 20260 12912
rect 20312 12900 20318 12912
rect 20312 12872 20576 12900
rect 20312 12860 20318 12872
rect 19797 12835 19855 12841
rect 19797 12832 19809 12835
rect 19306 12804 19809 12832
rect 19797 12801 19809 12804
rect 19843 12801 19855 12835
rect 19797 12795 19855 12801
rect 20064 12835 20122 12841
rect 20064 12801 20076 12835
rect 20110 12832 20122 12835
rect 20438 12832 20444 12844
rect 20110 12804 20444 12832
rect 20110 12801 20122 12804
rect 20064 12795 20122 12801
rect 20438 12792 20444 12804
rect 20496 12792 20502 12844
rect 20548 12832 20576 12872
rect 21082 12860 21088 12912
rect 21140 12900 21146 12912
rect 21453 12903 21511 12909
rect 21453 12900 21465 12903
rect 21140 12872 21465 12900
rect 21140 12860 21146 12872
rect 21453 12869 21465 12872
rect 21499 12869 21511 12903
rect 23198 12900 23204 12912
rect 21453 12863 21511 12869
rect 22066 12872 23204 12900
rect 22066 12832 22094 12872
rect 22848 12841 22876 12872
rect 23198 12860 23204 12872
rect 23256 12860 23262 12912
rect 20548 12804 22094 12832
rect 22189 12835 22247 12841
rect 22189 12801 22201 12835
rect 22235 12832 22247 12835
rect 22833 12835 22891 12841
rect 22235 12804 22508 12832
rect 22235 12801 22247 12804
rect 22189 12795 22247 12801
rect 22480 12776 22508 12804
rect 22833 12801 22845 12835
rect 22879 12801 22891 12835
rect 22833 12795 22891 12801
rect 22925 12835 22983 12841
rect 22925 12801 22937 12835
rect 22971 12832 22983 12835
rect 23474 12832 23480 12844
rect 22971 12804 23480 12832
rect 22971 12801 22983 12804
rect 22925 12795 22983 12801
rect 23474 12792 23480 12804
rect 23532 12792 23538 12844
rect 11256 12736 11652 12764
rect 4522 12656 4528 12708
rect 4580 12696 4586 12708
rect 4985 12699 5043 12705
rect 4985 12696 4997 12699
rect 4580 12668 4997 12696
rect 4580 12656 4586 12668
rect 4985 12665 4997 12668
rect 5031 12665 5043 12699
rect 8478 12696 8484 12708
rect 4985 12659 5043 12665
rect 7944 12668 8484 12696
rect 7944 12628 7972 12668
rect 8478 12656 8484 12668
rect 8536 12656 8542 12708
rect 11624 12705 11652 12736
rect 14660 12736 14872 12764
rect 21269 12767 21327 12773
rect 14660 12705 14688 12736
rect 21269 12733 21281 12767
rect 21315 12764 21327 12767
rect 21634 12764 21640 12776
rect 21315 12736 21640 12764
rect 21315 12733 21327 12736
rect 21269 12727 21327 12733
rect 21634 12724 21640 12736
rect 21692 12764 21698 12776
rect 21913 12767 21971 12773
rect 21913 12764 21925 12767
rect 21692 12736 21925 12764
rect 21692 12724 21698 12736
rect 21913 12733 21925 12736
rect 21959 12733 21971 12767
rect 21913 12727 21971 12733
rect 22462 12724 22468 12776
rect 22520 12724 22526 12776
rect 23198 12724 23204 12776
rect 23256 12764 23262 12776
rect 23382 12764 23388 12776
rect 23256 12736 23388 12764
rect 23256 12724 23262 12736
rect 23382 12724 23388 12736
rect 23440 12724 23446 12776
rect 11609 12699 11667 12705
rect 11609 12665 11621 12699
rect 11655 12665 11667 12699
rect 11609 12659 11667 12665
rect 14645 12699 14703 12705
rect 14645 12665 14657 12699
rect 14691 12665 14703 12699
rect 16114 12696 16120 12708
rect 16027 12668 16120 12696
rect 14645 12659 14703 12665
rect 16114 12656 16120 12668
rect 16172 12696 16178 12708
rect 16172 12668 17172 12696
rect 16172 12656 16178 12668
rect 4448 12600 7972 12628
rect 3329 12591 3387 12597
rect 9674 12588 9680 12640
rect 9732 12628 9738 12640
rect 9953 12631 10011 12637
rect 9953 12628 9965 12631
rect 9732 12600 9965 12628
rect 9732 12588 9738 12600
rect 9953 12597 9965 12600
rect 9999 12597 10011 12631
rect 9953 12591 10011 12597
rect 16574 12588 16580 12640
rect 16632 12628 16638 12640
rect 16669 12631 16727 12637
rect 16669 12628 16681 12631
rect 16632 12600 16681 12628
rect 16632 12588 16638 12600
rect 16669 12597 16681 12600
rect 16715 12597 16727 12631
rect 17144 12628 17172 12668
rect 19242 12628 19248 12640
rect 17144 12600 19248 12628
rect 16669 12591 16727 12597
rect 19242 12588 19248 12600
rect 19300 12588 19306 12640
rect 19705 12631 19763 12637
rect 19705 12597 19717 12631
rect 19751 12628 19763 12631
rect 21082 12628 21088 12640
rect 19751 12600 21088 12628
rect 19751 12597 19763 12600
rect 19705 12591 19763 12597
rect 21082 12588 21088 12600
rect 21140 12588 21146 12640
rect 22094 12588 22100 12640
rect 22152 12628 22158 12640
rect 22649 12631 22707 12637
rect 22649 12628 22661 12631
rect 22152 12600 22661 12628
rect 22152 12588 22158 12600
rect 22649 12597 22661 12600
rect 22695 12597 22707 12631
rect 22649 12591 22707 12597
rect 1104 12538 23460 12560
rect 1104 12486 3749 12538
rect 3801 12486 3813 12538
rect 3865 12486 3877 12538
rect 3929 12486 3941 12538
rect 3993 12486 4005 12538
rect 4057 12486 9347 12538
rect 9399 12486 9411 12538
rect 9463 12486 9475 12538
rect 9527 12486 9539 12538
rect 9591 12486 9603 12538
rect 9655 12486 14945 12538
rect 14997 12486 15009 12538
rect 15061 12486 15073 12538
rect 15125 12486 15137 12538
rect 15189 12486 15201 12538
rect 15253 12486 20543 12538
rect 20595 12486 20607 12538
rect 20659 12486 20671 12538
rect 20723 12486 20735 12538
rect 20787 12486 20799 12538
rect 20851 12486 23460 12538
rect 1104 12464 23460 12486
rect 1762 12384 1768 12436
rect 1820 12424 1826 12436
rect 2041 12427 2099 12433
rect 2041 12424 2053 12427
rect 1820 12396 2053 12424
rect 1820 12384 1826 12396
rect 2041 12393 2053 12396
rect 2087 12393 2099 12427
rect 2041 12387 2099 12393
rect 2866 12384 2872 12436
rect 2924 12424 2930 12436
rect 3789 12427 3847 12433
rect 3789 12424 3801 12427
rect 2924 12396 3801 12424
rect 2924 12384 2930 12396
rect 3789 12393 3801 12396
rect 3835 12393 3847 12427
rect 5902 12424 5908 12436
rect 3789 12387 3847 12393
rect 4540 12396 5908 12424
rect 2682 12288 2688 12300
rect 2643 12260 2688 12288
rect 2682 12248 2688 12260
rect 2740 12248 2746 12300
rect 3053 12291 3111 12297
rect 3053 12257 3065 12291
rect 3099 12288 3111 12291
rect 3602 12288 3608 12300
rect 3099 12260 3608 12288
rect 3099 12257 3111 12260
rect 3053 12251 3111 12257
rect 3602 12248 3608 12260
rect 3660 12248 3666 12300
rect 3510 12180 3516 12232
rect 3568 12220 3574 12232
rect 3973 12223 4031 12229
rect 3973 12220 3985 12223
rect 3568 12192 3985 12220
rect 3568 12180 3574 12192
rect 3973 12189 3985 12192
rect 4019 12189 4031 12223
rect 4540 12220 4568 12396
rect 5902 12384 5908 12396
rect 5960 12384 5966 12436
rect 16574 12384 16580 12436
rect 16632 12424 16638 12436
rect 18506 12424 18512 12436
rect 16632 12396 17816 12424
rect 18467 12396 18512 12424
rect 16632 12384 16638 12396
rect 17681 12359 17739 12365
rect 17681 12325 17693 12359
rect 17727 12325 17739 12359
rect 17788 12356 17816 12396
rect 18506 12384 18512 12396
rect 18564 12384 18570 12436
rect 20714 12424 20720 12436
rect 18607 12396 20720 12424
rect 18607 12356 18635 12396
rect 20714 12384 20720 12396
rect 20772 12384 20778 12436
rect 20806 12384 20812 12436
rect 20864 12424 20870 12436
rect 20864 12396 21312 12424
rect 20864 12384 20870 12396
rect 18782 12356 18788 12368
rect 17788 12328 18635 12356
rect 18743 12328 18788 12356
rect 17681 12319 17739 12325
rect 4709 12291 4767 12297
rect 4709 12257 4721 12291
rect 4755 12288 4767 12291
rect 4798 12288 4804 12300
rect 4755 12260 4804 12288
rect 4755 12257 4767 12260
rect 4709 12251 4767 12257
rect 4798 12248 4804 12260
rect 4856 12248 4862 12300
rect 9674 12248 9680 12300
rect 9732 12288 9738 12300
rect 14185 12291 14243 12297
rect 9732 12260 10180 12288
rect 9732 12248 9738 12260
rect 3973 12183 4031 12189
rect 4448 12192 4568 12220
rect 4893 12223 4951 12229
rect 2409 12155 2467 12161
rect 2409 12121 2421 12155
rect 2455 12152 2467 12155
rect 2866 12152 2872 12164
rect 2455 12124 2872 12152
rect 2455 12121 2467 12124
rect 2409 12115 2467 12121
rect 2866 12112 2872 12124
rect 2924 12112 2930 12164
rect 3237 12155 3295 12161
rect 3237 12121 3249 12155
rect 3283 12152 3295 12155
rect 4448 12152 4476 12192
rect 4893 12189 4905 12223
rect 4939 12220 4951 12223
rect 6362 12220 6368 12232
rect 4939 12192 6368 12220
rect 4939 12189 4951 12192
rect 4893 12183 4951 12189
rect 6362 12180 6368 12192
rect 6420 12180 6426 12232
rect 9858 12180 9864 12232
rect 9916 12220 9922 12232
rect 10045 12223 10103 12229
rect 10045 12220 10057 12223
rect 9916 12192 10057 12220
rect 9916 12180 9922 12192
rect 10045 12189 10057 12192
rect 10091 12189 10103 12223
rect 10045 12183 10103 12189
rect 3283 12124 4476 12152
rect 4525 12155 4583 12161
rect 3283 12121 3295 12124
rect 3237 12115 3295 12121
rect 4525 12121 4537 12155
rect 4571 12152 4583 12155
rect 5160 12155 5218 12161
rect 5160 12152 5172 12155
rect 4571 12124 5172 12152
rect 4571 12121 4583 12124
rect 4525 12115 4583 12121
rect 5160 12121 5172 12124
rect 5206 12152 5218 12155
rect 5258 12152 5264 12164
rect 5206 12124 5264 12152
rect 5206 12121 5218 12124
rect 5160 12115 5218 12121
rect 5258 12112 5264 12124
rect 5316 12112 5322 12164
rect 6178 12112 6184 12164
rect 6236 12152 6242 12164
rect 6610 12155 6668 12161
rect 6610 12152 6622 12155
rect 6236 12124 6622 12152
rect 6236 12112 6242 12124
rect 6610 12121 6622 12124
rect 6656 12121 6668 12155
rect 9306 12152 9312 12164
rect 6610 12115 6668 12121
rect 7760 12124 9312 12152
rect 2498 12044 2504 12096
rect 2556 12084 2562 12096
rect 3145 12087 3203 12093
rect 2556 12056 2601 12084
rect 2556 12044 2562 12056
rect 3145 12053 3157 12087
rect 3191 12084 3203 12087
rect 3326 12084 3332 12096
rect 3191 12056 3332 12084
rect 3191 12053 3203 12056
rect 3145 12047 3203 12053
rect 3326 12044 3332 12056
rect 3384 12044 3390 12096
rect 3602 12084 3608 12096
rect 3563 12056 3608 12084
rect 3602 12044 3608 12056
rect 3660 12044 3666 12096
rect 4062 12084 4068 12096
rect 4023 12056 4068 12084
rect 4062 12044 4068 12056
rect 4120 12044 4126 12096
rect 4433 12087 4491 12093
rect 4433 12053 4445 12087
rect 4479 12084 4491 12087
rect 6270 12084 6276 12096
rect 4479 12056 6276 12084
rect 4479 12053 4491 12056
rect 4433 12047 4491 12053
rect 6270 12044 6276 12056
rect 6328 12044 6334 12096
rect 6454 12044 6460 12096
rect 6512 12084 6518 12096
rect 7760 12093 7788 12124
rect 9306 12112 9312 12124
rect 9364 12112 9370 12164
rect 7745 12087 7803 12093
rect 7745 12084 7757 12087
rect 6512 12056 7757 12084
rect 6512 12044 6518 12056
rect 7745 12053 7757 12056
rect 7791 12053 7803 12087
rect 7745 12047 7803 12053
rect 7834 12044 7840 12096
rect 7892 12084 7898 12096
rect 8481 12087 8539 12093
rect 8481 12084 8493 12087
rect 7892 12056 8493 12084
rect 7892 12044 7898 12056
rect 8481 12053 8493 12056
rect 8527 12084 8539 12087
rect 9217 12087 9275 12093
rect 9217 12084 9229 12087
rect 8527 12056 9229 12084
rect 8527 12053 8539 12056
rect 8481 12047 8539 12053
rect 9217 12053 9229 12056
rect 9263 12084 9275 12087
rect 9861 12087 9919 12093
rect 9861 12084 9873 12087
rect 9263 12056 9873 12084
rect 9263 12053 9275 12056
rect 9217 12047 9275 12053
rect 9861 12053 9873 12056
rect 9907 12084 9919 12087
rect 10060 12084 10088 12183
rect 10152 12152 10180 12260
rect 14185 12257 14197 12291
rect 14231 12288 14243 12291
rect 14829 12291 14887 12297
rect 14829 12288 14841 12291
rect 14231 12260 14841 12288
rect 14231 12257 14243 12260
rect 14185 12251 14243 12257
rect 14829 12257 14841 12260
rect 14875 12288 14887 12291
rect 16206 12288 16212 12300
rect 14875 12260 16212 12288
rect 14875 12257 14887 12260
rect 14829 12251 14887 12257
rect 12529 12223 12587 12229
rect 12529 12220 12541 12223
rect 12406 12192 12541 12220
rect 10318 12161 10324 12164
rect 10312 12152 10324 12161
rect 10152 12124 10324 12152
rect 10312 12115 10324 12124
rect 10318 12112 10324 12115
rect 10376 12112 10382 12164
rect 11517 12155 11575 12161
rect 11517 12152 11529 12155
rect 10428 12124 11529 12152
rect 10428 12084 10456 12124
rect 11517 12121 11529 12124
rect 11563 12152 11575 12155
rect 11701 12155 11759 12161
rect 11701 12152 11713 12155
rect 11563 12124 11713 12152
rect 11563 12121 11575 12124
rect 11517 12115 11575 12121
rect 11701 12121 11713 12124
rect 11747 12152 11759 12155
rect 12406 12152 12434 12192
rect 12529 12189 12541 12192
rect 12575 12220 12587 12223
rect 13078 12220 13084 12232
rect 12575 12192 13084 12220
rect 12575 12189 12587 12192
rect 12529 12183 12587 12189
rect 13078 12180 13084 12192
rect 13136 12220 13142 12232
rect 14200 12220 14228 12251
rect 16206 12248 16212 12260
rect 16264 12288 16270 12300
rect 16301 12291 16359 12297
rect 16301 12288 16313 12291
rect 16264 12260 16313 12288
rect 16264 12248 16270 12260
rect 16301 12257 16313 12260
rect 16347 12257 16359 12291
rect 17696 12288 17724 12319
rect 18782 12316 18788 12328
rect 18840 12316 18846 12368
rect 19058 12356 19064 12368
rect 19019 12328 19064 12356
rect 19058 12316 19064 12328
rect 19116 12316 19122 12368
rect 20732 12328 21220 12356
rect 17696 12260 19104 12288
rect 16301 12251 16359 12257
rect 16574 12229 16580 12232
rect 16568 12220 16580 12229
rect 13136 12192 14228 12220
rect 16535 12192 16580 12220
rect 13136 12180 13142 12192
rect 16568 12183 16580 12192
rect 16574 12180 16580 12183
rect 16632 12180 16638 12232
rect 18325 12223 18383 12229
rect 18325 12189 18337 12223
rect 18371 12220 18383 12223
rect 18601 12223 18659 12229
rect 18601 12220 18613 12223
rect 18371 12192 18613 12220
rect 18371 12189 18383 12192
rect 18325 12183 18383 12189
rect 18601 12189 18613 12192
rect 18647 12189 18659 12223
rect 18874 12220 18880 12232
rect 18835 12192 18880 12220
rect 18601 12183 18659 12189
rect 11747 12124 12434 12152
rect 12796 12155 12854 12161
rect 11747 12121 11759 12124
rect 11701 12115 11759 12121
rect 12796 12121 12808 12155
rect 12842 12152 12854 12155
rect 14090 12152 14096 12164
rect 12842 12124 14096 12152
rect 12842 12121 12854 12124
rect 12796 12115 12854 12121
rect 14090 12112 14096 12124
rect 14148 12112 14154 12164
rect 17865 12155 17923 12161
rect 17865 12121 17877 12155
rect 17911 12152 17923 12155
rect 18141 12155 18199 12161
rect 18141 12152 18153 12155
rect 17911 12124 18153 12152
rect 17911 12121 17923 12124
rect 17865 12115 17923 12121
rect 18141 12121 18153 12124
rect 18187 12152 18199 12155
rect 18506 12152 18512 12164
rect 18187 12124 18512 12152
rect 18187 12121 18199 12124
rect 18141 12115 18199 12121
rect 18506 12112 18512 12124
rect 18564 12112 18570 12164
rect 18616 12152 18644 12183
rect 18874 12180 18880 12192
rect 18932 12180 18938 12232
rect 19076 12220 19104 12260
rect 19150 12248 19156 12300
rect 19208 12288 19214 12300
rect 19245 12291 19303 12297
rect 19245 12288 19257 12291
rect 19208 12260 19257 12288
rect 19208 12248 19214 12260
rect 19245 12257 19257 12260
rect 19291 12257 19303 12291
rect 19245 12251 19303 12257
rect 19501 12223 19559 12229
rect 19501 12220 19513 12223
rect 19076 12192 19513 12220
rect 19501 12189 19513 12192
rect 19547 12220 19559 12223
rect 20732 12220 20760 12328
rect 20806 12248 20812 12300
rect 20864 12288 20870 12300
rect 20864 12260 20909 12288
rect 20864 12248 20870 12260
rect 19547 12192 20760 12220
rect 19547 12189 19559 12192
rect 19501 12183 19559 12189
rect 20898 12180 20904 12232
rect 20956 12220 20962 12232
rect 21085 12223 21143 12229
rect 21085 12220 21097 12223
rect 20956 12192 21097 12220
rect 20956 12180 20962 12192
rect 21085 12189 21097 12192
rect 21131 12189 21143 12223
rect 21192 12220 21220 12328
rect 21284 12288 21312 12396
rect 21358 12316 21364 12368
rect 21416 12356 21422 12368
rect 21416 12328 22968 12356
rect 21416 12316 21422 12328
rect 21634 12288 21640 12300
rect 21284 12260 21640 12288
rect 21634 12248 21640 12260
rect 21692 12248 21698 12300
rect 22830 12288 22836 12300
rect 22791 12260 22836 12288
rect 22830 12248 22836 12260
rect 22888 12248 22894 12300
rect 22940 12297 22968 12328
rect 22925 12291 22983 12297
rect 22925 12257 22937 12291
rect 22971 12257 22983 12291
rect 22925 12251 22983 12257
rect 21913 12223 21971 12229
rect 21913 12220 21925 12223
rect 21192 12192 21925 12220
rect 21085 12183 21143 12189
rect 21913 12189 21925 12192
rect 21959 12189 21971 12223
rect 21913 12183 21971 12189
rect 22646 12180 22652 12232
rect 22704 12220 22710 12232
rect 22741 12223 22799 12229
rect 22741 12220 22753 12223
rect 22704 12192 22753 12220
rect 22704 12180 22710 12192
rect 22741 12189 22753 12192
rect 22787 12189 22799 12223
rect 22741 12183 22799 12189
rect 19334 12152 19340 12164
rect 18616 12124 19340 12152
rect 19334 12112 19340 12124
rect 19392 12112 19398 12164
rect 19610 12112 19616 12164
rect 19668 12152 19674 12164
rect 20993 12155 21051 12161
rect 20993 12152 21005 12155
rect 19668 12124 21005 12152
rect 19668 12112 19674 12124
rect 20993 12121 21005 12124
rect 21039 12121 21051 12155
rect 21821 12155 21879 12161
rect 21821 12152 21833 12155
rect 20993 12115 21051 12121
rect 21100 12124 21833 12152
rect 9907 12056 10456 12084
rect 9907 12053 9919 12056
rect 9861 12047 9919 12053
rect 11330 12044 11336 12096
rect 11388 12084 11394 12096
rect 11425 12087 11483 12093
rect 11425 12084 11437 12087
rect 11388 12056 11437 12084
rect 11388 12044 11394 12056
rect 11425 12053 11437 12056
rect 11471 12053 11483 12087
rect 13906 12084 13912 12096
rect 13819 12056 13912 12084
rect 11425 12047 11483 12053
rect 13906 12044 13912 12056
rect 13964 12084 13970 12096
rect 19702 12084 19708 12096
rect 13964 12056 19708 12084
rect 13964 12044 13970 12056
rect 19702 12044 19708 12056
rect 19760 12044 19766 12096
rect 20622 12084 20628 12096
rect 20583 12056 20628 12084
rect 20622 12044 20628 12056
rect 20680 12044 20686 12096
rect 20714 12044 20720 12096
rect 20772 12084 20778 12096
rect 21100 12084 21128 12124
rect 21821 12121 21833 12124
rect 21867 12121 21879 12155
rect 21821 12115 21879 12121
rect 21450 12084 21456 12096
rect 20772 12056 21128 12084
rect 21411 12056 21456 12084
rect 20772 12044 20778 12056
rect 21450 12044 21456 12056
rect 21508 12044 21514 12096
rect 22278 12084 22284 12096
rect 22239 12056 22284 12084
rect 22278 12044 22284 12056
rect 22336 12044 22342 12096
rect 22373 12087 22431 12093
rect 22373 12053 22385 12087
rect 22419 12084 22431 12087
rect 23474 12084 23480 12096
rect 22419 12056 23480 12084
rect 22419 12053 22431 12056
rect 22373 12047 22431 12053
rect 23474 12044 23480 12056
rect 23532 12044 23538 12096
rect 1104 11994 23460 12016
rect 1104 11942 6548 11994
rect 6600 11942 6612 11994
rect 6664 11942 6676 11994
rect 6728 11942 6740 11994
rect 6792 11942 6804 11994
rect 6856 11942 12146 11994
rect 12198 11942 12210 11994
rect 12262 11942 12274 11994
rect 12326 11942 12338 11994
rect 12390 11942 12402 11994
rect 12454 11942 17744 11994
rect 17796 11942 17808 11994
rect 17860 11942 17872 11994
rect 17924 11942 17936 11994
rect 17988 11942 18000 11994
rect 18052 11942 23460 11994
rect 1104 11920 23460 11942
rect 2590 11880 2596 11892
rect 2551 11852 2596 11880
rect 2590 11840 2596 11852
rect 2648 11840 2654 11892
rect 2869 11883 2927 11889
rect 2869 11849 2881 11883
rect 2915 11880 2927 11883
rect 3050 11880 3056 11892
rect 2915 11852 3056 11880
rect 2915 11849 2927 11852
rect 2869 11843 2927 11849
rect 3050 11840 3056 11852
rect 3108 11840 3114 11892
rect 3605 11883 3663 11889
rect 3605 11849 3617 11883
rect 3651 11880 3663 11883
rect 3973 11883 4031 11889
rect 3973 11880 3985 11883
rect 3651 11852 3985 11880
rect 3651 11849 3663 11852
rect 3605 11843 3663 11849
rect 3973 11849 3985 11852
rect 4019 11849 4031 11883
rect 6362 11880 6368 11892
rect 6323 11852 6368 11880
rect 3973 11843 4031 11849
rect 6362 11840 6368 11852
rect 6420 11840 6426 11892
rect 10597 11883 10655 11889
rect 10597 11880 10609 11883
rect 6748 11852 10609 11880
rect 3513 11815 3571 11821
rect 3513 11781 3525 11815
rect 3559 11812 3571 11815
rect 4062 11812 4068 11824
rect 3559 11784 4068 11812
rect 3559 11781 3571 11784
rect 3513 11775 3571 11781
rect 4062 11772 4068 11784
rect 4120 11772 4126 11824
rect 4264 11784 6132 11812
rect 2774 11704 2780 11756
rect 2832 11744 2838 11756
rect 3053 11747 3111 11753
rect 2832 11716 2877 11744
rect 2832 11704 2838 11716
rect 3053 11713 3065 11747
rect 3099 11744 3111 11747
rect 3099 11716 3188 11744
rect 3099 11713 3111 11716
rect 3053 11707 3111 11713
rect 3160 11617 3188 11716
rect 3326 11704 3332 11756
rect 3384 11744 3390 11756
rect 4264 11744 4292 11784
rect 3384 11716 4292 11744
rect 4341 11747 4399 11753
rect 3384 11704 3390 11716
rect 4341 11713 4353 11747
rect 4387 11744 4399 11747
rect 4706 11744 4712 11756
rect 4387 11716 4712 11744
rect 4387 11713 4399 11716
rect 4341 11707 4399 11713
rect 4706 11704 4712 11716
rect 4764 11704 4770 11756
rect 5902 11704 5908 11756
rect 5960 11753 5966 11756
rect 5960 11744 5972 11753
rect 5960 11716 6005 11744
rect 5960 11707 5972 11716
rect 5960 11704 5966 11707
rect 3418 11636 3424 11688
rect 3476 11676 3482 11688
rect 3697 11679 3755 11685
rect 3697 11676 3709 11679
rect 3476 11648 3709 11676
rect 3476 11636 3482 11648
rect 3697 11645 3709 11648
rect 3743 11645 3755 11679
rect 3697 11639 3755 11645
rect 4433 11679 4491 11685
rect 4433 11645 4445 11679
rect 4479 11645 4491 11679
rect 4433 11639 4491 11645
rect 4617 11679 4675 11685
rect 4617 11645 4629 11679
rect 4663 11676 4675 11679
rect 4798 11676 4804 11688
rect 4663 11648 4804 11676
rect 4663 11645 4675 11648
rect 4617 11639 4675 11645
rect 3145 11611 3203 11617
rect 3145 11577 3157 11611
rect 3191 11577 3203 11611
rect 4448 11608 4476 11639
rect 4798 11636 4804 11648
rect 4856 11636 4862 11688
rect 6104 11676 6132 11784
rect 6181 11747 6239 11753
rect 6181 11713 6193 11747
rect 6227 11744 6239 11747
rect 6380 11744 6408 11840
rect 6549 11747 6607 11753
rect 6549 11744 6561 11747
rect 6227 11716 6561 11744
rect 6227 11713 6239 11716
rect 6181 11707 6239 11713
rect 6549 11713 6561 11716
rect 6595 11713 6607 11747
rect 6549 11707 6607 11713
rect 6748 11676 6776 11852
rect 10597 11849 10609 11852
rect 10643 11880 10655 11883
rect 11514 11880 11520 11892
rect 10643 11852 11520 11880
rect 10643 11849 10655 11852
rect 10597 11843 10655 11849
rect 11514 11840 11520 11852
rect 11572 11840 11578 11892
rect 12434 11840 12440 11892
rect 12492 11880 12498 11892
rect 12710 11880 12716 11892
rect 12492 11852 12716 11880
rect 12492 11840 12498 11852
rect 12710 11840 12716 11852
rect 12768 11880 12774 11892
rect 12897 11883 12955 11889
rect 12897 11880 12909 11883
rect 12768 11852 12909 11880
rect 12768 11840 12774 11852
rect 12897 11849 12909 11852
rect 12943 11849 12955 11883
rect 12897 11843 12955 11849
rect 17037 11883 17095 11889
rect 17037 11849 17049 11883
rect 17083 11880 17095 11883
rect 18874 11880 18880 11892
rect 17083 11852 18880 11880
rect 17083 11849 17095 11852
rect 17037 11843 17095 11849
rect 18874 11840 18880 11852
rect 18932 11840 18938 11892
rect 20438 11880 20444 11892
rect 20399 11852 20444 11880
rect 20438 11840 20444 11852
rect 20496 11880 20502 11892
rect 20901 11883 20959 11889
rect 20901 11880 20913 11883
rect 20496 11852 20913 11880
rect 20496 11840 20502 11852
rect 20901 11849 20913 11852
rect 20947 11849 20959 11883
rect 20901 11843 20959 11849
rect 21450 11840 21456 11892
rect 21508 11880 21514 11892
rect 22189 11883 22247 11889
rect 22189 11880 22201 11883
rect 21508 11852 22201 11880
rect 21508 11840 21514 11852
rect 22189 11849 22201 11852
rect 22235 11849 22247 11883
rect 22189 11843 22247 11849
rect 9232 11784 10548 11812
rect 7834 11704 7840 11756
rect 7892 11704 7898 11756
rect 8012 11747 8070 11753
rect 8012 11713 8024 11747
rect 8058 11744 8070 11747
rect 9030 11744 9036 11756
rect 8058 11716 9036 11744
rect 8058 11713 8070 11716
rect 8012 11707 8070 11713
rect 9030 11704 9036 11716
rect 9088 11704 9094 11756
rect 9232 11753 9260 11784
rect 9217 11747 9275 11753
rect 9217 11713 9229 11747
rect 9263 11713 9275 11747
rect 9217 11707 9275 11713
rect 9306 11704 9312 11756
rect 9364 11744 9370 11756
rect 9473 11747 9531 11753
rect 9473 11744 9485 11747
rect 9364 11716 9485 11744
rect 9364 11704 9370 11716
rect 9473 11713 9485 11716
rect 9519 11713 9531 11747
rect 9473 11707 9531 11713
rect 6104 11648 6776 11676
rect 6822 11636 6828 11688
rect 6880 11676 6886 11688
rect 7745 11679 7803 11685
rect 7745 11676 7757 11679
rect 6880 11648 7757 11676
rect 6880 11636 6886 11648
rect 7745 11645 7757 11648
rect 7791 11676 7803 11679
rect 7852 11676 7880 11704
rect 10520 11688 10548 11784
rect 11606 11772 11612 11824
rect 11664 11812 11670 11824
rect 11762 11815 11820 11821
rect 11762 11812 11774 11815
rect 11664 11784 11774 11812
rect 11664 11772 11670 11784
rect 11762 11781 11774 11784
rect 11808 11781 11820 11815
rect 11762 11775 11820 11781
rect 16853 11815 16911 11821
rect 16853 11781 16865 11815
rect 16899 11812 16911 11815
rect 19328 11815 19386 11821
rect 16899 11784 18828 11812
rect 16899 11781 16911 11784
rect 16853 11775 16911 11781
rect 10778 11704 10784 11756
rect 10836 11744 10842 11756
rect 12618 11744 12624 11756
rect 10836 11716 12624 11744
rect 10836 11704 10842 11716
rect 12618 11704 12624 11716
rect 12676 11704 12682 11756
rect 15746 11704 15752 11756
rect 15804 11753 15810 11756
rect 15804 11744 15816 11753
rect 15804 11716 15849 11744
rect 15804 11707 15816 11716
rect 15804 11704 15810 11707
rect 18230 11704 18236 11756
rect 18288 11753 18294 11756
rect 18800 11753 18828 11784
rect 19328 11781 19340 11815
rect 19374 11812 19386 11815
rect 20622 11812 20628 11824
rect 19374 11784 20628 11812
rect 19374 11781 19386 11784
rect 19328 11775 19386 11781
rect 20622 11772 20628 11784
rect 20680 11812 20686 11824
rect 20809 11815 20867 11821
rect 20809 11812 20821 11815
rect 20680 11784 20821 11812
rect 20680 11772 20686 11784
rect 20809 11781 20821 11784
rect 20855 11781 20867 11815
rect 20809 11775 20867 11781
rect 21545 11815 21603 11821
rect 21545 11781 21557 11815
rect 21591 11812 21603 11815
rect 21910 11812 21916 11824
rect 21591 11784 21916 11812
rect 21591 11781 21603 11784
rect 21545 11775 21603 11781
rect 21910 11772 21916 11784
rect 21968 11772 21974 11824
rect 22462 11812 22468 11824
rect 22066 11784 22468 11812
rect 18288 11744 18300 11753
rect 18785 11747 18843 11753
rect 18288 11716 18333 11744
rect 18288 11707 18300 11716
rect 18785 11713 18797 11747
rect 18831 11744 18843 11747
rect 19610 11744 19616 11756
rect 18831 11716 19616 11744
rect 18831 11713 18843 11716
rect 18785 11707 18843 11713
rect 18288 11704 18294 11707
rect 19610 11704 19616 11716
rect 19668 11704 19674 11756
rect 19702 11704 19708 11756
rect 19760 11744 19766 11756
rect 22066 11744 22094 11784
rect 22462 11772 22468 11784
rect 22520 11772 22526 11824
rect 19760 11716 22094 11744
rect 19760 11704 19766 11716
rect 22186 11704 22192 11756
rect 22244 11744 22250 11756
rect 22281 11747 22339 11753
rect 22281 11744 22293 11747
rect 22244 11716 22293 11744
rect 22244 11704 22250 11716
rect 22281 11713 22293 11716
rect 22327 11713 22339 11747
rect 22281 11707 22339 11713
rect 22833 11747 22891 11753
rect 22833 11713 22845 11747
rect 22879 11744 22891 11747
rect 22922 11744 22928 11756
rect 22879 11716 22928 11744
rect 22879 11713 22891 11716
rect 22833 11707 22891 11713
rect 22922 11704 22928 11716
rect 22980 11704 22986 11756
rect 23109 11747 23167 11753
rect 23109 11713 23121 11747
rect 23155 11744 23167 11747
rect 23198 11744 23204 11756
rect 23155 11716 23204 11744
rect 23155 11713 23167 11716
rect 23109 11707 23167 11713
rect 23198 11704 23204 11716
rect 23256 11704 23262 11756
rect 7791 11648 7880 11676
rect 7791 11645 7803 11648
rect 7745 11639 7803 11645
rect 10502 11636 10508 11688
rect 10560 11676 10566 11688
rect 10689 11679 10747 11685
rect 10689 11676 10701 11679
rect 10560 11648 10701 11676
rect 10560 11636 10566 11648
rect 10689 11645 10701 11648
rect 10735 11676 10747 11679
rect 11517 11679 11575 11685
rect 11517 11676 11529 11679
rect 10735 11648 11529 11676
rect 10735 11645 10747 11648
rect 10689 11639 10747 11645
rect 11517 11645 11529 11648
rect 11563 11645 11575 11679
rect 11517 11639 11575 11645
rect 16025 11679 16083 11685
rect 16025 11645 16037 11679
rect 16071 11676 16083 11679
rect 16071 11648 16160 11676
rect 16071 11645 16083 11648
rect 16025 11639 16083 11645
rect 4448 11580 4844 11608
rect 3145 11571 3203 11577
rect 4816 11549 4844 11580
rect 16132 11552 16160 11648
rect 18506 11636 18512 11688
rect 18564 11676 18570 11688
rect 19061 11679 19119 11685
rect 19061 11676 19073 11679
rect 18564 11648 19073 11676
rect 18564 11636 18570 11648
rect 16390 11568 16396 11620
rect 16448 11608 16454 11620
rect 16448 11580 17632 11608
rect 16448 11568 16454 11580
rect 4801 11543 4859 11549
rect 4801 11509 4813 11543
rect 4847 11540 4859 11543
rect 5810 11540 5816 11552
rect 4847 11512 5816 11540
rect 4847 11509 4859 11512
rect 4801 11503 4859 11509
rect 5810 11500 5816 11512
rect 5868 11500 5874 11552
rect 9125 11543 9183 11549
rect 9125 11509 9137 11543
rect 9171 11540 9183 11543
rect 10410 11540 10416 11552
rect 9171 11512 10416 11540
rect 9171 11509 9183 11512
rect 9125 11503 9183 11509
rect 10410 11500 10416 11512
rect 10468 11540 10474 11552
rect 10778 11540 10784 11552
rect 10468 11512 10784 11540
rect 10468 11500 10474 11512
rect 10778 11500 10784 11512
rect 10836 11500 10842 11552
rect 13078 11540 13084 11552
rect 13039 11512 13084 11540
rect 13078 11500 13084 11512
rect 13136 11540 13142 11552
rect 13173 11543 13231 11549
rect 13173 11540 13185 11543
rect 13136 11512 13185 11540
rect 13136 11500 13142 11512
rect 13173 11509 13185 11512
rect 13219 11509 13231 11543
rect 13173 11503 13231 11509
rect 14645 11543 14703 11549
rect 14645 11509 14657 11543
rect 14691 11540 14703 11543
rect 15286 11540 15292 11552
rect 14691 11512 15292 11540
rect 14691 11509 14703 11512
rect 14645 11503 14703 11509
rect 15286 11500 15292 11512
rect 15344 11500 15350 11552
rect 16114 11540 16120 11552
rect 16075 11512 16120 11540
rect 16114 11500 16120 11512
rect 16172 11500 16178 11552
rect 16482 11540 16488 11552
rect 16443 11512 16488 11540
rect 16482 11500 16488 11512
rect 16540 11500 16546 11552
rect 17126 11540 17132 11552
rect 17087 11512 17132 11540
rect 17126 11500 17132 11512
rect 17184 11500 17190 11552
rect 17604 11540 17632 11580
rect 18892 11552 18920 11648
rect 19061 11645 19073 11648
rect 19107 11645 19119 11679
rect 19061 11639 19119 11645
rect 20717 11679 20775 11685
rect 20717 11645 20729 11679
rect 20763 11676 20775 11679
rect 20806 11676 20812 11688
rect 20763 11648 20812 11676
rect 20763 11645 20775 11648
rect 20717 11639 20775 11645
rect 20806 11636 20812 11648
rect 20864 11636 20870 11688
rect 22370 11676 22376 11688
rect 22331 11648 22376 11676
rect 22370 11636 22376 11648
rect 22428 11636 22434 11688
rect 21358 11608 21364 11620
rect 21319 11580 21364 11608
rect 21358 11568 21364 11580
rect 21416 11568 21422 11620
rect 22462 11568 22468 11620
rect 22520 11608 22526 11620
rect 22925 11611 22983 11617
rect 22925 11608 22937 11611
rect 22520 11580 22937 11608
rect 22520 11568 22526 11580
rect 22925 11577 22937 11580
rect 22971 11577 22983 11611
rect 22925 11571 22983 11577
rect 18322 11540 18328 11552
rect 17604 11512 18328 11540
rect 18322 11500 18328 11512
rect 18380 11500 18386 11552
rect 18693 11543 18751 11549
rect 18693 11509 18705 11543
rect 18739 11540 18751 11543
rect 18874 11540 18880 11552
rect 18739 11512 18880 11540
rect 18739 11509 18751 11512
rect 18693 11503 18751 11509
rect 18874 11500 18880 11512
rect 18932 11500 18938 11552
rect 18969 11543 19027 11549
rect 18969 11509 18981 11543
rect 19015 11540 19027 11543
rect 20990 11540 20996 11552
rect 19015 11512 20996 11540
rect 19015 11509 19027 11512
rect 18969 11503 19027 11509
rect 20990 11500 20996 11512
rect 21048 11500 21054 11552
rect 21266 11540 21272 11552
rect 21227 11512 21272 11540
rect 21266 11500 21272 11512
rect 21324 11500 21330 11552
rect 21818 11540 21824 11552
rect 21779 11512 21824 11540
rect 21818 11500 21824 11512
rect 21876 11500 21882 11552
rect 22646 11540 22652 11552
rect 22607 11512 22652 11540
rect 22646 11500 22652 11512
rect 22704 11500 22710 11552
rect 1104 11450 23460 11472
rect 1104 11398 3749 11450
rect 3801 11398 3813 11450
rect 3865 11398 3877 11450
rect 3929 11398 3941 11450
rect 3993 11398 4005 11450
rect 4057 11398 9347 11450
rect 9399 11398 9411 11450
rect 9463 11398 9475 11450
rect 9527 11398 9539 11450
rect 9591 11398 9603 11450
rect 9655 11398 14945 11450
rect 14997 11398 15009 11450
rect 15061 11398 15073 11450
rect 15125 11398 15137 11450
rect 15189 11398 15201 11450
rect 15253 11398 20543 11450
rect 20595 11398 20607 11450
rect 20659 11398 20671 11450
rect 20723 11398 20735 11450
rect 20787 11398 20799 11450
rect 20851 11398 23460 11450
rect 1104 11376 23460 11398
rect 3510 11296 3516 11348
rect 3568 11336 3574 11348
rect 3605 11339 3663 11345
rect 3605 11336 3617 11339
rect 3568 11308 3617 11336
rect 3568 11296 3574 11308
rect 3605 11305 3617 11308
rect 3651 11305 3663 11339
rect 4246 11336 4252 11348
rect 4207 11308 4252 11336
rect 3605 11299 3663 11305
rect 4246 11296 4252 11308
rect 4304 11296 4310 11348
rect 5258 11336 5264 11348
rect 5219 11308 5264 11336
rect 5258 11296 5264 11308
rect 5316 11296 5322 11348
rect 9030 11336 9036 11348
rect 8943 11308 9036 11336
rect 9030 11296 9036 11308
rect 9088 11336 9094 11348
rect 10042 11336 10048 11348
rect 9088 11308 10048 11336
rect 9088 11296 9094 11308
rect 10042 11296 10048 11308
rect 10100 11296 10106 11348
rect 12437 11339 12495 11345
rect 12437 11305 12449 11339
rect 12483 11336 12495 11339
rect 12526 11336 12532 11348
rect 12483 11308 12532 11336
rect 12483 11305 12495 11308
rect 12437 11299 12495 11305
rect 12526 11296 12532 11308
rect 12584 11296 12590 11348
rect 13909 11339 13967 11345
rect 13909 11305 13921 11339
rect 13955 11336 13967 11339
rect 16390 11336 16396 11348
rect 13955 11308 16396 11336
rect 13955 11305 13967 11308
rect 13909 11299 13967 11305
rect 16390 11296 16396 11308
rect 16448 11296 16454 11348
rect 16482 11296 16488 11348
rect 16540 11336 16546 11348
rect 19061 11339 19119 11345
rect 16540 11308 18920 11336
rect 16540 11296 16546 11308
rect 3418 11268 3424 11280
rect 3068 11240 3424 11268
rect 3068 11209 3096 11240
rect 3418 11228 3424 11240
rect 3476 11268 3482 11280
rect 4982 11268 4988 11280
rect 3476 11240 4988 11268
rect 3476 11228 3482 11240
rect 4982 11228 4988 11240
rect 5040 11228 5046 11280
rect 6733 11271 6791 11277
rect 6733 11237 6745 11271
rect 6779 11237 6791 11271
rect 6733 11231 6791 11237
rect 18417 11271 18475 11277
rect 18417 11237 18429 11271
rect 18463 11268 18475 11271
rect 18506 11268 18512 11280
rect 18463 11240 18512 11268
rect 18463 11237 18475 11240
rect 18417 11231 18475 11237
rect 3053 11203 3111 11209
rect 3053 11169 3065 11203
rect 3099 11169 3111 11203
rect 4798 11200 4804 11212
rect 4759 11172 4804 11200
rect 3053 11163 3111 11169
rect 4798 11160 4804 11172
rect 4856 11160 4862 11212
rect 6748 11200 6776 11231
rect 18506 11228 18512 11240
rect 18564 11228 18570 11280
rect 6564 11172 6776 11200
rect 18892 11200 18920 11308
rect 19061 11305 19073 11339
rect 19107 11336 19119 11339
rect 19426 11336 19432 11348
rect 19107 11308 19432 11336
rect 19107 11305 19119 11308
rect 19061 11299 19119 11305
rect 19426 11296 19432 11308
rect 19484 11296 19490 11348
rect 22738 11296 22744 11348
rect 22796 11336 22802 11348
rect 23017 11339 23075 11345
rect 23017 11336 23029 11339
rect 22796 11308 23029 11336
rect 22796 11296 22802 11308
rect 23017 11305 23029 11308
rect 23063 11305 23075 11339
rect 23017 11299 23075 11305
rect 20346 11228 20352 11280
rect 20404 11268 20410 11280
rect 20625 11271 20683 11277
rect 20625 11268 20637 11271
rect 20404 11240 20637 11268
rect 20404 11228 20410 11240
rect 20625 11237 20637 11240
rect 20671 11237 20683 11271
rect 20625 11231 20683 11237
rect 20717 11271 20775 11277
rect 20717 11237 20729 11271
rect 20763 11268 20775 11271
rect 20898 11268 20904 11280
rect 20763 11240 20904 11268
rect 20763 11237 20775 11240
rect 20717 11231 20775 11237
rect 18892 11172 19380 11200
rect 3237 11135 3295 11141
rect 3237 11101 3249 11135
rect 3283 11132 3295 11135
rect 3602 11132 3608 11144
rect 3283 11104 3608 11132
rect 3283 11101 3295 11104
rect 3237 11095 3295 11101
rect 3602 11092 3608 11104
rect 3660 11092 3666 11144
rect 4617 11135 4675 11141
rect 4617 11101 4629 11135
rect 4663 11132 4675 11135
rect 5902 11132 5908 11144
rect 4663 11104 5908 11132
rect 4663 11101 4675 11104
rect 4617 11095 4675 11101
rect 5902 11092 5908 11104
rect 5960 11132 5966 11144
rect 6564 11132 6592 11172
rect 5960 11104 6592 11132
rect 6641 11135 6699 11141
rect 5960 11092 5966 11104
rect 6641 11101 6653 11135
rect 6687 11132 6699 11135
rect 6822 11132 6828 11144
rect 6687 11104 6828 11132
rect 6687 11101 6699 11104
rect 6641 11095 6699 11101
rect 6822 11092 6828 11104
rect 6880 11132 6886 11144
rect 8113 11135 8171 11141
rect 8113 11132 8125 11135
rect 6880 11104 8125 11132
rect 6880 11092 6886 11104
rect 8113 11101 8125 11104
rect 8159 11132 8171 11135
rect 10413 11135 10471 11141
rect 8159 11104 8340 11132
rect 8159 11101 8171 11104
rect 8113 11095 8171 11101
rect 4709 11067 4767 11073
rect 4709 11033 4721 11067
rect 4755 11064 4767 11067
rect 4755 11036 5488 11064
rect 4755 11033 4767 11036
rect 4709 11027 4767 11033
rect 3142 10996 3148 11008
rect 3103 10968 3148 10996
rect 3142 10956 3148 10968
rect 3200 10956 3206 11008
rect 5460 10996 5488 11036
rect 5534 11024 5540 11076
rect 5592 11064 5598 11076
rect 6374 11067 6432 11073
rect 6374 11064 6386 11067
rect 5592 11036 6386 11064
rect 5592 11024 5598 11036
rect 6374 11033 6386 11036
rect 6420 11033 6432 11067
rect 7846 11067 7904 11073
rect 7846 11064 7858 11067
rect 6374 11027 6432 11033
rect 6472 11036 7858 11064
rect 6472 10996 6500 11036
rect 7846 11033 7858 11036
rect 7892 11064 7904 11067
rect 8018 11064 8024 11076
rect 7892 11036 8024 11064
rect 7892 11033 7904 11036
rect 7846 11027 7904 11033
rect 8018 11024 8024 11036
rect 8076 11024 8082 11076
rect 8312 11005 8340 11104
rect 10413 11101 10425 11135
rect 10459 11132 10471 11135
rect 11057 11135 11115 11141
rect 11057 11132 11069 11135
rect 10459 11104 11069 11132
rect 10459 11101 10471 11104
rect 10413 11095 10471 11101
rect 9950 11024 9956 11076
rect 10008 11064 10014 11076
rect 10146 11067 10204 11073
rect 10146 11064 10158 11067
rect 10008 11036 10158 11064
rect 10008 11024 10014 11036
rect 10146 11033 10158 11036
rect 10192 11033 10204 11067
rect 10146 11027 10204 11033
rect 10520 11008 10548 11104
rect 11057 11101 11069 11104
rect 11103 11132 11115 11135
rect 12529 11135 12587 11141
rect 12529 11132 12541 11135
rect 11103 11104 12541 11132
rect 11103 11101 11115 11104
rect 11057 11095 11115 11101
rect 12529 11101 12541 11104
rect 12575 11132 12587 11135
rect 13078 11132 13084 11144
rect 12575 11104 13084 11132
rect 12575 11101 12587 11104
rect 12529 11095 12587 11101
rect 13078 11092 13084 11104
rect 13136 11132 13142 11144
rect 14093 11135 14151 11141
rect 14093 11132 14105 11135
rect 13136 11104 14105 11132
rect 13136 11092 13142 11104
rect 14093 11101 14105 11104
rect 14139 11132 14151 11135
rect 14829 11135 14887 11141
rect 14829 11132 14841 11135
rect 14139 11104 14841 11132
rect 14139 11101 14151 11104
rect 14093 11095 14151 11101
rect 14829 11101 14841 11104
rect 14875 11132 14887 11135
rect 15010 11132 15016 11144
rect 14875 11104 15016 11132
rect 14875 11101 14887 11104
rect 14829 11095 14887 11101
rect 15010 11092 15016 11104
rect 15068 11132 15074 11144
rect 16114 11132 16120 11144
rect 15068 11104 16120 11132
rect 15068 11092 15074 11104
rect 16114 11092 16120 11104
rect 16172 11132 16178 11144
rect 16485 11135 16543 11141
rect 16485 11132 16497 11135
rect 16172 11104 16497 11132
rect 16172 11092 16178 11104
rect 16485 11101 16497 11104
rect 16531 11132 16543 11135
rect 16669 11135 16727 11141
rect 16669 11132 16681 11135
rect 16531 11104 16681 11132
rect 16531 11101 16543 11104
rect 16485 11095 16543 11101
rect 16669 11101 16681 11104
rect 16715 11132 16727 11135
rect 16853 11135 16911 11141
rect 16853 11132 16865 11135
rect 16715 11104 16865 11132
rect 16715 11101 16727 11104
rect 16669 11095 16727 11101
rect 16853 11101 16865 11104
rect 16899 11132 16911 11135
rect 17037 11135 17095 11141
rect 17037 11132 17049 11135
rect 16899 11104 17049 11132
rect 16899 11101 16911 11104
rect 16853 11095 16911 11101
rect 17037 11101 17049 11104
rect 17083 11101 17095 11135
rect 18690 11132 18696 11144
rect 17037 11095 17095 11101
rect 17236 11104 18696 11132
rect 11324 11067 11382 11073
rect 11324 11033 11336 11067
rect 11370 11064 11382 11067
rect 12434 11064 12440 11076
rect 11370 11036 12440 11064
rect 11370 11033 11382 11036
rect 11324 11027 11382 11033
rect 12434 11024 12440 11036
rect 12492 11024 12498 11076
rect 12618 11024 12624 11076
rect 12676 11064 12682 11076
rect 12774 11067 12832 11073
rect 12774 11064 12786 11067
rect 12676 11036 12786 11064
rect 12676 11024 12682 11036
rect 12774 11033 12786 11036
rect 12820 11033 12832 11067
rect 12774 11027 12832 11033
rect 15280 11067 15338 11073
rect 15280 11033 15292 11067
rect 15326 11064 15338 11067
rect 17236 11064 17264 11104
rect 18690 11092 18696 11104
rect 18748 11092 18754 11144
rect 18892 11141 18920 11172
rect 19352 11144 19380 11172
rect 18877 11135 18935 11141
rect 18877 11101 18889 11135
rect 18923 11101 18935 11135
rect 18877 11095 18935 11101
rect 19245 11135 19303 11141
rect 19245 11101 19257 11135
rect 19291 11101 19303 11135
rect 19245 11095 19303 11101
rect 15326 11036 17264 11064
rect 17304 11067 17362 11073
rect 15326 11033 15338 11036
rect 15280 11027 15338 11033
rect 17304 11033 17316 11067
rect 17350 11033 17362 11067
rect 19260 11064 19288 11095
rect 19334 11092 19340 11144
rect 19392 11092 19398 11144
rect 19512 11135 19570 11141
rect 19512 11101 19524 11135
rect 19558 11132 19570 11135
rect 20732 11132 20760 11231
rect 20898 11228 20904 11240
rect 20956 11228 20962 11280
rect 22756 11268 22784 11296
rect 22922 11268 22928 11280
rect 22112 11240 22784 11268
rect 22883 11240 22928 11268
rect 22112 11209 22140 11240
rect 22922 11228 22928 11240
rect 22980 11228 22986 11280
rect 22097 11203 22155 11209
rect 22097 11169 22109 11203
rect 22143 11169 22155 11203
rect 22370 11200 22376 11212
rect 22331 11172 22376 11200
rect 22097 11163 22155 11169
rect 22370 11160 22376 11172
rect 22428 11160 22434 11212
rect 19558 11104 20760 11132
rect 19558 11101 19570 11104
rect 19512 11095 19570 11101
rect 21266 11092 21272 11144
rect 21324 11132 21330 11144
rect 22557 11135 22615 11141
rect 22557 11132 22569 11135
rect 21324 11104 22569 11132
rect 21324 11092 21330 11104
rect 22557 11101 22569 11104
rect 22603 11101 22615 11135
rect 22557 11095 22615 11101
rect 17304 11027 17362 11033
rect 18892 11036 19288 11064
rect 5460 10968 6500 10996
rect 8297 10999 8355 11005
rect 8297 10965 8309 10999
rect 8343 10996 8355 10999
rect 8386 10996 8392 11008
rect 8343 10968 8392 10996
rect 8343 10965 8355 10968
rect 8297 10959 8355 10965
rect 8386 10956 8392 10968
rect 8444 10956 8450 11008
rect 10502 10996 10508 11008
rect 10463 10968 10508 10996
rect 10502 10956 10508 10968
rect 10560 10956 10566 11008
rect 16390 10996 16396 11008
rect 16351 10968 16396 10996
rect 16390 10956 16396 10968
rect 16448 10956 16454 11008
rect 17034 10956 17040 11008
rect 17092 10996 17098 11008
rect 17328 10996 17356 11027
rect 18892 11008 18920 11036
rect 21082 11024 21088 11076
rect 21140 11064 21146 11076
rect 21450 11064 21456 11076
rect 21140 11036 21456 11064
rect 21140 11024 21146 11036
rect 21450 11024 21456 11036
rect 21508 11064 21514 11076
rect 21830 11067 21888 11073
rect 21830 11064 21842 11067
rect 21508 11036 21842 11064
rect 21508 11024 21514 11036
rect 21830 11033 21842 11036
rect 21876 11033 21888 11067
rect 21830 11027 21888 11033
rect 22278 11024 22284 11076
rect 22336 11064 22342 11076
rect 22465 11067 22523 11073
rect 22465 11064 22477 11067
rect 22336 11036 22477 11064
rect 22336 11024 22342 11036
rect 22465 11033 22477 11036
rect 22511 11033 22523 11067
rect 22465 11027 22523 11033
rect 17092 10968 17356 10996
rect 18693 10999 18751 11005
rect 17092 10956 17098 10968
rect 18693 10965 18705 10999
rect 18739 10996 18751 10999
rect 18874 10996 18880 11008
rect 18739 10968 18880 10996
rect 18739 10965 18751 10968
rect 18693 10959 18751 10965
rect 18874 10956 18880 10968
rect 18932 10956 18938 11008
rect 1104 10906 23460 10928
rect 1104 10854 6548 10906
rect 6600 10854 6612 10906
rect 6664 10854 6676 10906
rect 6728 10854 6740 10906
rect 6792 10854 6804 10906
rect 6856 10854 12146 10906
rect 12198 10854 12210 10906
rect 12262 10854 12274 10906
rect 12326 10854 12338 10906
rect 12390 10854 12402 10906
rect 12454 10854 17744 10906
rect 17796 10854 17808 10906
rect 17860 10854 17872 10906
rect 17924 10854 17936 10906
rect 17988 10854 18000 10906
rect 18052 10854 23460 10906
rect 1104 10832 23460 10854
rect 2866 10752 2872 10804
rect 2924 10792 2930 10804
rect 3053 10795 3111 10801
rect 3053 10792 3065 10795
rect 2924 10764 3065 10792
rect 2924 10752 2930 10764
rect 3053 10761 3065 10764
rect 3099 10761 3111 10795
rect 3053 10755 3111 10761
rect 3142 10752 3148 10804
rect 3200 10792 3206 10804
rect 3881 10795 3939 10801
rect 3881 10792 3893 10795
rect 3200 10764 3893 10792
rect 3200 10752 3206 10764
rect 3881 10761 3893 10764
rect 3927 10761 3939 10795
rect 3881 10755 3939 10761
rect 5445 10795 5503 10801
rect 5445 10761 5457 10795
rect 5491 10792 5503 10795
rect 5534 10792 5540 10804
rect 5491 10764 5540 10792
rect 5491 10761 5503 10764
rect 5445 10755 5503 10761
rect 5534 10752 5540 10764
rect 5592 10752 5598 10804
rect 6178 10792 6184 10804
rect 6139 10764 6184 10792
rect 6178 10752 6184 10764
rect 6236 10752 6242 10804
rect 6362 10752 6368 10804
rect 6420 10792 6426 10804
rect 6733 10795 6791 10801
rect 6733 10792 6745 10795
rect 6420 10764 6745 10792
rect 6420 10752 6426 10764
rect 6733 10761 6745 10764
rect 6779 10761 6791 10795
rect 13538 10792 13544 10804
rect 13499 10764 13544 10792
rect 6733 10755 6791 10761
rect 13538 10752 13544 10764
rect 13596 10752 13602 10804
rect 22094 10792 22100 10804
rect 20824 10764 22100 10792
rect 4249 10727 4307 10733
rect 4249 10693 4261 10727
rect 4295 10724 4307 10727
rect 6454 10724 6460 10736
rect 4295 10696 6460 10724
rect 4295 10693 4307 10696
rect 4249 10687 4307 10693
rect 6454 10684 6460 10696
rect 6512 10684 6518 10736
rect 8478 10684 8484 10736
rect 8536 10724 8542 10736
rect 11146 10733 11152 10736
rect 9594 10727 9652 10733
rect 9594 10724 9606 10727
rect 8536 10696 9606 10724
rect 8536 10684 8542 10696
rect 9594 10693 9606 10696
rect 9640 10693 9652 10727
rect 9594 10687 9652 10693
rect 11088 10727 11152 10733
rect 11088 10693 11100 10727
rect 11134 10693 11152 10727
rect 11088 10687 11152 10693
rect 11146 10684 11152 10687
rect 11204 10684 11210 10736
rect 12428 10727 12486 10733
rect 12428 10693 12440 10727
rect 12474 10724 12486 10727
rect 12526 10724 12532 10736
rect 12474 10696 12532 10724
rect 12474 10693 12486 10696
rect 12428 10687 12486 10693
rect 12526 10684 12532 10696
rect 12584 10684 12590 10736
rect 14768 10727 14826 10733
rect 14768 10693 14780 10727
rect 14814 10724 14826 10727
rect 14814 10696 15148 10724
rect 14814 10693 14826 10696
rect 14768 10687 14826 10693
rect 2774 10616 2780 10668
rect 2832 10656 2838 10668
rect 3237 10659 3295 10665
rect 3237 10656 3249 10659
rect 2832 10628 3249 10656
rect 2832 10616 2838 10628
rect 3237 10625 3249 10628
rect 3283 10625 3295 10659
rect 3237 10619 3295 10625
rect 4341 10659 4399 10665
rect 4341 10625 4353 10659
rect 4387 10656 4399 10659
rect 5442 10656 5448 10668
rect 4387 10628 5448 10656
rect 4387 10625 4399 10628
rect 4341 10619 4399 10625
rect 5442 10616 5448 10628
rect 5500 10656 5506 10668
rect 5537 10659 5595 10665
rect 5537 10656 5549 10659
rect 5500 10628 5549 10656
rect 5500 10616 5506 10628
rect 5537 10625 5549 10628
rect 5583 10625 5595 10659
rect 5537 10619 5595 10625
rect 8133 10659 8191 10665
rect 8133 10625 8145 10659
rect 8179 10656 8191 10659
rect 8846 10656 8852 10668
rect 8179 10628 8852 10656
rect 8179 10625 8191 10628
rect 8133 10619 8191 10625
rect 8846 10616 8852 10628
rect 8904 10616 8910 10668
rect 10502 10656 10508 10668
rect 9876 10628 10508 10656
rect 4522 10588 4528 10600
rect 4483 10560 4528 10588
rect 4522 10548 4528 10560
rect 4580 10548 4586 10600
rect 4706 10548 4712 10600
rect 4764 10588 4770 10600
rect 4801 10591 4859 10597
rect 4801 10588 4813 10591
rect 4764 10560 4813 10588
rect 4764 10548 4770 10560
rect 4801 10557 4813 10560
rect 4847 10557 4859 10591
rect 8386 10588 8392 10600
rect 8347 10560 8392 10588
rect 4801 10551 4859 10557
rect 8386 10548 8392 10560
rect 8444 10548 8450 10600
rect 9876 10597 9904 10628
rect 10502 10616 10508 10628
rect 10560 10656 10566 10668
rect 15010 10656 15016 10668
rect 10560 10628 11376 10656
rect 14971 10628 15016 10656
rect 10560 10616 10566 10628
rect 11348 10597 11376 10628
rect 15010 10616 15016 10628
rect 15068 10616 15074 10668
rect 9861 10591 9919 10597
rect 9861 10557 9873 10591
rect 9907 10557 9919 10591
rect 9861 10551 9919 10557
rect 11333 10591 11391 10597
rect 11333 10557 11345 10591
rect 11379 10588 11391 10591
rect 12161 10591 12219 10597
rect 12161 10588 12173 10591
rect 11379 10560 12173 10588
rect 11379 10557 11391 10560
rect 11333 10551 11391 10557
rect 8481 10523 8539 10529
rect 8481 10489 8493 10523
rect 8527 10489 8539 10523
rect 8481 10483 8539 10489
rect 6454 10412 6460 10464
rect 6512 10452 6518 10464
rect 7009 10455 7067 10461
rect 7009 10452 7021 10455
rect 6512 10424 7021 10452
rect 6512 10412 6518 10424
rect 7009 10421 7021 10424
rect 7055 10421 7067 10455
rect 7009 10415 7067 10421
rect 8018 10412 8024 10464
rect 8076 10452 8082 10464
rect 8496 10452 8524 10483
rect 11532 10464 11560 10560
rect 12161 10557 12173 10560
rect 12207 10557 12219 10591
rect 12161 10551 12219 10557
rect 9950 10452 9956 10464
rect 8076 10424 8524 10452
rect 9911 10424 9956 10452
rect 8076 10412 8082 10424
rect 9950 10412 9956 10424
rect 10008 10412 10014 10464
rect 11514 10452 11520 10464
rect 11475 10424 11520 10452
rect 11514 10412 11520 10424
rect 11572 10452 11578 10464
rect 11701 10455 11759 10461
rect 11701 10452 11713 10455
rect 11572 10424 11713 10452
rect 11572 10412 11578 10424
rect 11701 10421 11713 10424
rect 11747 10421 11759 10455
rect 13630 10452 13636 10464
rect 13591 10424 13636 10452
rect 11701 10415 11759 10421
rect 13630 10412 13636 10424
rect 13688 10412 13694 10464
rect 15120 10461 15148 10696
rect 16114 10684 16120 10736
rect 16172 10724 16178 10736
rect 16172 10696 16528 10724
rect 16172 10684 16178 10696
rect 16500 10665 16528 10696
rect 17034 10684 17040 10736
rect 17092 10724 17098 10736
rect 20824 10733 20852 10764
rect 22094 10752 22100 10764
rect 22152 10752 22158 10804
rect 22462 10792 22468 10804
rect 22423 10764 22468 10792
rect 22462 10752 22468 10764
rect 22520 10752 22526 10804
rect 22557 10795 22615 10801
rect 22557 10761 22569 10795
rect 22603 10792 22615 10795
rect 22646 10792 22652 10804
rect 22603 10764 22652 10792
rect 22603 10761 22615 10764
rect 22557 10755 22615 10761
rect 22646 10752 22652 10764
rect 22704 10752 22710 10804
rect 20809 10727 20867 10733
rect 17092 10696 20760 10724
rect 17092 10684 17098 10696
rect 16229 10659 16287 10665
rect 16229 10625 16241 10659
rect 16275 10656 16287 10659
rect 16485 10659 16543 10665
rect 16275 10628 16436 10656
rect 16275 10625 16287 10628
rect 16229 10619 16287 10625
rect 16408 10588 16436 10628
rect 16485 10625 16497 10659
rect 16531 10656 16543 10659
rect 16669 10659 16727 10665
rect 16669 10656 16681 10659
rect 16531 10628 16681 10656
rect 16531 10625 16543 10628
rect 16485 10619 16543 10625
rect 16669 10625 16681 10628
rect 16715 10625 16727 10659
rect 16669 10619 16727 10625
rect 16758 10616 16764 10668
rect 16816 10656 16822 10668
rect 16925 10659 16983 10665
rect 16925 10656 16937 10659
rect 16816 10628 16937 10656
rect 16816 10616 16822 10628
rect 16925 10625 16937 10628
rect 16971 10625 16983 10659
rect 18322 10656 18328 10668
rect 18283 10628 18328 10656
rect 16925 10619 16983 10625
rect 18322 10616 18328 10628
rect 18380 10616 18386 10668
rect 19144 10659 19202 10665
rect 19144 10656 19156 10659
rect 18616 10628 19156 10656
rect 18616 10588 18644 10628
rect 19144 10625 19156 10628
rect 19190 10656 19202 10659
rect 20625 10659 20683 10665
rect 20625 10656 20637 10659
rect 19190 10628 20637 10656
rect 19190 10625 19202 10628
rect 19144 10619 19202 10625
rect 20625 10625 20637 10628
rect 20671 10625 20683 10659
rect 20625 10619 20683 10625
rect 18782 10588 18788 10600
rect 16408 10560 16712 10588
rect 15105 10455 15163 10461
rect 15105 10421 15117 10455
rect 15151 10452 15163 10455
rect 16574 10452 16580 10464
rect 15151 10424 16580 10452
rect 15151 10421 15163 10424
rect 15105 10415 15163 10421
rect 16574 10412 16580 10424
rect 16632 10412 16638 10464
rect 16684 10452 16712 10560
rect 18064 10560 18644 10588
rect 18743 10560 18788 10588
rect 18064 10529 18092 10560
rect 18782 10548 18788 10560
rect 18840 10548 18846 10600
rect 18874 10548 18880 10600
rect 18932 10588 18938 10600
rect 18932 10560 18977 10588
rect 18932 10548 18938 10560
rect 18049 10523 18107 10529
rect 18049 10489 18061 10523
rect 18095 10489 18107 10523
rect 18049 10483 18107 10489
rect 18233 10523 18291 10529
rect 18233 10489 18245 10523
rect 18279 10520 18291 10523
rect 18892 10520 18920 10548
rect 18279 10492 18920 10520
rect 18279 10489 18291 10492
rect 18233 10483 18291 10489
rect 19886 10480 19892 10532
rect 19944 10520 19950 10532
rect 20441 10523 20499 10529
rect 20441 10520 20453 10523
rect 19944 10492 20453 10520
rect 19944 10480 19950 10492
rect 20441 10489 20453 10492
rect 20487 10489 20499 10523
rect 20732 10520 20760 10696
rect 20809 10693 20821 10727
rect 20855 10693 20867 10727
rect 20809 10687 20867 10693
rect 21269 10727 21327 10733
rect 21269 10693 21281 10727
rect 21315 10724 21327 10727
rect 22278 10724 22284 10736
rect 21315 10696 22284 10724
rect 21315 10693 21327 10696
rect 21269 10687 21327 10693
rect 22278 10684 22284 10696
rect 22336 10684 22342 10736
rect 21818 10656 21824 10668
rect 21779 10628 21824 10656
rect 21818 10616 21824 10628
rect 21876 10616 21882 10668
rect 23109 10659 23167 10665
rect 23109 10625 23121 10659
rect 23155 10656 23167 10659
rect 23290 10656 23296 10668
rect 23155 10628 23296 10656
rect 23155 10625 23167 10628
rect 23109 10619 23167 10625
rect 23290 10616 23296 10628
rect 23348 10616 23354 10668
rect 21358 10588 21364 10600
rect 21319 10560 21364 10588
rect 21358 10548 21364 10560
rect 21416 10548 21422 10600
rect 21450 10548 21456 10600
rect 21508 10588 21514 10600
rect 21508 10560 21553 10588
rect 21508 10548 21514 10560
rect 22186 10548 22192 10600
rect 22244 10588 22250 10600
rect 22649 10591 22707 10597
rect 22649 10588 22661 10591
rect 22244 10560 22661 10588
rect 22244 10548 22250 10560
rect 22649 10557 22661 10560
rect 22695 10557 22707 10591
rect 22649 10551 22707 10557
rect 21818 10520 21824 10532
rect 20732 10492 21824 10520
rect 20441 10483 20499 10489
rect 21818 10480 21824 10492
rect 21876 10480 21882 10532
rect 17402 10452 17408 10464
rect 16684 10424 17408 10452
rect 17402 10412 17408 10424
rect 17460 10412 17466 10464
rect 18509 10455 18567 10461
rect 18509 10421 18521 10455
rect 18555 10452 18567 10455
rect 19242 10452 19248 10464
rect 18555 10424 19248 10452
rect 18555 10421 18567 10424
rect 18509 10415 18567 10421
rect 19242 10412 19248 10424
rect 19300 10412 19306 10464
rect 20254 10452 20260 10464
rect 20215 10424 20260 10452
rect 20254 10412 20260 10424
rect 20312 10412 20318 10464
rect 20901 10455 20959 10461
rect 20901 10421 20913 10455
rect 20947 10452 20959 10455
rect 21174 10452 21180 10464
rect 20947 10424 21180 10452
rect 20947 10421 20959 10424
rect 20901 10415 20959 10421
rect 21174 10412 21180 10424
rect 21232 10412 21238 10464
rect 22002 10452 22008 10464
rect 21963 10424 22008 10452
rect 22002 10412 22008 10424
rect 22060 10412 22066 10464
rect 22094 10412 22100 10464
rect 22152 10452 22158 10464
rect 22152 10424 22197 10452
rect 22152 10412 22158 10424
rect 22370 10412 22376 10464
rect 22428 10452 22434 10464
rect 22925 10455 22983 10461
rect 22925 10452 22937 10455
rect 22428 10424 22937 10452
rect 22428 10412 22434 10424
rect 22925 10421 22937 10424
rect 22971 10421 22983 10455
rect 22925 10415 22983 10421
rect 1104 10362 23460 10384
rect 1104 10310 3749 10362
rect 3801 10310 3813 10362
rect 3865 10310 3877 10362
rect 3929 10310 3941 10362
rect 3993 10310 4005 10362
rect 4057 10310 9347 10362
rect 9399 10310 9411 10362
rect 9463 10310 9475 10362
rect 9527 10310 9539 10362
rect 9591 10310 9603 10362
rect 9655 10310 14945 10362
rect 14997 10310 15009 10362
rect 15061 10310 15073 10362
rect 15125 10310 15137 10362
rect 15189 10310 15201 10362
rect 15253 10310 20543 10362
rect 20595 10310 20607 10362
rect 20659 10310 20671 10362
rect 20723 10310 20735 10362
rect 20787 10310 20799 10362
rect 20851 10310 23460 10362
rect 1104 10288 23460 10310
rect 2498 10248 2504 10260
rect 2459 10220 2504 10248
rect 2498 10208 2504 10220
rect 2556 10208 2562 10260
rect 2777 10251 2835 10257
rect 2777 10217 2789 10251
rect 2823 10248 2835 10251
rect 2958 10248 2964 10260
rect 2823 10220 2964 10248
rect 2823 10217 2835 10220
rect 2777 10211 2835 10217
rect 2958 10208 2964 10220
rect 3016 10208 3022 10260
rect 5077 10251 5135 10257
rect 5077 10217 5089 10251
rect 5123 10248 5135 10251
rect 6362 10248 6368 10260
rect 5123 10220 6368 10248
rect 5123 10217 5135 10220
rect 5077 10211 5135 10217
rect 6362 10208 6368 10220
rect 6420 10248 6426 10260
rect 6420 10220 6776 10248
rect 6420 10208 6426 10220
rect 2869 10183 2927 10189
rect 2869 10180 2881 10183
rect 2746 10152 2881 10180
rect 2314 10044 2320 10056
rect 2275 10016 2320 10044
rect 2314 10004 2320 10016
rect 2372 10004 2378 10056
rect 2593 10047 2651 10053
rect 2593 10013 2605 10047
rect 2639 10044 2651 10047
rect 2746 10044 2774 10152
rect 2869 10149 2881 10152
rect 2915 10149 2927 10183
rect 2869 10143 2927 10149
rect 4706 10140 4712 10192
rect 4764 10180 4770 10192
rect 5353 10183 5411 10189
rect 5353 10180 5365 10183
rect 4764 10152 5365 10180
rect 4764 10140 4770 10152
rect 5353 10149 5365 10152
rect 5399 10149 5411 10183
rect 5353 10143 5411 10149
rect 3050 10072 3056 10124
rect 3108 10112 3114 10124
rect 3418 10112 3424 10124
rect 3108 10084 3424 10112
rect 3108 10072 3114 10084
rect 3418 10072 3424 10084
rect 3476 10072 3482 10124
rect 4433 10115 4491 10121
rect 4433 10081 4445 10115
rect 4479 10112 4491 10115
rect 4522 10112 4528 10124
rect 4479 10084 4528 10112
rect 4479 10081 4491 10084
rect 4433 10075 4491 10081
rect 4522 10072 4528 10084
rect 4580 10112 4586 10124
rect 6748 10121 6776 10220
rect 8846 10208 8852 10260
rect 8904 10248 8910 10260
rect 8941 10251 8999 10257
rect 8941 10248 8953 10251
rect 8904 10220 8953 10248
rect 8904 10208 8910 10220
rect 8941 10217 8953 10220
rect 8987 10217 8999 10251
rect 17221 10251 17279 10257
rect 17221 10248 17233 10251
rect 8941 10211 8999 10217
rect 15672 10220 17233 10248
rect 15672 10121 15700 10220
rect 17221 10217 17233 10220
rect 17267 10248 17279 10251
rect 17405 10251 17463 10257
rect 17405 10248 17417 10251
rect 17267 10220 17417 10248
rect 17267 10217 17279 10220
rect 17221 10211 17279 10217
rect 17405 10217 17417 10220
rect 17451 10248 17463 10251
rect 17681 10251 17739 10257
rect 17681 10248 17693 10251
rect 17451 10220 17693 10248
rect 17451 10217 17463 10220
rect 17405 10211 17463 10217
rect 17681 10217 17693 10220
rect 17727 10248 17739 10251
rect 18874 10248 18880 10260
rect 17727 10220 18880 10248
rect 17727 10217 17739 10220
rect 17681 10211 17739 10217
rect 18874 10208 18880 10220
rect 18932 10248 18938 10260
rect 18932 10220 20668 10248
rect 18932 10208 18938 10220
rect 17034 10180 17040 10192
rect 16995 10152 17040 10180
rect 17034 10140 17040 10152
rect 17092 10140 17098 10192
rect 17957 10183 18015 10189
rect 17957 10149 17969 10183
rect 18003 10180 18015 10183
rect 19610 10180 19616 10192
rect 18003 10152 19616 10180
rect 18003 10149 18015 10152
rect 17957 10143 18015 10149
rect 19610 10140 19616 10152
rect 19668 10140 19674 10192
rect 6733 10115 6791 10121
rect 4580 10084 4844 10112
rect 4580 10072 4586 10084
rect 2639 10016 2774 10044
rect 4249 10047 4307 10053
rect 2639 10013 2651 10016
rect 2593 10007 2651 10013
rect 4249 10013 4261 10047
rect 4295 10044 4307 10047
rect 4706 10044 4712 10056
rect 4295 10016 4712 10044
rect 4295 10013 4307 10016
rect 4249 10007 4307 10013
rect 4706 10004 4712 10016
rect 4764 10004 4770 10056
rect 4816 10053 4844 10084
rect 6733 10081 6745 10115
rect 6779 10112 6791 10115
rect 6825 10115 6883 10121
rect 6825 10112 6837 10115
rect 6779 10084 6837 10112
rect 6779 10081 6791 10084
rect 6733 10075 6791 10081
rect 6825 10081 6837 10084
rect 6871 10081 6883 10115
rect 6825 10075 6883 10081
rect 15565 10115 15623 10121
rect 15565 10081 15577 10115
rect 15611 10112 15623 10115
rect 15657 10115 15715 10121
rect 15657 10112 15669 10115
rect 15611 10084 15669 10112
rect 15611 10081 15623 10084
rect 15565 10075 15623 10081
rect 15657 10081 15669 10084
rect 15703 10081 15715 10115
rect 18230 10112 18236 10124
rect 15657 10075 15715 10081
rect 18064 10084 18236 10112
rect 4801 10047 4859 10053
rect 4801 10013 4813 10047
rect 4847 10013 4859 10047
rect 4801 10007 4859 10013
rect 4890 10004 4896 10056
rect 4948 10044 4954 10056
rect 9493 10047 9551 10053
rect 9493 10044 9505 10047
rect 4948 10016 9505 10044
rect 4948 10004 4954 10016
rect 4157 9979 4215 9985
rect 4157 9945 4169 9979
rect 4203 9976 4215 9979
rect 4203 9948 4844 9976
rect 4203 9945 4215 9948
rect 4157 9939 4215 9945
rect 2866 9868 2872 9920
rect 2924 9908 2930 9920
rect 3237 9911 3295 9917
rect 3237 9908 3249 9911
rect 2924 9880 3249 9908
rect 2924 9868 2930 9880
rect 3237 9877 3249 9880
rect 3283 9877 3295 9911
rect 3237 9871 3295 9877
rect 3329 9911 3387 9917
rect 3329 9877 3341 9911
rect 3375 9908 3387 9911
rect 3789 9911 3847 9917
rect 3789 9908 3801 9911
rect 3375 9880 3801 9908
rect 3375 9877 3387 9880
rect 3329 9871 3387 9877
rect 3789 9877 3801 9880
rect 3835 9877 3847 9911
rect 4706 9908 4712 9920
rect 4667 9880 4712 9908
rect 3789 9871 3847 9877
rect 4706 9868 4712 9880
rect 4764 9868 4770 9920
rect 4816 9908 4844 9948
rect 5810 9936 5816 9988
rect 5868 9976 5874 9988
rect 7098 9985 7104 9988
rect 6466 9979 6524 9985
rect 6466 9976 6478 9979
rect 5868 9948 6478 9976
rect 5868 9936 5874 9948
rect 6466 9945 6478 9948
rect 6512 9945 6524 9979
rect 7092 9976 7104 9985
rect 7059 9948 7104 9976
rect 6466 9939 6524 9945
rect 7092 9939 7104 9948
rect 7098 9936 7104 9939
rect 7156 9936 7162 9988
rect 6546 9908 6552 9920
rect 4816 9880 6552 9908
rect 6546 9868 6552 9880
rect 6604 9868 6610 9920
rect 8220 9917 8248 10016
rect 9493 10013 9505 10016
rect 9539 10013 9551 10047
rect 11514 10044 11520 10056
rect 9493 10007 9551 10013
rect 9968 10016 11520 10044
rect 9968 9985 9996 10016
rect 11514 10004 11520 10016
rect 11572 10044 11578 10056
rect 11609 10047 11667 10053
rect 11609 10044 11621 10047
rect 11572 10016 11621 10044
rect 11572 10004 11578 10016
rect 11609 10013 11621 10016
rect 11655 10044 11667 10047
rect 12894 10044 12900 10056
rect 11655 10016 12900 10044
rect 11655 10013 11667 10016
rect 11609 10007 11667 10013
rect 12894 10004 12900 10016
rect 12952 10044 12958 10056
rect 13081 10047 13139 10053
rect 13081 10044 13093 10047
rect 12952 10016 13093 10044
rect 12952 10004 12958 10016
rect 13081 10013 13093 10016
rect 13127 10044 13139 10047
rect 13633 10047 13691 10053
rect 13633 10044 13645 10047
rect 13127 10016 13645 10044
rect 13127 10013 13139 10016
rect 13081 10007 13139 10013
rect 13633 10013 13645 10016
rect 13679 10013 13691 10047
rect 13633 10007 13691 10013
rect 15309 10047 15367 10053
rect 15309 10013 15321 10047
rect 15355 10044 15367 10047
rect 17586 10044 17592 10056
rect 15355 10016 17592 10044
rect 15355 10013 15367 10016
rect 15309 10007 15367 10013
rect 17586 10004 17592 10016
rect 17644 10004 17650 10056
rect 18064 10053 18092 10084
rect 18230 10072 18236 10084
rect 18288 10112 18294 10124
rect 18877 10115 18935 10121
rect 18288 10084 18736 10112
rect 18288 10072 18294 10084
rect 17773 10047 17831 10053
rect 17773 10013 17785 10047
rect 17819 10013 17831 10047
rect 17773 10007 17831 10013
rect 18049 10047 18107 10053
rect 18049 10013 18061 10047
rect 18095 10013 18107 10047
rect 18601 10047 18659 10053
rect 18601 10044 18613 10047
rect 18049 10007 18107 10013
rect 18432 10016 18613 10044
rect 9953 9979 10011 9985
rect 9953 9976 9965 9979
rect 8496 9948 9965 9976
rect 8205 9911 8263 9917
rect 8205 9877 8217 9911
rect 8251 9877 8263 9911
rect 8386 9908 8392 9920
rect 8347 9880 8392 9908
rect 8205 9871 8263 9877
rect 8386 9868 8392 9880
rect 8444 9908 8450 9920
rect 8496 9917 8524 9948
rect 9953 9945 9965 9948
rect 9999 9945 10011 9979
rect 9953 9939 10011 9945
rect 10226 9936 10232 9988
rect 10284 9976 10290 9988
rect 11250 9979 11308 9985
rect 11250 9976 11262 9979
rect 10284 9948 11262 9976
rect 10284 9936 10290 9948
rect 11250 9945 11262 9948
rect 11296 9945 11308 9979
rect 11854 9979 11912 9985
rect 11854 9976 11866 9979
rect 11250 9939 11308 9945
rect 11348 9948 11866 9976
rect 11348 9920 11376 9948
rect 11854 9945 11866 9948
rect 11900 9945 11912 9979
rect 11854 9939 11912 9945
rect 15924 9979 15982 9985
rect 15924 9945 15936 9979
rect 15970 9976 15982 9979
rect 16390 9976 16396 9988
rect 15970 9948 16396 9976
rect 15970 9945 15982 9948
rect 15924 9939 15982 9945
rect 16390 9936 16396 9948
rect 16448 9936 16454 9988
rect 17788 9976 17816 10007
rect 18138 9976 18144 9988
rect 17788 9948 18144 9976
rect 18138 9936 18144 9948
rect 18196 9936 18202 9988
rect 8481 9911 8539 9917
rect 8481 9908 8493 9911
rect 8444 9880 8493 9908
rect 8444 9868 8450 9880
rect 8481 9877 8493 9880
rect 8527 9877 8539 9911
rect 8481 9871 8539 9877
rect 8570 9868 8576 9920
rect 8628 9908 8634 9920
rect 10137 9911 10195 9917
rect 10137 9908 10149 9911
rect 8628 9880 10149 9908
rect 8628 9868 8634 9880
rect 10137 9877 10149 9880
rect 10183 9877 10195 9911
rect 10137 9871 10195 9877
rect 11330 9868 11336 9920
rect 11388 9868 11394 9920
rect 12986 9908 12992 9920
rect 12947 9880 12992 9908
rect 12986 9868 12992 9880
rect 13044 9868 13050 9920
rect 14182 9908 14188 9920
rect 14095 9880 14188 9908
rect 14182 9868 14188 9880
rect 14240 9908 14246 9920
rect 17310 9908 17316 9920
rect 14240 9880 17316 9908
rect 14240 9868 14246 9880
rect 17310 9868 17316 9880
rect 17368 9868 17374 9920
rect 18046 9868 18052 9920
rect 18104 9908 18110 9920
rect 18233 9911 18291 9917
rect 18233 9908 18245 9911
rect 18104 9880 18245 9908
rect 18104 9868 18110 9880
rect 18233 9877 18245 9880
rect 18279 9877 18291 9911
rect 18432 9908 18460 10016
rect 18601 10013 18613 10016
rect 18647 10013 18659 10047
rect 18708 10044 18736 10084
rect 18877 10081 18889 10115
rect 18923 10112 18935 10115
rect 18966 10112 18972 10124
rect 18923 10084 18972 10112
rect 18923 10081 18935 10084
rect 18877 10075 18935 10081
rect 18966 10072 18972 10084
rect 19024 10072 19030 10124
rect 20640 10121 20668 10220
rect 20806 10208 20812 10260
rect 20864 10248 20870 10260
rect 21910 10248 21916 10260
rect 20864 10220 21916 10248
rect 20864 10208 20870 10220
rect 21910 10208 21916 10220
rect 21968 10208 21974 10260
rect 21726 10140 21732 10192
rect 21784 10180 21790 10192
rect 21784 10152 23152 10180
rect 21784 10140 21790 10152
rect 20625 10115 20683 10121
rect 20625 10081 20637 10115
rect 20671 10081 20683 10115
rect 21266 10112 21272 10124
rect 21227 10084 21272 10112
rect 20625 10075 20683 10081
rect 21266 10072 21272 10084
rect 21324 10072 21330 10124
rect 21542 10072 21548 10124
rect 21600 10112 21606 10124
rect 21913 10115 21971 10121
rect 21913 10112 21925 10115
rect 21600 10084 21925 10112
rect 21600 10072 21606 10084
rect 21913 10081 21925 10084
rect 21959 10081 21971 10115
rect 22186 10112 22192 10124
rect 22147 10084 22192 10112
rect 21913 10075 21971 10081
rect 22186 10072 22192 10084
rect 22244 10072 22250 10124
rect 22370 10112 22376 10124
rect 22331 10084 22376 10112
rect 22370 10072 22376 10084
rect 22428 10072 22434 10124
rect 19150 10044 19156 10056
rect 18708 10016 19156 10044
rect 18601 10007 18659 10013
rect 19150 10004 19156 10016
rect 19208 10004 19214 10056
rect 21082 10044 21088 10056
rect 20272 10016 21088 10044
rect 18509 9979 18567 9985
rect 18509 9945 18521 9979
rect 18555 9976 18567 9979
rect 20272 9976 20300 10016
rect 21082 10004 21088 10016
rect 21140 10004 21146 10056
rect 22002 10004 22008 10056
rect 22060 10044 22066 10056
rect 23124 10053 23152 10152
rect 22465 10047 22523 10053
rect 22465 10044 22477 10047
rect 22060 10016 22477 10044
rect 22060 10004 22066 10016
rect 22465 10013 22477 10016
rect 22511 10013 22523 10047
rect 22465 10007 22523 10013
rect 23109 10047 23167 10053
rect 23109 10013 23121 10047
rect 23155 10013 23167 10047
rect 23109 10007 23167 10013
rect 18555 9948 20300 9976
rect 20358 9979 20416 9985
rect 18555 9945 18567 9948
rect 18509 9939 18567 9945
rect 20358 9945 20370 9979
rect 20404 9945 20416 9979
rect 20358 9939 20416 9945
rect 18598 9908 18604 9920
rect 18432 9880 18604 9908
rect 18233 9871 18291 9877
rect 18598 9868 18604 9880
rect 18656 9868 18662 9920
rect 18690 9868 18696 9920
rect 18748 9908 18754 9920
rect 19245 9911 19303 9917
rect 19245 9908 19257 9911
rect 18748 9880 19257 9908
rect 18748 9868 18754 9880
rect 19245 9877 19257 9880
rect 19291 9877 19303 9911
rect 19245 9871 19303 9877
rect 20070 9868 20076 9920
rect 20128 9908 20134 9920
rect 20364 9908 20392 9939
rect 20990 9936 20996 9988
rect 21048 9976 21054 9988
rect 21545 9979 21603 9985
rect 21545 9976 21557 9979
rect 21048 9948 21557 9976
rect 21048 9936 21054 9948
rect 21545 9945 21557 9948
rect 21591 9945 21603 9979
rect 21545 9939 21603 9945
rect 21634 9936 21640 9988
rect 21692 9976 21698 9988
rect 21729 9979 21787 9985
rect 21729 9976 21741 9979
rect 21692 9948 21741 9976
rect 21692 9936 21698 9948
rect 21729 9945 21741 9948
rect 21775 9945 21787 9979
rect 21729 9939 21787 9945
rect 20714 9908 20720 9920
rect 20128 9880 20392 9908
rect 20675 9880 20720 9908
rect 20128 9868 20134 9880
rect 20714 9868 20720 9880
rect 20772 9868 20778 9920
rect 20806 9868 20812 9920
rect 20864 9908 20870 9920
rect 21085 9911 21143 9917
rect 21085 9908 21097 9911
rect 20864 9880 21097 9908
rect 20864 9868 20870 9880
rect 21085 9877 21097 9880
rect 21131 9877 21143 9911
rect 21085 9871 21143 9877
rect 21177 9911 21235 9917
rect 21177 9877 21189 9911
rect 21223 9908 21235 9911
rect 21450 9908 21456 9920
rect 21223 9880 21456 9908
rect 21223 9877 21235 9880
rect 21177 9871 21235 9877
rect 21450 9868 21456 9880
rect 21508 9868 21514 9920
rect 22830 9908 22836 9920
rect 22791 9880 22836 9908
rect 22830 9868 22836 9880
rect 22888 9868 22894 9920
rect 22922 9868 22928 9920
rect 22980 9908 22986 9920
rect 22980 9880 23025 9908
rect 22980 9868 22986 9880
rect 1104 9818 23460 9840
rect 1104 9766 6548 9818
rect 6600 9766 6612 9818
rect 6664 9766 6676 9818
rect 6728 9766 6740 9818
rect 6792 9766 6804 9818
rect 6856 9766 12146 9818
rect 12198 9766 12210 9818
rect 12262 9766 12274 9818
rect 12326 9766 12338 9818
rect 12390 9766 12402 9818
rect 12454 9766 17744 9818
rect 17796 9766 17808 9818
rect 17860 9766 17872 9818
rect 17924 9766 17936 9818
rect 17988 9766 18000 9818
rect 18052 9766 23460 9818
rect 1104 9744 23460 9766
rect 4522 9704 4528 9716
rect 2884 9676 4528 9704
rect 2884 9636 2912 9676
rect 4522 9664 4528 9676
rect 4580 9664 4586 9716
rect 4709 9707 4767 9713
rect 4709 9673 4721 9707
rect 4755 9673 4767 9707
rect 6362 9704 6368 9716
rect 6323 9676 6368 9704
rect 4709 9667 4767 9673
rect 2792 9608 2912 9636
rect 2961 9639 3019 9645
rect 1394 9568 1400 9580
rect 1355 9540 1400 9568
rect 1394 9528 1400 9540
rect 1452 9568 1458 9580
rect 1673 9571 1731 9577
rect 1673 9568 1685 9571
rect 1452 9540 1685 9568
rect 1452 9528 1458 9540
rect 1673 9537 1685 9540
rect 1719 9537 1731 9571
rect 1673 9531 1731 9537
rect 2792 9500 2820 9608
rect 2961 9605 2973 9639
rect 3007 9636 3019 9639
rect 4724 9636 4752 9667
rect 6362 9664 6368 9676
rect 6420 9704 6426 9716
rect 6638 9704 6644 9716
rect 6420 9676 6644 9704
rect 6420 9664 6426 9676
rect 6638 9664 6644 9676
rect 6696 9664 6702 9716
rect 11238 9704 11244 9716
rect 11164 9676 11244 9704
rect 6380 9636 6408 9664
rect 10505 9639 10563 9645
rect 10505 9636 10517 9639
rect 3007 9608 4752 9636
rect 3007 9605 3019 9608
rect 2961 9599 3019 9605
rect 2869 9571 2927 9577
rect 2869 9537 2881 9571
rect 2915 9568 2927 9571
rect 3142 9568 3148 9580
rect 2915 9540 3148 9568
rect 2915 9537 2927 9540
rect 2869 9531 2927 9537
rect 3142 9528 3148 9540
rect 3200 9528 3206 9580
rect 3585 9571 3643 9577
rect 3585 9568 3597 9571
rect 3252 9540 3597 9568
rect 3252 9512 3280 9540
rect 3585 9537 3597 9540
rect 3631 9537 3643 9571
rect 3585 9531 3643 9537
rect 3878 9528 3884 9580
rect 3936 9568 3942 9580
rect 3936 9540 4660 9568
rect 3936 9528 3942 9540
rect 3053 9503 3111 9509
rect 3053 9500 3065 9503
rect 2792 9472 3065 9500
rect 3053 9469 3065 9472
rect 3099 9469 3111 9503
rect 3053 9463 3111 9469
rect 3234 9460 3240 9512
rect 3292 9460 3298 9512
rect 3336 9503 3394 9509
rect 3336 9469 3348 9503
rect 3382 9469 3394 9503
rect 3336 9463 3394 9469
rect 1581 9435 1639 9441
rect 1581 9401 1593 9435
rect 1627 9432 1639 9435
rect 3142 9432 3148 9444
rect 1627 9404 3148 9432
rect 1627 9401 1639 9404
rect 1581 9395 1639 9401
rect 3142 9392 3148 9404
rect 3200 9392 3206 9444
rect 2406 9324 2412 9376
rect 2464 9364 2470 9376
rect 2501 9367 2559 9373
rect 2501 9364 2513 9367
rect 2464 9336 2513 9364
rect 2464 9324 2470 9336
rect 2501 9333 2513 9336
rect 2547 9333 2559 9367
rect 3344 9364 3372 9463
rect 4430 9364 4436 9376
rect 3344 9336 4436 9364
rect 2501 9327 2559 9333
rect 4430 9324 4436 9336
rect 4488 9324 4494 9376
rect 4632 9364 4660 9540
rect 4724 9500 4752 9608
rect 4816 9608 6408 9636
rect 9048 9608 10517 9636
rect 4816 9577 4844 9608
rect 4801 9571 4859 9577
rect 4801 9537 4813 9571
rect 4847 9537 4859 9571
rect 5057 9571 5115 9577
rect 5057 9568 5069 9571
rect 4801 9531 4859 9537
rect 4908 9540 5069 9568
rect 4908 9500 4936 9540
rect 5057 9537 5069 9540
rect 5103 9537 5115 9571
rect 5057 9531 5115 9537
rect 6638 9528 6644 9580
rect 6696 9568 6702 9580
rect 7561 9571 7619 9577
rect 7561 9568 7573 9571
rect 6696 9540 7573 9568
rect 6696 9528 6702 9540
rect 7561 9537 7573 9540
rect 7607 9537 7619 9571
rect 7561 9531 7619 9537
rect 7828 9571 7886 9577
rect 7828 9537 7840 9571
rect 7874 9568 7886 9571
rect 8846 9568 8852 9580
rect 7874 9540 8852 9568
rect 7874 9537 7886 9540
rect 7828 9531 7886 9537
rect 8846 9528 8852 9540
rect 8904 9528 8910 9580
rect 9048 9512 9076 9608
rect 10505 9605 10517 9608
rect 10551 9605 10563 9639
rect 10505 9599 10563 9605
rect 9300 9571 9358 9577
rect 9300 9537 9312 9571
rect 9346 9568 9358 9571
rect 10134 9568 10140 9580
rect 9346 9540 10140 9568
rect 9346 9537 9358 9540
rect 9300 9531 9358 9537
rect 10134 9528 10140 9540
rect 10192 9568 10198 9580
rect 11164 9568 11192 9676
rect 11238 9664 11244 9676
rect 11296 9664 11302 9716
rect 12618 9664 12624 9716
rect 12676 9704 12682 9716
rect 13630 9704 13636 9716
rect 12676 9676 13636 9704
rect 12676 9664 12682 9676
rect 13630 9664 13636 9676
rect 13688 9704 13694 9716
rect 13688 9676 14504 9704
rect 13688 9664 13694 9676
rect 12802 9636 12808 9648
rect 10192 9540 11192 9568
rect 11256 9608 12808 9636
rect 10192 9528 10198 9540
rect 6914 9500 6920 9512
rect 4724 9472 4936 9500
rect 6875 9472 6920 9500
rect 6914 9460 6920 9472
rect 6972 9460 6978 9512
rect 9030 9500 9036 9512
rect 8991 9472 9036 9500
rect 9030 9460 9036 9472
rect 9088 9460 9094 9512
rect 6181 9367 6239 9373
rect 6181 9364 6193 9367
rect 4632 9336 6193 9364
rect 6181 9333 6193 9336
rect 6227 9364 6239 9367
rect 7098 9364 7104 9376
rect 6227 9336 7104 9364
rect 6227 9333 6239 9336
rect 6181 9327 6239 9333
rect 7098 9324 7104 9336
rect 7156 9324 7162 9376
rect 7466 9364 7472 9376
rect 7427 9336 7472 9364
rect 7466 9324 7472 9336
rect 7524 9324 7530 9376
rect 8941 9367 8999 9373
rect 8941 9333 8953 9367
rect 8987 9364 8999 9367
rect 9214 9364 9220 9376
rect 8987 9336 9220 9364
rect 8987 9333 8999 9336
rect 8941 9327 8999 9333
rect 9214 9324 9220 9336
rect 9272 9324 9278 9376
rect 10226 9324 10232 9376
rect 10284 9364 10290 9376
rect 10413 9367 10471 9373
rect 10413 9364 10425 9367
rect 10284 9336 10425 9364
rect 10284 9324 10290 9336
rect 10413 9333 10425 9336
rect 10459 9333 10471 9367
rect 10686 9364 10692 9376
rect 10647 9336 10692 9364
rect 10413 9327 10471 9333
rect 10686 9324 10692 9336
rect 10744 9324 10750 9376
rect 10778 9324 10784 9376
rect 10836 9364 10842 9376
rect 11256 9364 11284 9608
rect 12802 9596 12808 9608
rect 12860 9596 12866 9648
rect 14476 9636 14504 9676
rect 17494 9664 17500 9716
rect 17552 9704 17558 9716
rect 18046 9704 18052 9716
rect 17552 9676 18052 9704
rect 17552 9664 17558 9676
rect 18046 9664 18052 9676
rect 18104 9664 18110 9716
rect 18690 9664 18696 9716
rect 18748 9704 18754 9716
rect 20990 9704 20996 9716
rect 18748 9676 20996 9704
rect 18748 9664 18754 9676
rect 20990 9664 20996 9676
rect 21048 9664 21054 9716
rect 21358 9704 21364 9716
rect 21319 9676 21364 9704
rect 21358 9664 21364 9676
rect 21416 9664 21422 9716
rect 22186 9664 22192 9716
rect 22244 9704 22250 9716
rect 22649 9707 22707 9713
rect 22649 9704 22661 9707
rect 22244 9676 22661 9704
rect 22244 9664 22250 9676
rect 22649 9673 22661 9676
rect 22695 9673 22707 9707
rect 22649 9667 22707 9673
rect 22830 9664 22836 9716
rect 22888 9664 22894 9716
rect 22281 9639 22339 9645
rect 12912 9608 14412 9636
rect 14476 9608 20668 9636
rect 12912 9580 12940 9608
rect 12618 9528 12624 9580
rect 12676 9577 12682 9580
rect 12676 9568 12688 9577
rect 12894 9568 12900 9580
rect 12676 9540 12721 9568
rect 12855 9540 12900 9568
rect 12676 9531 12688 9540
rect 12676 9528 12682 9531
rect 12894 9528 12900 9540
rect 12952 9528 12958 9580
rect 12986 9528 12992 9580
rect 13044 9568 13050 9580
rect 14384 9577 14412 9608
rect 15378 9577 15384 9580
rect 14102 9571 14160 9577
rect 14102 9568 14114 9571
rect 13044 9540 14114 9568
rect 13044 9528 13050 9540
rect 14102 9537 14114 9540
rect 14148 9537 14160 9571
rect 14102 9531 14160 9537
rect 14369 9571 14427 9577
rect 14369 9537 14381 9571
rect 14415 9568 14427 9571
rect 14461 9571 14519 9577
rect 14461 9568 14473 9571
rect 14415 9540 14473 9568
rect 14415 9537 14427 9540
rect 14369 9531 14427 9537
rect 14461 9537 14473 9540
rect 14507 9568 14519 9571
rect 15105 9571 15163 9577
rect 15105 9568 15117 9571
rect 14507 9540 15117 9568
rect 14507 9537 14519 9540
rect 14461 9531 14519 9537
rect 15105 9537 15117 9540
rect 15151 9537 15163 9571
rect 15372 9568 15384 9577
rect 15339 9540 15384 9568
rect 15105 9531 15163 9537
rect 15372 9531 15384 9540
rect 15378 9528 15384 9531
rect 15436 9528 15442 9580
rect 17129 9571 17187 9577
rect 17129 9537 17141 9571
rect 17175 9568 17187 9571
rect 18230 9568 18236 9580
rect 17175 9540 18236 9568
rect 17175 9537 17187 9540
rect 17129 9531 17187 9537
rect 18230 9528 18236 9540
rect 18288 9528 18294 9580
rect 18506 9528 18512 9580
rect 18564 9577 18570 9580
rect 18564 9568 18576 9577
rect 18564 9540 18609 9568
rect 18564 9531 18576 9540
rect 18564 9528 18570 9531
rect 18966 9528 18972 9580
rect 19024 9568 19030 9580
rect 19133 9571 19191 9577
rect 19133 9568 19145 9571
rect 19024 9540 19145 9568
rect 19024 9528 19030 9540
rect 19133 9537 19145 9540
rect 19179 9537 19191 9571
rect 19133 9531 19191 9537
rect 19426 9528 19432 9580
rect 19484 9568 19490 9580
rect 19484 9540 20576 9568
rect 19484 9528 19490 9540
rect 11333 9503 11391 9509
rect 11333 9469 11345 9503
rect 11379 9469 11391 9503
rect 18782 9500 18788 9512
rect 18743 9472 18788 9500
rect 11333 9463 11391 9469
rect 11348 9432 11376 9463
rect 18782 9460 18788 9472
rect 18840 9500 18846 9512
rect 18877 9503 18935 9509
rect 18877 9500 18889 9503
rect 18840 9472 18889 9500
rect 18840 9460 18846 9472
rect 18877 9469 18889 9472
rect 18923 9469 18935 9503
rect 18877 9463 18935 9469
rect 11348 9404 11836 9432
rect 11517 9367 11575 9373
rect 11517 9364 11529 9367
rect 10836 9336 11529 9364
rect 10836 9324 10842 9336
rect 11517 9333 11529 9336
rect 11563 9333 11575 9367
rect 11808 9364 11836 9404
rect 16298 9392 16304 9444
rect 16356 9432 16362 9444
rect 16669 9435 16727 9441
rect 16669 9432 16681 9435
rect 16356 9404 16681 9432
rect 16356 9392 16362 9404
rect 16669 9401 16681 9404
rect 16715 9432 16727 9435
rect 16853 9435 16911 9441
rect 16853 9432 16865 9435
rect 16715 9404 16865 9432
rect 16715 9401 16727 9404
rect 16669 9395 16727 9401
rect 16853 9401 16865 9404
rect 16899 9432 16911 9435
rect 17221 9435 17279 9441
rect 17221 9432 17233 9435
rect 16899 9404 17233 9432
rect 16899 9401 16911 9404
rect 16853 9395 16911 9401
rect 17221 9401 17233 9404
rect 17267 9401 17279 9435
rect 20548 9432 20576 9540
rect 20640 9509 20668 9608
rect 22281 9605 22293 9639
rect 22327 9636 22339 9639
rect 22848 9636 22876 9664
rect 22327 9608 23152 9636
rect 22327 9605 22339 9608
rect 22281 9599 22339 9605
rect 20714 9528 20720 9580
rect 20772 9568 20778 9580
rect 20809 9571 20867 9577
rect 20809 9568 20821 9571
rect 20772 9540 20821 9568
rect 20772 9528 20778 9540
rect 20809 9537 20821 9540
rect 20855 9537 20867 9571
rect 20809 9531 20867 9537
rect 20901 9571 20959 9577
rect 20901 9537 20913 9571
rect 20947 9537 20959 9571
rect 20901 9531 20959 9537
rect 21545 9571 21603 9577
rect 21545 9537 21557 9571
rect 21591 9568 21603 9571
rect 21591 9540 21864 9568
rect 21591 9537 21603 9540
rect 21545 9531 21603 9537
rect 20625 9503 20683 9509
rect 20625 9469 20637 9503
rect 20671 9469 20683 9503
rect 20916 9500 20944 9531
rect 21726 9500 21732 9512
rect 20916 9472 21732 9500
rect 20625 9463 20683 9469
rect 21726 9460 21732 9472
rect 21784 9460 21790 9512
rect 21836 9441 21864 9540
rect 22094 9528 22100 9580
rect 22152 9568 22158 9580
rect 22189 9571 22247 9577
rect 22189 9568 22201 9571
rect 22152 9540 22201 9568
rect 22152 9528 22158 9540
rect 22189 9537 22201 9540
rect 22235 9568 22247 9571
rect 22833 9571 22891 9577
rect 22235 9540 22324 9568
rect 22235 9537 22247 9540
rect 22189 9531 22247 9537
rect 21821 9435 21879 9441
rect 20548 9404 21404 9432
rect 17221 9395 17279 9401
rect 12618 9364 12624 9376
rect 11808 9336 12624 9364
rect 11517 9327 11575 9333
rect 12618 9324 12624 9336
rect 12676 9324 12682 9376
rect 12710 9324 12716 9376
rect 12768 9364 12774 9376
rect 12989 9367 13047 9373
rect 12989 9364 13001 9367
rect 12768 9336 13001 9364
rect 12768 9324 12774 9336
rect 12989 9333 13001 9336
rect 13035 9333 13047 9367
rect 12989 9327 13047 9333
rect 16485 9367 16543 9373
rect 16485 9333 16497 9367
rect 16531 9364 16543 9367
rect 16574 9364 16580 9376
rect 16531 9336 16580 9364
rect 16531 9333 16543 9336
rect 16485 9327 16543 9333
rect 16574 9324 16580 9336
rect 16632 9324 16638 9376
rect 17402 9364 17408 9376
rect 17315 9336 17408 9364
rect 17402 9324 17408 9336
rect 17460 9364 17466 9376
rect 20070 9364 20076 9376
rect 17460 9336 20076 9364
rect 17460 9324 17466 9336
rect 20070 9324 20076 9336
rect 20128 9324 20134 9376
rect 20162 9324 20168 9376
rect 20220 9364 20226 9376
rect 20257 9367 20315 9373
rect 20257 9364 20269 9367
rect 20220 9336 20269 9364
rect 20220 9324 20226 9336
rect 20257 9333 20269 9336
rect 20303 9333 20315 9367
rect 20438 9364 20444 9376
rect 20399 9336 20444 9364
rect 20257 9327 20315 9333
rect 20438 9324 20444 9336
rect 20496 9324 20502 9376
rect 21266 9364 21272 9376
rect 21227 9336 21272 9364
rect 21266 9324 21272 9336
rect 21324 9324 21330 9376
rect 21376 9364 21404 9404
rect 21821 9401 21833 9435
rect 21867 9401 21879 9435
rect 22296 9432 22324 9540
rect 22833 9537 22845 9571
rect 22879 9568 22891 9571
rect 23014 9568 23020 9580
rect 22879 9540 23020 9568
rect 22879 9537 22891 9540
rect 22833 9531 22891 9537
rect 23014 9528 23020 9540
rect 23072 9528 23078 9580
rect 23124 9577 23152 9608
rect 23109 9571 23167 9577
rect 23109 9537 23121 9571
rect 23155 9537 23167 9571
rect 23109 9531 23167 9537
rect 22465 9503 22523 9509
rect 22465 9469 22477 9503
rect 22511 9500 22523 9503
rect 22922 9500 22928 9512
rect 22511 9472 22928 9500
rect 22511 9469 22523 9472
rect 22465 9463 22523 9469
rect 22922 9460 22928 9472
rect 22980 9460 22986 9512
rect 23198 9432 23204 9444
rect 22296 9404 23204 9432
rect 21821 9395 21879 9401
rect 23198 9392 23204 9404
rect 23256 9392 23262 9444
rect 22186 9364 22192 9376
rect 21376 9336 22192 9364
rect 22186 9324 22192 9336
rect 22244 9324 22250 9376
rect 22278 9324 22284 9376
rect 22336 9364 22342 9376
rect 22925 9367 22983 9373
rect 22925 9364 22937 9367
rect 22336 9336 22937 9364
rect 22336 9324 22342 9336
rect 22925 9333 22937 9336
rect 22971 9333 22983 9367
rect 22925 9327 22983 9333
rect 1104 9274 23460 9296
rect 1104 9222 3749 9274
rect 3801 9222 3813 9274
rect 3865 9222 3877 9274
rect 3929 9222 3941 9274
rect 3993 9222 4005 9274
rect 4057 9222 9347 9274
rect 9399 9222 9411 9274
rect 9463 9222 9475 9274
rect 9527 9222 9539 9274
rect 9591 9222 9603 9274
rect 9655 9222 14945 9274
rect 14997 9222 15009 9274
rect 15061 9222 15073 9274
rect 15125 9222 15137 9274
rect 15189 9222 15201 9274
rect 15253 9222 20543 9274
rect 20595 9222 20607 9274
rect 20659 9222 20671 9274
rect 20723 9222 20735 9274
rect 20787 9222 20799 9274
rect 20851 9222 23460 9274
rect 1104 9200 23460 9222
rect 2774 9120 2780 9172
rect 2832 9160 2838 9172
rect 4706 9160 4712 9172
rect 2832 9132 2877 9160
rect 3620 9132 4712 9160
rect 2832 9120 2838 9132
rect 2866 9092 2872 9104
rect 2827 9064 2872 9092
rect 2866 9052 2872 9064
rect 2924 9052 2930 9104
rect 3142 9052 3148 9104
rect 3200 9092 3206 9104
rect 3510 9092 3516 9104
rect 3200 9064 3516 9092
rect 3200 9052 3206 9064
rect 3510 9052 3516 9064
rect 3568 9052 3574 9104
rect 2225 9027 2283 9033
rect 2225 8993 2237 9027
rect 2271 9024 2283 9027
rect 3050 9024 3056 9036
rect 2271 8996 3056 9024
rect 2271 8993 2283 8996
rect 2225 8987 2283 8993
rect 3050 8984 3056 8996
rect 3108 8984 3114 9036
rect 3234 8984 3240 9036
rect 3292 9024 3298 9036
rect 3421 9027 3479 9033
rect 3421 9024 3433 9027
rect 3292 8996 3433 9024
rect 3292 8984 3298 8996
rect 3421 8993 3433 8996
rect 3467 9024 3479 9027
rect 3620 9024 3648 9132
rect 4706 9120 4712 9132
rect 4764 9120 4770 9172
rect 5442 9160 5448 9172
rect 5403 9132 5448 9160
rect 5442 9120 5448 9132
rect 5500 9120 5506 9172
rect 6638 9120 6644 9172
rect 6696 9160 6702 9172
rect 7009 9163 7067 9169
rect 7009 9160 7021 9163
rect 6696 9132 7021 9160
rect 6696 9120 6702 9132
rect 6932 9033 6960 9132
rect 7009 9129 7021 9132
rect 7055 9160 7067 9163
rect 7193 9163 7251 9169
rect 7193 9160 7205 9163
rect 7055 9132 7205 9160
rect 7055 9129 7067 9132
rect 7009 9123 7067 9129
rect 7193 9129 7205 9132
rect 7239 9129 7251 9163
rect 7193 9123 7251 9129
rect 8386 9120 8392 9172
rect 8444 9160 8450 9172
rect 9030 9160 9036 9172
rect 8444 9132 9036 9160
rect 8444 9120 8450 9132
rect 9030 9120 9036 9132
rect 9088 9120 9094 9172
rect 12894 9120 12900 9172
rect 12952 9160 12958 9172
rect 13173 9163 13231 9169
rect 13173 9160 13185 9163
rect 12952 9132 13185 9160
rect 12952 9120 12958 9132
rect 3467 8996 3648 9024
rect 6917 9027 6975 9033
rect 3467 8993 3479 8996
rect 3421 8987 3479 8993
rect 6917 8993 6929 9027
rect 6963 9024 6975 9027
rect 7377 9027 7435 9033
rect 7377 9024 7389 9027
rect 6963 8996 7389 9024
rect 6963 8993 6975 8996
rect 6917 8987 6975 8993
rect 7377 8993 7389 8996
rect 7423 8993 7435 9027
rect 9048 9024 9076 9120
rect 13096 9033 13124 9132
rect 13173 9129 13185 9132
rect 13219 9160 13231 9163
rect 13357 9163 13415 9169
rect 13357 9160 13369 9163
rect 13219 9132 13369 9160
rect 13219 9129 13231 9132
rect 13173 9123 13231 9129
rect 13357 9129 13369 9132
rect 13403 9129 13415 9163
rect 13357 9123 13415 9129
rect 17586 9120 17592 9172
rect 17644 9160 17650 9172
rect 17644 9132 18276 9160
rect 17644 9120 17650 9132
rect 18248 9092 18276 9132
rect 18322 9120 18328 9172
rect 18380 9160 18386 9172
rect 19061 9163 19119 9169
rect 19061 9160 19073 9163
rect 18380 9132 19073 9160
rect 18380 9120 18386 9132
rect 19061 9129 19073 9132
rect 19107 9160 19119 9163
rect 19242 9160 19248 9172
rect 19107 9132 19248 9160
rect 19107 9129 19119 9132
rect 19061 9123 19119 9129
rect 19242 9120 19248 9132
rect 19300 9120 19306 9172
rect 21450 9160 21456 9172
rect 19720 9132 21312 9160
rect 21411 9132 21456 9160
rect 18874 9092 18880 9104
rect 18248 9064 18880 9092
rect 18874 9052 18880 9064
rect 18932 9052 18938 9104
rect 18966 9052 18972 9104
rect 19024 9092 19030 9104
rect 19720 9092 19748 9132
rect 19024 9064 19748 9092
rect 21284 9092 21312 9132
rect 21450 9120 21456 9132
rect 21508 9120 21514 9172
rect 21634 9120 21640 9172
rect 21692 9120 21698 9172
rect 22373 9163 22431 9169
rect 22373 9129 22385 9163
rect 22419 9160 22431 9163
rect 23566 9160 23572 9172
rect 22419 9132 23572 9160
rect 22419 9129 22431 9132
rect 22373 9123 22431 9129
rect 23566 9120 23572 9132
rect 23624 9160 23630 9172
rect 23842 9160 23848 9172
rect 23624 9132 23848 9160
rect 23624 9120 23630 9132
rect 23842 9120 23848 9132
rect 23900 9120 23906 9172
rect 21652 9092 21680 9120
rect 21284 9064 21680 9092
rect 19024 9052 19030 9064
rect 22186 9052 22192 9104
rect 22244 9092 22250 9104
rect 23658 9092 23664 9104
rect 22244 9064 23664 9092
rect 22244 9052 22250 9064
rect 23658 9052 23664 9064
rect 23716 9052 23722 9104
rect 10045 9027 10103 9033
rect 10045 9024 10057 9027
rect 9048 8996 10057 9024
rect 7377 8987 7435 8993
rect 10045 8993 10057 8996
rect 10091 8993 10103 9027
rect 10045 8987 10103 8993
rect 13081 9027 13139 9033
rect 13081 8993 13093 9027
rect 13127 8993 13139 9027
rect 13081 8987 13139 8993
rect 17773 9027 17831 9033
rect 17773 8993 17785 9027
rect 17819 9024 17831 9027
rect 18693 9027 18751 9033
rect 18693 9024 18705 9027
rect 17819 8996 18705 9024
rect 17819 8993 17831 8996
rect 17773 8987 17831 8993
rect 18693 8993 18705 8996
rect 18739 9024 18751 9027
rect 18782 9024 18788 9036
rect 18739 8996 18788 9024
rect 18739 8993 18751 8996
rect 18693 8987 18751 8993
rect 18782 8984 18788 8996
rect 18840 9024 18846 9036
rect 19150 9024 19156 9036
rect 18840 8996 19156 9024
rect 18840 8984 18846 8996
rect 19150 8984 19156 8996
rect 19208 8984 19214 9036
rect 20901 9027 20959 9033
rect 20901 8993 20913 9027
rect 20947 9024 20959 9027
rect 20990 9024 20996 9036
rect 20947 8996 20996 9024
rect 20947 8993 20959 8996
rect 20901 8987 20959 8993
rect 20990 8984 20996 8996
rect 21048 8984 21054 9036
rect 21637 9027 21695 9033
rect 21637 9024 21649 9027
rect 21192 8996 21649 9024
rect 2406 8956 2412 8968
rect 2367 8928 2412 8956
rect 2406 8916 2412 8928
rect 2464 8916 2470 8968
rect 4065 8959 4123 8965
rect 4065 8925 4077 8959
rect 4111 8956 4123 8959
rect 4111 8928 4476 8956
rect 4111 8925 4123 8928
rect 4065 8919 4123 8925
rect 4448 8900 4476 8928
rect 7466 8916 7472 8968
rect 7524 8956 7530 8968
rect 7633 8959 7691 8965
rect 7633 8956 7645 8959
rect 7524 8928 7645 8956
rect 7524 8916 7530 8928
rect 7633 8925 7645 8928
rect 7679 8925 7691 8959
rect 7633 8919 7691 8925
rect 9401 8959 9459 8965
rect 9401 8925 9413 8959
rect 9447 8956 9459 8959
rect 9766 8956 9772 8968
rect 9447 8928 9772 8956
rect 9447 8925 9459 8928
rect 9401 8919 9459 8925
rect 9766 8916 9772 8928
rect 9824 8916 9830 8968
rect 16298 8956 16304 8968
rect 16259 8928 16304 8956
rect 16298 8916 16304 8928
rect 16356 8916 16362 8968
rect 16390 8916 16396 8968
rect 16448 8956 16454 8968
rect 18049 8959 18107 8965
rect 16448 8928 17632 8956
rect 16448 8916 16454 8928
rect 2317 8891 2375 8897
rect 2317 8857 2329 8891
rect 2363 8888 2375 8891
rect 2866 8888 2872 8900
rect 2363 8860 2872 8888
rect 2363 8857 2375 8860
rect 2317 8851 2375 8857
rect 2866 8848 2872 8860
rect 2924 8848 2930 8900
rect 4338 8897 4344 8900
rect 3237 8891 3295 8897
rect 3237 8857 3249 8891
rect 3283 8888 3295 8891
rect 4332 8888 4344 8897
rect 3283 8860 4344 8888
rect 3283 8857 3295 8860
rect 3237 8851 3295 8857
rect 4332 8851 4344 8860
rect 4338 8848 4344 8851
rect 4396 8848 4402 8900
rect 4430 8848 4436 8900
rect 4488 8848 4494 8900
rect 6454 8848 6460 8900
rect 6512 8888 6518 8900
rect 6650 8891 6708 8897
rect 6650 8888 6662 8891
rect 6512 8860 6662 8888
rect 6512 8848 6518 8860
rect 6650 8857 6662 8860
rect 6696 8857 6708 8891
rect 6650 8851 6708 8857
rect 9953 8891 10011 8897
rect 9953 8857 9965 8891
rect 9999 8888 10011 8891
rect 10290 8891 10348 8897
rect 10290 8888 10302 8891
rect 9999 8860 10302 8888
rect 9999 8857 10011 8860
rect 9953 8851 10011 8857
rect 10290 8857 10302 8860
rect 10336 8857 10348 8891
rect 10290 8851 10348 8857
rect 12710 8848 12716 8900
rect 12768 8888 12774 8900
rect 12814 8891 12872 8897
rect 12814 8888 12826 8891
rect 12768 8860 12826 8888
rect 12768 8848 12774 8860
rect 12814 8857 12826 8860
rect 12860 8857 12872 8891
rect 12814 8851 12872 8857
rect 15930 8848 15936 8900
rect 15988 8888 15994 8900
rect 16034 8891 16092 8897
rect 16034 8888 16046 8891
rect 15988 8860 16046 8888
rect 15988 8848 15994 8860
rect 16034 8857 16046 8860
rect 16080 8857 16092 8891
rect 17494 8888 17500 8900
rect 17552 8897 17558 8900
rect 16034 8851 16092 8857
rect 16132 8860 16528 8888
rect 17464 8860 17500 8888
rect 3329 8823 3387 8829
rect 3329 8789 3341 8823
rect 3375 8820 3387 8823
rect 5534 8820 5540 8832
rect 3375 8792 5540 8820
rect 3375 8789 3387 8792
rect 3329 8783 3387 8789
rect 5534 8780 5540 8792
rect 5592 8780 5598 8832
rect 8757 8823 8815 8829
rect 8757 8789 8769 8823
rect 8803 8820 8815 8823
rect 8846 8820 8852 8832
rect 8803 8792 8852 8820
rect 8803 8789 8815 8792
rect 8757 8783 8815 8789
rect 8846 8780 8852 8792
rect 8904 8780 8910 8832
rect 11146 8780 11152 8832
rect 11204 8820 11210 8832
rect 11425 8823 11483 8829
rect 11425 8820 11437 8823
rect 11204 8792 11437 8820
rect 11204 8780 11210 8792
rect 11425 8789 11437 8792
rect 11471 8789 11483 8823
rect 11425 8783 11483 8789
rect 11514 8780 11520 8832
rect 11572 8820 11578 8832
rect 11701 8823 11759 8829
rect 11572 8792 11617 8820
rect 11572 8780 11578 8792
rect 11701 8789 11713 8823
rect 11747 8820 11759 8823
rect 12618 8820 12624 8832
rect 11747 8792 12624 8820
rect 11747 8789 11759 8792
rect 11701 8783 11759 8789
rect 12618 8780 12624 8792
rect 12676 8780 12682 8832
rect 14921 8823 14979 8829
rect 14921 8789 14933 8823
rect 14967 8820 14979 8823
rect 15378 8820 15384 8832
rect 14967 8792 15384 8820
rect 14967 8789 14979 8792
rect 14921 8783 14979 8789
rect 15378 8780 15384 8792
rect 15436 8820 15442 8832
rect 16132 8820 16160 8860
rect 16390 8820 16396 8832
rect 15436 8792 16160 8820
rect 16351 8792 16396 8820
rect 15436 8780 15442 8792
rect 16390 8780 16396 8792
rect 16448 8780 16454 8832
rect 16500 8820 16528 8860
rect 17494 8848 17500 8860
rect 17552 8851 17564 8897
rect 17604 8888 17632 8928
rect 18049 8925 18061 8959
rect 18095 8956 18107 8959
rect 18230 8956 18236 8968
rect 18095 8928 18236 8956
rect 18095 8925 18107 8928
rect 18049 8919 18107 8925
rect 18230 8916 18236 8928
rect 18288 8956 18294 8968
rect 18598 8956 18604 8968
rect 18288 8928 18604 8956
rect 18288 8916 18294 8928
rect 18598 8916 18604 8928
rect 18656 8956 18662 8968
rect 19334 8956 19340 8968
rect 18656 8928 19340 8956
rect 18656 8916 18662 8928
rect 19334 8916 19340 8928
rect 19392 8916 19398 8968
rect 19610 8916 19616 8968
rect 19668 8956 19674 8968
rect 20530 8956 20536 8968
rect 19668 8928 20536 8956
rect 19668 8916 19674 8928
rect 20530 8916 20536 8928
rect 20588 8956 20594 8968
rect 20625 8959 20683 8965
rect 20625 8956 20637 8959
rect 20588 8928 20637 8956
rect 20588 8916 20594 8928
rect 20625 8925 20637 8928
rect 20671 8925 20683 8959
rect 21082 8956 21088 8968
rect 21043 8928 21088 8956
rect 20625 8919 20683 8925
rect 21082 8916 21088 8928
rect 21140 8916 21146 8968
rect 17604 8860 20107 8888
rect 17552 8848 17558 8851
rect 18782 8820 18788 8832
rect 16500 8792 18788 8820
rect 18782 8780 18788 8792
rect 18840 8780 18846 8832
rect 19245 8823 19303 8829
rect 19245 8789 19257 8823
rect 19291 8820 19303 8823
rect 19978 8820 19984 8832
rect 19291 8792 19984 8820
rect 19291 8789 19303 8792
rect 19245 8783 19303 8789
rect 19978 8780 19984 8792
rect 20036 8780 20042 8832
rect 20079 8820 20107 8860
rect 20346 8848 20352 8900
rect 20404 8897 20410 8900
rect 20404 8888 20416 8897
rect 21192 8888 21220 8996
rect 21637 8993 21649 8996
rect 21683 8993 21695 9027
rect 21637 8987 21695 8993
rect 21818 8984 21824 9036
rect 21876 9024 21882 9036
rect 22925 9027 22983 9033
rect 22925 9024 22937 9027
rect 21876 8996 22937 9024
rect 21876 8984 21882 8996
rect 22925 8993 22937 8996
rect 22971 8993 22983 9027
rect 22925 8987 22983 8993
rect 21450 8916 21456 8968
rect 21508 8956 21514 8968
rect 21913 8959 21971 8965
rect 21913 8956 21925 8959
rect 21508 8928 21925 8956
rect 21508 8916 21514 8928
rect 21913 8925 21925 8928
rect 21959 8925 21971 8959
rect 22738 8956 22744 8968
rect 22699 8928 22744 8956
rect 21913 8919 21971 8925
rect 22738 8916 22744 8928
rect 22796 8916 22802 8968
rect 20404 8860 20449 8888
rect 20916 8860 21220 8888
rect 21821 8891 21879 8897
rect 20404 8851 20416 8860
rect 20404 8848 20410 8851
rect 20916 8820 20944 8860
rect 21821 8857 21833 8891
rect 21867 8888 21879 8891
rect 22186 8888 22192 8900
rect 21867 8860 22192 8888
rect 21867 8857 21879 8860
rect 21821 8851 21879 8857
rect 22186 8848 22192 8860
rect 22244 8848 22250 8900
rect 22833 8891 22891 8897
rect 22833 8888 22845 8891
rect 22296 8860 22845 8888
rect 20079 8792 20944 8820
rect 20993 8823 21051 8829
rect 20993 8789 21005 8823
rect 21039 8820 21051 8823
rect 21634 8820 21640 8832
rect 21039 8792 21640 8820
rect 21039 8789 21051 8792
rect 20993 8783 21051 8789
rect 21634 8780 21640 8792
rect 21692 8780 21698 8832
rect 22296 8829 22324 8860
rect 22833 8857 22845 8860
rect 22879 8857 22891 8891
rect 22833 8851 22891 8857
rect 22281 8823 22339 8829
rect 22281 8789 22293 8823
rect 22327 8789 22339 8823
rect 22281 8783 22339 8789
rect 1104 8730 23460 8752
rect 1104 8678 6548 8730
rect 6600 8678 6612 8730
rect 6664 8678 6676 8730
rect 6728 8678 6740 8730
rect 6792 8678 6804 8730
rect 6856 8678 12146 8730
rect 12198 8678 12210 8730
rect 12262 8678 12274 8730
rect 12326 8678 12338 8730
rect 12390 8678 12402 8730
rect 12454 8678 17744 8730
rect 17796 8678 17808 8730
rect 17860 8678 17872 8730
rect 17924 8678 17936 8730
rect 17988 8678 18000 8730
rect 18052 8678 23460 8730
rect 1104 8656 23460 8678
rect 1949 8619 2007 8625
rect 1949 8585 1961 8619
rect 1995 8616 2007 8619
rect 2501 8619 2559 8625
rect 2501 8616 2513 8619
rect 1995 8588 2513 8616
rect 1995 8585 2007 8588
rect 1949 8579 2007 8585
rect 2501 8585 2513 8588
rect 2547 8585 2559 8619
rect 3326 8616 3332 8628
rect 3287 8588 3332 8616
rect 2501 8579 2559 8585
rect 3326 8576 3332 8588
rect 3384 8576 3390 8628
rect 6178 8616 6184 8628
rect 4356 8588 6184 8616
rect 2958 8548 2964 8560
rect 2919 8520 2964 8548
rect 2958 8508 2964 8520
rect 3016 8508 3022 8560
rect 2038 8480 2044 8492
rect 1999 8452 2044 8480
rect 2038 8440 2044 8452
rect 2096 8440 2102 8492
rect 2869 8483 2927 8489
rect 2869 8449 2881 8483
rect 2915 8480 2927 8483
rect 4356 8480 4384 8588
rect 6178 8576 6184 8588
rect 6236 8576 6242 8628
rect 14277 8619 14335 8625
rect 14277 8585 14289 8619
rect 14323 8616 14335 8619
rect 15746 8616 15752 8628
rect 14323 8588 15752 8616
rect 14323 8585 14335 8588
rect 14277 8579 14335 8585
rect 15746 8576 15752 8588
rect 15804 8616 15810 8628
rect 16206 8616 16212 8628
rect 15804 8588 16212 8616
rect 15804 8576 15810 8588
rect 16206 8576 16212 8588
rect 16264 8576 16270 8628
rect 17497 8619 17555 8625
rect 17497 8585 17509 8619
rect 17543 8616 17555 8619
rect 18230 8616 18236 8628
rect 17543 8588 18236 8616
rect 17543 8585 17555 8588
rect 17497 8579 17555 8585
rect 18230 8576 18236 8588
rect 18288 8576 18294 8628
rect 19306 8588 20484 8616
rect 4798 8508 4804 8560
rect 4856 8508 4862 8560
rect 8144 8551 8202 8557
rect 8144 8517 8156 8551
rect 8190 8548 8202 8551
rect 8294 8548 8300 8560
rect 8190 8520 8300 8548
rect 8190 8517 8202 8520
rect 8144 8511 8202 8517
rect 8294 8508 8300 8520
rect 8352 8548 8358 8560
rect 8570 8548 8576 8560
rect 8352 8520 8576 8548
rect 8352 8508 8358 8520
rect 8570 8508 8576 8520
rect 8628 8508 8634 8560
rect 11514 8548 11520 8560
rect 9048 8520 11520 8548
rect 2915 8452 4384 8480
rect 4453 8483 4511 8489
rect 2915 8449 2927 8452
rect 2869 8443 2927 8449
rect 4453 8449 4465 8483
rect 4499 8480 4511 8483
rect 4816 8480 4844 8508
rect 4499 8452 4844 8480
rect 4499 8449 4511 8452
rect 4453 8443 4511 8449
rect 4890 8440 4896 8492
rect 4948 8480 4954 8492
rect 5057 8483 5115 8489
rect 5057 8480 5069 8483
rect 4948 8452 5069 8480
rect 4948 8440 4954 8452
rect 5057 8449 5069 8452
rect 5103 8480 5115 8483
rect 5810 8480 5816 8492
rect 5103 8452 5816 8480
rect 5103 8449 5115 8452
rect 5057 8443 5115 8449
rect 5810 8440 5816 8452
rect 5868 8440 5874 8492
rect 9048 8480 9076 8520
rect 6840 8452 9076 8480
rect 1857 8415 1915 8421
rect 1857 8381 1869 8415
rect 1903 8412 1915 8415
rect 3050 8412 3056 8424
rect 1903 8384 3056 8412
rect 1903 8381 1915 8384
rect 1857 8375 1915 8381
rect 3050 8372 3056 8384
rect 3108 8372 3114 8424
rect 3145 8415 3203 8421
rect 3145 8381 3157 8415
rect 3191 8412 3203 8415
rect 3234 8412 3240 8424
rect 3191 8384 3240 8412
rect 3191 8381 3203 8384
rect 3145 8375 3203 8381
rect 3234 8372 3240 8384
rect 3292 8372 3298 8424
rect 4709 8415 4767 8421
rect 4709 8381 4721 8415
rect 4755 8412 4767 8415
rect 4801 8415 4859 8421
rect 4801 8412 4813 8415
rect 4755 8384 4813 8412
rect 4755 8381 4767 8384
rect 4709 8375 4767 8381
rect 4801 8381 4813 8384
rect 4847 8381 4859 8415
rect 4801 8375 4859 8381
rect 2314 8304 2320 8356
rect 2372 8344 2378 8356
rect 2409 8347 2467 8353
rect 2409 8344 2421 8347
rect 2372 8316 2421 8344
rect 2372 8304 2378 8316
rect 2409 8313 2421 8316
rect 2455 8313 2467 8347
rect 2409 8307 2467 8313
rect 4430 8236 4436 8288
rect 4488 8276 4494 8288
rect 4724 8276 4752 8375
rect 5994 8304 6000 8356
rect 6052 8344 6058 8356
rect 6840 8353 6868 8452
rect 8404 8424 8432 8452
rect 9122 8440 9128 8492
rect 9180 8480 9186 8492
rect 9876 8489 9904 8520
rect 11514 8508 11520 8520
rect 11572 8548 11578 8560
rect 11572 8520 13216 8548
rect 11572 8508 11578 8520
rect 9594 8483 9652 8489
rect 9594 8480 9606 8483
rect 9180 8452 9606 8480
rect 9180 8440 9186 8452
rect 9594 8449 9606 8452
rect 9640 8449 9652 8483
rect 9594 8443 9652 8449
rect 9861 8483 9919 8489
rect 9861 8449 9873 8483
rect 9907 8480 9919 8483
rect 9953 8483 10011 8489
rect 9953 8480 9965 8483
rect 9907 8452 9965 8480
rect 9907 8449 9919 8452
rect 9861 8443 9919 8449
rect 9953 8449 9965 8452
rect 9999 8449 10011 8483
rect 9953 8443 10011 8449
rect 10220 8483 10278 8489
rect 10220 8449 10232 8483
rect 10266 8480 10278 8483
rect 10686 8480 10692 8492
rect 10266 8452 10692 8480
rect 10266 8449 10278 8452
rect 10220 8443 10278 8449
rect 10686 8440 10692 8452
rect 10744 8440 10750 8492
rect 12526 8440 12532 8492
rect 12584 8480 12590 8492
rect 13188 8489 13216 8520
rect 18138 8508 18144 8560
rect 18196 8548 18202 8560
rect 19306 8548 19334 8588
rect 19518 8557 19524 8560
rect 19512 8548 19524 8557
rect 18196 8520 19334 8548
rect 19479 8520 19524 8548
rect 18196 8508 18202 8520
rect 19512 8511 19524 8520
rect 19518 8508 19524 8511
rect 19576 8508 19582 8560
rect 20456 8548 20484 8588
rect 20530 8576 20536 8628
rect 20588 8616 20594 8628
rect 21545 8619 21603 8625
rect 21545 8616 21557 8619
rect 20588 8588 21557 8616
rect 20588 8576 20594 8588
rect 21545 8585 21557 8588
rect 21591 8585 21603 8619
rect 21545 8579 21603 8585
rect 21726 8576 21732 8628
rect 21784 8616 21790 8628
rect 21821 8619 21879 8625
rect 21821 8616 21833 8619
rect 21784 8588 21833 8616
rect 21784 8576 21790 8588
rect 21821 8585 21833 8588
rect 21867 8585 21879 8619
rect 21821 8579 21879 8585
rect 22373 8551 22431 8557
rect 22373 8548 22385 8551
rect 20456 8520 22385 8548
rect 22373 8517 22385 8520
rect 22419 8517 22431 8551
rect 22373 8511 22431 8517
rect 22462 8508 22468 8560
rect 22520 8548 22526 8560
rect 22925 8551 22983 8557
rect 22925 8548 22937 8551
rect 22520 8520 22937 8548
rect 22520 8508 22526 8520
rect 22925 8517 22937 8520
rect 22971 8517 22983 8551
rect 22925 8511 22983 8517
rect 12906 8483 12964 8489
rect 12906 8480 12918 8483
rect 12584 8452 12918 8480
rect 12584 8440 12590 8452
rect 12906 8449 12918 8452
rect 12952 8449 12964 8483
rect 12906 8443 12964 8449
rect 13173 8483 13231 8489
rect 13173 8449 13185 8483
rect 13219 8480 13231 8483
rect 13265 8483 13323 8489
rect 13265 8480 13277 8483
rect 13219 8452 13277 8480
rect 13219 8449 13231 8452
rect 13173 8443 13231 8449
rect 13265 8449 13277 8452
rect 13311 8449 13323 8483
rect 13265 8443 13323 8449
rect 15401 8483 15459 8489
rect 15401 8449 15413 8483
rect 15447 8480 15459 8483
rect 16482 8480 16488 8492
rect 15447 8452 16488 8480
rect 15447 8449 15459 8452
rect 15401 8443 15459 8449
rect 16482 8440 16488 8452
rect 16540 8440 16546 8492
rect 16574 8440 16580 8492
rect 16632 8480 16638 8492
rect 18322 8480 18328 8492
rect 16632 8452 18328 8480
rect 16632 8440 16638 8452
rect 18322 8440 18328 8452
rect 18380 8440 18386 8492
rect 18897 8483 18955 8489
rect 18897 8449 18909 8483
rect 18943 8480 18955 8483
rect 19058 8480 19064 8492
rect 18943 8452 19064 8480
rect 18943 8449 18955 8452
rect 18897 8443 18955 8449
rect 19058 8440 19064 8452
rect 19116 8440 19122 8492
rect 20438 8440 20444 8492
rect 20496 8480 20502 8492
rect 20898 8480 20904 8492
rect 20496 8452 20904 8480
rect 20496 8440 20502 8452
rect 20898 8440 20904 8452
rect 20956 8440 20962 8492
rect 21082 8480 21088 8492
rect 21043 8452 21088 8480
rect 21082 8440 21088 8452
rect 21140 8440 21146 8492
rect 21174 8440 21180 8492
rect 21232 8480 21238 8492
rect 21232 8452 21277 8480
rect 21232 8440 21238 8452
rect 21726 8440 21732 8492
rect 21784 8480 21790 8492
rect 22646 8480 22652 8492
rect 21784 8452 22094 8480
rect 22607 8452 22652 8480
rect 21784 8440 21790 8452
rect 8386 8372 8392 8424
rect 8444 8412 8450 8424
rect 15657 8415 15715 8421
rect 8444 8384 8537 8412
rect 8444 8372 8450 8384
rect 15657 8381 15669 8415
rect 15703 8381 15715 8415
rect 15657 8375 15715 8381
rect 6365 8347 6423 8353
rect 6365 8344 6377 8347
rect 6052 8316 6377 8344
rect 6052 8304 6058 8316
rect 6365 8313 6377 8316
rect 6411 8344 6423 8347
rect 6549 8347 6607 8353
rect 6549 8344 6561 8347
rect 6411 8316 6561 8344
rect 6411 8313 6423 8316
rect 6365 8307 6423 8313
rect 6549 8313 6561 8316
rect 6595 8344 6607 8347
rect 6825 8347 6883 8353
rect 6825 8344 6837 8347
rect 6595 8316 6837 8344
rect 6595 8313 6607 8316
rect 6549 8307 6607 8313
rect 6825 8313 6837 8316
rect 6871 8313 6883 8347
rect 6825 8307 6883 8313
rect 11793 8347 11851 8353
rect 11793 8313 11805 8347
rect 11839 8344 11851 8347
rect 12066 8344 12072 8356
rect 11839 8316 12072 8344
rect 11839 8313 11851 8316
rect 11793 8307 11851 8313
rect 12066 8304 12072 8316
rect 12124 8304 12130 8356
rect 15672 8344 15700 8375
rect 19150 8372 19156 8424
rect 19208 8412 19214 8424
rect 19245 8415 19303 8421
rect 19245 8412 19257 8415
rect 19208 8384 19257 8412
rect 19208 8372 19214 8384
rect 19245 8381 19257 8384
rect 19291 8381 19303 8415
rect 19245 8375 19303 8381
rect 15841 8347 15899 8353
rect 15841 8344 15853 8347
rect 15672 8316 15853 8344
rect 15841 8313 15853 8316
rect 15887 8344 15899 8347
rect 16022 8344 16028 8356
rect 15887 8316 16028 8344
rect 15887 8313 15899 8316
rect 15841 8307 15899 8313
rect 16022 8304 16028 8316
rect 16080 8344 16086 8356
rect 16298 8344 16304 8356
rect 16080 8316 16304 8344
rect 16080 8304 16086 8316
rect 16298 8304 16304 8316
rect 16356 8344 16362 8356
rect 16485 8347 16543 8353
rect 16485 8344 16497 8347
rect 16356 8316 16497 8344
rect 16356 8304 16362 8316
rect 16485 8313 16497 8316
rect 16531 8344 16543 8347
rect 16761 8347 16819 8353
rect 16761 8344 16773 8347
rect 16531 8316 16773 8344
rect 16531 8313 16543 8316
rect 16485 8307 16543 8313
rect 16761 8313 16773 8316
rect 16807 8344 16819 8347
rect 16945 8347 17003 8353
rect 16945 8344 16957 8347
rect 16807 8316 16957 8344
rect 16807 8313 16819 8316
rect 16761 8307 16819 8313
rect 16945 8313 16957 8316
rect 16991 8344 17003 8347
rect 17129 8347 17187 8353
rect 17129 8344 17141 8347
rect 16991 8316 17141 8344
rect 16991 8313 17003 8316
rect 16945 8307 17003 8313
rect 17129 8313 17141 8316
rect 17175 8344 17187 8347
rect 17313 8347 17371 8353
rect 17313 8344 17325 8347
rect 17175 8316 17325 8344
rect 17175 8313 17187 8316
rect 17129 8307 17187 8313
rect 17313 8313 17325 8316
rect 17359 8344 17371 8347
rect 17681 8347 17739 8353
rect 17681 8344 17693 8347
rect 17359 8316 17693 8344
rect 17359 8313 17371 8316
rect 17313 8307 17371 8313
rect 17681 8313 17693 8316
rect 17727 8344 17739 8347
rect 17727 8316 18000 8344
rect 17727 8313 17739 8316
rect 17681 8307 17739 8313
rect 7006 8276 7012 8288
rect 4488 8248 4752 8276
rect 6967 8248 7012 8276
rect 4488 8236 4494 8248
rect 7006 8236 7012 8248
rect 7064 8236 7070 8288
rect 8481 8279 8539 8285
rect 8481 8245 8493 8279
rect 8527 8276 8539 8279
rect 8662 8276 8668 8288
rect 8527 8248 8668 8276
rect 8527 8245 8539 8248
rect 8481 8239 8539 8245
rect 8662 8236 8668 8248
rect 8720 8236 8726 8288
rect 11333 8279 11391 8285
rect 11333 8245 11345 8279
rect 11379 8276 11391 8279
rect 11514 8276 11520 8288
rect 11379 8248 11520 8276
rect 11379 8245 11391 8248
rect 11333 8239 11391 8245
rect 11514 8236 11520 8248
rect 11572 8236 11578 8288
rect 11882 8236 11888 8288
rect 11940 8276 11946 8288
rect 16390 8276 16396 8288
rect 11940 8248 16396 8276
rect 11940 8236 11946 8248
rect 16390 8236 16396 8248
rect 16448 8236 16454 8288
rect 17586 8236 17592 8288
rect 17644 8276 17650 8288
rect 17773 8279 17831 8285
rect 17773 8276 17785 8279
rect 17644 8248 17785 8276
rect 17644 8236 17650 8248
rect 17773 8245 17785 8248
rect 17819 8245 17831 8279
rect 17972 8276 18000 8316
rect 19260 8276 19288 8375
rect 20806 8372 20812 8424
rect 20864 8412 20870 8424
rect 21269 8415 21327 8421
rect 21269 8412 21281 8415
rect 20864 8384 21281 8412
rect 20864 8372 20870 8384
rect 21269 8381 21281 8384
rect 21315 8381 21327 8415
rect 22066 8412 22094 8452
rect 22646 8440 22652 8452
rect 22704 8440 22710 8492
rect 22554 8412 22560 8424
rect 22066 8384 22560 8412
rect 21269 8375 21327 8381
rect 22554 8372 22560 8384
rect 22612 8372 22618 8424
rect 20717 8347 20775 8353
rect 20717 8313 20729 8347
rect 20763 8344 20775 8347
rect 20990 8344 20996 8356
rect 20763 8316 20996 8344
rect 20763 8313 20775 8316
rect 20717 8307 20775 8313
rect 20990 8304 20996 8316
rect 21048 8304 21054 8356
rect 22462 8304 22468 8356
rect 22520 8344 22526 8356
rect 22741 8347 22799 8353
rect 22741 8344 22753 8347
rect 22520 8316 22753 8344
rect 22520 8304 22526 8316
rect 22741 8313 22753 8316
rect 22787 8313 22799 8347
rect 22741 8307 22799 8313
rect 19610 8276 19616 8288
rect 17972 8248 19616 8276
rect 17773 8239 17831 8245
rect 19610 8236 19616 8248
rect 19668 8236 19674 8288
rect 20438 8236 20444 8288
rect 20496 8276 20502 8288
rect 20625 8279 20683 8285
rect 20625 8276 20637 8279
rect 20496 8248 20637 8276
rect 20496 8236 20502 8248
rect 20625 8245 20637 8248
rect 20671 8245 20683 8279
rect 20625 8239 20683 8245
rect 20806 8236 20812 8288
rect 20864 8276 20870 8288
rect 22554 8276 22560 8288
rect 20864 8248 22560 8276
rect 20864 8236 20870 8248
rect 22554 8236 22560 8248
rect 22612 8236 22618 8288
rect 1104 8186 23460 8208
rect 1104 8134 3749 8186
rect 3801 8134 3813 8186
rect 3865 8134 3877 8186
rect 3929 8134 3941 8186
rect 3993 8134 4005 8186
rect 4057 8134 9347 8186
rect 9399 8134 9411 8186
rect 9463 8134 9475 8186
rect 9527 8134 9539 8186
rect 9591 8134 9603 8186
rect 9655 8134 14945 8186
rect 14997 8134 15009 8186
rect 15061 8134 15073 8186
rect 15125 8134 15137 8186
rect 15189 8134 15201 8186
rect 15253 8134 20543 8186
rect 20595 8134 20607 8186
rect 20659 8134 20671 8186
rect 20723 8134 20735 8186
rect 20787 8134 20799 8186
rect 20851 8134 23460 8186
rect 1104 8112 23460 8134
rect 2038 8072 2044 8084
rect 1999 8044 2044 8072
rect 2038 8032 2044 8044
rect 2096 8032 2102 8084
rect 2866 8072 2872 8084
rect 2827 8044 2872 8072
rect 2866 8032 2872 8044
rect 2924 8032 2930 8084
rect 5810 8072 5816 8084
rect 5771 8044 5816 8072
rect 5810 8032 5816 8044
rect 5868 8032 5874 8084
rect 6914 8032 6920 8084
rect 6972 8072 6978 8084
rect 7377 8075 7435 8081
rect 7377 8072 7389 8075
rect 6972 8044 7389 8072
rect 6972 8032 6978 8044
rect 7377 8041 7389 8044
rect 7423 8072 7435 8075
rect 7466 8072 7472 8084
rect 7423 8044 7472 8072
rect 7423 8041 7435 8044
rect 7377 8035 7435 8041
rect 7466 8032 7472 8044
rect 7524 8032 7530 8084
rect 11238 8032 11244 8084
rect 11296 8072 11302 8084
rect 18601 8075 18659 8081
rect 18601 8072 18613 8075
rect 11296 8044 18613 8072
rect 11296 8032 11302 8044
rect 18601 8041 18613 8044
rect 18647 8041 18659 8075
rect 22830 8072 22836 8084
rect 18601 8035 18659 8041
rect 19536 8044 22836 8072
rect 18417 8007 18475 8013
rect 18417 8004 18429 8007
rect 18064 7976 18429 8004
rect 2685 7939 2743 7945
rect 2685 7905 2697 7939
rect 2731 7936 2743 7939
rect 3234 7936 3240 7948
rect 2731 7908 3240 7936
rect 2731 7905 2743 7908
rect 2685 7899 2743 7905
rect 3234 7896 3240 7908
rect 3292 7936 3298 7948
rect 3421 7939 3479 7945
rect 3421 7936 3433 7939
rect 3292 7908 3433 7936
rect 3292 7896 3298 7908
rect 3421 7905 3433 7908
rect 3467 7905 3479 7939
rect 3421 7899 3479 7905
rect 2501 7871 2559 7877
rect 2501 7837 2513 7871
rect 2547 7868 2559 7871
rect 3142 7868 3148 7880
rect 2547 7840 3148 7868
rect 2547 7837 2559 7840
rect 2501 7831 2559 7837
rect 3142 7828 3148 7840
rect 3200 7828 3206 7880
rect 3326 7828 3332 7880
rect 3384 7868 3390 7880
rect 4430 7868 4436 7880
rect 3384 7840 4436 7868
rect 3384 7828 3390 7840
rect 4430 7828 4436 7840
rect 4488 7868 4494 7880
rect 5905 7871 5963 7877
rect 5905 7868 5917 7871
rect 4488 7840 5917 7868
rect 4488 7828 4494 7840
rect 5905 7837 5917 7840
rect 5951 7868 5963 7871
rect 5994 7868 6000 7880
rect 5951 7840 6000 7868
rect 5951 7837 5963 7840
rect 5905 7831 5963 7837
rect 5994 7828 6000 7840
rect 6052 7828 6058 7880
rect 8757 7871 8815 7877
rect 8757 7868 8769 7871
rect 8404 7840 8769 7868
rect 8404 7812 8432 7840
rect 8757 7837 8769 7840
rect 8803 7868 8815 7871
rect 8941 7871 8999 7877
rect 8941 7868 8953 7871
rect 8803 7840 8953 7868
rect 8803 7837 8815 7840
rect 8757 7831 8815 7837
rect 8941 7837 8953 7840
rect 8987 7868 8999 7871
rect 9125 7871 9183 7877
rect 9125 7868 9137 7871
rect 8987 7840 9137 7868
rect 8987 7837 8999 7840
rect 8941 7831 8999 7837
rect 9125 7837 9137 7840
rect 9171 7868 9183 7871
rect 9309 7871 9367 7877
rect 9309 7868 9321 7871
rect 9171 7840 9321 7868
rect 9171 7837 9183 7840
rect 9125 7831 9183 7837
rect 9309 7837 9321 7840
rect 9355 7868 9367 7871
rect 9493 7871 9551 7877
rect 9493 7868 9505 7871
rect 9355 7840 9505 7868
rect 9355 7837 9367 7840
rect 9309 7831 9367 7837
rect 9493 7837 9505 7840
rect 9539 7868 9551 7871
rect 10686 7868 10692 7880
rect 9539 7840 10692 7868
rect 9539 7837 9551 7840
rect 9493 7831 9551 7837
rect 10686 7828 10692 7840
rect 10744 7868 10750 7880
rect 10965 7871 11023 7877
rect 10965 7868 10977 7871
rect 10744 7840 10977 7868
rect 10744 7828 10750 7840
rect 10965 7837 10977 7840
rect 11011 7868 11023 7871
rect 12437 7871 12495 7877
rect 12437 7868 12449 7871
rect 11011 7840 12449 7868
rect 11011 7837 11023 7840
rect 10965 7831 11023 7837
rect 12437 7837 12449 7840
rect 12483 7868 12495 7871
rect 14093 7871 14151 7877
rect 14093 7868 14105 7871
rect 12483 7840 14105 7868
rect 12483 7837 12495 7840
rect 12437 7831 12495 7837
rect 14093 7837 14105 7840
rect 14139 7868 14151 7871
rect 15565 7871 15623 7877
rect 15565 7868 15577 7871
rect 14139 7840 15577 7868
rect 14139 7837 14151 7840
rect 14093 7831 14151 7837
rect 15565 7837 15577 7840
rect 15611 7868 15623 7871
rect 16298 7868 16304 7880
rect 15611 7840 16304 7868
rect 15611 7837 15623 7840
rect 15565 7831 15623 7837
rect 16298 7828 16304 7840
rect 16356 7868 16362 7880
rect 17037 7871 17095 7877
rect 17037 7868 17049 7871
rect 16356 7840 17049 7868
rect 16356 7828 16362 7840
rect 17037 7837 17049 7840
rect 17083 7837 17095 7871
rect 18064 7868 18092 7976
rect 18417 7973 18429 7976
rect 18463 8004 18475 8007
rect 19536 8004 19564 8044
rect 22830 8032 22836 8044
rect 22888 8032 22894 8084
rect 18463 7976 19564 8004
rect 18463 7973 18475 7976
rect 18417 7967 18475 7973
rect 22186 7964 22192 8016
rect 22244 8004 22250 8016
rect 22557 8007 22615 8013
rect 22557 8004 22569 8007
rect 22244 7976 22569 8004
rect 22244 7964 22250 7976
rect 22557 7973 22569 7976
rect 22603 8004 22615 8007
rect 23290 8004 23296 8016
rect 22603 7976 23296 8004
rect 22603 7973 22615 7976
rect 22557 7967 22615 7973
rect 23290 7964 23296 7976
rect 23348 7964 23354 8016
rect 21180 7939 21238 7945
rect 21180 7905 21192 7939
rect 21226 7936 21238 7939
rect 21266 7936 21272 7948
rect 21226 7908 21272 7936
rect 21226 7905 21238 7908
rect 21180 7899 21238 7905
rect 21266 7896 21272 7908
rect 21324 7896 21330 7948
rect 21453 7939 21511 7945
rect 21453 7905 21465 7939
rect 21499 7936 21511 7939
rect 21910 7936 21916 7948
rect 21499 7908 21916 7936
rect 21499 7905 21511 7908
rect 21453 7899 21511 7905
rect 21910 7896 21916 7908
rect 21968 7896 21974 7948
rect 17037 7831 17095 7837
rect 17420 7840 18092 7868
rect 17420 7812 17448 7840
rect 18414 7828 18420 7880
rect 18472 7868 18478 7880
rect 18785 7871 18843 7877
rect 18785 7868 18797 7871
rect 18472 7840 18797 7868
rect 18472 7828 18478 7840
rect 18785 7837 18797 7840
rect 18831 7837 18843 7871
rect 18785 7831 18843 7837
rect 18877 7871 18935 7877
rect 18877 7837 18889 7871
rect 18923 7868 18935 7871
rect 19886 7868 19892 7880
rect 18923 7840 19892 7868
rect 18923 7837 18935 7840
rect 18877 7831 18935 7837
rect 19886 7828 19892 7840
rect 19944 7828 19950 7880
rect 20622 7868 20628 7880
rect 20583 7840 20628 7868
rect 20622 7828 20628 7840
rect 20680 7828 20686 7880
rect 20717 7871 20775 7877
rect 20717 7837 20729 7871
rect 20763 7868 20775 7871
rect 21542 7868 21548 7880
rect 20763 7840 21548 7868
rect 20763 7837 20775 7840
rect 20717 7831 20775 7837
rect 21542 7828 21548 7840
rect 21600 7828 21606 7880
rect 21818 7828 21824 7880
rect 21876 7868 21882 7880
rect 23014 7868 23020 7880
rect 21876 7840 23020 7868
rect 21876 7828 21882 7840
rect 23014 7828 23020 7840
rect 23072 7828 23078 7880
rect 3237 7803 3295 7809
rect 3237 7769 3249 7803
rect 3283 7800 3295 7803
rect 3418 7800 3424 7812
rect 3283 7772 3424 7800
rect 3283 7769 3295 7772
rect 3237 7763 3295 7769
rect 3418 7760 3424 7772
rect 3476 7760 3482 7812
rect 3510 7760 3516 7812
rect 3568 7800 3574 7812
rect 4678 7803 4736 7809
rect 4678 7800 4690 7803
rect 3568 7772 4690 7800
rect 3568 7760 3574 7772
rect 4678 7769 4690 7772
rect 4724 7769 4736 7803
rect 4678 7763 4736 7769
rect 6172 7803 6230 7809
rect 6172 7769 6184 7803
rect 6218 7800 6230 7803
rect 7190 7800 7196 7812
rect 6218 7772 7196 7800
rect 6218 7769 6230 7772
rect 6172 7763 6230 7769
rect 7190 7760 7196 7772
rect 7248 7760 7254 7812
rect 7558 7800 7564 7812
rect 7300 7772 7564 7800
rect 2406 7732 2412 7744
rect 2367 7704 2412 7732
rect 2406 7692 2412 7704
rect 2464 7692 2470 7744
rect 3329 7735 3387 7741
rect 3329 7701 3341 7735
rect 3375 7732 3387 7735
rect 4798 7732 4804 7744
rect 3375 7704 4804 7732
rect 3375 7701 3387 7704
rect 3329 7695 3387 7701
rect 4798 7692 4804 7704
rect 4856 7692 4862 7744
rect 7300 7741 7328 7772
rect 7558 7760 7564 7772
rect 7616 7800 7622 7812
rect 7616 7772 7788 7800
rect 7616 7760 7622 7772
rect 7285 7735 7343 7741
rect 7285 7701 7297 7735
rect 7331 7701 7343 7735
rect 7760 7732 7788 7772
rect 8386 7760 8392 7812
rect 8444 7760 8450 7812
rect 8490 7803 8548 7809
rect 8490 7769 8502 7803
rect 8536 7769 8548 7803
rect 8490 7763 8548 7769
rect 9760 7803 9818 7809
rect 9760 7769 9772 7803
rect 9806 7800 9818 7803
rect 11232 7803 11290 7809
rect 9806 7772 11192 7800
rect 9806 7769 9818 7772
rect 9760 7763 9818 7769
rect 8496 7732 8524 7763
rect 7760 7704 8524 7732
rect 10873 7735 10931 7741
rect 7285 7695 7343 7701
rect 10873 7701 10885 7735
rect 10919 7732 10931 7735
rect 11054 7732 11060 7744
rect 10919 7704 11060 7732
rect 10919 7701 10931 7704
rect 10873 7695 10931 7701
rect 11054 7692 11060 7704
rect 11112 7692 11118 7744
rect 11164 7732 11192 7772
rect 11232 7769 11244 7803
rect 11278 7800 11290 7803
rect 11514 7800 11520 7812
rect 11278 7772 11520 7800
rect 11278 7769 11290 7772
rect 11232 7763 11290 7769
rect 11514 7760 11520 7772
rect 11572 7760 11578 7812
rect 11606 7760 11612 7812
rect 11664 7800 11670 7812
rect 12682 7803 12740 7809
rect 12682 7800 12694 7803
rect 11664 7772 12694 7800
rect 11664 7760 11670 7772
rect 12682 7769 12694 7772
rect 12728 7769 12740 7803
rect 12682 7763 12740 7769
rect 13354 7760 13360 7812
rect 13412 7800 13418 7812
rect 14338 7803 14396 7809
rect 14338 7800 14350 7803
rect 13412 7772 14350 7800
rect 13412 7760 13418 7772
rect 14338 7769 14350 7772
rect 14384 7769 14396 7803
rect 15810 7803 15868 7809
rect 15810 7800 15822 7803
rect 14338 7763 14396 7769
rect 14476 7772 15822 7800
rect 11882 7732 11888 7744
rect 11164 7704 11888 7732
rect 11882 7692 11888 7704
rect 11940 7692 11946 7744
rect 12345 7735 12403 7741
rect 12345 7701 12357 7735
rect 12391 7732 12403 7735
rect 12526 7732 12532 7744
rect 12391 7704 12532 7732
rect 12391 7701 12403 7704
rect 12345 7695 12403 7701
rect 12526 7692 12532 7704
rect 12584 7692 12590 7744
rect 13814 7732 13820 7744
rect 13727 7704 13820 7732
rect 13814 7692 13820 7704
rect 13872 7732 13878 7744
rect 14476 7732 14504 7772
rect 15810 7769 15822 7772
rect 15856 7769 15868 7803
rect 17282 7803 17340 7809
rect 17282 7800 17294 7803
rect 15810 7763 15868 7769
rect 16960 7772 17294 7800
rect 13872 7704 14504 7732
rect 13872 7692 13878 7704
rect 14734 7692 14740 7744
rect 14792 7732 14798 7744
rect 15473 7735 15531 7741
rect 15473 7732 15485 7735
rect 14792 7704 15485 7732
rect 14792 7692 14798 7704
rect 15473 7701 15485 7704
rect 15519 7701 15531 7735
rect 15473 7695 15531 7701
rect 16666 7692 16672 7744
rect 16724 7732 16730 7744
rect 16960 7741 16988 7772
rect 17282 7769 17294 7772
rect 17328 7769 17340 7803
rect 17282 7763 17340 7769
rect 17402 7760 17408 7812
rect 17460 7760 17466 7812
rect 20162 7800 20168 7812
rect 19076 7772 20168 7800
rect 19076 7741 19104 7772
rect 20162 7760 20168 7772
rect 20220 7760 20226 7812
rect 20254 7760 20260 7812
rect 20312 7800 20318 7812
rect 20358 7803 20416 7809
rect 20358 7800 20370 7803
rect 20312 7772 20370 7800
rect 20312 7760 20318 7772
rect 20358 7769 20370 7772
rect 20404 7769 20416 7803
rect 20358 7763 20416 7769
rect 16945 7735 17003 7741
rect 16945 7732 16957 7735
rect 16724 7704 16957 7732
rect 16724 7692 16730 7704
rect 16945 7701 16957 7704
rect 16991 7701 17003 7735
rect 16945 7695 17003 7701
rect 19061 7735 19119 7741
rect 19061 7701 19073 7735
rect 19107 7701 19119 7735
rect 19061 7695 19119 7701
rect 19245 7735 19303 7741
rect 19245 7701 19257 7735
rect 19291 7732 19303 7735
rect 19518 7732 19524 7744
rect 19291 7704 19524 7732
rect 19291 7701 19303 7704
rect 19245 7695 19303 7701
rect 19518 7692 19524 7704
rect 19576 7692 19582 7744
rect 21174 7732 21180 7744
rect 21232 7741 21238 7744
rect 21141 7704 21180 7732
rect 21174 7692 21180 7704
rect 21232 7695 21241 7741
rect 22646 7732 22652 7744
rect 22607 7704 22652 7732
rect 21232 7692 21238 7695
rect 22646 7692 22652 7704
rect 22704 7692 22710 7744
rect 22925 7735 22983 7741
rect 22925 7701 22937 7735
rect 22971 7732 22983 7735
rect 23566 7732 23572 7744
rect 22971 7704 23572 7732
rect 22971 7701 22983 7704
rect 22925 7695 22983 7701
rect 23566 7692 23572 7704
rect 23624 7692 23630 7744
rect 1104 7642 23460 7664
rect 1104 7590 6548 7642
rect 6600 7590 6612 7642
rect 6664 7590 6676 7642
rect 6728 7590 6740 7642
rect 6792 7590 6804 7642
rect 6856 7590 12146 7642
rect 12198 7590 12210 7642
rect 12262 7590 12274 7642
rect 12326 7590 12338 7642
rect 12390 7590 12402 7642
rect 12454 7590 17744 7642
rect 17796 7590 17808 7642
rect 17860 7590 17872 7642
rect 17924 7590 17936 7642
rect 17988 7590 18000 7642
rect 18052 7590 23460 7642
rect 1104 7568 23460 7590
rect 4338 7488 4344 7540
rect 4396 7528 4402 7540
rect 4801 7531 4859 7537
rect 4801 7528 4813 7531
rect 4396 7500 4813 7528
rect 4396 7488 4402 7500
rect 4801 7497 4813 7500
rect 4847 7497 4859 7531
rect 4801 7491 4859 7497
rect 9214 7488 9220 7540
rect 9272 7528 9278 7540
rect 9861 7531 9919 7537
rect 9861 7528 9873 7531
rect 9272 7500 9873 7528
rect 9272 7488 9278 7500
rect 9861 7497 9873 7500
rect 9907 7497 9919 7531
rect 9861 7491 9919 7497
rect 10042 7488 10048 7540
rect 10100 7528 10106 7540
rect 10321 7531 10379 7537
rect 10321 7528 10333 7531
rect 10100 7500 10333 7528
rect 10100 7488 10106 7500
rect 10321 7497 10333 7500
rect 10367 7497 10379 7531
rect 10686 7528 10692 7540
rect 10647 7500 10692 7528
rect 10321 7491 10379 7497
rect 10686 7488 10692 7500
rect 10744 7528 10750 7540
rect 10965 7531 11023 7537
rect 10965 7528 10977 7531
rect 10744 7500 10977 7528
rect 10744 7488 10750 7500
rect 10965 7497 10977 7500
rect 11011 7528 11023 7531
rect 11793 7531 11851 7537
rect 11793 7528 11805 7531
rect 11011 7500 11805 7528
rect 11011 7497 11023 7500
rect 10965 7491 11023 7497
rect 11793 7497 11805 7500
rect 11839 7497 11851 7531
rect 13354 7528 13360 7540
rect 13315 7500 13360 7528
rect 11793 7491 11851 7497
rect 3142 7420 3148 7472
rect 3200 7460 3206 7472
rect 3200 7432 3464 7460
rect 3200 7420 3206 7432
rect 3326 7392 3332 7404
rect 3287 7364 3332 7392
rect 3326 7352 3332 7364
rect 3384 7352 3390 7404
rect 3436 7392 3464 7432
rect 5534 7420 5540 7472
rect 5592 7460 5598 7472
rect 5914 7463 5972 7469
rect 5914 7460 5926 7463
rect 5592 7432 5926 7460
rect 5592 7420 5598 7432
rect 5914 7429 5926 7432
rect 5960 7429 5972 7463
rect 5914 7423 5972 7429
rect 10229 7463 10287 7469
rect 10229 7429 10241 7463
rect 10275 7460 10287 7463
rect 10410 7460 10416 7472
rect 10275 7432 10416 7460
rect 10275 7429 10287 7432
rect 10229 7423 10287 7429
rect 10410 7420 10416 7432
rect 10468 7420 10474 7472
rect 11054 7420 11060 7472
rect 11112 7460 11118 7472
rect 11606 7460 11612 7472
rect 11112 7432 11612 7460
rect 11112 7420 11118 7432
rect 11606 7420 11612 7432
rect 11664 7420 11670 7472
rect 3596 7395 3654 7401
rect 3596 7392 3608 7395
rect 3436 7364 3608 7392
rect 3596 7361 3608 7364
rect 3642 7392 3654 7395
rect 5074 7392 5080 7404
rect 3642 7364 5080 7392
rect 3642 7361 3654 7364
rect 3596 7355 3654 7361
rect 5074 7352 5080 7364
rect 5132 7352 5138 7404
rect 6086 7352 6092 7404
rect 6144 7392 6150 7404
rect 6181 7395 6239 7401
rect 6181 7392 6193 7395
rect 6144 7364 6193 7392
rect 6144 7352 6150 7364
rect 6181 7361 6193 7364
rect 6227 7392 6239 7395
rect 6365 7395 6423 7401
rect 6365 7392 6377 7395
rect 6227 7364 6377 7392
rect 6227 7361 6239 7364
rect 6181 7355 6239 7361
rect 6365 7361 6377 7364
rect 6411 7392 6423 7395
rect 6549 7395 6607 7401
rect 6549 7392 6561 7395
rect 6411 7364 6561 7392
rect 6411 7361 6423 7364
rect 6365 7355 6423 7361
rect 6549 7361 6561 7364
rect 6595 7392 6607 7395
rect 6638 7392 6644 7404
rect 6595 7364 6644 7392
rect 6595 7361 6607 7364
rect 6549 7355 6607 7361
rect 6638 7352 6644 7364
rect 6696 7392 6702 7404
rect 6733 7395 6791 7401
rect 6733 7392 6745 7395
rect 6696 7364 6745 7392
rect 6696 7352 6702 7364
rect 6733 7361 6745 7364
rect 6779 7392 6791 7395
rect 6917 7395 6975 7401
rect 6917 7392 6929 7395
rect 6779 7364 6929 7392
rect 6779 7361 6791 7364
rect 6733 7355 6791 7361
rect 6917 7361 6929 7364
rect 6963 7361 6975 7395
rect 6917 7355 6975 7361
rect 7006 7352 7012 7404
rect 7064 7392 7070 7404
rect 7184 7395 7242 7401
rect 7184 7392 7196 7395
rect 7064 7364 7196 7392
rect 7064 7352 7070 7364
rect 7184 7361 7196 7364
rect 7230 7392 7242 7395
rect 7650 7392 7656 7404
rect 7230 7364 7656 7392
rect 7230 7361 7242 7364
rect 7184 7355 7242 7361
rect 7650 7352 7656 7364
rect 7708 7352 7714 7404
rect 8386 7392 8392 7404
rect 8347 7364 8392 7392
rect 8386 7352 8392 7364
rect 8444 7352 8450 7404
rect 8662 7401 8668 7404
rect 8656 7392 8668 7401
rect 8623 7364 8668 7392
rect 8656 7355 8668 7364
rect 8662 7352 8668 7355
rect 8720 7352 8726 7404
rect 11808 7392 11836 7491
rect 13354 7488 13360 7500
rect 13412 7488 13418 7540
rect 16022 7528 16028 7540
rect 15983 7500 16028 7528
rect 16022 7488 16028 7500
rect 16080 7488 16086 7540
rect 19518 7528 19524 7540
rect 18064 7500 19524 7528
rect 12066 7420 12072 7472
rect 12124 7460 12130 7472
rect 12222 7463 12280 7469
rect 12222 7460 12234 7463
rect 12124 7432 12234 7460
rect 12124 7420 12130 7432
rect 12222 7429 12234 7432
rect 12268 7429 12280 7463
rect 12222 7423 12280 7429
rect 14001 7463 14059 7469
rect 14001 7429 14013 7463
rect 14047 7460 14059 7463
rect 14185 7463 14243 7469
rect 14185 7460 14197 7463
rect 14047 7432 14197 7460
rect 14047 7429 14059 7432
rect 14001 7423 14059 7429
rect 14185 7429 14197 7432
rect 14231 7460 14243 7463
rect 16040 7460 16068 7488
rect 14231 7432 16068 7460
rect 16936 7463 16994 7469
rect 14231 7429 14243 7432
rect 14185 7423 14243 7429
rect 11977 7395 12035 7401
rect 11977 7392 11989 7395
rect 11808 7364 11989 7392
rect 11977 7361 11989 7364
rect 12023 7361 12035 7395
rect 11977 7355 12035 7361
rect 13633 7395 13691 7401
rect 13633 7361 13645 7395
rect 13679 7392 13691 7395
rect 13722 7392 13728 7404
rect 13679 7364 13728 7392
rect 13679 7361 13691 7364
rect 13633 7355 13691 7361
rect 13722 7352 13728 7364
rect 13780 7352 13786 7404
rect 14476 7401 14504 7432
rect 16936 7429 16948 7463
rect 16982 7460 16994 7463
rect 18064 7460 18092 7500
rect 19518 7488 19524 7500
rect 19576 7488 19582 7540
rect 21082 7528 21088 7540
rect 19904 7500 20944 7528
rect 21043 7500 21088 7528
rect 16982 7432 18092 7460
rect 16982 7429 16994 7432
rect 16936 7423 16994 7429
rect 18690 7420 18696 7472
rect 18748 7460 18754 7472
rect 19904 7460 19932 7500
rect 18748 7432 19932 7460
rect 18748 7420 18754 7432
rect 19978 7420 19984 7472
rect 20036 7460 20042 7472
rect 20916 7460 20944 7500
rect 21082 7488 21088 7500
rect 21140 7488 21146 7540
rect 23014 7528 23020 7540
rect 22975 7500 23020 7528
rect 23014 7488 23020 7500
rect 23072 7488 23078 7540
rect 21450 7460 21456 7472
rect 20036 7432 20852 7460
rect 20916 7432 21456 7460
rect 20036 7420 20042 7432
rect 14734 7401 14740 7404
rect 14461 7395 14519 7401
rect 14461 7361 14473 7395
rect 14507 7361 14519 7395
rect 14728 7392 14740 7401
rect 14695 7364 14740 7392
rect 14461 7355 14519 7361
rect 14728 7355 14740 7364
rect 14734 7352 14740 7355
rect 14792 7352 14798 7404
rect 16298 7392 16304 7404
rect 16259 7364 16304 7392
rect 16298 7352 16304 7364
rect 16356 7352 16362 7404
rect 18141 7395 18199 7401
rect 18141 7392 18153 7395
rect 16684 7364 18153 7392
rect 10410 7284 10416 7336
rect 10468 7324 10474 7336
rect 10468 7296 10513 7324
rect 10468 7284 10474 7296
rect 16022 7284 16028 7336
rect 16080 7324 16086 7336
rect 16684 7333 16712 7364
rect 18141 7361 18153 7364
rect 18187 7361 18199 7395
rect 18397 7395 18455 7401
rect 18397 7392 18409 7395
rect 18141 7355 18199 7361
rect 18248 7364 18409 7392
rect 16669 7327 16727 7333
rect 16669 7324 16681 7327
rect 16080 7296 16681 7324
rect 16080 7284 16086 7296
rect 16669 7293 16681 7296
rect 16715 7293 16727 7327
rect 18248 7324 18276 7364
rect 18397 7361 18409 7364
rect 18443 7361 18455 7395
rect 18397 7355 18455 7361
rect 19880 7395 19938 7401
rect 19880 7361 19892 7395
rect 19926 7392 19938 7395
rect 20438 7392 20444 7404
rect 19926 7364 20444 7392
rect 19926 7361 19938 7364
rect 19880 7355 19938 7361
rect 20438 7352 20444 7364
rect 20496 7352 20502 7404
rect 20824 7392 20852 7432
rect 21450 7420 21456 7432
rect 21508 7420 21514 7472
rect 21542 7392 21548 7404
rect 20824 7364 21404 7392
rect 21503 7364 21548 7392
rect 19610 7324 19616 7336
rect 16669 7287 16727 7293
rect 18156 7296 18276 7324
rect 19523 7296 19616 7324
rect 9766 7256 9772 7268
rect 4724 7228 5304 7256
rect 9727 7228 9772 7256
rect 2406 7148 2412 7200
rect 2464 7188 2470 7200
rect 4724 7197 4752 7228
rect 4709 7191 4767 7197
rect 4709 7188 4721 7191
rect 2464 7160 4721 7188
rect 2464 7148 2470 7160
rect 4709 7157 4721 7160
rect 4755 7157 4767 7191
rect 5276 7188 5304 7228
rect 9766 7216 9772 7228
rect 9824 7216 9830 7268
rect 15396 7228 16252 7256
rect 5902 7188 5908 7200
rect 5276 7160 5908 7188
rect 4709 7151 4767 7157
rect 5902 7148 5908 7160
rect 5960 7148 5966 7200
rect 8297 7191 8355 7197
rect 8297 7157 8309 7191
rect 8343 7188 8355 7191
rect 8570 7188 8576 7200
rect 8343 7160 8576 7188
rect 8343 7157 8355 7160
rect 8297 7151 8355 7157
rect 8570 7148 8576 7160
rect 8628 7148 8634 7200
rect 10042 7148 10048 7200
rect 10100 7188 10106 7200
rect 13446 7188 13452 7200
rect 10100 7160 13452 7188
rect 10100 7148 10106 7160
rect 13446 7148 13452 7160
rect 13504 7148 13510 7200
rect 13538 7148 13544 7200
rect 13596 7188 13602 7200
rect 13596 7160 13641 7188
rect 13596 7148 13602 7160
rect 13722 7148 13728 7200
rect 13780 7188 13786 7200
rect 15396 7188 15424 7228
rect 15838 7188 15844 7200
rect 13780 7160 15424 7188
rect 15799 7160 15844 7188
rect 13780 7148 13786 7160
rect 15838 7148 15844 7160
rect 15896 7148 15902 7200
rect 16224 7197 16252 7228
rect 18156 7200 18184 7296
rect 19610 7284 19616 7296
rect 19668 7284 19674 7336
rect 21376 7324 21404 7364
rect 21542 7352 21548 7364
rect 21600 7352 21606 7404
rect 22186 7392 22192 7404
rect 22147 7364 22192 7392
rect 22186 7352 22192 7364
rect 22244 7352 22250 7404
rect 22833 7395 22891 7401
rect 22833 7361 22845 7395
rect 22879 7392 22891 7395
rect 22922 7392 22928 7404
rect 22879 7364 22928 7392
rect 22879 7361 22891 7364
rect 22833 7355 22891 7361
rect 22922 7352 22928 7364
rect 22980 7352 22986 7404
rect 21913 7327 21971 7333
rect 21913 7324 21925 7327
rect 21376 7296 21925 7324
rect 21913 7293 21925 7296
rect 21959 7293 21971 7327
rect 21913 7287 21971 7293
rect 22094 7284 22100 7336
rect 22152 7324 22158 7336
rect 22152 7296 22197 7324
rect 22152 7284 22158 7296
rect 16209 7191 16267 7197
rect 16209 7157 16221 7191
rect 16255 7188 16267 7191
rect 17954 7188 17960 7200
rect 16255 7160 17960 7188
rect 16255 7157 16267 7160
rect 16209 7151 16267 7157
rect 17954 7148 17960 7160
rect 18012 7148 18018 7200
rect 18049 7191 18107 7197
rect 18049 7157 18061 7191
rect 18095 7188 18107 7191
rect 18138 7188 18144 7200
rect 18095 7160 18144 7188
rect 18095 7157 18107 7160
rect 18049 7151 18107 7157
rect 18138 7148 18144 7160
rect 18196 7148 18202 7200
rect 19426 7148 19432 7200
rect 19484 7188 19490 7200
rect 19521 7191 19579 7197
rect 19521 7188 19533 7191
rect 19484 7160 19533 7188
rect 19484 7148 19490 7160
rect 19521 7157 19533 7160
rect 19567 7157 19579 7191
rect 19628 7188 19656 7284
rect 20993 7259 21051 7265
rect 20993 7225 21005 7259
rect 21039 7256 21051 7259
rect 21266 7256 21272 7268
rect 21039 7228 21272 7256
rect 21039 7225 21051 7228
rect 20993 7219 21051 7225
rect 21266 7216 21272 7228
rect 21324 7216 21330 7268
rect 22554 7256 22560 7268
rect 22515 7228 22560 7256
rect 22554 7216 22560 7228
rect 22612 7216 22618 7268
rect 20346 7188 20352 7200
rect 19628 7160 20352 7188
rect 19521 7151 19579 7157
rect 20346 7148 20352 7160
rect 20404 7188 20410 7200
rect 20622 7188 20628 7200
rect 20404 7160 20628 7188
rect 20404 7148 20410 7160
rect 20622 7148 20628 7160
rect 20680 7148 20686 7200
rect 21082 7148 21088 7200
rect 21140 7188 21146 7200
rect 21361 7191 21419 7197
rect 21361 7188 21373 7191
rect 21140 7160 21373 7188
rect 21140 7148 21146 7160
rect 21361 7157 21373 7160
rect 21407 7157 21419 7191
rect 22646 7188 22652 7200
rect 22607 7160 22652 7188
rect 21361 7151 21419 7157
rect 22646 7148 22652 7160
rect 22704 7148 22710 7200
rect 1104 7098 23460 7120
rect 1104 7046 3749 7098
rect 3801 7046 3813 7098
rect 3865 7046 3877 7098
rect 3929 7046 3941 7098
rect 3993 7046 4005 7098
rect 4057 7046 9347 7098
rect 9399 7046 9411 7098
rect 9463 7046 9475 7098
rect 9527 7046 9539 7098
rect 9591 7046 9603 7098
rect 9655 7046 14945 7098
rect 14997 7046 15009 7098
rect 15061 7046 15073 7098
rect 15125 7046 15137 7098
rect 15189 7046 15201 7098
rect 15253 7046 20543 7098
rect 20595 7046 20607 7098
rect 20659 7046 20671 7098
rect 20723 7046 20735 7098
rect 20787 7046 20799 7098
rect 20851 7046 23460 7098
rect 1104 7024 23460 7046
rect 3326 6944 3332 6996
rect 3384 6984 3390 6996
rect 4801 6987 4859 6993
rect 4801 6984 4813 6987
rect 3384 6956 4813 6984
rect 3384 6944 3390 6956
rect 4801 6953 4813 6956
rect 4847 6953 4859 6987
rect 5074 6984 5080 6996
rect 5035 6956 5080 6984
rect 4801 6947 4859 6953
rect 5074 6944 5080 6956
rect 5132 6944 5138 6996
rect 6638 6984 6644 6996
rect 6599 6956 6644 6984
rect 6638 6944 6644 6956
rect 6696 6984 6702 6996
rect 7101 6987 7159 6993
rect 7101 6984 7113 6987
rect 6696 6956 7113 6984
rect 6696 6944 6702 6956
rect 7101 6953 7113 6956
rect 7147 6953 7159 6987
rect 7101 6947 7159 6953
rect 7190 6944 7196 6996
rect 7248 6984 7254 6996
rect 7285 6987 7343 6993
rect 7285 6984 7297 6987
rect 7248 6956 7297 6984
rect 7248 6944 7254 6956
rect 7285 6953 7297 6956
rect 7331 6953 7343 6987
rect 7285 6947 7343 6953
rect 8386 6944 8392 6996
rect 8444 6984 8450 6996
rect 8941 6987 8999 6993
rect 8941 6984 8953 6987
rect 8444 6956 8953 6984
rect 8444 6944 8450 6956
rect 6454 6808 6460 6860
rect 6512 6848 6518 6860
rect 6656 6848 6684 6944
rect 8680 6857 8708 6956
rect 8941 6953 8953 6956
rect 8987 6953 8999 6987
rect 8941 6947 8999 6953
rect 13446 6944 13452 6996
rect 13504 6984 13510 6996
rect 22462 6984 22468 6996
rect 13504 6956 22468 6984
rect 13504 6944 13510 6956
rect 22462 6944 22468 6956
rect 22520 6944 22526 6996
rect 10428 6888 11376 6916
rect 10428 6860 10456 6888
rect 6512 6820 6684 6848
rect 8665 6851 8723 6857
rect 6512 6808 6518 6820
rect 8665 6817 8677 6851
rect 8711 6817 8723 6851
rect 10137 6851 10195 6857
rect 10137 6848 10149 6851
rect 8665 6811 8723 6817
rect 9416 6820 10149 6848
rect 6178 6740 6184 6792
rect 6236 6789 6242 6792
rect 6236 6780 6248 6789
rect 6236 6752 6281 6780
rect 6236 6743 6248 6752
rect 6236 6740 6242 6743
rect 2130 6672 2136 6724
rect 2188 6712 2194 6724
rect 8202 6712 8208 6724
rect 2188 6684 8208 6712
rect 2188 6672 2194 6684
rect 8202 6672 8208 6684
rect 8260 6672 8266 6724
rect 8420 6715 8478 6721
rect 8420 6681 8432 6715
rect 8466 6712 8478 6715
rect 8570 6712 8576 6724
rect 8466 6684 8576 6712
rect 8466 6681 8478 6684
rect 8420 6675 8478 6681
rect 8570 6672 8576 6684
rect 8628 6672 8634 6724
rect 8754 6672 8760 6724
rect 8812 6712 8818 6724
rect 9416 6721 9444 6820
rect 10137 6817 10149 6820
rect 10183 6848 10195 6851
rect 10410 6848 10416 6860
rect 10183 6820 10416 6848
rect 10183 6817 10195 6820
rect 10137 6811 10195 6817
rect 10410 6808 10416 6820
rect 10468 6808 10474 6860
rect 11057 6851 11115 6857
rect 11057 6817 11069 6851
rect 11103 6848 11115 6851
rect 11238 6848 11244 6860
rect 11103 6820 11244 6848
rect 11103 6817 11115 6820
rect 11057 6811 11115 6817
rect 11238 6808 11244 6820
rect 11296 6808 11302 6860
rect 11348 6848 11376 6888
rect 13004 6888 13768 6916
rect 11517 6851 11575 6857
rect 11517 6848 11529 6851
rect 11348 6820 11529 6848
rect 11517 6817 11529 6820
rect 11563 6817 11575 6851
rect 11517 6811 11575 6817
rect 12526 6808 12532 6860
rect 12584 6848 12590 6860
rect 13004 6857 13032 6888
rect 13740 6860 13768 6888
rect 17954 6876 17960 6928
rect 18012 6916 18018 6928
rect 18230 6916 18236 6928
rect 18012 6888 18236 6916
rect 18012 6876 18018 6888
rect 18230 6876 18236 6888
rect 18288 6876 18294 6928
rect 20806 6876 20812 6928
rect 20864 6916 20870 6928
rect 21266 6916 21272 6928
rect 20864 6888 21272 6916
rect 20864 6876 20870 6888
rect 21266 6876 21272 6888
rect 21324 6876 21330 6928
rect 21453 6919 21511 6925
rect 21453 6885 21465 6919
rect 21499 6885 21511 6919
rect 21453 6879 21511 6885
rect 12805 6851 12863 6857
rect 12805 6848 12817 6851
rect 12584 6820 12817 6848
rect 12584 6808 12590 6820
rect 12805 6817 12817 6820
rect 12851 6817 12863 6851
rect 12805 6811 12863 6817
rect 12989 6851 13047 6857
rect 12989 6817 13001 6851
rect 13035 6817 13047 6851
rect 12989 6811 13047 6817
rect 13354 6808 13360 6860
rect 13412 6848 13418 6860
rect 13633 6851 13691 6857
rect 13633 6848 13645 6851
rect 13412 6820 13645 6848
rect 13412 6808 13418 6820
rect 13633 6817 13645 6820
rect 13679 6817 13691 6851
rect 13633 6811 13691 6817
rect 13722 6808 13728 6860
rect 13780 6848 13786 6860
rect 13780 6820 13825 6848
rect 13780 6808 13786 6820
rect 16022 6808 16028 6860
rect 16080 6848 16086 6860
rect 16117 6851 16175 6857
rect 16117 6848 16129 6851
rect 16080 6820 16129 6848
rect 16080 6808 16086 6820
rect 16117 6817 16129 6820
rect 16163 6817 16175 6851
rect 17773 6851 17831 6857
rect 17773 6848 17785 6851
rect 16117 6811 16175 6817
rect 17144 6820 17785 6848
rect 9950 6740 9956 6792
rect 10008 6780 10014 6792
rect 10781 6783 10839 6789
rect 10781 6780 10793 6783
rect 10008 6752 10793 6780
rect 10008 6740 10014 6752
rect 10781 6749 10793 6752
rect 10827 6749 10839 6783
rect 10781 6743 10839 6749
rect 10873 6783 10931 6789
rect 10873 6749 10885 6783
rect 10919 6780 10931 6783
rect 11146 6780 11152 6792
rect 10919 6752 11152 6780
rect 10919 6749 10931 6752
rect 10873 6743 10931 6749
rect 11146 6740 11152 6752
rect 11204 6740 11210 6792
rect 12066 6740 12072 6792
rect 12124 6780 12130 6792
rect 12713 6783 12771 6789
rect 12713 6780 12725 6783
rect 12124 6752 12725 6780
rect 12124 6740 12130 6752
rect 12713 6749 12725 6752
rect 12759 6749 12771 6783
rect 12713 6743 12771 6749
rect 14369 6783 14427 6789
rect 14369 6749 14381 6783
rect 14415 6780 14427 6783
rect 14553 6783 14611 6789
rect 14553 6780 14565 6783
rect 14415 6752 14565 6780
rect 14415 6749 14427 6752
rect 14369 6743 14427 6749
rect 14553 6749 14565 6752
rect 14599 6780 14611 6783
rect 14645 6783 14703 6789
rect 14645 6780 14657 6783
rect 14599 6752 14657 6780
rect 14599 6749 14611 6752
rect 14553 6743 14611 6749
rect 14645 6749 14657 6752
rect 14691 6780 14703 6783
rect 16040 6780 16068 6808
rect 17144 6780 17172 6820
rect 17773 6817 17785 6820
rect 17819 6848 17831 6851
rect 19061 6851 19119 6857
rect 17819 6820 18000 6848
rect 17819 6817 17831 6820
rect 17773 6811 17831 6817
rect 17865 6783 17923 6789
rect 17865 6780 17877 6783
rect 14691 6752 16068 6780
rect 16224 6752 17172 6780
rect 17512 6752 17877 6780
rect 14691 6749 14703 6752
rect 14645 6743 14703 6749
rect 9401 6715 9459 6721
rect 9401 6712 9413 6715
rect 8812 6684 9413 6712
rect 8812 6672 8818 6684
rect 9401 6681 9413 6684
rect 9447 6681 9459 6715
rect 10226 6712 10232 6724
rect 9401 6675 9459 6681
rect 9968 6684 10232 6712
rect 9306 6644 9312 6656
rect 9267 6616 9312 6644
rect 9306 6604 9312 6616
rect 9364 6604 9370 6656
rect 9585 6647 9643 6653
rect 9585 6613 9597 6647
rect 9631 6644 9643 6647
rect 9674 6644 9680 6656
rect 9631 6616 9680 6644
rect 9631 6613 9643 6616
rect 9585 6607 9643 6613
rect 9674 6604 9680 6616
rect 9732 6604 9738 6656
rect 9968 6653 9996 6684
rect 10226 6672 10232 6684
rect 10284 6672 10290 6724
rect 11790 6672 11796 6724
rect 11848 6712 11854 6724
rect 13541 6715 13599 6721
rect 11848 6684 13492 6712
rect 11848 6672 11854 6684
rect 9953 6647 10011 6653
rect 9953 6613 9965 6647
rect 9999 6613 10011 6647
rect 9953 6607 10011 6613
rect 10045 6647 10103 6653
rect 10045 6613 10057 6647
rect 10091 6644 10103 6647
rect 10134 6644 10140 6656
rect 10091 6616 10140 6644
rect 10091 6613 10103 6616
rect 10045 6607 10103 6613
rect 10134 6604 10140 6616
rect 10192 6604 10198 6656
rect 10410 6644 10416 6656
rect 10371 6616 10416 6644
rect 10410 6604 10416 6616
rect 10468 6604 10474 6656
rect 12066 6604 12072 6656
rect 12124 6644 12130 6656
rect 12345 6647 12403 6653
rect 12345 6644 12357 6647
rect 12124 6616 12357 6644
rect 12124 6604 12130 6616
rect 12345 6613 12357 6616
rect 12391 6613 12403 6647
rect 13170 6644 13176 6656
rect 13131 6616 13176 6644
rect 12345 6607 12403 6613
rect 13170 6604 13176 6616
rect 13228 6604 13234 6656
rect 13464 6644 13492 6684
rect 13541 6681 13553 6715
rect 13587 6712 13599 6715
rect 14734 6712 14740 6724
rect 13587 6684 14740 6712
rect 13587 6681 13599 6684
rect 13541 6675 13599 6681
rect 14734 6672 14740 6684
rect 14792 6672 14798 6724
rect 14912 6715 14970 6721
rect 14912 6681 14924 6715
rect 14958 6712 14970 6715
rect 15746 6712 15752 6724
rect 14958 6684 15752 6712
rect 14958 6681 14970 6684
rect 14912 6675 14970 6681
rect 15746 6672 15752 6684
rect 15804 6672 15810 6724
rect 16224 6712 16252 6752
rect 16390 6721 16396 6724
rect 16384 6712 16396 6721
rect 15856 6684 16252 6712
rect 16351 6684 16396 6712
rect 15856 6644 15884 6684
rect 16384 6675 16396 6684
rect 16390 6672 16396 6675
rect 16448 6672 16454 6724
rect 16482 6672 16488 6724
rect 16540 6712 16546 6724
rect 17512 6712 17540 6752
rect 17865 6749 17877 6752
rect 17911 6749 17923 6783
rect 17972 6780 18000 6820
rect 19061 6817 19073 6851
rect 19107 6848 19119 6851
rect 19242 6848 19248 6860
rect 19107 6820 19248 6848
rect 19107 6817 19119 6820
rect 19061 6811 19119 6817
rect 19242 6808 19248 6820
rect 19300 6808 19306 6860
rect 20622 6848 20628 6860
rect 20583 6820 20628 6848
rect 20622 6808 20628 6820
rect 20680 6808 20686 6860
rect 20898 6848 20904 6860
rect 20859 6820 20904 6848
rect 20898 6808 20904 6820
rect 20956 6808 20962 6860
rect 21468 6848 21496 6879
rect 22094 6848 22100 6860
rect 21468 6820 22100 6848
rect 22094 6808 22100 6820
rect 22152 6808 22158 6860
rect 22189 6851 22247 6857
rect 22189 6817 22201 6851
rect 22235 6817 22247 6851
rect 22189 6811 22247 6817
rect 19886 6780 19892 6792
rect 17972 6752 19892 6780
rect 17865 6743 17923 6749
rect 19886 6740 19892 6752
rect 19944 6740 19950 6792
rect 20714 6780 20720 6792
rect 19996 6752 20720 6780
rect 16540 6684 17540 6712
rect 16540 6672 16546 6684
rect 17586 6672 17592 6724
rect 17644 6712 17650 6724
rect 17957 6715 18015 6721
rect 17957 6712 17969 6715
rect 17644 6684 17969 6712
rect 17644 6672 17650 6684
rect 17957 6681 17969 6684
rect 18003 6681 18015 6715
rect 18874 6712 18880 6724
rect 17957 6675 18015 6681
rect 18340 6684 18880 6712
rect 13464 6616 15884 6644
rect 15930 6604 15936 6656
rect 15988 6644 15994 6656
rect 16025 6647 16083 6653
rect 16025 6644 16037 6647
rect 15988 6616 16037 6644
rect 15988 6604 15994 6616
rect 16025 6613 16037 6616
rect 16071 6613 16083 6647
rect 17494 6644 17500 6656
rect 17455 6616 17500 6644
rect 16025 6607 16083 6613
rect 17494 6604 17500 6616
rect 17552 6604 17558 6656
rect 18340 6653 18368 6684
rect 18874 6672 18880 6684
rect 18932 6672 18938 6724
rect 19150 6672 19156 6724
rect 19208 6712 19214 6724
rect 19996 6712 20024 6752
rect 20714 6740 20720 6752
rect 20772 6740 20778 6792
rect 22204 6780 22232 6811
rect 22462 6780 22468 6792
rect 20824 6752 22232 6780
rect 22423 6752 22468 6780
rect 19208 6684 20024 6712
rect 20380 6715 20438 6721
rect 19208 6672 19214 6684
rect 20380 6681 20392 6715
rect 20426 6712 20438 6715
rect 20530 6712 20536 6724
rect 20426 6684 20536 6712
rect 20426 6681 20438 6684
rect 20380 6675 20438 6681
rect 20530 6672 20536 6684
rect 20588 6672 20594 6724
rect 18325 6647 18383 6653
rect 18325 6613 18337 6647
rect 18371 6613 18383 6647
rect 18325 6607 18383 6613
rect 18414 6604 18420 6656
rect 18472 6644 18478 6656
rect 18690 6644 18696 6656
rect 18472 6616 18517 6644
rect 18651 6616 18696 6644
rect 18472 6604 18478 6616
rect 18690 6604 18696 6616
rect 18748 6604 18754 6656
rect 19058 6604 19064 6656
rect 19116 6644 19122 6656
rect 19245 6647 19303 6653
rect 19245 6644 19257 6647
rect 19116 6616 19257 6644
rect 19116 6604 19122 6616
rect 19245 6613 19257 6616
rect 19291 6644 19303 6647
rect 20824 6644 20852 6752
rect 22462 6740 22468 6752
rect 22520 6740 22526 6792
rect 22830 6780 22836 6792
rect 22791 6752 22836 6780
rect 22830 6740 22836 6752
rect 22888 6740 22894 6792
rect 20898 6672 20904 6724
rect 20956 6712 20962 6724
rect 21085 6715 21143 6721
rect 21085 6712 21097 6715
rect 20956 6684 21097 6712
rect 20956 6672 20962 6684
rect 21085 6681 21097 6684
rect 21131 6681 21143 6715
rect 21085 6675 21143 6681
rect 21450 6672 21456 6724
rect 21508 6712 21514 6724
rect 22097 6715 22155 6721
rect 22097 6712 22109 6715
rect 21508 6684 22109 6712
rect 21508 6672 21514 6684
rect 22097 6681 22109 6684
rect 22143 6681 22155 6715
rect 22097 6675 22155 6681
rect 20990 6644 20996 6656
rect 19291 6616 20852 6644
rect 20951 6616 20996 6644
rect 19291 6613 19303 6616
rect 19245 6607 19303 6613
rect 20990 6604 20996 6616
rect 21048 6604 21054 6656
rect 21266 6604 21272 6656
rect 21324 6644 21330 6656
rect 21637 6647 21695 6653
rect 21637 6644 21649 6647
rect 21324 6616 21649 6644
rect 21324 6604 21330 6616
rect 21637 6613 21649 6616
rect 21683 6613 21695 6647
rect 22002 6644 22008 6656
rect 21963 6616 22008 6644
rect 21637 6607 21695 6613
rect 22002 6604 22008 6616
rect 22060 6604 22066 6656
rect 22649 6647 22707 6653
rect 22649 6613 22661 6647
rect 22695 6644 22707 6647
rect 22830 6644 22836 6656
rect 22695 6616 22836 6644
rect 22695 6613 22707 6616
rect 22649 6607 22707 6613
rect 22830 6604 22836 6616
rect 22888 6604 22894 6656
rect 23014 6644 23020 6656
rect 22975 6616 23020 6644
rect 23014 6604 23020 6616
rect 23072 6604 23078 6656
rect 1104 6554 23460 6576
rect 1104 6502 6548 6554
rect 6600 6502 6612 6554
rect 6664 6502 6676 6554
rect 6728 6502 6740 6554
rect 6792 6502 6804 6554
rect 6856 6502 12146 6554
rect 12198 6502 12210 6554
rect 12262 6502 12274 6554
rect 12326 6502 12338 6554
rect 12390 6502 12402 6554
rect 12454 6502 17744 6554
rect 17796 6502 17808 6554
rect 17860 6502 17872 6554
rect 17924 6502 17936 6554
rect 17988 6502 18000 6554
rect 18052 6502 23460 6554
rect 1104 6480 23460 6502
rect 4798 6440 4804 6452
rect 4759 6412 4804 6440
rect 4798 6400 4804 6412
rect 4856 6400 4862 6452
rect 6454 6440 6460 6452
rect 6415 6412 6460 6440
rect 6454 6400 6460 6412
rect 6512 6400 6518 6452
rect 7558 6440 7564 6452
rect 7519 6412 7564 6440
rect 7558 6400 7564 6412
rect 7616 6400 7622 6452
rect 7650 6400 7656 6452
rect 7708 6440 7714 6452
rect 8481 6443 8539 6449
rect 8481 6440 8493 6443
rect 7708 6412 8493 6440
rect 7708 6400 7714 6412
rect 8481 6409 8493 6412
rect 8527 6409 8539 6443
rect 8481 6403 8539 6409
rect 9214 6400 9220 6452
rect 9272 6440 9278 6452
rect 9309 6443 9367 6449
rect 9309 6440 9321 6443
rect 9272 6412 9321 6440
rect 9272 6400 9278 6412
rect 9309 6409 9321 6412
rect 9355 6409 9367 6443
rect 9309 6403 9367 6409
rect 10045 6443 10103 6449
rect 10045 6409 10057 6443
rect 10091 6440 10103 6443
rect 10318 6440 10324 6452
rect 10091 6412 10324 6440
rect 10091 6409 10103 6412
rect 10045 6403 10103 6409
rect 10318 6400 10324 6412
rect 10376 6400 10382 6452
rect 10873 6443 10931 6449
rect 10873 6409 10885 6443
rect 10919 6440 10931 6443
rect 12345 6443 12403 6449
rect 12345 6440 12357 6443
rect 10919 6412 12357 6440
rect 10919 6409 10931 6412
rect 10873 6403 10931 6409
rect 12345 6409 12357 6412
rect 12391 6409 12403 6443
rect 12710 6440 12716 6452
rect 12671 6412 12716 6440
rect 12345 6403 12403 6409
rect 12710 6400 12716 6412
rect 12768 6400 12774 6452
rect 12805 6443 12863 6449
rect 12805 6409 12817 6443
rect 12851 6440 12863 6443
rect 12986 6440 12992 6452
rect 12851 6412 12992 6440
rect 12851 6409 12863 6412
rect 12805 6403 12863 6409
rect 12986 6400 12992 6412
rect 13044 6400 13050 6452
rect 13265 6443 13323 6449
rect 13265 6409 13277 6443
rect 13311 6440 13323 6443
rect 15746 6440 15752 6452
rect 13311 6412 15752 6440
rect 13311 6409 13323 6412
rect 13265 6403 13323 6409
rect 5902 6332 5908 6384
rect 5960 6381 5966 6384
rect 5960 6372 5972 6381
rect 5960 6344 6005 6372
rect 5960 6335 5972 6344
rect 5960 6332 5966 6335
rect 6181 6307 6239 6313
rect 6181 6273 6193 6307
rect 6227 6304 6239 6307
rect 6472 6304 6500 6400
rect 8294 6332 8300 6384
rect 8352 6372 8358 6384
rect 8573 6375 8631 6381
rect 8573 6372 8585 6375
rect 8352 6344 8585 6372
rect 8352 6332 8358 6344
rect 8573 6341 8585 6344
rect 8619 6341 8631 6375
rect 10410 6372 10416 6384
rect 8573 6335 8631 6341
rect 9232 6344 10416 6372
rect 6227 6276 6500 6304
rect 6227 6273 6239 6276
rect 6181 6267 6239 6273
rect 7466 6264 7472 6316
rect 7524 6304 7530 6316
rect 9232 6313 9260 6344
rect 10410 6332 10416 6344
rect 10468 6332 10474 6384
rect 11330 6372 11336 6384
rect 10796 6344 11336 6372
rect 7653 6307 7711 6313
rect 7653 6304 7665 6307
rect 7524 6276 7665 6304
rect 7524 6264 7530 6276
rect 7653 6273 7665 6276
rect 7699 6273 7711 6307
rect 9217 6307 9275 6313
rect 7653 6267 7711 6273
rect 8496 6276 9168 6304
rect 7374 6236 7380 6248
rect 7287 6208 7380 6236
rect 7374 6196 7380 6208
rect 7432 6236 7438 6248
rect 8496 6236 8524 6276
rect 8754 6236 8760 6248
rect 7432 6208 8524 6236
rect 8715 6208 8760 6236
rect 7432 6196 7438 6208
rect 8754 6196 8760 6208
rect 8812 6196 8818 6248
rect 9033 6239 9091 6245
rect 9033 6205 9045 6239
rect 9079 6205 9091 6239
rect 9140 6236 9168 6276
rect 9217 6273 9229 6307
rect 9263 6273 9275 6307
rect 9217 6267 9275 6273
rect 10137 6307 10195 6313
rect 10137 6273 10149 6307
rect 10183 6304 10195 6307
rect 10796 6304 10824 6344
rect 11330 6332 11336 6344
rect 11388 6332 11394 6384
rect 11422 6332 11428 6384
rect 11480 6372 11486 6384
rect 11793 6375 11851 6381
rect 11793 6372 11805 6375
rect 11480 6344 11805 6372
rect 11480 6332 11486 6344
rect 11793 6341 11805 6344
rect 11839 6372 11851 6375
rect 13280 6372 13308 6403
rect 15746 6400 15752 6412
rect 15804 6400 15810 6452
rect 15930 6400 15936 6452
rect 15988 6440 15994 6452
rect 16025 6443 16083 6449
rect 16025 6440 16037 6443
rect 15988 6412 16037 6440
rect 15988 6400 15994 6412
rect 16025 6409 16037 6412
rect 16071 6409 16083 6443
rect 16025 6403 16083 6409
rect 16393 6443 16451 6449
rect 16393 6409 16405 6443
rect 16439 6440 16451 6443
rect 16482 6440 16488 6452
rect 16439 6412 16488 6440
rect 16439 6409 16451 6412
rect 16393 6403 16451 6409
rect 16482 6400 16488 6412
rect 16540 6400 16546 6452
rect 17405 6443 17463 6449
rect 17405 6409 17417 6443
rect 17451 6440 17463 6443
rect 17957 6443 18015 6449
rect 17957 6440 17969 6443
rect 17451 6412 17969 6440
rect 17451 6409 17463 6412
rect 17405 6403 17463 6409
rect 17957 6409 17969 6412
rect 18003 6409 18015 6443
rect 17957 6403 18015 6409
rect 18785 6443 18843 6449
rect 18785 6409 18797 6443
rect 18831 6440 18843 6443
rect 19426 6440 19432 6452
rect 18831 6412 19432 6440
rect 18831 6409 18843 6412
rect 18785 6403 18843 6409
rect 19426 6400 19432 6412
rect 19484 6400 19490 6452
rect 20530 6400 20536 6452
rect 20588 6440 20594 6452
rect 20625 6443 20683 6449
rect 20625 6440 20637 6443
rect 20588 6412 20637 6440
rect 20588 6400 20594 6412
rect 20625 6409 20637 6412
rect 20671 6409 20683 6443
rect 20625 6403 20683 6409
rect 20714 6400 20720 6452
rect 20772 6440 20778 6452
rect 20993 6443 21051 6449
rect 20993 6440 21005 6443
rect 20772 6412 21005 6440
rect 20772 6400 20778 6412
rect 20993 6409 21005 6412
rect 21039 6409 21051 6443
rect 21450 6440 21456 6452
rect 21411 6412 21456 6440
rect 20993 6403 21051 6409
rect 21450 6400 21456 6412
rect 21508 6400 21514 6452
rect 21634 6400 21640 6452
rect 21692 6440 21698 6452
rect 21821 6443 21879 6449
rect 21821 6440 21833 6443
rect 21692 6412 21833 6440
rect 21692 6400 21698 6412
rect 21821 6409 21833 6412
rect 21867 6409 21879 6443
rect 21821 6403 21879 6409
rect 11839 6344 13308 6372
rect 15197 6375 15255 6381
rect 11839 6341 11851 6344
rect 11793 6335 11851 6341
rect 15197 6341 15209 6375
rect 15243 6372 15255 6375
rect 15378 6372 15384 6384
rect 15243 6344 15384 6372
rect 15243 6341 15255 6344
rect 15197 6335 15255 6341
rect 15378 6332 15384 6344
rect 15436 6332 15442 6384
rect 16758 6332 16764 6384
rect 16816 6372 16822 6384
rect 17037 6375 17095 6381
rect 17037 6372 17049 6375
rect 16816 6344 17049 6372
rect 16816 6332 16822 6344
rect 17037 6341 17049 6344
rect 17083 6372 17095 6375
rect 18877 6375 18935 6381
rect 17083 6344 18635 6372
rect 17083 6341 17095 6344
rect 17037 6335 17095 6341
rect 10962 6304 10968 6316
rect 10183 6276 10824 6304
rect 10923 6276 10968 6304
rect 10183 6273 10195 6276
rect 10137 6267 10195 6273
rect 10962 6264 10968 6276
rect 11020 6264 11026 6316
rect 11882 6304 11888 6316
rect 11843 6276 11888 6304
rect 11882 6264 11888 6276
rect 11940 6264 11946 6316
rect 14001 6307 14059 6313
rect 14001 6273 14013 6307
rect 14047 6304 14059 6307
rect 14461 6307 14519 6313
rect 14461 6304 14473 6307
rect 14047 6276 14473 6304
rect 14047 6273 14059 6276
rect 14001 6267 14059 6273
rect 14461 6273 14473 6276
rect 14507 6273 14519 6307
rect 14461 6267 14519 6273
rect 15289 6307 15347 6313
rect 15289 6273 15301 6307
rect 15335 6304 15347 6307
rect 15654 6304 15660 6316
rect 15335 6276 15660 6304
rect 15335 6273 15347 6276
rect 15289 6267 15347 6273
rect 15654 6264 15660 6276
rect 15712 6264 15718 6316
rect 15838 6264 15844 6316
rect 15896 6304 15902 6316
rect 15933 6307 15991 6313
rect 15933 6304 15945 6307
rect 15896 6276 15945 6304
rect 15896 6264 15902 6276
rect 15933 6273 15945 6276
rect 15979 6273 15991 6307
rect 15933 6267 15991 6273
rect 17865 6307 17923 6313
rect 17865 6273 17877 6307
rect 17911 6304 17923 6307
rect 18506 6304 18512 6316
rect 17911 6276 18512 6304
rect 17911 6273 17923 6276
rect 17865 6267 17923 6273
rect 18506 6264 18512 6276
rect 18564 6264 18570 6316
rect 18607 6304 18635 6344
rect 18877 6341 18889 6375
rect 18923 6372 18935 6375
rect 19512 6375 19570 6381
rect 18923 6344 19380 6372
rect 18923 6341 18935 6344
rect 18877 6335 18935 6341
rect 19150 6304 19156 6316
rect 18607 6276 19156 6304
rect 19150 6264 19156 6276
rect 19208 6264 19214 6316
rect 19352 6304 19380 6344
rect 19512 6341 19524 6375
rect 19558 6372 19570 6375
rect 19610 6372 19616 6384
rect 19558 6344 19616 6372
rect 19558 6341 19570 6344
rect 19512 6335 19570 6341
rect 19610 6332 19616 6344
rect 19668 6332 19674 6384
rect 19794 6304 19800 6316
rect 19352 6276 19800 6304
rect 19794 6264 19800 6276
rect 19852 6264 19858 6316
rect 19886 6264 19892 6316
rect 19944 6304 19950 6316
rect 20898 6304 20904 6316
rect 19944 6276 20904 6304
rect 19944 6264 19950 6276
rect 20898 6264 20904 6276
rect 20956 6264 20962 6316
rect 21085 6307 21143 6313
rect 21085 6273 21097 6307
rect 21131 6304 21143 6307
rect 21266 6304 21272 6316
rect 21131 6276 21272 6304
rect 21131 6273 21143 6276
rect 21085 6267 21143 6273
rect 21266 6264 21272 6276
rect 21324 6264 21330 6316
rect 22189 6307 22247 6313
rect 22189 6273 22201 6307
rect 22235 6304 22247 6307
rect 22462 6304 22468 6316
rect 22235 6276 22468 6304
rect 22235 6273 22247 6276
rect 22189 6267 22247 6273
rect 22462 6264 22468 6276
rect 22520 6264 22526 6316
rect 22833 6307 22891 6313
rect 22833 6273 22845 6307
rect 22879 6304 22891 6307
rect 23382 6304 23388 6316
rect 22879 6276 23388 6304
rect 22879 6273 22891 6276
rect 22833 6267 22891 6273
rect 23382 6264 23388 6276
rect 23440 6264 23446 6316
rect 9306 6236 9312 6248
rect 9140 6208 9312 6236
rect 9033 6199 9091 6205
rect 8021 6171 8079 6177
rect 8021 6137 8033 6171
rect 8067 6168 8079 6171
rect 8478 6168 8484 6180
rect 8067 6140 8484 6168
rect 8067 6137 8079 6140
rect 8021 6131 8079 6137
rect 8478 6128 8484 6140
rect 8536 6128 8542 6180
rect 9048 6168 9076 6199
rect 9306 6196 9312 6208
rect 9364 6196 9370 6248
rect 9950 6236 9956 6248
rect 9911 6208 9956 6236
rect 9950 6196 9956 6208
rect 10008 6196 10014 6248
rect 10781 6239 10839 6245
rect 10781 6205 10793 6239
rect 10827 6236 10839 6239
rect 11146 6236 11152 6248
rect 10827 6208 11152 6236
rect 10827 6205 10839 6208
rect 10781 6199 10839 6205
rect 11146 6196 11152 6208
rect 11204 6196 11210 6248
rect 11606 6236 11612 6248
rect 11567 6208 11612 6236
rect 11606 6196 11612 6208
rect 11664 6196 11670 6248
rect 12710 6196 12716 6248
rect 12768 6236 12774 6248
rect 12989 6239 13047 6245
rect 12989 6236 13001 6239
rect 12768 6208 13001 6236
rect 12768 6196 12774 6208
rect 12989 6205 13001 6208
rect 13035 6236 13047 6239
rect 13538 6236 13544 6248
rect 13035 6208 13544 6236
rect 13035 6205 13047 6208
rect 12989 6199 13047 6205
rect 13538 6196 13544 6208
rect 13596 6196 13602 6248
rect 13814 6236 13820 6248
rect 13775 6208 13820 6236
rect 13814 6196 13820 6208
rect 13872 6196 13878 6248
rect 13909 6239 13967 6245
rect 13909 6205 13921 6239
rect 13955 6205 13967 6239
rect 13909 6199 13967 6205
rect 15381 6239 15439 6245
rect 15381 6205 15393 6239
rect 15427 6205 15439 6239
rect 15381 6199 15439 6205
rect 15749 6239 15807 6245
rect 15749 6205 15761 6239
rect 15795 6236 15807 6239
rect 16298 6236 16304 6248
rect 15795 6208 16304 6236
rect 15795 6205 15807 6208
rect 15749 6199 15807 6205
rect 10042 6168 10048 6180
rect 9048 6140 10048 6168
rect 10042 6128 10048 6140
rect 10100 6128 10106 6180
rect 12253 6171 12311 6177
rect 12253 6137 12265 6171
rect 12299 6168 12311 6171
rect 13924 6168 13952 6199
rect 14366 6168 14372 6180
rect 12299 6140 13952 6168
rect 14327 6140 14372 6168
rect 12299 6137 12311 6140
rect 12253 6131 12311 6137
rect 14366 6128 14372 6140
rect 14424 6128 14430 6180
rect 15286 6128 15292 6180
rect 15344 6168 15350 6180
rect 15396 6168 15424 6199
rect 16298 6196 16304 6208
rect 16356 6196 16362 6248
rect 16666 6196 16672 6248
rect 16724 6236 16730 6248
rect 16761 6239 16819 6245
rect 16761 6236 16773 6239
rect 16724 6208 16773 6236
rect 16724 6196 16730 6208
rect 16761 6205 16773 6208
rect 16807 6205 16819 6239
rect 16761 6199 16819 6205
rect 16942 6196 16948 6248
rect 17000 6236 17006 6248
rect 17770 6236 17776 6248
rect 17000 6208 17776 6236
rect 17000 6196 17006 6208
rect 17770 6196 17776 6208
rect 17828 6196 17834 6248
rect 18049 6239 18107 6245
rect 18049 6236 18061 6239
rect 17880 6208 18061 6236
rect 15344 6140 15424 6168
rect 15344 6128 15350 6140
rect 17402 6128 17408 6180
rect 17460 6168 17466 6180
rect 17880 6168 17908 6208
rect 18049 6205 18061 6208
rect 18095 6205 18107 6239
rect 18966 6236 18972 6248
rect 18927 6208 18972 6236
rect 18049 6199 18107 6205
rect 18966 6196 18972 6208
rect 19024 6196 19030 6248
rect 19245 6239 19303 6245
rect 19245 6205 19257 6239
rect 19291 6205 19303 6239
rect 19245 6199 19303 6205
rect 17460 6140 17908 6168
rect 17460 6128 17466 6140
rect 17954 6128 17960 6180
rect 18012 6168 18018 6180
rect 18782 6168 18788 6180
rect 18012 6140 18788 6168
rect 18012 6128 18018 6140
rect 18782 6128 18788 6140
rect 18840 6128 18846 6180
rect 8113 6103 8171 6109
rect 8113 6069 8125 6103
rect 8159 6100 8171 6103
rect 8386 6100 8392 6112
rect 8159 6072 8392 6100
rect 8159 6069 8171 6072
rect 8113 6063 8171 6069
rect 8386 6060 8392 6072
rect 8444 6060 8450 6112
rect 9677 6103 9735 6109
rect 9677 6069 9689 6103
rect 9723 6100 9735 6103
rect 10410 6100 10416 6112
rect 9723 6072 10416 6100
rect 9723 6069 9735 6072
rect 9677 6063 9735 6069
rect 10410 6060 10416 6072
rect 10468 6060 10474 6112
rect 10505 6103 10563 6109
rect 10505 6069 10517 6103
rect 10551 6100 10563 6103
rect 11238 6100 11244 6112
rect 10551 6072 11244 6100
rect 10551 6069 10563 6072
rect 10505 6063 10563 6069
rect 11238 6060 11244 6072
rect 11296 6060 11302 6112
rect 11330 6060 11336 6112
rect 11388 6100 11394 6112
rect 11388 6072 11433 6100
rect 11388 6060 11394 6072
rect 14642 6060 14648 6112
rect 14700 6100 14706 6112
rect 14829 6103 14887 6109
rect 14829 6100 14841 6103
rect 14700 6072 14841 6100
rect 14700 6060 14706 6072
rect 14829 6069 14841 6072
rect 14875 6069 14887 6103
rect 14829 6063 14887 6069
rect 17034 6060 17040 6112
rect 17092 6100 17098 6112
rect 17497 6103 17555 6109
rect 17497 6100 17509 6103
rect 17092 6072 17509 6100
rect 17092 6060 17098 6072
rect 17497 6069 17509 6072
rect 17543 6069 17555 6103
rect 17497 6063 17555 6069
rect 17678 6060 17684 6112
rect 17736 6100 17742 6112
rect 18417 6103 18475 6109
rect 18417 6100 18429 6103
rect 17736 6072 18429 6100
rect 17736 6060 17742 6072
rect 18417 6069 18429 6072
rect 18463 6069 18475 6103
rect 19260 6100 19288 6199
rect 20530 6196 20536 6248
rect 20588 6236 20594 6248
rect 20809 6239 20867 6245
rect 20809 6236 20821 6239
rect 20588 6208 20821 6236
rect 20588 6196 20594 6208
rect 20809 6205 20821 6208
rect 20855 6205 20867 6239
rect 22278 6236 22284 6248
rect 22239 6208 22284 6236
rect 20809 6199 20867 6205
rect 22278 6196 22284 6208
rect 22336 6196 22342 6248
rect 22370 6196 22376 6248
rect 22428 6236 22434 6248
rect 22428 6208 22473 6236
rect 22428 6196 22434 6208
rect 21545 6171 21603 6177
rect 21545 6168 21557 6171
rect 20640 6140 21557 6168
rect 20640 6112 20668 6140
rect 21545 6137 21557 6140
rect 21591 6168 21603 6171
rect 22646 6168 22652 6180
rect 21591 6140 22652 6168
rect 21591 6137 21603 6140
rect 21545 6131 21603 6137
rect 22646 6128 22652 6140
rect 22704 6128 22710 6180
rect 20346 6100 20352 6112
rect 19260 6072 20352 6100
rect 18417 6063 18475 6069
rect 20346 6060 20352 6072
rect 20404 6100 20410 6112
rect 20622 6100 20628 6112
rect 20404 6072 20628 6100
rect 20404 6060 20410 6072
rect 20622 6060 20628 6072
rect 20680 6060 20686 6112
rect 21910 6060 21916 6112
rect 21968 6100 21974 6112
rect 22830 6100 22836 6112
rect 21968 6072 22836 6100
rect 21968 6060 21974 6072
rect 22830 6060 22836 6072
rect 22888 6060 22894 6112
rect 23014 6100 23020 6112
rect 22975 6072 23020 6100
rect 23014 6060 23020 6072
rect 23072 6060 23078 6112
rect 1104 6010 23460 6032
rect 1104 5958 3749 6010
rect 3801 5958 3813 6010
rect 3865 5958 3877 6010
rect 3929 5958 3941 6010
rect 3993 5958 4005 6010
rect 4057 5958 9347 6010
rect 9399 5958 9411 6010
rect 9463 5958 9475 6010
rect 9527 5958 9539 6010
rect 9591 5958 9603 6010
rect 9655 5958 14945 6010
rect 14997 5958 15009 6010
rect 15061 5958 15073 6010
rect 15125 5958 15137 6010
rect 15189 5958 15201 6010
rect 15253 5958 20543 6010
rect 20595 5958 20607 6010
rect 20659 5958 20671 6010
rect 20723 5958 20735 6010
rect 20787 5958 20799 6010
rect 20851 5958 23460 6010
rect 1104 5936 23460 5958
rect 9861 5899 9919 5905
rect 9861 5896 9873 5899
rect 8588 5868 9873 5896
rect 7929 5831 7987 5837
rect 7929 5797 7941 5831
rect 7975 5828 7987 5831
rect 8294 5828 8300 5840
rect 7975 5800 8300 5828
rect 7975 5797 7987 5800
rect 7929 5791 7987 5797
rect 8294 5788 8300 5800
rect 8352 5788 8358 5840
rect 7374 5760 7380 5772
rect 7335 5732 7380 5760
rect 7374 5720 7380 5732
rect 7432 5720 7438 5772
rect 8205 5763 8263 5769
rect 8205 5729 8217 5763
rect 8251 5760 8263 5763
rect 8588 5760 8616 5868
rect 9861 5865 9873 5868
rect 9907 5896 9919 5899
rect 10042 5896 10048 5908
rect 9907 5868 10048 5896
rect 9907 5865 9919 5868
rect 9861 5859 9919 5865
rect 10042 5856 10048 5868
rect 10100 5856 10106 5908
rect 10962 5856 10968 5908
rect 11020 5896 11026 5908
rect 12069 5899 12127 5905
rect 12069 5896 12081 5899
rect 11020 5868 12081 5896
rect 11020 5856 11026 5868
rect 12069 5865 12081 5868
rect 12115 5865 12127 5899
rect 12069 5859 12127 5865
rect 13909 5899 13967 5905
rect 13909 5865 13921 5899
rect 13955 5896 13967 5899
rect 13955 5868 16344 5896
rect 13955 5865 13967 5868
rect 13909 5859 13967 5865
rect 8757 5831 8815 5837
rect 8757 5797 8769 5831
rect 8803 5828 8815 5831
rect 8803 5800 9904 5828
rect 8803 5797 8815 5800
rect 8757 5791 8815 5797
rect 8251 5732 8616 5760
rect 8251 5729 8263 5732
rect 8205 5723 8263 5729
rect 8662 5720 8668 5772
rect 8720 5760 8726 5772
rect 9401 5763 9459 5769
rect 9401 5760 9413 5763
rect 8720 5732 9413 5760
rect 8720 5720 8726 5732
rect 9401 5729 9413 5732
rect 9447 5729 9459 5763
rect 9401 5723 9459 5729
rect 9490 5720 9496 5772
rect 9548 5760 9554 5772
rect 9548 5732 9593 5760
rect 9548 5720 9554 5732
rect 7190 5652 7196 5704
rect 7248 5692 7254 5704
rect 7561 5695 7619 5701
rect 7561 5692 7573 5695
rect 7248 5664 7573 5692
rect 7248 5652 7254 5664
rect 7561 5661 7573 5664
rect 7607 5661 7619 5695
rect 8386 5692 8392 5704
rect 8347 5664 8392 5692
rect 7561 5655 7619 5661
rect 8386 5652 8392 5664
rect 8444 5652 8450 5704
rect 9309 5695 9367 5701
rect 9309 5661 9321 5695
rect 9355 5692 9367 5695
rect 9766 5692 9772 5704
rect 9355 5664 9772 5692
rect 9355 5661 9367 5664
rect 9309 5655 9367 5661
rect 9766 5652 9772 5664
rect 9824 5652 9830 5704
rect 7469 5627 7527 5633
rect 7469 5593 7481 5627
rect 7515 5624 7527 5627
rect 8570 5624 8576 5636
rect 7515 5596 8576 5624
rect 7515 5593 7527 5596
rect 7469 5587 7527 5593
rect 8570 5584 8576 5596
rect 8628 5584 8634 5636
rect 9582 5624 9588 5636
rect 8680 5596 9588 5624
rect 8297 5559 8355 5565
rect 8297 5525 8309 5559
rect 8343 5556 8355 5559
rect 8680 5556 8708 5596
rect 9582 5584 9588 5596
rect 9640 5584 9646 5636
rect 9876 5624 9904 5800
rect 9950 5788 9956 5840
rect 10008 5828 10014 5840
rect 10008 5800 12756 5828
rect 10008 5788 10014 5800
rect 10612 5769 10640 5800
rect 12728 5772 12756 5800
rect 10597 5763 10655 5769
rect 10597 5729 10609 5763
rect 10643 5729 10655 5763
rect 10597 5723 10655 5729
rect 10686 5720 10692 5772
rect 10744 5760 10750 5772
rect 10744 5732 10789 5760
rect 10744 5720 10750 5732
rect 11146 5720 11152 5772
rect 11204 5760 11210 5772
rect 11333 5763 11391 5769
rect 11333 5760 11345 5763
rect 11204 5732 11345 5760
rect 11204 5720 11210 5732
rect 11333 5729 11345 5732
rect 11379 5729 11391 5763
rect 12710 5760 12716 5772
rect 12671 5732 12716 5760
rect 11333 5723 11391 5729
rect 12710 5720 12716 5732
rect 12768 5720 12774 5772
rect 14556 5763 14614 5769
rect 14556 5729 14568 5763
rect 14602 5760 14614 5763
rect 14642 5760 14648 5772
rect 14602 5732 14648 5760
rect 14602 5729 14614 5732
rect 14556 5723 14614 5729
rect 14642 5720 14648 5732
rect 14700 5720 14706 5772
rect 14752 5732 16068 5760
rect 10781 5695 10839 5701
rect 10781 5661 10793 5695
rect 10827 5692 10839 5695
rect 10870 5692 10876 5704
rect 10827 5664 10876 5692
rect 10827 5661 10839 5664
rect 10781 5655 10839 5661
rect 10870 5652 10876 5664
rect 10928 5652 10934 5704
rect 11238 5652 11244 5704
rect 11296 5692 11302 5704
rect 11609 5695 11667 5701
rect 11609 5692 11621 5695
rect 11296 5664 11621 5692
rect 11296 5652 11302 5664
rect 11609 5661 11621 5664
rect 11655 5661 11667 5695
rect 13725 5695 13783 5701
rect 13725 5692 13737 5695
rect 11609 5655 11667 5661
rect 11716 5664 13737 5692
rect 11716 5624 11744 5664
rect 13725 5661 13737 5664
rect 13771 5661 13783 5695
rect 13725 5655 13783 5661
rect 14093 5695 14151 5701
rect 14093 5661 14105 5695
rect 14139 5692 14151 5695
rect 14752 5692 14780 5732
rect 14139 5664 14780 5692
rect 14829 5695 14887 5701
rect 14139 5661 14151 5664
rect 14093 5655 14151 5661
rect 14829 5661 14841 5695
rect 14875 5692 14887 5695
rect 15102 5692 15108 5704
rect 14875 5664 15108 5692
rect 14875 5661 14887 5664
rect 14829 5655 14887 5661
rect 15102 5652 15108 5664
rect 15160 5652 15166 5704
rect 12437 5627 12495 5633
rect 12437 5624 12449 5627
rect 9876 5596 11744 5624
rect 11808 5596 12449 5624
rect 8938 5556 8944 5568
rect 8343 5528 8708 5556
rect 8899 5528 8944 5556
rect 8343 5525 8355 5528
rect 8297 5519 8355 5525
rect 8938 5516 8944 5528
rect 8996 5516 9002 5568
rect 11149 5559 11207 5565
rect 11149 5525 11161 5559
rect 11195 5556 11207 5559
rect 11517 5559 11575 5565
rect 11517 5556 11529 5559
rect 11195 5528 11529 5556
rect 11195 5525 11207 5528
rect 11149 5519 11207 5525
rect 11517 5525 11529 5528
rect 11563 5525 11575 5559
rect 11517 5519 11575 5525
rect 11606 5516 11612 5568
rect 11664 5556 11670 5568
rect 11808 5556 11836 5596
rect 12437 5593 12449 5596
rect 12483 5593 12495 5627
rect 12437 5587 12495 5593
rect 12529 5627 12587 5633
rect 12529 5593 12541 5627
rect 12575 5624 12587 5627
rect 12618 5624 12624 5636
rect 12575 5596 12624 5624
rect 12575 5593 12587 5596
rect 12529 5587 12587 5593
rect 12618 5584 12624 5596
rect 12676 5584 12682 5636
rect 16040 5624 16068 5732
rect 16114 5720 16120 5772
rect 16172 5760 16178 5772
rect 16316 5769 16344 5868
rect 17586 5856 17592 5908
rect 17644 5896 17650 5908
rect 17681 5899 17739 5905
rect 17681 5896 17693 5899
rect 17644 5868 17693 5896
rect 17644 5856 17650 5868
rect 17681 5865 17693 5868
rect 17727 5865 17739 5899
rect 17681 5859 17739 5865
rect 17770 5856 17776 5908
rect 17828 5896 17834 5908
rect 20901 5899 20959 5905
rect 20901 5896 20913 5899
rect 17828 5868 20913 5896
rect 17828 5856 17834 5868
rect 20901 5865 20913 5868
rect 20947 5865 20959 5899
rect 20901 5859 20959 5865
rect 21542 5856 21548 5908
rect 21600 5896 21606 5908
rect 21729 5899 21787 5905
rect 21729 5896 21741 5899
rect 21600 5868 21741 5896
rect 21600 5856 21606 5868
rect 21729 5865 21741 5868
rect 21775 5865 21787 5899
rect 22646 5896 22652 5908
rect 22607 5868 22652 5896
rect 21729 5859 21787 5865
rect 22646 5856 22652 5868
rect 22704 5856 22710 5908
rect 16761 5831 16819 5837
rect 16761 5797 16773 5831
rect 16807 5828 16819 5831
rect 20806 5828 20812 5840
rect 16807 5800 20812 5828
rect 16807 5797 16819 5800
rect 16761 5791 16819 5797
rect 20806 5788 20812 5800
rect 20864 5788 20870 5840
rect 22094 5788 22100 5840
rect 22152 5828 22158 5840
rect 22281 5831 22339 5837
rect 22281 5828 22293 5831
rect 22152 5800 22293 5828
rect 22152 5788 22158 5800
rect 22281 5797 22293 5800
rect 22327 5797 22339 5831
rect 23474 5828 23480 5840
rect 22281 5791 22339 5797
rect 22388 5800 23480 5828
rect 16301 5763 16359 5769
rect 16172 5732 16217 5760
rect 16172 5720 16178 5732
rect 16301 5729 16313 5763
rect 16347 5729 16359 5763
rect 16301 5723 16359 5729
rect 16574 5720 16580 5772
rect 16632 5760 16638 5772
rect 16945 5763 17003 5769
rect 16945 5760 16957 5763
rect 16632 5732 16957 5760
rect 16632 5720 16638 5732
rect 16945 5729 16957 5732
rect 16991 5729 17003 5763
rect 18230 5760 18236 5772
rect 18191 5732 18236 5760
rect 16945 5723 17003 5729
rect 18230 5720 18236 5732
rect 18288 5720 18294 5772
rect 18506 5760 18512 5772
rect 18467 5732 18512 5760
rect 18506 5720 18512 5732
rect 18564 5720 18570 5772
rect 19794 5760 19800 5772
rect 19755 5732 19800 5760
rect 19794 5720 19800 5732
rect 19852 5720 19858 5772
rect 20070 5720 20076 5772
rect 20128 5760 20134 5772
rect 20165 5763 20223 5769
rect 20165 5760 20177 5763
rect 20128 5732 20177 5760
rect 20128 5720 20134 5732
rect 20165 5729 20177 5732
rect 20211 5729 20223 5763
rect 20165 5723 20223 5729
rect 21450 5720 21456 5772
rect 21508 5760 21514 5772
rect 22388 5760 22416 5800
rect 23474 5788 23480 5800
rect 23532 5788 23538 5840
rect 23198 5760 23204 5772
rect 21508 5732 21553 5760
rect 21836 5732 22416 5760
rect 22480 5732 23204 5760
rect 21508 5720 21514 5732
rect 16390 5692 16396 5704
rect 16351 5664 16396 5692
rect 16390 5652 16396 5664
rect 16448 5652 16454 5704
rect 17221 5695 17279 5701
rect 17221 5661 17233 5695
rect 17267 5692 17279 5695
rect 18414 5692 18420 5704
rect 17267 5664 18420 5692
rect 17267 5661 17279 5664
rect 17221 5655 17279 5661
rect 18414 5652 18420 5664
rect 18472 5652 18478 5704
rect 19334 5652 19340 5704
rect 19392 5692 19398 5704
rect 21361 5695 21419 5701
rect 19392 5664 19748 5692
rect 19392 5652 19398 5664
rect 17310 5624 17316 5636
rect 16040 5596 17316 5624
rect 17310 5584 17316 5596
rect 17368 5584 17374 5636
rect 18049 5627 18107 5633
rect 18049 5593 18061 5627
rect 18095 5624 18107 5627
rect 18322 5624 18328 5636
rect 18095 5596 18328 5624
rect 18095 5593 18107 5596
rect 18049 5587 18107 5593
rect 18322 5584 18328 5596
rect 18380 5584 18386 5636
rect 19061 5627 19119 5633
rect 19061 5593 19073 5627
rect 19107 5624 19119 5627
rect 19613 5627 19671 5633
rect 19613 5624 19625 5627
rect 19107 5596 19625 5624
rect 19107 5593 19119 5596
rect 19061 5587 19119 5593
rect 19613 5593 19625 5596
rect 19659 5593 19671 5627
rect 19720 5624 19748 5664
rect 21361 5661 21373 5695
rect 21407 5692 21419 5695
rect 21836 5692 21864 5732
rect 21407 5664 21864 5692
rect 21913 5695 21971 5701
rect 21407 5661 21419 5664
rect 21361 5655 21419 5661
rect 21913 5661 21925 5695
rect 21959 5692 21971 5695
rect 22480 5692 22508 5732
rect 23198 5720 23204 5732
rect 23256 5720 23262 5772
rect 21959 5664 22508 5692
rect 21959 5661 21971 5664
rect 21913 5655 21971 5661
rect 22554 5652 22560 5704
rect 22612 5692 22618 5704
rect 22833 5695 22891 5701
rect 22833 5692 22845 5695
rect 22612 5664 22845 5692
rect 22612 5652 22618 5664
rect 22833 5661 22845 5664
rect 22879 5661 22891 5695
rect 22833 5655 22891 5661
rect 20349 5627 20407 5633
rect 20349 5624 20361 5627
rect 19720 5596 20361 5624
rect 19613 5587 19671 5593
rect 20349 5593 20361 5596
rect 20395 5593 20407 5627
rect 20349 5587 20407 5593
rect 21269 5627 21327 5633
rect 21269 5593 21281 5627
rect 21315 5624 21327 5627
rect 22005 5627 22063 5633
rect 22005 5624 22017 5627
rect 21315 5596 22017 5624
rect 21315 5593 21327 5596
rect 21269 5587 21327 5593
rect 22005 5593 22017 5596
rect 22051 5593 22063 5627
rect 22005 5587 22063 5593
rect 22465 5627 22523 5633
rect 22465 5593 22477 5627
rect 22511 5624 22523 5627
rect 23106 5624 23112 5636
rect 22511 5596 23112 5624
rect 22511 5593 22523 5596
rect 22465 5587 22523 5593
rect 23106 5584 23112 5596
rect 23164 5584 23170 5636
rect 11974 5556 11980 5568
rect 11664 5528 11836 5556
rect 11935 5528 11980 5556
rect 11664 5516 11670 5528
rect 11974 5516 11980 5528
rect 12032 5516 12038 5568
rect 13633 5559 13691 5565
rect 13633 5525 13645 5559
rect 13679 5556 13691 5559
rect 13814 5556 13820 5568
rect 13679 5528 13820 5556
rect 13679 5525 13691 5528
rect 13633 5519 13691 5525
rect 13814 5516 13820 5528
rect 13872 5556 13878 5568
rect 14550 5556 14556 5568
rect 14608 5565 14614 5568
rect 13872 5528 14556 5556
rect 13872 5516 13878 5528
rect 14550 5516 14556 5528
rect 14608 5556 14617 5565
rect 15933 5559 15991 5565
rect 14608 5528 14653 5556
rect 14608 5519 14617 5528
rect 15933 5525 15945 5559
rect 15979 5556 15991 5559
rect 16666 5556 16672 5568
rect 15979 5528 16672 5556
rect 15979 5525 15991 5528
rect 15933 5519 15991 5525
rect 14608 5516 14614 5519
rect 16666 5516 16672 5528
rect 16724 5516 16730 5568
rect 17126 5556 17132 5568
rect 17087 5528 17132 5556
rect 17126 5516 17132 5528
rect 17184 5516 17190 5568
rect 17218 5516 17224 5568
rect 17276 5556 17282 5568
rect 17589 5559 17647 5565
rect 17589 5556 17601 5559
rect 17276 5528 17601 5556
rect 17276 5516 17282 5528
rect 17589 5525 17601 5528
rect 17635 5525 17647 5559
rect 17589 5519 17647 5525
rect 17954 5516 17960 5568
rect 18012 5556 18018 5568
rect 18141 5559 18199 5565
rect 18141 5556 18153 5559
rect 18012 5528 18153 5556
rect 18012 5516 18018 5528
rect 18141 5525 18153 5528
rect 18187 5525 18199 5559
rect 18141 5519 18199 5525
rect 18230 5516 18236 5568
rect 18288 5556 18294 5568
rect 19245 5559 19303 5565
rect 19245 5556 19257 5559
rect 18288 5528 19257 5556
rect 18288 5516 18294 5528
rect 19245 5525 19257 5528
rect 19291 5525 19303 5559
rect 19702 5556 19708 5568
rect 19663 5528 19708 5556
rect 19245 5519 19303 5525
rect 19702 5516 19708 5528
rect 19760 5516 19766 5568
rect 20438 5516 20444 5568
rect 20496 5556 20502 5568
rect 20809 5559 20867 5565
rect 20496 5528 20541 5556
rect 20496 5516 20502 5528
rect 20809 5525 20821 5559
rect 20855 5556 20867 5559
rect 21726 5556 21732 5568
rect 20855 5528 21732 5556
rect 20855 5525 20867 5528
rect 20809 5519 20867 5525
rect 21726 5516 21732 5528
rect 21784 5556 21790 5568
rect 22646 5556 22652 5568
rect 21784 5528 22652 5556
rect 21784 5516 21790 5528
rect 22646 5516 22652 5528
rect 22704 5516 22710 5568
rect 23014 5556 23020 5568
rect 22975 5528 23020 5556
rect 23014 5516 23020 5528
rect 23072 5516 23078 5568
rect 1104 5466 23460 5488
rect 1104 5414 6548 5466
rect 6600 5414 6612 5466
rect 6664 5414 6676 5466
rect 6728 5414 6740 5466
rect 6792 5414 6804 5466
rect 6856 5414 12146 5466
rect 12198 5414 12210 5466
rect 12262 5414 12274 5466
rect 12326 5414 12338 5466
rect 12390 5414 12402 5466
rect 12454 5414 17744 5466
rect 17796 5414 17808 5466
rect 17860 5414 17872 5466
rect 17924 5414 17936 5466
rect 17988 5414 18000 5466
rect 18052 5414 23460 5466
rect 1104 5392 23460 5414
rect 8205 5355 8263 5361
rect 8205 5321 8217 5355
rect 8251 5352 8263 5355
rect 8757 5355 8815 5361
rect 8757 5352 8769 5355
rect 8251 5324 8769 5352
rect 8251 5321 8263 5324
rect 8205 5315 8263 5321
rect 8757 5321 8769 5324
rect 8803 5321 8815 5355
rect 9122 5352 9128 5364
rect 9083 5324 9128 5352
rect 8757 5315 8815 5321
rect 9122 5312 9128 5324
rect 9180 5312 9186 5364
rect 9677 5355 9735 5361
rect 9677 5321 9689 5355
rect 9723 5352 9735 5355
rect 10042 5352 10048 5364
rect 9723 5324 10048 5352
rect 9723 5321 9735 5324
rect 9677 5315 9735 5321
rect 10042 5312 10048 5324
rect 10100 5312 10106 5364
rect 12066 5312 12072 5364
rect 12124 5352 12130 5364
rect 12253 5355 12311 5361
rect 12253 5352 12265 5355
rect 12124 5324 12265 5352
rect 12124 5312 12130 5324
rect 12253 5321 12265 5324
rect 12299 5321 12311 5355
rect 12253 5315 12311 5321
rect 12345 5355 12403 5361
rect 12345 5321 12357 5355
rect 12391 5352 12403 5355
rect 13170 5352 13176 5364
rect 12391 5324 13176 5352
rect 12391 5321 12403 5324
rect 12345 5315 12403 5321
rect 13170 5312 13176 5324
rect 13228 5312 13234 5364
rect 15013 5355 15071 5361
rect 15013 5321 15025 5355
rect 15059 5321 15071 5355
rect 15378 5352 15384 5364
rect 15339 5324 15384 5352
rect 15013 5315 15071 5321
rect 8297 5287 8355 5293
rect 8297 5253 8309 5287
rect 8343 5284 8355 5287
rect 8938 5284 8944 5296
rect 8343 5256 8944 5284
rect 8343 5253 8355 5256
rect 8297 5247 8355 5253
rect 8938 5244 8944 5256
rect 8996 5244 9002 5296
rect 14369 5287 14427 5293
rect 14369 5253 14381 5287
rect 14415 5284 14427 5287
rect 14550 5284 14556 5296
rect 14415 5256 14556 5284
rect 14415 5253 14427 5256
rect 14369 5247 14427 5253
rect 14550 5244 14556 5256
rect 14608 5244 14614 5296
rect 15028 5284 15056 5315
rect 15378 5312 15384 5324
rect 15436 5312 15442 5364
rect 15654 5352 15660 5364
rect 15615 5324 15660 5352
rect 15654 5312 15660 5324
rect 15712 5312 15718 5364
rect 16942 5312 16948 5364
rect 17000 5352 17006 5364
rect 17037 5355 17095 5361
rect 17037 5352 17049 5355
rect 17000 5324 17049 5352
rect 17000 5312 17006 5324
rect 17037 5321 17049 5324
rect 17083 5321 17095 5355
rect 17037 5315 17095 5321
rect 17126 5312 17132 5364
rect 17184 5352 17190 5364
rect 17405 5355 17463 5361
rect 17405 5352 17417 5355
rect 17184 5324 17417 5352
rect 17184 5312 17190 5324
rect 17405 5321 17417 5324
rect 17451 5321 17463 5355
rect 17405 5315 17463 5321
rect 17586 5312 17592 5364
rect 17644 5352 17650 5364
rect 17957 5355 18015 5361
rect 17957 5352 17969 5355
rect 17644 5324 17969 5352
rect 17644 5312 17650 5324
rect 17957 5321 17969 5324
rect 18003 5321 18015 5355
rect 17957 5315 18015 5321
rect 19153 5355 19211 5361
rect 19153 5321 19165 5355
rect 19199 5352 19211 5355
rect 19334 5352 19340 5364
rect 19199 5324 19340 5352
rect 19199 5321 19211 5324
rect 19153 5315 19211 5321
rect 19334 5312 19340 5324
rect 19392 5312 19398 5364
rect 19702 5312 19708 5364
rect 19760 5352 19766 5364
rect 20073 5355 20131 5361
rect 20073 5352 20085 5355
rect 19760 5324 20085 5352
rect 19760 5312 19766 5324
rect 20073 5321 20085 5324
rect 20119 5321 20131 5355
rect 22189 5355 22247 5361
rect 22189 5352 22201 5355
rect 20073 5315 20131 5321
rect 20180 5324 22201 5352
rect 16390 5284 16396 5296
rect 15028 5256 16396 5284
rect 16390 5244 16396 5256
rect 16448 5244 16454 5296
rect 16574 5244 16580 5296
rect 16632 5284 16638 5296
rect 17494 5284 17500 5296
rect 16632 5256 17500 5284
rect 16632 5244 16638 5256
rect 17494 5244 17500 5256
rect 17552 5244 17558 5296
rect 17865 5287 17923 5293
rect 17865 5253 17877 5287
rect 17911 5284 17923 5287
rect 18690 5284 18696 5296
rect 17911 5256 18696 5284
rect 17911 5253 17923 5256
rect 17865 5247 17923 5253
rect 18690 5244 18696 5256
rect 18748 5244 18754 5296
rect 19058 5244 19064 5296
rect 19116 5284 19122 5296
rect 20180 5284 20208 5324
rect 22189 5321 22201 5324
rect 22235 5321 22247 5355
rect 22738 5352 22744 5364
rect 22699 5324 22744 5352
rect 22189 5315 22247 5321
rect 22738 5312 22744 5324
rect 22796 5312 22802 5364
rect 19116 5256 20208 5284
rect 19116 5244 19122 5256
rect 20254 5244 20260 5296
rect 20312 5284 20318 5296
rect 20312 5256 20668 5284
rect 20312 5244 20318 5256
rect 8846 5176 8852 5228
rect 8904 5216 8910 5228
rect 9217 5219 9275 5225
rect 9217 5216 9229 5219
rect 8904 5188 9229 5216
rect 8904 5176 8910 5188
rect 9217 5185 9229 5188
rect 9263 5185 9275 5219
rect 14826 5216 14832 5228
rect 14787 5188 14832 5216
rect 9217 5179 9275 5185
rect 14826 5176 14832 5188
rect 14884 5176 14890 5228
rect 15105 5219 15163 5225
rect 15105 5185 15117 5219
rect 15151 5185 15163 5219
rect 15105 5179 15163 5185
rect 8110 5148 8116 5160
rect 8071 5120 8116 5148
rect 8110 5108 8116 5120
rect 8168 5108 8174 5160
rect 9306 5108 9312 5160
rect 9364 5148 9370 5160
rect 9364 5120 9409 5148
rect 9364 5108 9370 5120
rect 11146 5108 11152 5160
rect 11204 5148 11210 5160
rect 11790 5148 11796 5160
rect 11204 5120 11796 5148
rect 11204 5108 11210 5120
rect 11790 5108 11796 5120
rect 11848 5148 11854 5160
rect 12069 5151 12127 5157
rect 12069 5148 12081 5151
rect 11848 5120 12081 5148
rect 11848 5108 11854 5120
rect 12069 5117 12081 5120
rect 12115 5117 12127 5151
rect 12069 5111 12127 5117
rect 8665 5083 8723 5089
rect 8665 5049 8677 5083
rect 8711 5080 8723 5083
rect 15120 5080 15148 5179
rect 15194 5176 15200 5228
rect 15252 5216 15258 5228
rect 16022 5216 16028 5228
rect 15252 5188 16028 5216
rect 15252 5176 15258 5188
rect 16022 5176 16028 5188
rect 16080 5176 16086 5228
rect 16117 5219 16175 5225
rect 16117 5185 16129 5219
rect 16163 5216 16175 5219
rect 16776 5216 16896 5220
rect 18230 5216 18236 5228
rect 16163 5192 18236 5216
rect 16163 5188 16804 5192
rect 16868 5188 18236 5192
rect 16163 5185 16175 5188
rect 16117 5179 16175 5185
rect 18230 5176 18236 5188
rect 18288 5176 18294 5228
rect 18782 5216 18788 5228
rect 18743 5188 18788 5216
rect 18782 5176 18788 5188
rect 18840 5176 18846 5228
rect 18966 5176 18972 5228
rect 19024 5216 19030 5228
rect 19613 5219 19671 5225
rect 19613 5216 19625 5219
rect 19024 5188 19625 5216
rect 19024 5176 19030 5188
rect 19613 5185 19625 5188
rect 19659 5185 19671 5219
rect 19613 5179 19671 5185
rect 19886 5176 19892 5228
rect 19944 5216 19950 5228
rect 20441 5219 20499 5225
rect 20441 5216 20453 5219
rect 19944 5188 20453 5216
rect 19944 5176 19950 5188
rect 20441 5185 20453 5188
rect 20487 5185 20499 5219
rect 20441 5179 20499 5185
rect 16206 5148 16212 5160
rect 16167 5120 16212 5148
rect 16206 5108 16212 5120
rect 16264 5108 16270 5160
rect 16574 5108 16580 5160
rect 16632 5148 16638 5160
rect 16761 5151 16819 5157
rect 16761 5148 16773 5151
rect 16632 5120 16773 5148
rect 16632 5108 16638 5120
rect 16761 5117 16773 5120
rect 16807 5117 16819 5151
rect 16761 5111 16819 5117
rect 16850 5108 16856 5160
rect 16908 5148 16914 5160
rect 16945 5151 17003 5157
rect 16945 5148 16957 5151
rect 16908 5120 16957 5148
rect 16908 5108 16914 5120
rect 16945 5117 16957 5120
rect 16991 5117 17003 5151
rect 16945 5111 17003 5117
rect 17402 5108 17408 5160
rect 17460 5148 17466 5160
rect 18049 5151 18107 5157
rect 18049 5148 18061 5151
rect 17460 5120 18061 5148
rect 17460 5108 17466 5120
rect 18049 5117 18061 5120
rect 18095 5117 18107 5151
rect 18598 5148 18604 5160
rect 18559 5120 18604 5148
rect 18049 5111 18107 5117
rect 18598 5108 18604 5120
rect 18656 5108 18662 5160
rect 18693 5151 18751 5157
rect 18693 5117 18705 5151
rect 18739 5117 18751 5151
rect 19426 5148 19432 5160
rect 19387 5120 19432 5148
rect 18693 5111 18751 5117
rect 17126 5080 17132 5092
rect 8711 5052 15148 5080
rect 15212 5052 17132 5080
rect 8711 5049 8723 5052
rect 8665 5043 8723 5049
rect 12713 5015 12771 5021
rect 12713 4981 12725 5015
rect 12759 5012 12771 5015
rect 14182 5012 14188 5024
rect 12759 4984 14188 5012
rect 12759 4981 12771 4984
rect 12713 4975 12771 4981
rect 14182 4972 14188 4984
rect 14240 4972 14246 5024
rect 14645 5015 14703 5021
rect 14645 4981 14657 5015
rect 14691 5012 14703 5015
rect 15212 5012 15240 5052
rect 17126 5040 17132 5052
rect 17184 5040 17190 5092
rect 18708 5080 18736 5111
rect 19426 5108 19432 5120
rect 19484 5108 19490 5160
rect 19518 5108 19524 5160
rect 19576 5148 19582 5160
rect 20640 5157 20668 5256
rect 20806 5244 20812 5296
rect 20864 5284 20870 5296
rect 22281 5287 22339 5293
rect 22281 5284 22293 5287
rect 20864 5256 22293 5284
rect 20864 5244 20870 5256
rect 22281 5253 22293 5256
rect 22327 5253 22339 5287
rect 22281 5247 22339 5253
rect 21266 5216 21272 5228
rect 21227 5188 21272 5216
rect 21266 5176 21272 5188
rect 21324 5176 21330 5228
rect 22830 5216 22836 5228
rect 22791 5188 22836 5216
rect 22830 5176 22836 5188
rect 22888 5176 22894 5228
rect 20533 5151 20591 5157
rect 20533 5148 20545 5151
rect 19576 5120 19621 5148
rect 19720 5120 20545 5148
rect 19576 5108 19582 5120
rect 17328 5052 18736 5080
rect 14691 4984 15240 5012
rect 15289 5015 15347 5021
rect 14691 4981 14703 4984
rect 14645 4975 14703 4981
rect 15289 4981 15301 5015
rect 15335 5012 15347 5015
rect 15654 5012 15660 5024
rect 15335 4984 15660 5012
rect 15335 4981 15347 4984
rect 15289 4975 15347 4981
rect 15654 4972 15660 4984
rect 15712 4972 15718 5024
rect 16022 4972 16028 5024
rect 16080 5012 16086 5024
rect 17328 5012 17356 5052
rect 17494 5012 17500 5024
rect 16080 4984 17356 5012
rect 17455 4984 17500 5012
rect 16080 4972 16086 4984
rect 17494 4972 17500 4984
rect 17552 4972 17558 5024
rect 18708 5012 18736 5052
rect 19334 5040 19340 5092
rect 19392 5080 19398 5092
rect 19720 5080 19748 5120
rect 20533 5117 20545 5120
rect 20579 5117 20591 5151
rect 20533 5111 20591 5117
rect 20625 5151 20683 5157
rect 20625 5117 20637 5151
rect 20671 5117 20683 5151
rect 20625 5111 20683 5117
rect 20898 5108 20904 5160
rect 20956 5148 20962 5160
rect 20993 5151 21051 5157
rect 20993 5148 21005 5151
rect 20956 5120 21005 5148
rect 20956 5108 20962 5120
rect 20993 5117 21005 5120
rect 21039 5117 21051 5151
rect 20993 5111 21051 5117
rect 21177 5151 21235 5157
rect 21177 5117 21189 5151
rect 21223 5117 21235 5151
rect 21177 5111 21235 5117
rect 19392 5052 19748 5080
rect 19812 5052 20107 5080
rect 19392 5040 19398 5052
rect 19812 5012 19840 5052
rect 19978 5012 19984 5024
rect 18708 4984 19840 5012
rect 19939 4984 19984 5012
rect 19978 4972 19984 4984
rect 20036 4972 20042 5024
rect 20079 5012 20107 5052
rect 20254 5040 20260 5092
rect 20312 5080 20318 5092
rect 21192 5080 21220 5111
rect 22370 5108 22376 5160
rect 22428 5148 22434 5160
rect 22428 5120 22473 5148
rect 22428 5108 22434 5120
rect 21634 5080 21640 5092
rect 20312 5052 21220 5080
rect 21595 5052 21640 5080
rect 20312 5040 20318 5052
rect 21634 5040 21640 5052
rect 21692 5080 21698 5092
rect 22554 5080 22560 5092
rect 21692 5052 22560 5080
rect 21692 5040 21698 5052
rect 22554 5040 22560 5052
rect 22612 5040 22618 5092
rect 21450 5012 21456 5024
rect 20079 4984 21456 5012
rect 21450 4972 21456 4984
rect 21508 4972 21514 5024
rect 21818 5012 21824 5024
rect 21779 4984 21824 5012
rect 21818 4972 21824 4984
rect 21876 4972 21882 5024
rect 23014 5012 23020 5024
rect 22975 4984 23020 5012
rect 23014 4972 23020 4984
rect 23072 4972 23078 5024
rect 1104 4922 23460 4944
rect 1104 4870 3749 4922
rect 3801 4870 3813 4922
rect 3865 4870 3877 4922
rect 3929 4870 3941 4922
rect 3993 4870 4005 4922
rect 4057 4870 9347 4922
rect 9399 4870 9411 4922
rect 9463 4870 9475 4922
rect 9527 4870 9539 4922
rect 9591 4870 9603 4922
rect 9655 4870 14945 4922
rect 14997 4870 15009 4922
rect 15061 4870 15073 4922
rect 15125 4870 15137 4922
rect 15189 4870 15201 4922
rect 15253 4870 20543 4922
rect 20595 4870 20607 4922
rect 20659 4870 20671 4922
rect 20723 4870 20735 4922
rect 20787 4870 20799 4922
rect 20851 4870 23460 4922
rect 1104 4848 23460 4870
rect 8757 4811 8815 4817
rect 8757 4777 8769 4811
rect 8803 4808 8815 4811
rect 14826 4808 14832 4820
rect 8803 4780 14832 4808
rect 8803 4777 8815 4780
rect 8757 4771 8815 4777
rect 14826 4768 14832 4780
rect 14884 4768 14890 4820
rect 18325 4811 18383 4817
rect 18325 4777 18337 4811
rect 18371 4808 18383 4811
rect 19518 4808 19524 4820
rect 18371 4780 19524 4808
rect 18371 4777 18383 4780
rect 18325 4771 18383 4777
rect 19518 4768 19524 4780
rect 19576 4768 19582 4820
rect 19981 4811 20039 4817
rect 19981 4777 19993 4811
rect 20027 4808 20039 4811
rect 20254 4808 20260 4820
rect 20027 4780 20260 4808
rect 20027 4777 20039 4780
rect 19981 4771 20039 4777
rect 20254 4768 20260 4780
rect 20312 4768 20318 4820
rect 20717 4811 20775 4817
rect 20717 4777 20729 4811
rect 20763 4808 20775 4811
rect 22370 4808 22376 4820
rect 20763 4780 22376 4808
rect 20763 4777 20775 4780
rect 20717 4771 20775 4777
rect 22370 4768 22376 4780
rect 22428 4768 22434 4820
rect 9033 4743 9091 4749
rect 9033 4740 9045 4743
rect 8159 4712 9045 4740
rect 8159 4684 8187 4712
rect 9033 4709 9045 4712
rect 9079 4740 9091 4743
rect 10042 4740 10048 4752
rect 9079 4712 10048 4740
rect 9079 4709 9091 4712
rect 9033 4703 9091 4709
rect 10042 4700 10048 4712
rect 10100 4700 10106 4752
rect 18782 4700 18788 4752
rect 18840 4740 18846 4752
rect 19061 4743 19119 4749
rect 19061 4740 19073 4743
rect 18840 4712 19073 4740
rect 18840 4700 18846 4712
rect 19061 4709 19073 4712
rect 19107 4740 19119 4743
rect 19107 4712 20576 4740
rect 19107 4709 19119 4712
rect 19061 4703 19119 4709
rect 8110 4672 8116 4684
rect 8023 4644 8116 4672
rect 8110 4632 8116 4644
rect 8168 4644 8187 4684
rect 8294 4672 8300 4684
rect 8255 4644 8300 4672
rect 8168 4632 8174 4644
rect 8294 4632 8300 4644
rect 8352 4632 8358 4684
rect 10410 4632 10416 4684
rect 10468 4672 10474 4684
rect 10468 4644 15424 4672
rect 10468 4632 10474 4644
rect 8389 4607 8447 4613
rect 8389 4573 8401 4607
rect 8435 4604 8447 4607
rect 8478 4604 8484 4616
rect 8435 4576 8484 4604
rect 8435 4573 8447 4576
rect 8389 4567 8447 4573
rect 8478 4564 8484 4576
rect 8536 4564 8542 4616
rect 11701 4607 11759 4613
rect 11701 4573 11713 4607
rect 11747 4573 11759 4607
rect 11701 4567 11759 4573
rect 12253 4607 12311 4613
rect 12253 4573 12265 4607
rect 12299 4604 12311 4607
rect 13814 4604 13820 4616
rect 12299 4576 13820 4604
rect 12299 4573 12311 4576
rect 12253 4567 12311 4573
rect 8202 4496 8208 4548
rect 8260 4536 8266 4548
rect 11716 4536 11744 4567
rect 13814 4564 13820 4576
rect 13872 4564 13878 4616
rect 15396 4613 15424 4644
rect 16666 4632 16672 4684
rect 16724 4672 16730 4684
rect 17034 4672 17040 4684
rect 16724 4644 16896 4672
rect 16995 4644 17040 4672
rect 16724 4632 16730 4644
rect 15381 4607 15439 4613
rect 15381 4573 15393 4607
rect 15427 4573 15439 4607
rect 16758 4604 16764 4616
rect 16719 4576 16764 4604
rect 15381 4567 15439 4573
rect 16758 4564 16764 4576
rect 16816 4564 16822 4616
rect 16868 4604 16896 4644
rect 17034 4632 17040 4644
rect 17092 4632 17098 4684
rect 17310 4632 17316 4684
rect 17368 4672 17374 4684
rect 17497 4675 17555 4681
rect 17497 4672 17509 4675
rect 17368 4644 17509 4672
rect 17368 4632 17374 4644
rect 17497 4641 17509 4644
rect 17543 4641 17555 4675
rect 17497 4635 17555 4641
rect 17773 4675 17831 4681
rect 17773 4641 17785 4675
rect 17819 4672 17831 4675
rect 18138 4672 18144 4684
rect 17819 4644 18144 4672
rect 17819 4641 17831 4644
rect 17773 4635 17831 4641
rect 18138 4632 18144 4644
rect 18196 4632 18202 4684
rect 18693 4675 18751 4681
rect 18693 4641 18705 4675
rect 18739 4672 18751 4675
rect 18966 4672 18972 4684
rect 18739 4644 18972 4672
rect 18739 4641 18751 4644
rect 18693 4635 18751 4641
rect 18966 4632 18972 4644
rect 19024 4632 19030 4684
rect 19429 4675 19487 4681
rect 19429 4641 19441 4675
rect 19475 4672 19487 4675
rect 20070 4672 20076 4684
rect 19475 4644 20076 4672
rect 19475 4641 19487 4644
rect 19429 4635 19487 4641
rect 20070 4632 20076 4644
rect 20128 4632 20134 4684
rect 20257 4675 20315 4681
rect 20257 4641 20269 4675
rect 20303 4672 20315 4675
rect 20438 4672 20444 4684
rect 20303 4644 20444 4672
rect 20303 4641 20315 4644
rect 20257 4635 20315 4641
rect 20438 4632 20444 4644
rect 20496 4632 20502 4684
rect 20548 4672 20576 4712
rect 21272 4675 21330 4681
rect 21272 4672 21284 4675
rect 20548 4644 21284 4672
rect 21272 4641 21284 4644
rect 21318 4641 21330 4675
rect 21272 4635 21330 4641
rect 21545 4675 21603 4681
rect 21545 4641 21557 4675
rect 21591 4672 21603 4675
rect 23290 4672 23296 4684
rect 21591 4644 23296 4672
rect 21591 4641 21603 4644
rect 21545 4635 21603 4641
rect 23290 4632 23296 4644
rect 23348 4632 23354 4684
rect 17402 4604 17408 4616
rect 16868 4576 17408 4604
rect 17402 4564 17408 4576
rect 17460 4564 17466 4616
rect 17957 4607 18015 4613
rect 17957 4573 17969 4607
rect 18003 4604 18015 4607
rect 18230 4604 18236 4616
rect 18003 4576 18236 4604
rect 18003 4573 18015 4576
rect 17957 4567 18015 4573
rect 18230 4564 18236 4576
rect 18288 4564 18294 4616
rect 18877 4607 18935 4613
rect 18877 4573 18889 4607
rect 18923 4604 18935 4607
rect 19058 4604 19064 4616
rect 18923 4576 19064 4604
rect 18923 4573 18935 4576
rect 18877 4567 18935 4573
rect 19058 4564 19064 4576
rect 19116 4564 19122 4616
rect 19521 4607 19579 4613
rect 19521 4573 19533 4607
rect 19567 4604 19579 4607
rect 19610 4604 19616 4616
rect 19567 4576 19616 4604
rect 19567 4573 19579 4576
rect 19521 4567 19579 4573
rect 19610 4564 19616 4576
rect 19668 4564 19674 4616
rect 20533 4607 20591 4613
rect 20533 4573 20545 4607
rect 20579 4573 20591 4607
rect 20806 4604 20812 4616
rect 20767 4576 20812 4604
rect 20533 4567 20591 4573
rect 12437 4539 12495 4545
rect 12437 4536 12449 4539
rect 8260 4508 12449 4536
rect 8260 4496 8266 4508
rect 12437 4505 12449 4508
rect 12483 4536 12495 4539
rect 13722 4536 13728 4548
rect 12483 4508 13728 4536
rect 12483 4505 12495 4508
rect 12437 4499 12495 4505
rect 13722 4496 13728 4508
rect 13780 4496 13786 4548
rect 17420 4536 17448 4564
rect 17865 4539 17923 4545
rect 17865 4536 17877 4539
rect 17420 4508 17877 4536
rect 17865 4505 17877 4508
rect 17911 4505 17923 4539
rect 20548 4536 20576 4567
rect 20806 4564 20812 4576
rect 20864 4564 20870 4616
rect 21358 4604 21364 4616
rect 20916 4576 21364 4604
rect 20916 4536 20944 4576
rect 21358 4564 21364 4576
rect 21416 4564 21422 4616
rect 21634 4564 21640 4616
rect 21692 4604 21698 4616
rect 22833 4607 22891 4613
rect 22833 4604 22845 4607
rect 21692 4576 22845 4604
rect 21692 4564 21698 4576
rect 22833 4573 22845 4576
rect 22879 4573 22891 4607
rect 22833 4567 22891 4573
rect 20548 4508 20944 4536
rect 17865 4499 17923 4505
rect 15562 4468 15568 4480
rect 15523 4440 15568 4468
rect 15562 4428 15568 4440
rect 15620 4428 15626 4480
rect 15657 4471 15715 4477
rect 15657 4437 15669 4471
rect 15703 4468 15715 4471
rect 16850 4468 16856 4480
rect 15703 4440 16856 4468
rect 15703 4437 15715 4440
rect 15657 4431 15715 4437
rect 16850 4428 16856 4440
rect 16908 4428 16914 4480
rect 17030 4471 17088 4477
rect 17030 4437 17042 4471
rect 17076 4468 17088 4471
rect 17126 4468 17132 4480
rect 17076 4440 17132 4468
rect 17076 4437 17088 4440
rect 17030 4431 17088 4437
rect 17126 4428 17132 4440
rect 17184 4428 17190 4480
rect 18782 4428 18788 4480
rect 18840 4468 18846 4480
rect 19150 4468 19156 4480
rect 18840 4440 19156 4468
rect 18840 4428 18846 4440
rect 19150 4428 19156 4440
rect 19208 4428 19214 4480
rect 19610 4468 19616 4480
rect 19571 4440 19616 4468
rect 19610 4428 19616 4440
rect 19668 4428 19674 4480
rect 20346 4468 20352 4480
rect 20307 4440 20352 4468
rect 20346 4428 20352 4440
rect 20404 4428 20410 4480
rect 20806 4428 20812 4480
rect 20864 4468 20870 4480
rect 21082 4468 21088 4480
rect 20864 4440 21088 4468
rect 20864 4428 20870 4440
rect 21082 4428 21088 4440
rect 21140 4428 21146 4480
rect 21174 4428 21180 4480
rect 21232 4468 21238 4480
rect 21275 4471 21333 4477
rect 21275 4468 21287 4471
rect 21232 4440 21287 4468
rect 21232 4428 21238 4440
rect 21275 4437 21287 4440
rect 21321 4437 21333 4471
rect 21275 4431 21333 4437
rect 21450 4428 21456 4480
rect 21508 4468 21514 4480
rect 22649 4471 22707 4477
rect 22649 4468 22661 4471
rect 21508 4440 22661 4468
rect 21508 4428 21514 4440
rect 22649 4437 22661 4440
rect 22695 4437 22707 4471
rect 23014 4468 23020 4480
rect 22975 4440 23020 4468
rect 22649 4431 22707 4437
rect 23014 4428 23020 4440
rect 23072 4428 23078 4480
rect 1104 4378 23460 4400
rect 1104 4326 6548 4378
rect 6600 4326 6612 4378
rect 6664 4326 6676 4378
rect 6728 4326 6740 4378
rect 6792 4326 6804 4378
rect 6856 4326 12146 4378
rect 12198 4326 12210 4378
rect 12262 4326 12274 4378
rect 12326 4326 12338 4378
rect 12390 4326 12402 4378
rect 12454 4326 17744 4378
rect 17796 4326 17808 4378
rect 17860 4326 17872 4378
rect 17924 4326 17936 4378
rect 17988 4326 18000 4378
rect 18052 4326 23460 4378
rect 1104 4304 23460 4326
rect 15562 4224 15568 4276
rect 15620 4264 15626 4276
rect 15749 4267 15807 4273
rect 15749 4264 15761 4267
rect 15620 4236 15761 4264
rect 15620 4224 15626 4236
rect 15749 4233 15761 4236
rect 15795 4233 15807 4267
rect 15749 4227 15807 4233
rect 16117 4267 16175 4273
rect 16117 4233 16129 4267
rect 16163 4264 16175 4267
rect 18966 4264 18972 4276
rect 16163 4236 18972 4264
rect 16163 4233 16175 4236
rect 16117 4227 16175 4233
rect 18966 4224 18972 4236
rect 19024 4224 19030 4276
rect 19061 4267 19119 4273
rect 19061 4233 19073 4267
rect 19107 4264 19119 4267
rect 19797 4267 19855 4273
rect 19797 4264 19809 4267
rect 19107 4236 19809 4264
rect 19107 4233 19119 4236
rect 19061 4227 19119 4233
rect 19797 4233 19809 4236
rect 19843 4233 19855 4267
rect 21266 4264 21272 4276
rect 21227 4236 21272 4264
rect 19797 4227 19855 4233
rect 21266 4224 21272 4236
rect 21324 4224 21330 4276
rect 22002 4264 22008 4276
rect 21963 4236 22008 4264
rect 22002 4224 22008 4236
rect 22060 4224 22066 4276
rect 22281 4267 22339 4273
rect 22281 4233 22293 4267
rect 22327 4264 22339 4267
rect 22370 4264 22376 4276
rect 22327 4236 22376 4264
rect 22327 4233 22339 4236
rect 22281 4227 22339 4233
rect 22370 4224 22376 4236
rect 22428 4224 22434 4276
rect 23750 4264 23756 4276
rect 22480 4236 23756 4264
rect 15654 4196 15660 4208
rect 15615 4168 15660 4196
rect 15654 4156 15660 4168
rect 15712 4156 15718 4208
rect 18524 4168 18736 4196
rect 11882 4088 11888 4140
rect 11940 4128 11946 4140
rect 16942 4128 16948 4140
rect 11940 4100 16948 4128
rect 11940 4088 11946 4100
rect 16942 4088 16948 4100
rect 17000 4088 17006 4140
rect 17494 4088 17500 4140
rect 17552 4128 17558 4140
rect 17678 4128 17684 4140
rect 17552 4100 17684 4128
rect 17552 4088 17558 4100
rect 17678 4088 17684 4100
rect 17736 4088 17742 4140
rect 18414 4128 18420 4140
rect 17788 4100 18420 4128
rect 15562 4060 15568 4072
rect 15523 4032 15568 4060
rect 15562 4020 15568 4032
rect 15620 4060 15626 4072
rect 16114 4060 16120 4072
rect 15620 4032 16120 4060
rect 15620 4020 15626 4032
rect 16114 4020 16120 4032
rect 16172 4020 16178 4072
rect 17788 4069 17816 4100
rect 18414 4088 18420 4100
rect 18472 4128 18478 4140
rect 18524 4128 18552 4168
rect 18472 4100 18552 4128
rect 18601 4131 18659 4137
rect 18472 4088 18478 4100
rect 18601 4097 18613 4131
rect 18647 4097 18659 4131
rect 18601 4091 18659 4097
rect 17773 4063 17831 4069
rect 17773 4029 17785 4063
rect 17819 4029 17831 4063
rect 17773 4023 17831 4029
rect 17954 4020 17960 4072
rect 18012 4060 18018 4072
rect 18046 4063 18104 4069
rect 18046 4060 18058 4063
rect 18012 4032 18058 4060
rect 18012 4020 18018 4032
rect 18046 4029 18058 4032
rect 18092 4029 18104 4063
rect 18046 4023 18104 4029
rect 18138 4020 18144 4072
rect 18196 4069 18202 4072
rect 18196 4063 18244 4069
rect 18196 4029 18198 4063
rect 18232 4029 18244 4063
rect 18506 4060 18512 4072
rect 18467 4032 18512 4060
rect 18196 4023 18244 4029
rect 18196 4020 18202 4023
rect 18506 4020 18512 4032
rect 18564 4020 18570 4072
rect 14182 3952 14188 4004
rect 14240 3992 14246 4004
rect 14240 3964 17172 3992
rect 14240 3952 14246 3964
rect 16666 3924 16672 3936
rect 16627 3896 16672 3924
rect 16666 3884 16672 3896
rect 16724 3884 16730 3936
rect 17144 3924 17172 3964
rect 18616 3924 18644 4091
rect 18708 4060 18736 4168
rect 19426 4156 19432 4208
rect 19484 4196 19490 4208
rect 20625 4199 20683 4205
rect 20625 4196 20637 4199
rect 19484 4168 20637 4196
rect 19484 4156 19490 4168
rect 20625 4165 20637 4168
rect 20671 4165 20683 4199
rect 22480 4196 22508 4236
rect 23750 4224 23756 4236
rect 23808 4224 23814 4276
rect 20625 4159 20683 4165
rect 22388 4168 22508 4196
rect 18874 4128 18880 4140
rect 18835 4100 18880 4128
rect 18874 4088 18880 4100
rect 18932 4088 18938 4140
rect 19150 4128 19156 4140
rect 19111 4100 19156 4128
rect 19150 4088 19156 4100
rect 19208 4088 19214 4140
rect 21361 4131 21419 4137
rect 19628 4100 20944 4128
rect 19518 4060 19524 4072
rect 18708 4032 19524 4060
rect 19518 4020 19524 4032
rect 19576 4020 19582 4072
rect 19628 4069 19656 4100
rect 20916 4069 20944 4100
rect 21361 4097 21373 4131
rect 21407 4128 21419 4131
rect 21818 4128 21824 4140
rect 21407 4100 21824 4128
rect 21407 4097 21419 4100
rect 21361 4091 21419 4097
rect 21818 4088 21824 4100
rect 21876 4088 21882 4140
rect 21910 4088 21916 4140
rect 21968 4128 21974 4140
rect 22388 4132 22416 4168
rect 22554 4156 22560 4208
rect 22612 4196 22618 4208
rect 22612 4168 22876 4196
rect 22612 4156 22618 4168
rect 22848 4137 22876 4168
rect 22465 4132 22523 4137
rect 22388 4131 22523 4132
rect 21968 4100 22013 4128
rect 22066 4100 22324 4128
rect 22388 4104 22477 4131
rect 21968 4088 21974 4100
rect 19613 4063 19671 4069
rect 19613 4029 19625 4063
rect 19659 4029 19671 4063
rect 19613 4023 19671 4029
rect 19705 4063 19763 4069
rect 19705 4029 19717 4063
rect 19751 4029 19763 4063
rect 20717 4063 20775 4069
rect 20717 4060 20729 4063
rect 19705 4023 19763 4029
rect 19904 4032 20729 4060
rect 18785 3995 18843 4001
rect 18785 3961 18797 3995
rect 18831 3992 18843 3995
rect 19720 3992 19748 4023
rect 18831 3964 19748 3992
rect 18831 3961 18843 3964
rect 18785 3955 18843 3961
rect 19334 3924 19340 3936
rect 17144 3896 18644 3924
rect 19295 3896 19340 3924
rect 19334 3884 19340 3896
rect 19392 3884 19398 3936
rect 19518 3884 19524 3936
rect 19576 3924 19582 3936
rect 19904 3924 19932 4032
rect 20717 4029 20729 4032
rect 20763 4029 20775 4063
rect 20717 4023 20775 4029
rect 20901 4063 20959 4069
rect 20901 4029 20913 4063
rect 20947 4060 20959 4063
rect 22066 4060 22094 4100
rect 20947 4032 22094 4060
rect 22296 4060 22324 4100
rect 22465 4097 22477 4104
rect 22511 4097 22523 4131
rect 22465 4091 22523 4097
rect 22741 4131 22799 4137
rect 22741 4097 22753 4131
rect 22787 4097 22799 4131
rect 22741 4091 22799 4097
rect 22833 4131 22891 4137
rect 22833 4097 22845 4131
rect 22879 4097 22891 4131
rect 22833 4091 22891 4097
rect 22296 4032 22600 4060
rect 20947 4029 20959 4032
rect 20901 4023 20959 4029
rect 21545 3995 21603 4001
rect 21545 3961 21557 3995
rect 21591 3992 21603 3995
rect 22278 3992 22284 4004
rect 21591 3964 22284 3992
rect 21591 3961 21603 3964
rect 21545 3955 21603 3961
rect 22278 3952 22284 3964
rect 22336 3952 22342 4004
rect 22572 4001 22600 4032
rect 22557 3995 22615 4001
rect 22557 3961 22569 3995
rect 22603 3961 22615 3995
rect 22557 3955 22615 3961
rect 20162 3924 20168 3936
rect 19576 3896 19932 3924
rect 20123 3896 20168 3924
rect 19576 3884 19582 3896
rect 20162 3884 20168 3896
rect 20220 3884 20226 3936
rect 20257 3927 20315 3933
rect 20257 3893 20269 3927
rect 20303 3924 20315 3927
rect 20438 3924 20444 3936
rect 20303 3896 20444 3924
rect 20303 3893 20315 3896
rect 20257 3887 20315 3893
rect 20438 3884 20444 3896
rect 20496 3884 20502 3936
rect 20530 3884 20536 3936
rect 20588 3924 20594 3936
rect 22756 3924 22784 4091
rect 23014 3924 23020 3936
rect 20588 3896 22784 3924
rect 22975 3896 23020 3924
rect 20588 3884 20594 3896
rect 23014 3884 23020 3896
rect 23072 3884 23078 3936
rect 1104 3834 23460 3856
rect 1104 3782 3749 3834
rect 3801 3782 3813 3834
rect 3865 3782 3877 3834
rect 3929 3782 3941 3834
rect 3993 3782 4005 3834
rect 4057 3782 9347 3834
rect 9399 3782 9411 3834
rect 9463 3782 9475 3834
rect 9527 3782 9539 3834
rect 9591 3782 9603 3834
rect 9655 3782 14945 3834
rect 14997 3782 15009 3834
rect 15061 3782 15073 3834
rect 15125 3782 15137 3834
rect 15189 3782 15201 3834
rect 15253 3782 20543 3834
rect 20595 3782 20607 3834
rect 20659 3782 20671 3834
rect 20723 3782 20735 3834
rect 20787 3782 20799 3834
rect 20851 3782 23460 3834
rect 1104 3760 23460 3782
rect 17310 3680 17316 3732
rect 17368 3720 17374 3732
rect 18049 3723 18107 3729
rect 18049 3720 18061 3723
rect 17368 3692 18061 3720
rect 17368 3680 17374 3692
rect 18049 3689 18061 3692
rect 18095 3689 18107 3723
rect 19426 3720 19432 3732
rect 19387 3692 19432 3720
rect 18049 3683 18107 3689
rect 19426 3680 19432 3692
rect 19484 3680 19490 3732
rect 19613 3723 19671 3729
rect 19613 3689 19625 3723
rect 19659 3720 19671 3723
rect 20346 3720 20352 3732
rect 19659 3692 20352 3720
rect 19659 3689 19671 3692
rect 19613 3683 19671 3689
rect 20346 3680 20352 3692
rect 20404 3680 20410 3732
rect 22462 3720 22468 3732
rect 22066 3692 22468 3720
rect 17957 3655 18015 3661
rect 17957 3621 17969 3655
rect 18003 3652 18015 3655
rect 18138 3652 18144 3664
rect 18003 3624 18144 3652
rect 18003 3621 18015 3624
rect 17957 3615 18015 3621
rect 18138 3612 18144 3624
rect 18196 3652 18202 3664
rect 18966 3652 18972 3664
rect 18196 3624 18972 3652
rect 18196 3612 18202 3624
rect 18966 3612 18972 3624
rect 19024 3612 19030 3664
rect 19061 3655 19119 3661
rect 19061 3621 19073 3655
rect 19107 3621 19119 3655
rect 19061 3615 19119 3621
rect 16850 3584 16856 3596
rect 16811 3556 16856 3584
rect 16850 3544 16856 3556
rect 16908 3544 16914 3596
rect 17034 3544 17040 3596
rect 17092 3584 17098 3596
rect 17126 3587 17184 3593
rect 17126 3584 17138 3587
rect 17092 3556 17138 3584
rect 17092 3544 17098 3556
rect 17126 3553 17138 3556
rect 17172 3553 17184 3587
rect 17126 3547 17184 3553
rect 17218 3544 17224 3596
rect 17276 3584 17282 3596
rect 17276 3556 17816 3584
rect 17276 3544 17282 3556
rect 1581 3519 1639 3525
rect 1581 3485 1593 3519
rect 1627 3516 1639 3519
rect 16206 3516 16212 3528
rect 1627 3488 16212 3516
rect 1627 3485 1639 3488
rect 1581 3479 1639 3485
rect 16206 3476 16212 3488
rect 16264 3476 16270 3528
rect 16574 3476 16580 3528
rect 16632 3516 16638 3528
rect 17310 3516 17316 3528
rect 16632 3488 17316 3516
rect 16632 3476 16638 3488
rect 17310 3476 17316 3488
rect 17368 3516 17374 3528
rect 17788 3525 17816 3556
rect 18322 3544 18328 3596
rect 18380 3584 18386 3596
rect 19076 3584 19104 3615
rect 19150 3612 19156 3664
rect 19208 3652 19214 3664
rect 19981 3655 20039 3661
rect 19981 3652 19993 3655
rect 19208 3624 19993 3652
rect 19208 3612 19214 3624
rect 19981 3621 19993 3624
rect 20027 3621 20039 3655
rect 19981 3615 20039 3621
rect 20254 3612 20260 3664
rect 20312 3652 20318 3664
rect 20993 3655 21051 3661
rect 20312 3624 20576 3652
rect 20312 3612 20318 3624
rect 19518 3584 19524 3596
rect 18380 3556 18920 3584
rect 19076 3556 19524 3584
rect 18380 3544 18386 3556
rect 17589 3519 17647 3525
rect 17589 3516 17601 3519
rect 17368 3488 17601 3516
rect 17368 3476 17374 3488
rect 17589 3485 17601 3488
rect 17635 3485 17647 3519
rect 17589 3479 17647 3485
rect 17773 3519 17831 3525
rect 17773 3485 17785 3519
rect 17819 3485 17831 3519
rect 17773 3479 17831 3485
rect 18233 3519 18291 3525
rect 18233 3485 18245 3519
rect 18279 3516 18291 3519
rect 18690 3516 18696 3528
rect 18279 3488 18696 3516
rect 18279 3485 18291 3488
rect 18233 3479 18291 3485
rect 18690 3476 18696 3488
rect 18748 3476 18754 3528
rect 18892 3525 18920 3556
rect 19518 3544 19524 3556
rect 19576 3544 19582 3596
rect 20438 3584 20444 3596
rect 19720 3556 20444 3584
rect 18785 3519 18843 3525
rect 18785 3485 18797 3519
rect 18831 3485 18843 3519
rect 18785 3479 18843 3485
rect 18877 3519 18935 3525
rect 18877 3485 18889 3519
rect 18923 3485 18935 3519
rect 18877 3479 18935 3485
rect 18800 3448 18828 3479
rect 19150 3476 19156 3528
rect 19208 3516 19214 3528
rect 19720 3525 19748 3556
rect 20438 3544 20444 3556
rect 20496 3544 20502 3596
rect 20548 3593 20576 3624
rect 20993 3621 21005 3655
rect 21039 3652 21051 3655
rect 22066 3652 22094 3692
rect 22462 3680 22468 3692
rect 22520 3680 22526 3732
rect 23566 3720 23572 3732
rect 22664 3692 23572 3720
rect 22554 3652 22560 3664
rect 21039 3624 22094 3652
rect 22515 3624 22560 3652
rect 21039 3621 21051 3624
rect 20993 3615 21051 3621
rect 22554 3612 22560 3624
rect 22612 3612 22618 3664
rect 20533 3587 20591 3593
rect 20533 3553 20545 3587
rect 20579 3553 20591 3587
rect 20533 3547 20591 3553
rect 21358 3544 21364 3596
rect 21416 3584 21422 3596
rect 21821 3587 21879 3593
rect 21821 3584 21833 3587
rect 21416 3556 21833 3584
rect 21416 3544 21422 3556
rect 21821 3553 21833 3556
rect 21867 3553 21879 3587
rect 22186 3584 22192 3596
rect 22147 3556 22192 3584
rect 21821 3547 21879 3553
rect 22186 3544 22192 3556
rect 22244 3544 22250 3596
rect 19245 3519 19303 3525
rect 19245 3516 19257 3519
rect 19208 3488 19257 3516
rect 19208 3476 19214 3488
rect 19245 3485 19257 3488
rect 19291 3485 19303 3519
rect 19245 3479 19303 3485
rect 19705 3519 19763 3525
rect 19705 3485 19717 3519
rect 19751 3485 19763 3519
rect 19705 3479 19763 3485
rect 20809 3519 20867 3525
rect 20809 3485 20821 3519
rect 20855 3516 20867 3519
rect 20898 3516 20904 3528
rect 20855 3488 20904 3516
rect 20855 3485 20867 3488
rect 20809 3479 20867 3485
rect 20898 3476 20904 3488
rect 20956 3476 20962 3528
rect 21450 3476 21456 3528
rect 21508 3516 21514 3528
rect 21545 3519 21603 3525
rect 21545 3516 21557 3519
rect 21508 3488 21557 3516
rect 21508 3476 21514 3488
rect 21545 3485 21557 3488
rect 21591 3516 21603 3519
rect 22281 3519 22339 3525
rect 22281 3516 22293 3519
rect 21591 3488 22293 3516
rect 21591 3485 21603 3488
rect 21545 3479 21603 3485
rect 22281 3485 22293 3488
rect 22327 3516 22339 3519
rect 22664 3516 22692 3692
rect 23566 3680 23572 3692
rect 23624 3680 23630 3732
rect 23658 3652 23664 3664
rect 22756 3624 23664 3652
rect 22756 3525 22784 3624
rect 23658 3612 23664 3624
rect 23716 3612 23722 3664
rect 22848 3525 22968 3532
rect 22327 3488 22692 3516
rect 22741 3519 22799 3525
rect 22327 3485 22339 3488
rect 22281 3479 22339 3485
rect 22741 3485 22753 3519
rect 22787 3485 22799 3519
rect 22741 3479 22799 3485
rect 22833 3519 22968 3525
rect 22833 3485 22845 3519
rect 22879 3516 22968 3519
rect 23106 3516 23112 3528
rect 22879 3504 23112 3516
rect 22879 3485 22891 3504
rect 22940 3488 23112 3504
rect 22833 3479 22891 3485
rect 23106 3476 23112 3488
rect 23164 3476 23170 3528
rect 20162 3448 20168 3460
rect 18800 3420 20168 3448
rect 20162 3408 20168 3420
rect 20220 3448 20226 3460
rect 20349 3451 20407 3457
rect 20349 3448 20361 3451
rect 20220 3420 20361 3448
rect 20220 3408 20226 3420
rect 20349 3417 20361 3420
rect 20395 3417 20407 3451
rect 22922 3448 22928 3460
rect 20349 3411 20407 3417
rect 22480 3420 22928 3448
rect 1394 3380 1400 3392
rect 1355 3352 1400 3380
rect 1394 3340 1400 3352
rect 1452 3340 1458 3392
rect 15746 3380 15752 3392
rect 15707 3352 15752 3380
rect 15746 3340 15752 3352
rect 15804 3340 15810 3392
rect 17126 3389 17132 3392
rect 17122 3380 17132 3389
rect 17087 3352 17132 3380
rect 17122 3343 17132 3352
rect 17126 3340 17132 3343
rect 17184 3340 17190 3392
rect 17218 3340 17224 3392
rect 17276 3380 17282 3392
rect 18601 3383 18659 3389
rect 18601 3380 18613 3383
rect 17276 3352 18613 3380
rect 17276 3340 17282 3352
rect 18601 3349 18613 3352
rect 18647 3380 18659 3383
rect 19610 3380 19616 3392
rect 18647 3352 19616 3380
rect 18647 3349 18659 3352
rect 18601 3343 18659 3349
rect 19610 3340 19616 3352
rect 19668 3340 19674 3392
rect 19886 3380 19892 3392
rect 19847 3352 19892 3380
rect 19886 3340 19892 3352
rect 19944 3340 19950 3392
rect 19978 3340 19984 3392
rect 20036 3380 20042 3392
rect 21634 3380 21640 3392
rect 20036 3352 21640 3380
rect 20036 3340 20042 3352
rect 21634 3340 21640 3352
rect 21692 3340 21698 3392
rect 22480 3389 22508 3420
rect 22922 3408 22928 3420
rect 22980 3408 22986 3460
rect 22465 3383 22523 3389
rect 22465 3349 22477 3383
rect 22511 3349 22523 3383
rect 23014 3380 23020 3392
rect 22975 3352 23020 3380
rect 22465 3343 22523 3349
rect 23014 3340 23020 3352
rect 23072 3340 23078 3392
rect 1104 3290 23460 3312
rect 1104 3238 6548 3290
rect 6600 3238 6612 3290
rect 6664 3238 6676 3290
rect 6728 3238 6740 3290
rect 6792 3238 6804 3290
rect 6856 3238 12146 3290
rect 12198 3238 12210 3290
rect 12262 3238 12274 3290
rect 12326 3238 12338 3290
rect 12390 3238 12402 3290
rect 12454 3238 17744 3290
rect 17796 3238 17808 3290
rect 17860 3238 17872 3290
rect 17924 3238 17936 3290
rect 17988 3238 18000 3290
rect 18052 3238 23460 3290
rect 1104 3216 23460 3238
rect 11330 3136 11336 3188
rect 11388 3176 11394 3188
rect 18966 3176 18972 3188
rect 11388 3148 18972 3176
rect 11388 3136 11394 3148
rect 18966 3136 18972 3148
rect 19024 3136 19030 3188
rect 19058 3136 19064 3188
rect 19116 3176 19122 3188
rect 19974 3179 20032 3185
rect 19974 3176 19986 3179
rect 19116 3148 19986 3176
rect 19116 3136 19122 3148
rect 19974 3145 19986 3148
rect 20020 3176 20032 3179
rect 21174 3176 21180 3188
rect 20020 3148 21180 3176
rect 20020 3145 20032 3148
rect 19974 3139 20032 3145
rect 21174 3136 21180 3148
rect 21232 3136 21238 3188
rect 22005 3179 22063 3185
rect 22005 3145 22017 3179
rect 22051 3176 22063 3179
rect 22738 3176 22744 3188
rect 22051 3148 22744 3176
rect 22051 3145 22063 3148
rect 22005 3139 22063 3145
rect 16206 3108 16212 3120
rect 16167 3080 16212 3108
rect 16206 3068 16212 3080
rect 16264 3068 16270 3120
rect 8573 3043 8631 3049
rect 8573 3009 8585 3043
rect 8619 3040 8631 3043
rect 16485 3043 16543 3049
rect 8619 3012 8800 3040
rect 8619 3009 8631 3012
rect 8573 3003 8631 3009
rect 8386 2836 8392 2848
rect 8347 2808 8392 2836
rect 8386 2796 8392 2808
rect 8444 2796 8450 2848
rect 8772 2845 8800 3012
rect 16485 3009 16497 3043
rect 16531 3040 16543 3043
rect 16758 3040 16764 3052
rect 16531 3012 16764 3040
rect 16531 3009 16543 3012
rect 16485 3003 16543 3009
rect 16758 3000 16764 3012
rect 16816 3040 16822 3052
rect 19242 3040 19248 3052
rect 16816 3012 19248 3040
rect 16816 3000 16822 3012
rect 19242 3000 19248 3012
rect 19300 3000 19306 3052
rect 19702 3040 19708 3052
rect 19663 3012 19708 3040
rect 19702 3000 19708 3012
rect 19760 3000 19766 3052
rect 21542 3040 21548 3052
rect 20364 3012 21548 3040
rect 19978 2993 20036 2999
rect 16574 2932 16580 2984
rect 16632 2972 16638 2984
rect 17034 2981 17040 2984
rect 16669 2975 16727 2981
rect 16669 2972 16681 2975
rect 16632 2944 16681 2972
rect 16632 2932 16638 2944
rect 16669 2941 16681 2944
rect 16715 2941 16727 2975
rect 16669 2935 16727 2941
rect 16992 2975 17040 2981
rect 16992 2941 17004 2975
rect 17038 2941 17040 2975
rect 16992 2935 17040 2941
rect 17034 2932 17040 2935
rect 17092 2932 17098 2984
rect 17132 2975 17190 2981
rect 17132 2941 17144 2975
rect 17178 2972 17190 2975
rect 17218 2972 17224 2984
rect 17178 2944 17224 2972
rect 17178 2941 17190 2944
rect 17132 2935 17190 2941
rect 17218 2932 17224 2944
rect 17276 2932 17282 2984
rect 17402 2972 17408 2984
rect 17363 2944 17408 2972
rect 17402 2932 17408 2944
rect 17460 2932 17466 2984
rect 18782 2972 18788 2984
rect 18616 2944 18788 2972
rect 8757 2839 8815 2845
rect 8757 2805 8769 2839
rect 8803 2836 8815 2839
rect 10778 2836 10784 2848
rect 8803 2808 10784 2836
rect 8803 2805 8815 2808
rect 8757 2799 8815 2805
rect 10778 2796 10784 2808
rect 10836 2796 10842 2848
rect 11974 2796 11980 2848
rect 12032 2836 12038 2848
rect 18322 2836 18328 2848
rect 12032 2808 18328 2836
rect 12032 2796 12038 2808
rect 18322 2796 18328 2808
rect 18380 2796 18386 2848
rect 18414 2796 18420 2848
rect 18472 2836 18478 2848
rect 18616 2845 18644 2944
rect 18782 2932 18788 2944
rect 18840 2932 18846 2984
rect 19978 2959 19990 2993
rect 20024 2972 20036 2993
rect 20364 2972 20392 3012
rect 21542 3000 21548 3012
rect 21600 3000 21606 3052
rect 22112 3049 22140 3148
rect 22738 3136 22744 3148
rect 22796 3136 22802 3188
rect 22646 3068 22652 3120
rect 22704 3108 22710 3120
rect 22704 3080 22876 3108
rect 22704 3068 22710 3080
rect 22848 3049 22876 3080
rect 22097 3043 22155 3049
rect 22097 3009 22109 3043
rect 22143 3009 22155 3043
rect 22097 3003 22155 3009
rect 22833 3043 22891 3049
rect 22833 3009 22845 3043
rect 22879 3009 22891 3043
rect 22833 3003 22891 3009
rect 20024 2959 20392 2972
rect 19978 2953 20392 2959
rect 19996 2944 20392 2953
rect 20441 2975 20499 2981
rect 20441 2941 20453 2975
rect 20487 2972 20499 2975
rect 21082 2972 21088 2984
rect 20487 2944 21088 2972
rect 20487 2941 20499 2944
rect 20441 2935 20499 2941
rect 18509 2839 18567 2845
rect 18509 2836 18521 2839
rect 18472 2808 18521 2836
rect 18472 2796 18478 2808
rect 18509 2805 18521 2808
rect 18555 2805 18567 2839
rect 18509 2799 18567 2805
rect 18601 2839 18659 2845
rect 18601 2805 18613 2839
rect 18647 2805 18659 2839
rect 18601 2799 18659 2805
rect 18690 2796 18696 2848
rect 18748 2836 18754 2848
rect 20456 2836 20484 2935
rect 21082 2932 21088 2944
rect 21140 2932 21146 2984
rect 22373 2975 22431 2981
rect 22373 2941 22385 2975
rect 22419 2972 22431 2975
rect 22646 2972 22652 2984
rect 22419 2944 22652 2972
rect 22419 2941 22431 2944
rect 22373 2935 22431 2941
rect 22646 2932 22652 2944
rect 22704 2932 22710 2984
rect 22741 2975 22799 2981
rect 22741 2941 22753 2975
rect 22787 2972 22799 2975
rect 23382 2972 23388 2984
rect 22787 2944 23388 2972
rect 22787 2941 22799 2944
rect 22741 2935 22799 2941
rect 23382 2932 23388 2944
rect 23440 2932 23446 2984
rect 23014 2836 23020 2848
rect 18748 2808 20484 2836
rect 22975 2808 23020 2836
rect 18748 2796 18754 2808
rect 23014 2796 23020 2808
rect 23072 2796 23078 2848
rect 23106 2796 23112 2848
rect 23164 2836 23170 2848
rect 23842 2836 23848 2848
rect 23164 2808 23848 2836
rect 23164 2796 23170 2808
rect 23842 2796 23848 2808
rect 23900 2796 23906 2848
rect 1104 2746 23460 2768
rect 1104 2694 3749 2746
rect 3801 2694 3813 2746
rect 3865 2694 3877 2746
rect 3929 2694 3941 2746
rect 3993 2694 4005 2746
rect 4057 2694 9347 2746
rect 9399 2694 9411 2746
rect 9463 2694 9475 2746
rect 9527 2694 9539 2746
rect 9591 2694 9603 2746
rect 9655 2694 14945 2746
rect 14997 2694 15009 2746
rect 15061 2694 15073 2746
rect 15125 2694 15137 2746
rect 15189 2694 15201 2746
rect 15253 2694 20543 2746
rect 20595 2694 20607 2746
rect 20659 2694 20671 2746
rect 20723 2694 20735 2746
rect 20787 2694 20799 2746
rect 20851 2694 23460 2746
rect 1104 2672 23460 2694
rect 10778 2632 10784 2644
rect 10691 2604 10784 2632
rect 10778 2592 10784 2604
rect 10836 2632 10842 2644
rect 15746 2632 15752 2644
rect 10836 2604 15752 2632
rect 10836 2592 10842 2604
rect 15746 2592 15752 2604
rect 15804 2592 15810 2644
rect 16758 2632 16764 2644
rect 16719 2604 16764 2632
rect 16758 2592 16764 2604
rect 16816 2592 16822 2644
rect 22833 2635 22891 2641
rect 22833 2601 22845 2635
rect 22879 2632 22891 2635
rect 23106 2632 23112 2644
rect 22879 2604 23112 2632
rect 22879 2601 22891 2604
rect 22833 2595 22891 2601
rect 23106 2592 23112 2604
rect 23164 2592 23170 2644
rect 8386 2496 8392 2508
rect 2516 2468 8392 2496
rect 2516 2437 2544 2468
rect 8386 2456 8392 2468
rect 8444 2456 8450 2508
rect 2501 2431 2559 2437
rect 2501 2397 2513 2431
rect 2547 2397 2559 2431
rect 2501 2391 2559 2397
rect 6178 2388 6184 2440
rect 6236 2428 6242 2440
rect 6365 2431 6423 2437
rect 6365 2428 6377 2431
rect 6236 2400 6377 2428
rect 6236 2388 6242 2400
rect 6365 2397 6377 2400
rect 6411 2397 6423 2431
rect 6365 2391 6423 2397
rect 10597 2431 10655 2437
rect 10597 2397 10609 2431
rect 10643 2428 10655 2431
rect 10796 2428 10824 2592
rect 22646 2428 22652 2440
rect 10643 2400 10824 2428
rect 22607 2400 22652 2428
rect 10643 2397 10655 2400
rect 10597 2391 10655 2397
rect 22646 2388 22652 2400
rect 22704 2388 22710 2440
rect 2130 2252 2136 2304
rect 2188 2292 2194 2304
rect 2317 2295 2375 2301
rect 2317 2292 2329 2295
rect 2188 2264 2329 2292
rect 2188 2252 2194 2264
rect 2317 2261 2329 2264
rect 2363 2261 2375 2295
rect 2317 2255 2375 2261
rect 10226 2252 10232 2304
rect 10284 2292 10290 2304
rect 10413 2295 10471 2301
rect 10413 2292 10425 2295
rect 10284 2264 10425 2292
rect 10284 2252 10290 2264
rect 10413 2261 10425 2264
rect 10459 2261 10471 2295
rect 10413 2255 10471 2261
rect 22370 2252 22376 2304
rect 22428 2292 22434 2304
rect 22465 2295 22523 2301
rect 22465 2292 22477 2295
rect 22428 2264 22477 2292
rect 22428 2252 22434 2264
rect 22465 2261 22477 2264
rect 22511 2261 22523 2295
rect 22465 2255 22523 2261
rect 1104 2202 23460 2224
rect 1104 2150 6548 2202
rect 6600 2150 6612 2202
rect 6664 2150 6676 2202
rect 6728 2150 6740 2202
rect 6792 2150 6804 2202
rect 6856 2150 12146 2202
rect 12198 2150 12210 2202
rect 12262 2150 12274 2202
rect 12326 2150 12338 2202
rect 12390 2150 12402 2202
rect 12454 2150 17744 2202
rect 17796 2150 17808 2202
rect 17860 2150 17872 2202
rect 17924 2150 17936 2202
rect 17988 2150 18000 2202
rect 18052 2150 23460 2202
rect 1104 2128 23460 2150
<< via1 >>
rect 11980 22788 12032 22840
rect 19064 22788 19116 22840
rect 9036 22720 9088 22772
rect 20168 22720 20220 22772
rect 7472 22652 7524 22704
rect 19708 22652 19760 22704
rect 5172 22584 5224 22636
rect 19340 22584 19392 22636
rect 14556 22516 14608 22568
rect 16304 22516 16356 22568
rect 14096 22448 14148 22500
rect 20996 22448 21048 22500
rect 13820 22380 13872 22432
rect 15568 22380 15620 22432
rect 3749 22278 3801 22330
rect 3813 22278 3865 22330
rect 3877 22278 3929 22330
rect 3941 22278 3993 22330
rect 4005 22278 4057 22330
rect 9347 22278 9399 22330
rect 9411 22278 9463 22330
rect 9475 22278 9527 22330
rect 9539 22278 9591 22330
rect 9603 22278 9655 22330
rect 14945 22278 14997 22330
rect 15009 22278 15061 22330
rect 15073 22278 15125 22330
rect 15137 22278 15189 22330
rect 15201 22278 15253 22330
rect 20543 22278 20595 22330
rect 20607 22278 20659 22330
rect 20671 22278 20723 22330
rect 20735 22278 20787 22330
rect 20799 22278 20851 22330
rect 5724 22176 5776 22228
rect 5448 22083 5500 22092
rect 5448 22049 5457 22083
rect 5457 22049 5491 22083
rect 5491 22049 5500 22083
rect 5448 22040 5500 22049
rect 2412 21972 2464 22024
rect 2964 21972 3016 22024
rect 3240 22015 3292 22024
rect 3240 21981 3249 22015
rect 3249 21981 3283 22015
rect 3283 21981 3292 22015
rect 3240 21972 3292 21981
rect 4160 21972 4212 22024
rect 3700 21904 3752 21956
rect 4988 21972 5040 22024
rect 6092 22040 6144 22092
rect 6460 22040 6512 22092
rect 7380 22040 7432 22092
rect 7656 22108 7708 22160
rect 6828 21972 6880 22024
rect 8024 21972 8076 22024
rect 9128 22108 9180 22160
rect 8484 22015 8536 22024
rect 8484 21981 8493 22015
rect 8493 21981 8527 22015
rect 8527 21981 8536 22015
rect 8484 21972 8536 21981
rect 9220 21972 9272 22024
rect 9956 21972 10008 22024
rect 10232 22015 10284 22024
rect 10232 21981 10241 22015
rect 10241 21981 10275 22015
rect 10275 21981 10284 22015
rect 10232 21972 10284 21981
rect 11060 22015 11112 22024
rect 1584 21836 1636 21888
rect 2228 21836 2280 21888
rect 2872 21836 2924 21888
rect 3516 21836 3568 21888
rect 4252 21836 4304 21888
rect 4620 21879 4672 21888
rect 4620 21845 4629 21879
rect 4629 21845 4663 21879
rect 4663 21845 4672 21879
rect 4620 21836 4672 21845
rect 4804 21836 4856 21888
rect 5816 21836 5868 21888
rect 6368 21879 6420 21888
rect 6368 21845 6377 21879
rect 6377 21845 6411 21879
rect 6411 21845 6420 21879
rect 6368 21836 6420 21845
rect 6460 21836 6512 21888
rect 6920 21836 6972 21888
rect 7564 21879 7616 21888
rect 7564 21845 7573 21879
rect 7573 21845 7607 21879
rect 7607 21845 7616 21879
rect 7564 21836 7616 21845
rect 7840 21879 7892 21888
rect 7840 21845 7849 21879
rect 7849 21845 7883 21879
rect 7883 21845 7892 21879
rect 7840 21836 7892 21845
rect 10600 21904 10652 21956
rect 11060 21981 11069 22015
rect 11069 21981 11103 22015
rect 11103 21981 11112 22015
rect 11060 21972 11112 21981
rect 11888 22040 11940 22092
rect 12440 22083 12492 22092
rect 11520 22015 11572 22024
rect 11520 21981 11529 22015
rect 11529 21981 11563 22015
rect 11563 21981 11572 22015
rect 11520 21972 11572 21981
rect 12440 22049 12449 22083
rect 12449 22049 12483 22083
rect 12483 22049 12492 22083
rect 12716 22083 12768 22092
rect 12440 22040 12492 22049
rect 12716 22049 12725 22083
rect 12725 22049 12759 22083
rect 12759 22049 12768 22083
rect 14464 22176 14516 22228
rect 16028 22176 16080 22228
rect 16304 22176 16356 22228
rect 22560 22176 22612 22228
rect 13636 22151 13688 22160
rect 13636 22117 13645 22151
rect 13645 22117 13679 22151
rect 13679 22117 13688 22151
rect 13636 22108 13688 22117
rect 14832 22108 14884 22160
rect 16120 22108 16172 22160
rect 16488 22108 16540 22160
rect 12716 22040 12768 22049
rect 12532 21972 12584 22024
rect 13176 21972 13228 22024
rect 13636 21972 13688 22024
rect 9220 21836 9272 21888
rect 9496 21879 9548 21888
rect 9496 21845 9505 21879
rect 9505 21845 9539 21879
rect 9539 21845 9548 21879
rect 9496 21836 9548 21845
rect 9772 21836 9824 21888
rect 10048 21879 10100 21888
rect 10048 21845 10057 21879
rect 10057 21845 10091 21879
rect 10091 21845 10100 21879
rect 10048 21836 10100 21845
rect 10876 21879 10928 21888
rect 10876 21845 10885 21879
rect 10885 21845 10919 21879
rect 10919 21845 10928 21879
rect 10876 21836 10928 21845
rect 11152 21879 11204 21888
rect 11152 21845 11161 21879
rect 11161 21845 11195 21879
rect 11195 21845 11204 21879
rect 11152 21836 11204 21845
rect 11704 21879 11756 21888
rect 11704 21845 11713 21879
rect 11713 21845 11747 21879
rect 11747 21845 11756 21879
rect 11704 21836 11756 21845
rect 11888 21879 11940 21888
rect 11888 21845 11897 21879
rect 11897 21845 11931 21879
rect 11931 21845 11940 21879
rect 11888 21836 11940 21845
rect 12072 21836 12124 21888
rect 12900 21879 12952 21888
rect 12900 21845 12909 21879
rect 12909 21845 12943 21879
rect 12943 21845 12952 21879
rect 12900 21836 12952 21845
rect 12992 21879 13044 21888
rect 12992 21845 13001 21879
rect 13001 21845 13035 21879
rect 13035 21845 13044 21879
rect 14372 21904 14424 21956
rect 15016 21904 15068 21956
rect 15476 22015 15528 22024
rect 15476 21981 15485 22015
rect 15485 21981 15519 22015
rect 15519 21981 15528 22015
rect 15752 22015 15804 22024
rect 15476 21972 15528 21981
rect 15752 21981 15761 22015
rect 15761 21981 15795 22015
rect 15795 21981 15804 22015
rect 15752 21972 15804 21981
rect 16028 22015 16080 22024
rect 16028 21981 16037 22015
rect 16037 21981 16071 22015
rect 16071 21981 16080 22015
rect 16028 21972 16080 21981
rect 16120 21972 16172 22024
rect 12992 21836 13044 21845
rect 13820 21836 13872 21888
rect 14740 21879 14792 21888
rect 14740 21845 14749 21879
rect 14749 21845 14783 21879
rect 14783 21845 14792 21879
rect 14740 21836 14792 21845
rect 15200 21836 15252 21888
rect 15384 21836 15436 21888
rect 15936 21904 15988 21956
rect 17316 22108 17368 22160
rect 16948 22083 17000 22092
rect 16948 22049 16957 22083
rect 16957 22049 16991 22083
rect 16991 22049 17000 22083
rect 16948 22040 17000 22049
rect 19156 22108 19208 22160
rect 17960 21972 18012 22024
rect 16120 21879 16172 21888
rect 16120 21845 16129 21879
rect 16129 21845 16163 21879
rect 16163 21845 16172 21879
rect 16120 21836 16172 21845
rect 16304 21836 16356 21888
rect 17592 21904 17644 21956
rect 18144 21904 18196 21956
rect 17132 21879 17184 21888
rect 17132 21845 17141 21879
rect 17141 21845 17175 21879
rect 17175 21845 17184 21879
rect 17132 21836 17184 21845
rect 17500 21879 17552 21888
rect 17500 21845 17509 21879
rect 17509 21845 17543 21879
rect 17543 21845 17552 21879
rect 17500 21836 17552 21845
rect 18236 21836 18288 21888
rect 18328 21879 18380 21888
rect 18328 21845 18337 21879
rect 18337 21845 18371 21879
rect 18371 21845 18380 21879
rect 18880 21972 18932 22024
rect 19340 22015 19392 22024
rect 19340 21981 19349 22015
rect 19349 21981 19383 22015
rect 19383 21981 19392 22015
rect 19340 21972 19392 21981
rect 19708 22015 19760 22024
rect 19708 21981 19717 22015
rect 19717 21981 19751 22015
rect 19751 21981 19760 22015
rect 19708 21972 19760 21981
rect 20168 22015 20220 22024
rect 20168 21981 20177 22015
rect 20177 21981 20211 22015
rect 20211 21981 20220 22015
rect 20168 21972 20220 21981
rect 24124 22040 24176 22092
rect 20996 21972 21048 22024
rect 21088 21972 21140 22024
rect 21456 21972 21508 22024
rect 21824 22015 21876 22024
rect 21824 21981 21833 22015
rect 21833 21981 21867 22015
rect 21867 21981 21876 22015
rect 21824 21972 21876 21981
rect 22468 21972 22520 22024
rect 18328 21836 18380 21845
rect 18696 21836 18748 21888
rect 19616 21836 19668 21888
rect 20260 21836 20312 21888
rect 20812 21879 20864 21888
rect 20812 21845 20821 21879
rect 20821 21845 20855 21879
rect 20855 21845 20864 21879
rect 20812 21836 20864 21845
rect 20904 21836 20956 21888
rect 21272 21879 21324 21888
rect 21272 21845 21281 21879
rect 21281 21845 21315 21879
rect 21315 21845 21324 21879
rect 21272 21836 21324 21845
rect 23204 21904 23256 21956
rect 21640 21836 21692 21888
rect 22192 21836 22244 21888
rect 22836 21836 22888 21888
rect 6548 21734 6600 21786
rect 6612 21734 6664 21786
rect 6676 21734 6728 21786
rect 6740 21734 6792 21786
rect 6804 21734 6856 21786
rect 12146 21734 12198 21786
rect 12210 21734 12262 21786
rect 12274 21734 12326 21786
rect 12338 21734 12390 21786
rect 12402 21734 12454 21786
rect 17744 21734 17796 21786
rect 17808 21734 17860 21786
rect 17872 21734 17924 21786
rect 17936 21734 17988 21786
rect 18000 21734 18052 21786
rect 296 21632 348 21684
rect 2412 21675 2464 21684
rect 2412 21641 2421 21675
rect 2421 21641 2455 21675
rect 2455 21641 2464 21675
rect 2412 21632 2464 21641
rect 2964 21675 3016 21684
rect 2964 21641 2973 21675
rect 2973 21641 3007 21675
rect 3007 21641 3016 21675
rect 2964 21632 3016 21641
rect 3240 21675 3292 21684
rect 3240 21641 3249 21675
rect 3249 21641 3283 21675
rect 3283 21641 3292 21675
rect 3240 21632 3292 21641
rect 3700 21675 3752 21684
rect 3700 21641 3709 21675
rect 3709 21641 3743 21675
rect 3743 21641 3752 21675
rect 3700 21632 3752 21641
rect 4988 21675 5040 21684
rect 4988 21641 4997 21675
rect 4997 21641 5031 21675
rect 5031 21641 5040 21675
rect 4988 21632 5040 21641
rect 5632 21632 5684 21684
rect 6460 21632 6512 21684
rect 7840 21632 7892 21684
rect 8484 21632 8536 21684
rect 9496 21632 9548 21684
rect 11520 21632 11572 21684
rect 12532 21675 12584 21684
rect 4252 21564 4304 21616
rect 5448 21564 5500 21616
rect 6368 21564 6420 21616
rect 940 21360 992 21412
rect 2780 21496 2832 21548
rect 2964 21496 3016 21548
rect 3148 21539 3200 21548
rect 3148 21505 3157 21539
rect 3157 21505 3191 21539
rect 3191 21505 3200 21539
rect 3148 21496 3200 21505
rect 3424 21539 3476 21548
rect 3424 21505 3433 21539
rect 3433 21505 3467 21539
rect 3467 21505 3476 21539
rect 3424 21496 3476 21505
rect 3608 21496 3660 21548
rect 3976 21539 4028 21548
rect 3976 21505 3985 21539
rect 3985 21505 4019 21539
rect 4019 21505 4028 21539
rect 3976 21496 4028 21505
rect 5172 21539 5224 21548
rect 3240 21428 3292 21480
rect 4804 21428 4856 21480
rect 5172 21505 5181 21539
rect 5181 21505 5215 21539
rect 5215 21505 5224 21539
rect 5172 21496 5224 21505
rect 5724 21496 5776 21548
rect 7564 21564 7616 21616
rect 11888 21564 11940 21616
rect 12532 21641 12541 21675
rect 12541 21641 12575 21675
rect 12575 21641 12584 21675
rect 12532 21632 12584 21641
rect 13360 21632 13412 21684
rect 13728 21632 13780 21684
rect 15292 21632 15344 21684
rect 15660 21632 15712 21684
rect 15936 21632 15988 21684
rect 16120 21564 16172 21616
rect 16948 21632 17000 21684
rect 17592 21632 17644 21684
rect 18880 21675 18932 21684
rect 7656 21428 7708 21480
rect 7840 21471 7892 21480
rect 7840 21437 7849 21471
rect 7849 21437 7883 21471
rect 7883 21437 7892 21471
rect 7840 21428 7892 21437
rect 1400 21292 1452 21344
rect 6092 21360 6144 21412
rect 9496 21496 9548 21548
rect 10968 21496 11020 21548
rect 11520 21539 11572 21548
rect 11520 21505 11529 21539
rect 11529 21505 11563 21539
rect 11563 21505 11572 21539
rect 11520 21496 11572 21505
rect 11796 21496 11848 21548
rect 8852 21471 8904 21480
rect 8852 21437 8861 21471
rect 8861 21437 8895 21471
rect 8895 21437 8904 21471
rect 8852 21428 8904 21437
rect 9036 21471 9088 21480
rect 9036 21437 9045 21471
rect 9045 21437 9079 21471
rect 9079 21437 9088 21471
rect 9036 21428 9088 21437
rect 9220 21428 9272 21480
rect 9864 21471 9916 21480
rect 9864 21437 9873 21471
rect 9873 21437 9907 21471
rect 9907 21437 9916 21471
rect 9864 21428 9916 21437
rect 10324 21428 10376 21480
rect 11152 21360 11204 21412
rect 11704 21428 11756 21480
rect 12716 21428 12768 21480
rect 13176 21428 13228 21480
rect 15108 21496 15160 21548
rect 17408 21496 17460 21548
rect 18880 21641 18889 21675
rect 18889 21641 18923 21675
rect 18923 21641 18932 21675
rect 18880 21632 18932 21641
rect 18236 21564 18288 21616
rect 19340 21632 19392 21684
rect 20536 21675 20588 21684
rect 20536 21641 20545 21675
rect 20545 21641 20579 21675
rect 20579 21641 20588 21675
rect 20536 21632 20588 21641
rect 20628 21632 20680 21684
rect 21364 21632 21416 21684
rect 21824 21564 21876 21616
rect 19064 21539 19116 21548
rect 4528 21292 4580 21344
rect 5724 21292 5776 21344
rect 6276 21292 6328 21344
rect 7380 21335 7432 21344
rect 7380 21301 7389 21335
rect 7389 21301 7423 21335
rect 7423 21301 7432 21335
rect 7380 21292 7432 21301
rect 8392 21335 8444 21344
rect 8392 21301 8401 21335
rect 8401 21301 8435 21335
rect 8435 21301 8444 21335
rect 8392 21292 8444 21301
rect 8484 21292 8536 21344
rect 8944 21292 8996 21344
rect 10508 21292 10560 21344
rect 14372 21428 14424 21480
rect 13636 21360 13688 21412
rect 14188 21360 14240 21412
rect 15016 21428 15068 21480
rect 15292 21428 15344 21480
rect 14004 21292 14056 21344
rect 15200 21292 15252 21344
rect 16120 21428 16172 21480
rect 16764 21471 16816 21480
rect 16764 21437 16773 21471
rect 16773 21437 16807 21471
rect 16807 21437 16816 21471
rect 16764 21428 16816 21437
rect 17408 21360 17460 21412
rect 19064 21505 19073 21539
rect 19073 21505 19107 21539
rect 19107 21505 19116 21539
rect 19064 21496 19116 21505
rect 19892 21539 19944 21548
rect 19892 21505 19901 21539
rect 19901 21505 19935 21539
rect 19935 21505 19944 21539
rect 19892 21496 19944 21505
rect 20352 21539 20404 21548
rect 20352 21505 20361 21539
rect 20361 21505 20395 21539
rect 20395 21505 20404 21539
rect 20352 21496 20404 21505
rect 21088 21539 21140 21548
rect 21088 21505 21097 21539
rect 21097 21505 21131 21539
rect 21131 21505 21140 21539
rect 21088 21496 21140 21505
rect 19524 21428 19576 21480
rect 20168 21428 20220 21480
rect 21180 21428 21232 21480
rect 19708 21360 19760 21412
rect 19800 21360 19852 21412
rect 22192 21539 22244 21548
rect 22192 21505 22201 21539
rect 22201 21505 22235 21539
rect 22235 21505 22244 21539
rect 22192 21496 22244 21505
rect 21732 21428 21784 21480
rect 16028 21292 16080 21344
rect 17868 21292 17920 21344
rect 20628 21292 20680 21344
rect 21364 21292 21416 21344
rect 22100 21292 22152 21344
rect 23020 21335 23072 21344
rect 23020 21301 23029 21335
rect 23029 21301 23063 21335
rect 23063 21301 23072 21335
rect 23020 21292 23072 21301
rect 3749 21190 3801 21242
rect 3813 21190 3865 21242
rect 3877 21190 3929 21242
rect 3941 21190 3993 21242
rect 4005 21190 4057 21242
rect 9347 21190 9399 21242
rect 9411 21190 9463 21242
rect 9475 21190 9527 21242
rect 9539 21190 9591 21242
rect 9603 21190 9655 21242
rect 14945 21190 14997 21242
rect 15009 21190 15061 21242
rect 15073 21190 15125 21242
rect 15137 21190 15189 21242
rect 15201 21190 15253 21242
rect 20543 21190 20595 21242
rect 20607 21190 20659 21242
rect 20671 21190 20723 21242
rect 20735 21190 20787 21242
rect 20799 21190 20851 21242
rect 4068 21088 4120 21140
rect 4344 21131 4396 21140
rect 4344 21097 4353 21131
rect 4353 21097 4387 21131
rect 4387 21097 4396 21131
rect 4344 21088 4396 21097
rect 2780 21063 2832 21072
rect 2780 21029 2789 21063
rect 2789 21029 2823 21063
rect 2823 21029 2832 21063
rect 2780 21020 2832 21029
rect 2964 21020 3016 21072
rect 7840 21088 7892 21140
rect 9772 21131 9824 21140
rect 9772 21097 9781 21131
rect 9781 21097 9815 21131
rect 9815 21097 9824 21131
rect 9772 21088 9824 21097
rect 10232 21088 10284 21140
rect 8484 21020 8536 21072
rect 8668 21020 8720 21072
rect 9864 21020 9916 21072
rect 5448 20952 5500 21004
rect 7288 20995 7340 21004
rect 7288 20961 7297 20995
rect 7297 20961 7331 20995
rect 7331 20961 7340 20995
rect 7288 20952 7340 20961
rect 3424 20884 3476 20936
rect 3700 20884 3752 20936
rect 4344 20884 4396 20936
rect 6184 20884 6236 20936
rect 8300 20952 8352 21004
rect 8576 20995 8628 21004
rect 8576 20961 8585 20995
rect 8585 20961 8619 20995
rect 8619 20961 8628 20995
rect 8576 20952 8628 20961
rect 3148 20816 3200 20868
rect 3608 20748 3660 20800
rect 3884 20791 3936 20800
rect 3884 20757 3893 20791
rect 3893 20757 3927 20791
rect 3927 20757 3936 20791
rect 3884 20748 3936 20757
rect 4344 20748 4396 20800
rect 4988 20791 5040 20800
rect 4988 20757 4997 20791
rect 4997 20757 5031 20791
rect 5031 20757 5040 20791
rect 5356 20791 5408 20800
rect 4988 20748 5040 20757
rect 5356 20757 5365 20791
rect 5365 20757 5399 20791
rect 5399 20757 5408 20791
rect 5356 20748 5408 20757
rect 5448 20791 5500 20800
rect 5448 20757 5457 20791
rect 5457 20757 5491 20791
rect 5491 20757 5500 20791
rect 6460 20816 6512 20868
rect 7840 20884 7892 20936
rect 10324 20952 10376 21004
rect 10600 20952 10652 21004
rect 8944 20816 8996 20868
rect 9956 20816 10008 20868
rect 7472 20791 7524 20800
rect 5448 20748 5500 20757
rect 7472 20757 7481 20791
rect 7481 20757 7515 20791
rect 7515 20757 7524 20791
rect 7472 20748 7524 20757
rect 7932 20791 7984 20800
rect 7932 20757 7941 20791
rect 7941 20757 7975 20791
rect 7975 20757 7984 20791
rect 7932 20748 7984 20757
rect 8300 20748 8352 20800
rect 8484 20791 8536 20800
rect 8484 20757 8493 20791
rect 8493 20757 8527 20791
rect 8527 20757 8536 20791
rect 8484 20748 8536 20757
rect 8760 20748 8812 20800
rect 9772 20748 9824 20800
rect 10508 20791 10560 20800
rect 10508 20757 10523 20791
rect 10523 20757 10557 20791
rect 10557 20757 10560 20791
rect 10508 20748 10560 20757
rect 10692 20748 10744 20800
rect 12072 21020 12124 21072
rect 13544 21088 13596 21140
rect 13728 21131 13780 21140
rect 13728 21097 13737 21131
rect 13737 21097 13771 21131
rect 13771 21097 13780 21131
rect 13728 21088 13780 21097
rect 14832 21088 14884 21140
rect 14924 21088 14976 21140
rect 15476 21088 15528 21140
rect 15752 21088 15804 21140
rect 12900 21020 12952 21072
rect 16948 21020 17000 21072
rect 17224 21063 17276 21072
rect 17224 21029 17233 21063
rect 17233 21029 17267 21063
rect 17267 21029 17276 21063
rect 18144 21088 18196 21140
rect 18604 21131 18656 21140
rect 18604 21097 18613 21131
rect 18613 21097 18647 21131
rect 18647 21097 18656 21131
rect 18604 21088 18656 21097
rect 18972 21088 19024 21140
rect 20444 21088 20496 21140
rect 22652 21131 22704 21140
rect 17224 21020 17276 21029
rect 12808 20884 12860 20936
rect 12072 20816 12124 20868
rect 13636 20952 13688 21004
rect 14924 20952 14976 21004
rect 16304 20952 16356 21004
rect 16856 20952 16908 21004
rect 17592 20952 17644 21004
rect 17868 20995 17920 21004
rect 17868 20961 17877 20995
rect 17877 20961 17911 20995
rect 17911 20961 17920 20995
rect 18328 21020 18380 21072
rect 22652 21097 22661 21131
rect 22661 21097 22695 21131
rect 22695 21097 22704 21131
rect 22652 21088 22704 21097
rect 23204 21020 23256 21072
rect 17868 20952 17920 20961
rect 13912 20927 13964 20936
rect 13912 20893 13921 20927
rect 13921 20893 13955 20927
rect 13955 20893 13964 20927
rect 13912 20884 13964 20893
rect 14280 20927 14332 20936
rect 14280 20893 14289 20927
rect 14289 20893 14323 20927
rect 14323 20893 14332 20927
rect 14280 20884 14332 20893
rect 15384 20884 15436 20936
rect 17500 20884 17552 20936
rect 18512 20927 18564 20936
rect 18512 20893 18521 20927
rect 18521 20893 18555 20927
rect 18555 20893 18564 20927
rect 18512 20884 18564 20893
rect 18604 20884 18656 20936
rect 18880 20884 18932 20936
rect 21088 20952 21140 21004
rect 20260 20927 20312 20936
rect 20260 20893 20269 20927
rect 20269 20893 20303 20927
rect 20303 20893 20312 20927
rect 20260 20884 20312 20893
rect 16120 20816 16172 20868
rect 12532 20748 12584 20800
rect 12900 20791 12952 20800
rect 12900 20757 12909 20791
rect 12909 20757 12943 20791
rect 12943 20757 12952 20791
rect 12900 20748 12952 20757
rect 13452 20748 13504 20800
rect 14832 20748 14884 20800
rect 15384 20748 15436 20800
rect 16028 20748 16080 20800
rect 16212 20748 16264 20800
rect 16488 20791 16540 20800
rect 16488 20757 16497 20791
rect 16497 20757 16531 20791
rect 16531 20757 16540 20791
rect 16764 20791 16816 20800
rect 16488 20748 16540 20757
rect 16764 20757 16773 20791
rect 16773 20757 16807 20791
rect 16807 20757 16816 20791
rect 16764 20748 16816 20757
rect 17500 20748 17552 20800
rect 17684 20791 17736 20800
rect 17684 20757 17693 20791
rect 17693 20757 17727 20791
rect 17727 20757 17736 20791
rect 19708 20816 19760 20868
rect 20996 20884 21048 20936
rect 22284 20884 22336 20936
rect 22560 20884 22612 20936
rect 23112 20816 23164 20868
rect 17684 20748 17736 20757
rect 20720 20748 20772 20800
rect 20812 20748 20864 20800
rect 21548 20748 21600 20800
rect 21640 20748 21692 20800
rect 23020 20791 23072 20800
rect 23020 20757 23029 20791
rect 23029 20757 23063 20791
rect 23063 20757 23072 20791
rect 23020 20748 23072 20757
rect 6548 20646 6600 20698
rect 6612 20646 6664 20698
rect 6676 20646 6728 20698
rect 6740 20646 6792 20698
rect 6804 20646 6856 20698
rect 12146 20646 12198 20698
rect 12210 20646 12262 20698
rect 12274 20646 12326 20698
rect 12338 20646 12390 20698
rect 12402 20646 12454 20698
rect 17744 20646 17796 20698
rect 17808 20646 17860 20698
rect 17872 20646 17924 20698
rect 17936 20646 17988 20698
rect 18000 20646 18052 20698
rect 4988 20544 5040 20596
rect 5356 20544 5408 20596
rect 7196 20476 7248 20528
rect 4712 20408 4764 20460
rect 7104 20408 7156 20460
rect 6184 20383 6236 20392
rect 6184 20349 6193 20383
rect 6193 20349 6227 20383
rect 6227 20349 6236 20383
rect 6184 20340 6236 20349
rect 7472 20544 7524 20596
rect 8484 20544 8536 20596
rect 9772 20544 9824 20596
rect 9956 20544 10008 20596
rect 10692 20587 10744 20596
rect 10692 20553 10701 20587
rect 10701 20553 10735 20587
rect 10735 20553 10744 20587
rect 10692 20544 10744 20553
rect 11060 20544 11112 20596
rect 12532 20544 12584 20596
rect 7748 20451 7800 20460
rect 7748 20417 7757 20451
rect 7757 20417 7791 20451
rect 7791 20417 7800 20451
rect 7748 20408 7800 20417
rect 7932 20408 7984 20460
rect 8944 20451 8996 20460
rect 8024 20383 8076 20392
rect 1584 20272 1636 20324
rect 4620 20272 4672 20324
rect 2136 20204 2188 20256
rect 4804 20247 4856 20256
rect 4804 20213 4813 20247
rect 4813 20213 4847 20247
rect 4847 20213 4856 20247
rect 4804 20204 4856 20213
rect 6828 20204 6880 20256
rect 8024 20349 8033 20383
rect 8033 20349 8067 20383
rect 8067 20349 8076 20383
rect 8024 20340 8076 20349
rect 8392 20340 8444 20392
rect 8944 20417 8953 20451
rect 8953 20417 8987 20451
rect 8987 20417 8996 20451
rect 8944 20408 8996 20417
rect 10600 20451 10652 20460
rect 10600 20417 10609 20451
rect 10609 20417 10643 20451
rect 10643 20417 10652 20451
rect 10600 20408 10652 20417
rect 12900 20476 12952 20528
rect 13912 20544 13964 20596
rect 14648 20544 14700 20596
rect 15292 20544 15344 20596
rect 15660 20544 15712 20596
rect 16764 20544 16816 20596
rect 17500 20544 17552 20596
rect 18144 20544 18196 20596
rect 19892 20544 19944 20596
rect 20720 20544 20772 20596
rect 20904 20544 20956 20596
rect 22008 20544 22060 20596
rect 14280 20476 14332 20528
rect 16212 20476 16264 20528
rect 11796 20451 11848 20460
rect 11796 20417 11805 20451
rect 11805 20417 11839 20451
rect 11839 20417 11848 20451
rect 11796 20408 11848 20417
rect 12440 20451 12492 20460
rect 12440 20417 12449 20451
rect 12449 20417 12483 20451
rect 12483 20417 12492 20451
rect 12440 20408 12492 20417
rect 13084 20408 13136 20460
rect 14372 20408 14424 20460
rect 15844 20408 15896 20460
rect 10784 20383 10836 20392
rect 10784 20349 10793 20383
rect 10793 20349 10827 20383
rect 10827 20349 10836 20383
rect 10784 20340 10836 20349
rect 12256 20340 12308 20392
rect 13176 20383 13228 20392
rect 13176 20349 13185 20383
rect 13185 20349 13219 20383
rect 13219 20349 13228 20383
rect 13176 20340 13228 20349
rect 15200 20383 15252 20392
rect 8760 20204 8812 20256
rect 8852 20204 8904 20256
rect 11520 20204 11572 20256
rect 13636 20272 13688 20324
rect 15200 20349 15209 20383
rect 15209 20349 15243 20383
rect 15243 20349 15252 20383
rect 15200 20340 15252 20349
rect 15384 20340 15436 20392
rect 16580 20408 16632 20460
rect 19984 20408 20036 20460
rect 21364 20451 21416 20460
rect 16672 20340 16724 20392
rect 16856 20340 16908 20392
rect 17224 20383 17276 20392
rect 17224 20349 17233 20383
rect 17233 20349 17267 20383
rect 17267 20349 17276 20383
rect 17224 20340 17276 20349
rect 17408 20340 17460 20392
rect 18328 20383 18380 20392
rect 18328 20349 18340 20383
rect 18340 20349 18374 20383
rect 18374 20349 18380 20383
rect 18328 20340 18380 20349
rect 18512 20340 18564 20392
rect 12992 20204 13044 20256
rect 13912 20204 13964 20256
rect 16304 20272 16356 20324
rect 21364 20417 21373 20451
rect 21373 20417 21407 20451
rect 21407 20417 21416 20451
rect 21364 20408 21416 20417
rect 22836 20451 22888 20460
rect 22836 20417 22845 20451
rect 22845 20417 22879 20451
rect 22879 20417 22888 20451
rect 22836 20408 22888 20417
rect 22284 20383 22336 20392
rect 22284 20349 22293 20383
rect 22293 20349 22327 20383
rect 22327 20349 22336 20383
rect 22284 20340 22336 20349
rect 22560 20340 22612 20392
rect 14464 20204 14516 20256
rect 16396 20247 16448 20256
rect 16396 20213 16405 20247
rect 16405 20213 16439 20247
rect 16439 20213 16448 20247
rect 16396 20204 16448 20213
rect 18144 20204 18196 20256
rect 21456 20272 21508 20324
rect 23480 20272 23532 20324
rect 21088 20204 21140 20256
rect 21824 20247 21876 20256
rect 21824 20213 21833 20247
rect 21833 20213 21867 20247
rect 21867 20213 21876 20247
rect 21824 20204 21876 20213
rect 22652 20247 22704 20256
rect 22652 20213 22661 20247
rect 22661 20213 22695 20247
rect 22695 20213 22704 20247
rect 22652 20204 22704 20213
rect 23020 20247 23072 20256
rect 23020 20213 23029 20247
rect 23029 20213 23063 20247
rect 23063 20213 23072 20247
rect 23020 20204 23072 20213
rect 3749 20102 3801 20154
rect 3813 20102 3865 20154
rect 3877 20102 3929 20154
rect 3941 20102 3993 20154
rect 4005 20102 4057 20154
rect 9347 20102 9399 20154
rect 9411 20102 9463 20154
rect 9475 20102 9527 20154
rect 9539 20102 9591 20154
rect 9603 20102 9655 20154
rect 14945 20102 14997 20154
rect 15009 20102 15061 20154
rect 15073 20102 15125 20154
rect 15137 20102 15189 20154
rect 15201 20102 15253 20154
rect 20543 20102 20595 20154
rect 20607 20102 20659 20154
rect 20671 20102 20723 20154
rect 20735 20102 20787 20154
rect 20799 20102 20851 20154
rect 3148 19932 3200 19984
rect 8392 19932 8444 19984
rect 9220 20000 9272 20052
rect 10876 20043 10928 20052
rect 10876 20009 10885 20043
rect 10885 20009 10919 20043
rect 10919 20009 10928 20043
rect 10876 20000 10928 20009
rect 11152 20000 11204 20052
rect 12256 20043 12308 20052
rect 12256 20009 12265 20043
rect 12265 20009 12299 20043
rect 12299 20009 12308 20043
rect 12256 20000 12308 20009
rect 2228 19796 2280 19848
rect 3516 19839 3568 19848
rect 3516 19805 3525 19839
rect 3525 19805 3559 19839
rect 3559 19805 3568 19839
rect 3516 19796 3568 19805
rect 6184 19796 6236 19848
rect 6828 19796 6880 19848
rect 7196 19796 7248 19848
rect 2504 19660 2556 19712
rect 5172 19771 5224 19780
rect 5172 19737 5190 19771
rect 5190 19737 5224 19771
rect 5172 19728 5224 19737
rect 3976 19703 4028 19712
rect 3976 19669 3985 19703
rect 3985 19669 4019 19703
rect 4019 19669 4028 19703
rect 3976 19660 4028 19669
rect 5908 19728 5960 19780
rect 7288 19728 7340 19780
rect 5632 19660 5684 19712
rect 6460 19660 6512 19712
rect 8300 19660 8352 19712
rect 10600 19932 10652 19984
rect 11244 19932 11296 19984
rect 11980 19975 12032 19984
rect 11980 19941 11989 19975
rect 11989 19941 12023 19975
rect 12023 19941 12032 19975
rect 11980 19932 12032 19941
rect 12164 19975 12216 19984
rect 12164 19941 12173 19975
rect 12173 19941 12207 19975
rect 12207 19941 12216 19975
rect 12164 19932 12216 19941
rect 9220 19907 9272 19916
rect 9220 19873 9229 19907
rect 9229 19873 9263 19907
rect 9263 19873 9272 19907
rect 9220 19864 9272 19873
rect 12624 19864 12676 19916
rect 12900 19907 12952 19916
rect 12900 19873 12909 19907
rect 12909 19873 12943 19907
rect 12943 19873 12952 19907
rect 12900 19864 12952 19873
rect 8852 19796 8904 19848
rect 14004 20000 14056 20052
rect 14372 20043 14424 20052
rect 14372 20009 14381 20043
rect 14381 20009 14415 20043
rect 14415 20009 14424 20043
rect 14372 20000 14424 20009
rect 15292 20000 15344 20052
rect 16856 20043 16908 20052
rect 16856 20009 16865 20043
rect 16865 20009 16899 20043
rect 16899 20009 16908 20043
rect 16856 20000 16908 20009
rect 17592 20000 17644 20052
rect 18788 20043 18840 20052
rect 18788 20009 18797 20043
rect 18797 20009 18831 20043
rect 18831 20009 18840 20043
rect 18788 20000 18840 20009
rect 13728 19932 13780 19984
rect 14096 19932 14148 19984
rect 14556 19932 14608 19984
rect 15476 19932 15528 19984
rect 13360 19796 13412 19848
rect 13544 19796 13596 19848
rect 9496 19771 9548 19780
rect 9496 19737 9505 19771
rect 9505 19737 9539 19771
rect 9539 19737 9548 19771
rect 9496 19728 9548 19737
rect 11428 19771 11480 19780
rect 11428 19737 11437 19771
rect 11437 19737 11471 19771
rect 11471 19737 11480 19771
rect 11428 19728 11480 19737
rect 14464 19796 14516 19848
rect 14556 19796 14608 19848
rect 15292 19864 15344 19916
rect 16120 19907 16172 19916
rect 16120 19873 16129 19907
rect 16129 19873 16163 19907
rect 16163 19873 16172 19907
rect 16120 19864 16172 19873
rect 17500 19907 17552 19916
rect 16488 19796 16540 19848
rect 9864 19660 9916 19712
rect 10324 19660 10376 19712
rect 11152 19703 11204 19712
rect 11152 19669 11161 19703
rect 11161 19669 11195 19703
rect 11195 19669 11204 19703
rect 11152 19660 11204 19669
rect 11520 19660 11572 19712
rect 11888 19660 11940 19712
rect 12624 19703 12676 19712
rect 12624 19669 12633 19703
rect 12633 19669 12667 19703
rect 12667 19669 12676 19703
rect 12624 19660 12676 19669
rect 12716 19703 12768 19712
rect 12716 19669 12725 19703
rect 12725 19669 12759 19703
rect 12759 19669 12768 19703
rect 12716 19660 12768 19669
rect 13636 19703 13688 19712
rect 13636 19669 13645 19703
rect 13645 19669 13679 19703
rect 13679 19669 13688 19703
rect 13636 19660 13688 19669
rect 14740 19703 14792 19712
rect 14740 19669 14749 19703
rect 14749 19669 14783 19703
rect 14783 19669 14792 19703
rect 14740 19660 14792 19669
rect 14832 19703 14884 19712
rect 14832 19669 14841 19703
rect 14841 19669 14875 19703
rect 14875 19669 14884 19703
rect 14832 19660 14884 19669
rect 15660 19703 15712 19712
rect 15660 19669 15669 19703
rect 15669 19669 15703 19703
rect 15703 19669 15712 19703
rect 15660 19660 15712 19669
rect 16028 19660 16080 19712
rect 17500 19873 17509 19907
rect 17509 19873 17543 19907
rect 17543 19873 17552 19907
rect 17500 19864 17552 19873
rect 18144 19907 18196 19916
rect 18144 19873 18153 19907
rect 18153 19873 18187 19907
rect 18187 19873 18196 19907
rect 18144 19864 18196 19873
rect 18052 19839 18104 19848
rect 17040 19728 17092 19780
rect 18052 19805 18061 19839
rect 18061 19805 18095 19839
rect 18095 19805 18104 19839
rect 18052 19796 18104 19805
rect 18328 19796 18380 19848
rect 18420 19796 18472 19848
rect 20444 20000 20496 20052
rect 20536 20000 20588 20052
rect 22008 20000 22060 20052
rect 22284 20000 22336 20052
rect 21272 19864 21324 19916
rect 21456 19864 21508 19916
rect 19248 19839 19300 19848
rect 19248 19805 19257 19839
rect 19257 19805 19291 19839
rect 19291 19805 19300 19839
rect 19248 19796 19300 19805
rect 20536 19796 20588 19848
rect 20904 19839 20956 19848
rect 20904 19805 20913 19839
rect 20913 19805 20947 19839
rect 20947 19805 20956 19839
rect 20904 19796 20956 19805
rect 18696 19728 18748 19780
rect 19156 19660 19208 19712
rect 19432 19660 19484 19712
rect 20168 19728 20220 19780
rect 20720 19660 20772 19712
rect 21732 19796 21784 19848
rect 22928 19796 22980 19848
rect 21548 19660 21600 19712
rect 23020 19703 23072 19712
rect 23020 19669 23029 19703
rect 23029 19669 23063 19703
rect 23063 19669 23072 19703
rect 23020 19660 23072 19669
rect 6548 19558 6600 19610
rect 6612 19558 6664 19610
rect 6676 19558 6728 19610
rect 6740 19558 6792 19610
rect 6804 19558 6856 19610
rect 12146 19558 12198 19610
rect 12210 19558 12262 19610
rect 12274 19558 12326 19610
rect 12338 19558 12390 19610
rect 12402 19558 12454 19610
rect 17744 19558 17796 19610
rect 17808 19558 17860 19610
rect 17872 19558 17924 19610
rect 17936 19558 17988 19610
rect 18000 19558 18052 19610
rect 2412 19456 2464 19508
rect 3976 19456 4028 19508
rect 4436 19499 4488 19508
rect 4436 19465 4445 19499
rect 4445 19465 4479 19499
rect 4479 19465 4488 19499
rect 4436 19456 4488 19465
rect 4712 19499 4764 19508
rect 4712 19465 4721 19499
rect 4721 19465 4755 19499
rect 4755 19465 4764 19499
rect 4712 19456 4764 19465
rect 7748 19499 7800 19508
rect 7748 19465 7757 19499
rect 7757 19465 7791 19499
rect 7791 19465 7800 19499
rect 7748 19456 7800 19465
rect 8576 19456 8628 19508
rect 2596 19388 2648 19440
rect 3424 19388 3476 19440
rect 2044 19320 2096 19372
rect 2688 19320 2740 19372
rect 3332 19363 3384 19372
rect 3332 19329 3341 19363
rect 3341 19329 3375 19363
rect 3375 19329 3384 19363
rect 3332 19320 3384 19329
rect 2780 19252 2832 19304
rect 3240 19252 3292 19304
rect 4436 19320 4488 19372
rect 5540 19320 5592 19372
rect 8852 19363 8904 19372
rect 8852 19329 8861 19363
rect 8861 19329 8895 19363
rect 8895 19329 8904 19363
rect 8852 19320 8904 19329
rect 9772 19320 9824 19372
rect 9864 19320 9916 19372
rect 10876 19456 10928 19508
rect 11612 19456 11664 19508
rect 14740 19456 14792 19508
rect 15844 19499 15896 19508
rect 15844 19465 15853 19499
rect 15853 19465 15887 19499
rect 15887 19465 15896 19499
rect 15844 19456 15896 19465
rect 12900 19388 12952 19440
rect 12992 19320 13044 19372
rect 13268 19320 13320 19372
rect 3608 19184 3660 19236
rect 5080 19252 5132 19304
rect 8116 19252 8168 19304
rect 14832 19388 14884 19440
rect 14556 19320 14608 19372
rect 15752 19363 15804 19372
rect 15752 19329 15761 19363
rect 15761 19329 15795 19363
rect 15795 19329 15804 19363
rect 16396 19456 16448 19508
rect 16580 19456 16632 19508
rect 16672 19499 16724 19508
rect 16672 19465 16681 19499
rect 16681 19465 16715 19499
rect 16715 19465 16724 19499
rect 17040 19499 17092 19508
rect 16672 19456 16724 19465
rect 17040 19465 17049 19499
rect 17049 19465 17083 19499
rect 17083 19465 17092 19499
rect 17040 19456 17092 19465
rect 18144 19456 18196 19508
rect 18512 19456 18564 19508
rect 19340 19456 19392 19508
rect 16304 19388 16356 19440
rect 20720 19388 20772 19440
rect 21088 19388 21140 19440
rect 15752 19320 15804 19329
rect 17408 19320 17460 19372
rect 19064 19320 19116 19372
rect 20076 19363 20128 19372
rect 20076 19329 20094 19363
rect 20094 19329 20128 19363
rect 20076 19320 20128 19329
rect 20536 19363 20588 19372
rect 9680 19227 9732 19236
rect 9680 19193 9689 19227
rect 9689 19193 9723 19227
rect 9723 19193 9732 19227
rect 9680 19184 9732 19193
rect 12900 19295 12952 19304
rect 12900 19261 12909 19295
rect 12909 19261 12943 19295
rect 12943 19261 12952 19295
rect 13544 19295 13596 19304
rect 12900 19252 12952 19261
rect 13544 19261 13553 19295
rect 13553 19261 13587 19295
rect 13587 19261 13596 19295
rect 13544 19252 13596 19261
rect 1952 19116 2004 19168
rect 6092 19116 6144 19168
rect 6184 19116 6236 19168
rect 11152 19159 11204 19168
rect 11152 19125 11161 19159
rect 11161 19125 11195 19159
rect 11195 19125 11204 19159
rect 11152 19116 11204 19125
rect 13084 19116 13136 19168
rect 13636 19116 13688 19168
rect 14280 19159 14332 19168
rect 14280 19125 14289 19159
rect 14289 19125 14323 19159
rect 14323 19125 14332 19159
rect 14280 19116 14332 19125
rect 14372 19116 14424 19168
rect 19248 19252 19300 19304
rect 20536 19329 20545 19363
rect 20545 19329 20579 19363
rect 20579 19329 20588 19363
rect 20536 19320 20588 19329
rect 20904 19320 20956 19372
rect 22100 19320 22152 19372
rect 22376 19320 22428 19372
rect 21732 19252 21784 19304
rect 21916 19252 21968 19304
rect 22468 19295 22520 19304
rect 22468 19261 22477 19295
rect 22477 19261 22511 19295
rect 22511 19261 22520 19295
rect 22468 19252 22520 19261
rect 18512 19116 18564 19168
rect 21180 19116 21232 19168
rect 22008 19184 22060 19236
rect 22836 19184 22888 19236
rect 22284 19116 22336 19168
rect 22744 19159 22796 19168
rect 22744 19125 22753 19159
rect 22753 19125 22787 19159
rect 22787 19125 22796 19159
rect 22744 19116 22796 19125
rect 23020 19159 23072 19168
rect 23020 19125 23029 19159
rect 23029 19125 23063 19159
rect 23063 19125 23072 19159
rect 23020 19116 23072 19125
rect 3749 19014 3801 19066
rect 3813 19014 3865 19066
rect 3877 19014 3929 19066
rect 3941 19014 3993 19066
rect 4005 19014 4057 19066
rect 9347 19014 9399 19066
rect 9411 19014 9463 19066
rect 9475 19014 9527 19066
rect 9539 19014 9591 19066
rect 9603 19014 9655 19066
rect 14945 19014 14997 19066
rect 15009 19014 15061 19066
rect 15073 19014 15125 19066
rect 15137 19014 15189 19066
rect 15201 19014 15253 19066
rect 20543 19014 20595 19066
rect 20607 19014 20659 19066
rect 20671 19014 20723 19066
rect 20735 19014 20787 19066
rect 20799 19014 20851 19066
rect 3516 18912 3568 18964
rect 4344 18844 4396 18896
rect 1952 18776 2004 18828
rect 5632 18912 5684 18964
rect 5908 18955 5960 18964
rect 5908 18921 5917 18955
rect 5917 18921 5951 18955
rect 5951 18921 5960 18955
rect 5908 18912 5960 18921
rect 4252 18708 4304 18760
rect 4804 18708 4856 18760
rect 6184 18708 6236 18760
rect 1952 18640 2004 18692
rect 4160 18683 4212 18692
rect 4160 18649 4169 18683
rect 4169 18649 4203 18683
rect 4203 18649 4212 18683
rect 4160 18640 4212 18649
rect 6920 18640 6972 18692
rect 8024 18912 8076 18964
rect 10876 18912 10928 18964
rect 12992 18955 13044 18964
rect 12992 18921 13001 18955
rect 13001 18921 13035 18955
rect 13035 18921 13044 18955
rect 12992 18912 13044 18921
rect 13636 18912 13688 18964
rect 13084 18844 13136 18896
rect 15292 18912 15344 18964
rect 15844 18912 15896 18964
rect 17316 18912 17368 18964
rect 22008 18912 22060 18964
rect 22100 18912 22152 18964
rect 19432 18844 19484 18896
rect 20812 18844 20864 18896
rect 9036 18776 9088 18828
rect 13820 18776 13872 18828
rect 15752 18776 15804 18828
rect 1676 18572 1728 18624
rect 2320 18615 2372 18624
rect 2320 18581 2329 18615
rect 2329 18581 2363 18615
rect 2363 18581 2372 18615
rect 2688 18615 2740 18624
rect 2320 18572 2372 18581
rect 2688 18581 2697 18615
rect 2697 18581 2731 18615
rect 2731 18581 2740 18615
rect 2688 18572 2740 18581
rect 3240 18615 3292 18624
rect 3240 18581 3249 18615
rect 3249 18581 3283 18615
rect 3283 18581 3292 18615
rect 3240 18572 3292 18581
rect 4436 18615 4488 18624
rect 4436 18581 4445 18615
rect 4445 18581 4479 18615
rect 4479 18581 4488 18615
rect 4436 18572 4488 18581
rect 5356 18572 5408 18624
rect 8116 18572 8168 18624
rect 8300 18572 8352 18624
rect 9588 18708 9640 18760
rect 11152 18751 11204 18760
rect 11152 18717 11161 18751
rect 11161 18717 11195 18751
rect 11195 18717 11204 18751
rect 11152 18708 11204 18717
rect 12900 18708 12952 18760
rect 13452 18708 13504 18760
rect 8852 18640 8904 18692
rect 13728 18640 13780 18692
rect 14280 18708 14332 18760
rect 22468 18776 22520 18828
rect 22652 18776 22704 18828
rect 18880 18751 18932 18760
rect 18880 18717 18889 18751
rect 18889 18717 18923 18751
rect 18923 18717 18932 18751
rect 18880 18708 18932 18717
rect 19248 18708 19300 18760
rect 20720 18708 20772 18760
rect 22376 18708 22428 18760
rect 15936 18640 15988 18692
rect 16948 18640 17000 18692
rect 17592 18683 17644 18692
rect 17592 18649 17626 18683
rect 17626 18649 17644 18683
rect 17592 18640 17644 18649
rect 14556 18572 14608 18624
rect 17224 18615 17276 18624
rect 17224 18581 17233 18615
rect 17233 18581 17267 18615
rect 17267 18581 17276 18615
rect 17224 18572 17276 18581
rect 17408 18572 17460 18624
rect 19800 18640 19852 18692
rect 20444 18640 20496 18692
rect 21916 18640 21968 18692
rect 19708 18572 19760 18624
rect 22468 18572 22520 18624
rect 6548 18470 6600 18522
rect 6612 18470 6664 18522
rect 6676 18470 6728 18522
rect 6740 18470 6792 18522
rect 6804 18470 6856 18522
rect 12146 18470 12198 18522
rect 12210 18470 12262 18522
rect 12274 18470 12326 18522
rect 12338 18470 12390 18522
rect 12402 18470 12454 18522
rect 17744 18470 17796 18522
rect 17808 18470 17860 18522
rect 17872 18470 17924 18522
rect 17936 18470 17988 18522
rect 18000 18470 18052 18522
rect 2320 18368 2372 18420
rect 5356 18368 5408 18420
rect 5448 18368 5500 18420
rect 7840 18368 7892 18420
rect 9588 18368 9640 18420
rect 1860 18275 1912 18284
rect 1860 18241 1869 18275
rect 1869 18241 1903 18275
rect 1903 18241 1912 18275
rect 1860 18232 1912 18241
rect 2412 18232 2464 18284
rect 4068 18232 4120 18284
rect 4160 18232 4212 18284
rect 4620 18232 4672 18284
rect 3516 18164 3568 18216
rect 2964 18028 3016 18080
rect 6184 18164 6236 18216
rect 5080 18028 5132 18080
rect 8300 18232 8352 18284
rect 9772 18368 9824 18420
rect 14280 18368 14332 18420
rect 14648 18368 14700 18420
rect 15752 18368 15804 18420
rect 13084 18300 13136 18352
rect 13636 18343 13688 18352
rect 13636 18309 13645 18343
rect 13645 18309 13679 18343
rect 13679 18309 13688 18343
rect 13636 18300 13688 18309
rect 14740 18300 14792 18352
rect 14648 18232 14700 18284
rect 15292 18232 15344 18284
rect 13728 18207 13780 18216
rect 13728 18173 13737 18207
rect 13737 18173 13771 18207
rect 13771 18173 13780 18207
rect 13728 18164 13780 18173
rect 13820 18207 13872 18216
rect 13820 18173 13829 18207
rect 13829 18173 13863 18207
rect 13863 18173 13872 18207
rect 17592 18368 17644 18420
rect 19432 18368 19484 18420
rect 19616 18368 19668 18420
rect 20628 18368 20680 18420
rect 22744 18411 22796 18420
rect 17224 18232 17276 18284
rect 18512 18300 18564 18352
rect 18972 18300 19024 18352
rect 20260 18300 20312 18352
rect 13820 18164 13872 18173
rect 19248 18232 19300 18284
rect 19708 18232 19760 18284
rect 21272 18300 21324 18352
rect 22744 18377 22753 18411
rect 22753 18377 22787 18411
rect 22787 18377 22796 18411
rect 22744 18368 22796 18377
rect 23020 18411 23072 18420
rect 23020 18377 23029 18411
rect 23029 18377 23063 18411
rect 23063 18377 23072 18411
rect 23020 18368 23072 18377
rect 21180 18275 21232 18284
rect 21180 18241 21189 18275
rect 21189 18241 21223 18275
rect 21223 18241 21232 18275
rect 21180 18232 21232 18241
rect 21456 18275 21508 18284
rect 21456 18241 21465 18275
rect 21465 18241 21499 18275
rect 21499 18241 21508 18275
rect 21456 18232 21508 18241
rect 22836 18275 22888 18284
rect 22836 18241 22845 18275
rect 22845 18241 22879 18275
rect 22879 18241 22888 18275
rect 22836 18232 22888 18241
rect 13176 18096 13228 18148
rect 13636 18096 13688 18148
rect 8576 18028 8628 18080
rect 9220 18028 9272 18080
rect 9680 18028 9732 18080
rect 13912 18028 13964 18080
rect 14280 18028 14332 18080
rect 14372 18028 14424 18080
rect 15936 18028 15988 18080
rect 22192 18164 22244 18216
rect 22376 18207 22428 18216
rect 22376 18173 22385 18207
rect 22385 18173 22419 18207
rect 22419 18173 22428 18207
rect 22376 18164 22428 18173
rect 20720 18096 20772 18148
rect 22468 18096 22520 18148
rect 20996 18071 21048 18080
rect 20996 18037 21005 18071
rect 21005 18037 21039 18071
rect 21039 18037 21048 18071
rect 20996 18028 21048 18037
rect 22100 18028 22152 18080
rect 22192 18028 22244 18080
rect 22560 18028 22612 18080
rect 3749 17926 3801 17978
rect 3813 17926 3865 17978
rect 3877 17926 3929 17978
rect 3941 17926 3993 17978
rect 4005 17926 4057 17978
rect 9347 17926 9399 17978
rect 9411 17926 9463 17978
rect 9475 17926 9527 17978
rect 9539 17926 9591 17978
rect 9603 17926 9655 17978
rect 14945 17926 14997 17978
rect 15009 17926 15061 17978
rect 15073 17926 15125 17978
rect 15137 17926 15189 17978
rect 15201 17926 15253 17978
rect 20543 17926 20595 17978
rect 20607 17926 20659 17978
rect 20671 17926 20723 17978
rect 20735 17926 20787 17978
rect 20799 17926 20851 17978
rect 1952 17867 2004 17876
rect 1952 17833 1961 17867
rect 1961 17833 1995 17867
rect 1995 17833 2004 17867
rect 1952 17824 2004 17833
rect 3332 17824 3384 17876
rect 3424 17824 3476 17876
rect 5540 17824 5592 17876
rect 7196 17824 7248 17876
rect 9036 17824 9088 17876
rect 10968 17867 11020 17876
rect 10968 17833 10977 17867
rect 10977 17833 11011 17867
rect 11011 17833 11020 17867
rect 10968 17824 11020 17833
rect 12532 17824 12584 17876
rect 13912 17867 13964 17876
rect 13912 17833 13921 17867
rect 13921 17833 13955 17867
rect 13955 17833 13964 17867
rect 13912 17824 13964 17833
rect 2136 17688 2188 17740
rect 4160 17756 4212 17808
rect 3516 17731 3568 17740
rect 3516 17697 3525 17731
rect 3525 17697 3559 17731
rect 3559 17697 3568 17731
rect 3516 17688 3568 17697
rect 4252 17731 4304 17740
rect 4252 17697 4261 17731
rect 4261 17697 4295 17731
rect 4295 17697 4304 17731
rect 4252 17688 4304 17697
rect 15200 17824 15252 17876
rect 15476 17867 15528 17876
rect 15476 17833 15485 17867
rect 15485 17833 15519 17867
rect 15519 17833 15528 17867
rect 15476 17824 15528 17833
rect 4528 17688 4580 17740
rect 13452 17688 13504 17740
rect 15752 17824 15804 17876
rect 16948 17867 17000 17876
rect 16948 17833 16957 17867
rect 16957 17833 16991 17867
rect 16991 17833 17000 17867
rect 16948 17824 17000 17833
rect 17040 17824 17092 17876
rect 20352 17824 20404 17876
rect 20444 17824 20496 17876
rect 21088 17824 21140 17876
rect 21732 17824 21784 17876
rect 19064 17799 19116 17808
rect 19064 17765 19073 17799
rect 19073 17765 19107 17799
rect 19107 17765 19116 17799
rect 19064 17756 19116 17765
rect 2228 17620 2280 17672
rect 4344 17620 4396 17672
rect 6184 17620 6236 17672
rect 10784 17620 10836 17672
rect 3148 17552 3200 17604
rect 2688 17484 2740 17536
rect 4436 17484 4488 17536
rect 6000 17527 6052 17536
rect 6000 17493 6009 17527
rect 6009 17493 6043 17527
rect 6043 17493 6052 17527
rect 6368 17595 6420 17604
rect 6368 17561 6402 17595
rect 6402 17561 6420 17595
rect 6368 17552 6420 17561
rect 14188 17620 14240 17672
rect 18420 17731 18472 17740
rect 18420 17697 18429 17731
rect 18429 17697 18463 17731
rect 18463 17697 18472 17731
rect 19248 17731 19300 17740
rect 18420 17688 18472 17697
rect 19248 17697 19257 17731
rect 19257 17697 19291 17731
rect 19291 17697 19300 17731
rect 19248 17688 19300 17697
rect 21548 17688 21600 17740
rect 22652 17688 22704 17740
rect 22928 17731 22980 17740
rect 22928 17697 22937 17731
rect 22937 17697 22971 17731
rect 22971 17697 22980 17731
rect 22928 17688 22980 17697
rect 15844 17663 15896 17672
rect 15844 17629 15878 17663
rect 15878 17629 15896 17663
rect 15844 17620 15896 17629
rect 18144 17663 18196 17672
rect 18144 17629 18162 17663
rect 18162 17629 18196 17663
rect 18144 17620 18196 17629
rect 18880 17663 18932 17672
rect 14004 17552 14056 17604
rect 15384 17552 15436 17604
rect 16028 17552 16080 17604
rect 18512 17552 18564 17604
rect 18880 17629 18889 17663
rect 18889 17629 18923 17663
rect 18923 17629 18932 17663
rect 18880 17620 18932 17629
rect 20996 17620 21048 17672
rect 21088 17663 21140 17672
rect 21088 17629 21097 17663
rect 21097 17629 21131 17663
rect 21131 17629 21140 17663
rect 21088 17620 21140 17629
rect 21272 17620 21324 17672
rect 19340 17552 19392 17604
rect 19800 17552 19852 17604
rect 6000 17484 6052 17493
rect 8300 17484 8352 17536
rect 8484 17527 8536 17536
rect 8484 17493 8493 17527
rect 8493 17493 8527 17527
rect 8527 17493 8536 17527
rect 8484 17484 8536 17493
rect 12532 17527 12584 17536
rect 12532 17493 12541 17527
rect 12541 17493 12575 17527
rect 12575 17493 12584 17527
rect 12532 17484 12584 17493
rect 13084 17527 13136 17536
rect 13084 17493 13093 17527
rect 13093 17493 13127 17527
rect 13127 17493 13136 17527
rect 13084 17484 13136 17493
rect 13360 17484 13412 17536
rect 14280 17484 14332 17536
rect 14648 17484 14700 17536
rect 15200 17484 15252 17536
rect 15568 17484 15620 17536
rect 17224 17484 17276 17536
rect 20720 17484 20772 17536
rect 22652 17484 22704 17536
rect 6548 17382 6600 17434
rect 6612 17382 6664 17434
rect 6676 17382 6728 17434
rect 6740 17382 6792 17434
rect 6804 17382 6856 17434
rect 12146 17382 12198 17434
rect 12210 17382 12262 17434
rect 12274 17382 12326 17434
rect 12338 17382 12390 17434
rect 12402 17382 12454 17434
rect 17744 17382 17796 17434
rect 17808 17382 17860 17434
rect 17872 17382 17924 17434
rect 17936 17382 17988 17434
rect 18000 17382 18052 17434
rect 1860 17280 1912 17332
rect 2136 17280 2188 17332
rect 2596 17280 2648 17332
rect 3240 17280 3292 17332
rect 5172 17280 5224 17332
rect 8852 17280 8904 17332
rect 10784 17280 10836 17332
rect 12072 17280 12124 17332
rect 12532 17323 12584 17332
rect 12532 17289 12541 17323
rect 12541 17289 12575 17323
rect 12575 17289 12584 17323
rect 14188 17323 14240 17332
rect 12532 17280 12584 17289
rect 4528 17212 4580 17264
rect 6276 17212 6328 17264
rect 8576 17212 8628 17264
rect 8760 17255 8812 17264
rect 8760 17221 8794 17255
rect 8794 17221 8812 17255
rect 8760 17212 8812 17221
rect 9128 17212 9180 17264
rect 10968 17212 11020 17264
rect 11336 17212 11388 17264
rect 2872 17187 2924 17196
rect 2872 17153 2881 17187
rect 2881 17153 2915 17187
rect 2915 17153 2924 17187
rect 2872 17144 2924 17153
rect 1860 17076 1912 17128
rect 2504 17119 2556 17128
rect 2504 17085 2513 17119
rect 2513 17085 2547 17119
rect 2547 17085 2556 17119
rect 2504 17076 2556 17085
rect 2596 17076 2648 17128
rect 3148 17144 3200 17196
rect 4344 17144 4396 17196
rect 10508 17144 10560 17196
rect 14188 17289 14197 17323
rect 14197 17289 14231 17323
rect 14231 17289 14240 17323
rect 14188 17280 14240 17289
rect 16028 17280 16080 17332
rect 13176 17212 13228 17264
rect 13636 17212 13688 17264
rect 17132 17280 17184 17332
rect 17316 17323 17368 17332
rect 17316 17289 17325 17323
rect 17325 17289 17359 17323
rect 17359 17289 17368 17323
rect 17316 17280 17368 17289
rect 17408 17280 17460 17332
rect 17960 17280 18012 17332
rect 18512 17280 18564 17332
rect 3516 17119 3568 17128
rect 3516 17085 3525 17119
rect 3525 17085 3559 17119
rect 3559 17085 3568 17119
rect 3516 17076 3568 17085
rect 8484 17119 8536 17128
rect 2780 17008 2832 17060
rect 4436 17008 4488 17060
rect 1768 16940 1820 16992
rect 4252 16940 4304 16992
rect 5172 16940 5224 16992
rect 8484 17085 8493 17119
rect 8493 17085 8527 17119
rect 8527 17085 8536 17119
rect 8484 17076 8536 17085
rect 9772 17076 9824 17128
rect 11796 17119 11848 17128
rect 11796 17085 11805 17119
rect 11805 17085 11839 17119
rect 11839 17085 11848 17119
rect 11796 17076 11848 17085
rect 6184 16940 6236 16992
rect 13728 17008 13780 17060
rect 16948 17144 17000 17196
rect 17592 17144 17644 17196
rect 17868 17144 17920 17196
rect 18420 17212 18472 17264
rect 20996 17212 21048 17264
rect 20720 17144 20772 17196
rect 20904 17076 20956 17128
rect 21088 17119 21140 17128
rect 21088 17085 21097 17119
rect 21097 17085 21131 17119
rect 21131 17085 21140 17119
rect 21088 17076 21140 17085
rect 21272 17187 21324 17196
rect 21272 17153 21281 17187
rect 21281 17153 21315 17187
rect 21315 17153 21324 17187
rect 21272 17144 21324 17153
rect 22376 17280 22428 17332
rect 22928 17280 22980 17332
rect 22192 17187 22244 17196
rect 22192 17153 22201 17187
rect 22201 17153 22235 17187
rect 22235 17153 22244 17187
rect 22192 17144 22244 17153
rect 22376 17076 22428 17128
rect 17408 17008 17460 17060
rect 22744 17076 22796 17128
rect 12808 16940 12860 16992
rect 14004 16983 14056 16992
rect 14004 16949 14013 16983
rect 14013 16949 14047 16983
rect 14047 16949 14056 16983
rect 14004 16940 14056 16949
rect 16764 16983 16816 16992
rect 16764 16949 16773 16983
rect 16773 16949 16807 16983
rect 16807 16949 16816 16983
rect 16764 16940 16816 16949
rect 17040 16983 17092 16992
rect 17040 16949 17049 16983
rect 17049 16949 17083 16983
rect 17083 16949 17092 16983
rect 17040 16940 17092 16949
rect 19340 16983 19392 16992
rect 19340 16949 19349 16983
rect 19349 16949 19383 16983
rect 19383 16949 19392 16983
rect 21640 16983 21692 16992
rect 19340 16940 19392 16949
rect 21640 16949 21649 16983
rect 21649 16949 21683 16983
rect 21683 16949 21692 16983
rect 21640 16940 21692 16949
rect 22560 16983 22612 16992
rect 22560 16949 22569 16983
rect 22569 16949 22603 16983
rect 22603 16949 22612 16983
rect 22560 16940 22612 16949
rect 3749 16838 3801 16890
rect 3813 16838 3865 16890
rect 3877 16838 3929 16890
rect 3941 16838 3993 16890
rect 4005 16838 4057 16890
rect 9347 16838 9399 16890
rect 9411 16838 9463 16890
rect 9475 16838 9527 16890
rect 9539 16838 9591 16890
rect 9603 16838 9655 16890
rect 14945 16838 14997 16890
rect 15009 16838 15061 16890
rect 15073 16838 15125 16890
rect 15137 16838 15189 16890
rect 15201 16838 15253 16890
rect 20543 16838 20595 16890
rect 20607 16838 20659 16890
rect 20671 16838 20723 16890
rect 20735 16838 20787 16890
rect 20799 16838 20851 16890
rect 2872 16736 2924 16788
rect 4988 16736 5040 16788
rect 5724 16736 5776 16788
rect 8760 16779 8812 16788
rect 8760 16745 8769 16779
rect 8769 16745 8803 16779
rect 8803 16745 8812 16779
rect 8760 16736 8812 16745
rect 17132 16736 17184 16788
rect 1952 16668 2004 16720
rect 2780 16600 2832 16652
rect 2964 16643 3016 16652
rect 2964 16609 2973 16643
rect 2973 16609 3007 16643
rect 3007 16609 3016 16643
rect 2964 16600 3016 16609
rect 3976 16668 4028 16720
rect 4252 16643 4304 16652
rect 4252 16609 4261 16643
rect 4261 16609 4295 16643
rect 4295 16609 4304 16643
rect 4252 16600 4304 16609
rect 4436 16643 4488 16652
rect 4436 16609 4445 16643
rect 4445 16609 4479 16643
rect 4479 16609 4488 16643
rect 4436 16600 4488 16609
rect 2320 16532 2372 16584
rect 3516 16532 3568 16584
rect 8484 16600 8536 16652
rect 11796 16600 11848 16652
rect 13544 16600 13596 16652
rect 18420 16736 18472 16788
rect 19340 16736 19392 16788
rect 21272 16736 21324 16788
rect 22192 16736 22244 16788
rect 22744 16779 22796 16788
rect 22744 16745 22753 16779
rect 22753 16745 22787 16779
rect 22787 16745 22796 16779
rect 22744 16736 22796 16745
rect 3700 16464 3752 16516
rect 5540 16464 5592 16516
rect 6000 16464 6052 16516
rect 6184 16464 6236 16516
rect 9772 16575 9824 16584
rect 9772 16541 9781 16575
rect 9781 16541 9815 16575
rect 9815 16541 9824 16575
rect 9772 16532 9824 16541
rect 15476 16532 15528 16584
rect 17500 16532 17552 16584
rect 18144 16532 18196 16584
rect 19432 16600 19484 16652
rect 20904 16668 20956 16720
rect 21824 16668 21876 16720
rect 7840 16464 7892 16516
rect 11060 16507 11112 16516
rect 11060 16473 11078 16507
rect 11078 16473 11112 16507
rect 11060 16464 11112 16473
rect 1492 16396 1544 16448
rect 2872 16396 2924 16448
rect 3608 16439 3660 16448
rect 3608 16405 3617 16439
rect 3617 16405 3651 16439
rect 3651 16405 3660 16439
rect 3608 16396 3660 16405
rect 4160 16439 4212 16448
rect 4160 16405 4169 16439
rect 4169 16405 4203 16439
rect 4203 16405 4212 16439
rect 4160 16396 4212 16405
rect 6276 16396 6328 16448
rect 11244 16396 11296 16448
rect 11796 16439 11848 16448
rect 11796 16405 11805 16439
rect 11805 16405 11839 16439
rect 11839 16405 11848 16439
rect 11796 16396 11848 16405
rect 12992 16396 13044 16448
rect 16672 16464 16724 16516
rect 16304 16439 16356 16448
rect 16304 16405 16313 16439
rect 16313 16405 16347 16439
rect 16347 16405 16356 16439
rect 16304 16396 16356 16405
rect 18604 16396 18656 16448
rect 21088 16600 21140 16652
rect 21640 16600 21692 16652
rect 20904 16532 20956 16584
rect 21732 16532 21784 16584
rect 22652 16575 22704 16584
rect 22652 16541 22661 16575
rect 22661 16541 22695 16575
rect 22695 16541 22704 16575
rect 22652 16532 22704 16541
rect 20352 16507 20404 16516
rect 20352 16473 20370 16507
rect 20370 16473 20404 16507
rect 20352 16464 20404 16473
rect 20536 16464 20588 16516
rect 23204 16532 23256 16584
rect 19892 16396 19944 16448
rect 21456 16396 21508 16448
rect 22008 16439 22060 16448
rect 22008 16405 22017 16439
rect 22017 16405 22051 16439
rect 22051 16405 22060 16439
rect 22008 16396 22060 16405
rect 23020 16396 23072 16448
rect 6548 16294 6600 16346
rect 6612 16294 6664 16346
rect 6676 16294 6728 16346
rect 6740 16294 6792 16346
rect 6804 16294 6856 16346
rect 12146 16294 12198 16346
rect 12210 16294 12262 16346
rect 12274 16294 12326 16346
rect 12338 16294 12390 16346
rect 12402 16294 12454 16346
rect 17744 16294 17796 16346
rect 17808 16294 17860 16346
rect 17872 16294 17924 16346
rect 17936 16294 17988 16346
rect 18000 16294 18052 16346
rect 1676 16235 1728 16244
rect 1676 16201 1685 16235
rect 1685 16201 1719 16235
rect 1719 16201 1728 16235
rect 1676 16192 1728 16201
rect 1952 16235 2004 16244
rect 1952 16201 1961 16235
rect 1961 16201 1995 16235
rect 1995 16201 2004 16235
rect 1952 16192 2004 16201
rect 2412 16235 2464 16244
rect 2412 16201 2421 16235
rect 2421 16201 2455 16235
rect 2455 16201 2464 16235
rect 2412 16192 2464 16201
rect 2872 16235 2924 16244
rect 2872 16201 2881 16235
rect 2881 16201 2915 16235
rect 2915 16201 2924 16235
rect 2872 16192 2924 16201
rect 3516 16192 3568 16244
rect 3700 16235 3752 16244
rect 3700 16201 3709 16235
rect 3709 16201 3743 16235
rect 3743 16201 3752 16235
rect 3700 16192 3752 16201
rect 4804 16235 4856 16244
rect 4804 16201 4813 16235
rect 4813 16201 4847 16235
rect 4847 16201 4856 16235
rect 4804 16192 4856 16201
rect 1492 16099 1544 16108
rect 1492 16065 1501 16099
rect 1501 16065 1535 16099
rect 1535 16065 1544 16099
rect 1492 16056 1544 16065
rect 1768 16099 1820 16108
rect 1768 16065 1777 16099
rect 1777 16065 1811 16099
rect 1811 16065 1820 16099
rect 1768 16056 1820 16065
rect 5724 16124 5776 16176
rect 9588 16192 9640 16244
rect 9864 16235 9916 16244
rect 9864 16201 9873 16235
rect 9873 16201 9907 16235
rect 9907 16201 9916 16235
rect 9864 16192 9916 16201
rect 11796 16192 11848 16244
rect 14832 16192 14884 16244
rect 4344 16056 4396 16108
rect 9772 16099 9824 16108
rect 9772 16065 9781 16099
rect 9781 16065 9815 16099
rect 9815 16065 9824 16099
rect 9772 16056 9824 16065
rect 11152 16056 11204 16108
rect 11980 16056 12032 16108
rect 12808 16056 12860 16108
rect 15292 16056 15344 16108
rect 16304 16192 16356 16244
rect 18420 16192 18472 16244
rect 18604 16192 18656 16244
rect 18144 16124 18196 16176
rect 20536 16192 20588 16244
rect 21916 16192 21968 16244
rect 19616 16056 19668 16108
rect 20168 16124 20220 16176
rect 21548 16167 21600 16176
rect 21548 16133 21557 16167
rect 21557 16133 21591 16167
rect 21591 16133 21600 16167
rect 21548 16124 21600 16133
rect 19892 16056 19944 16108
rect 20904 16056 20956 16108
rect 21456 16056 21508 16108
rect 23112 16099 23164 16108
rect 3332 16031 3384 16040
rect 3332 15997 3341 16031
rect 3341 15997 3375 16031
rect 3375 15997 3384 16031
rect 3332 15988 3384 15997
rect 3516 16031 3568 16040
rect 3516 15997 3525 16031
rect 3525 15997 3559 16031
rect 3559 15997 3568 16031
rect 3516 15988 3568 15997
rect 3976 15988 4028 16040
rect 4160 15920 4212 15972
rect 18512 15988 18564 16040
rect 21732 15988 21784 16040
rect 21272 15920 21324 15972
rect 23112 16065 23121 16099
rect 23121 16065 23155 16099
rect 23155 16065 23164 16099
rect 23112 16056 23164 16065
rect 22376 15920 22428 15972
rect 5540 15852 5592 15904
rect 6184 15852 6236 15904
rect 8392 15895 8444 15904
rect 8392 15861 8401 15895
rect 8401 15861 8435 15895
rect 8435 15861 8444 15895
rect 8392 15852 8444 15861
rect 14280 15852 14332 15904
rect 16120 15852 16172 15904
rect 18420 15852 18472 15904
rect 21088 15852 21140 15904
rect 22928 15895 22980 15904
rect 22928 15861 22937 15895
rect 22937 15861 22971 15895
rect 22971 15861 22980 15895
rect 22928 15852 22980 15861
rect 3749 15750 3801 15802
rect 3813 15750 3865 15802
rect 3877 15750 3929 15802
rect 3941 15750 3993 15802
rect 4005 15750 4057 15802
rect 9347 15750 9399 15802
rect 9411 15750 9463 15802
rect 9475 15750 9527 15802
rect 9539 15750 9591 15802
rect 9603 15750 9655 15802
rect 14945 15750 14997 15802
rect 15009 15750 15061 15802
rect 15073 15750 15125 15802
rect 15137 15750 15189 15802
rect 15201 15750 15253 15802
rect 20543 15750 20595 15802
rect 20607 15750 20659 15802
rect 20671 15750 20723 15802
rect 20735 15750 20787 15802
rect 20799 15750 20851 15802
rect 2044 15648 2096 15700
rect 4344 15648 4396 15700
rect 10508 15648 10560 15700
rect 11980 15691 12032 15700
rect 11980 15657 11989 15691
rect 11989 15657 12023 15691
rect 12023 15657 12032 15691
rect 11980 15648 12032 15657
rect 15292 15648 15344 15700
rect 18236 15648 18288 15700
rect 18604 15691 18656 15700
rect 18604 15657 18613 15691
rect 18613 15657 18647 15691
rect 18647 15657 18656 15691
rect 18604 15648 18656 15657
rect 2688 15555 2740 15564
rect 2688 15521 2697 15555
rect 2697 15521 2731 15555
rect 2731 15521 2740 15555
rect 2688 15512 2740 15521
rect 4068 15512 4120 15564
rect 1676 15487 1728 15496
rect 1676 15453 1685 15487
rect 1685 15453 1719 15487
rect 1719 15453 1728 15487
rect 1676 15444 1728 15453
rect 3240 15487 3292 15496
rect 1492 15351 1544 15360
rect 1492 15317 1501 15351
rect 1501 15317 1535 15351
rect 1535 15317 1544 15351
rect 1492 15308 1544 15317
rect 3240 15453 3249 15487
rect 3249 15453 3283 15487
rect 3283 15453 3292 15487
rect 3240 15444 3292 15453
rect 5816 15580 5868 15632
rect 17500 15580 17552 15632
rect 20168 15648 20220 15700
rect 20352 15648 20404 15700
rect 20812 15555 20864 15564
rect 4804 15444 4856 15496
rect 9864 15444 9916 15496
rect 11612 15487 11664 15496
rect 11612 15453 11630 15487
rect 11630 15453 11664 15487
rect 11612 15444 11664 15453
rect 20812 15521 20821 15555
rect 20821 15521 20855 15555
rect 20855 15521 20864 15555
rect 20812 15512 20864 15521
rect 22008 15648 22060 15700
rect 21088 15580 21140 15632
rect 18420 15444 18472 15496
rect 18880 15487 18932 15496
rect 18880 15453 18889 15487
rect 18889 15453 18923 15487
rect 18923 15453 18932 15487
rect 18880 15444 18932 15453
rect 19156 15444 19208 15496
rect 19340 15444 19392 15496
rect 19892 15444 19944 15496
rect 21548 15487 21600 15496
rect 21548 15453 21557 15487
rect 21557 15453 21591 15487
rect 21591 15453 21600 15487
rect 21548 15444 21600 15453
rect 2780 15376 2832 15428
rect 2412 15351 2464 15360
rect 2412 15317 2421 15351
rect 2421 15317 2455 15351
rect 2455 15317 2464 15351
rect 2412 15308 2464 15317
rect 2872 15351 2924 15360
rect 2872 15317 2881 15351
rect 2881 15317 2915 15351
rect 2915 15317 2924 15351
rect 2872 15308 2924 15317
rect 3608 15308 3660 15360
rect 5724 15351 5776 15360
rect 5724 15317 5733 15351
rect 5733 15317 5767 15351
rect 5767 15317 5776 15351
rect 5724 15308 5776 15317
rect 6184 15376 6236 15428
rect 6460 15376 6512 15428
rect 8392 15376 8444 15428
rect 12532 15376 12584 15428
rect 13084 15376 13136 15428
rect 14372 15419 14424 15428
rect 8668 15351 8720 15360
rect 8668 15317 8677 15351
rect 8677 15317 8711 15351
rect 8711 15317 8720 15351
rect 8668 15308 8720 15317
rect 11060 15308 11112 15360
rect 13268 15308 13320 15360
rect 14372 15385 14406 15419
rect 14406 15385 14424 15419
rect 14372 15376 14424 15385
rect 14556 15376 14608 15428
rect 16672 15376 16724 15428
rect 19984 15376 20036 15428
rect 22468 15512 22520 15564
rect 23296 15580 23348 15632
rect 23664 15512 23716 15564
rect 21640 15308 21692 15360
rect 22284 15351 22336 15360
rect 22284 15317 22293 15351
rect 22293 15317 22327 15351
rect 22327 15317 22336 15351
rect 22284 15308 22336 15317
rect 22376 15351 22428 15360
rect 22376 15317 22385 15351
rect 22385 15317 22419 15351
rect 22419 15317 22428 15351
rect 22376 15308 22428 15317
rect 22652 15308 22704 15360
rect 6548 15206 6600 15258
rect 6612 15206 6664 15258
rect 6676 15206 6728 15258
rect 6740 15206 6792 15258
rect 6804 15206 6856 15258
rect 12146 15206 12198 15258
rect 12210 15206 12262 15258
rect 12274 15206 12326 15258
rect 12338 15206 12390 15258
rect 12402 15206 12454 15258
rect 17744 15206 17796 15258
rect 17808 15206 17860 15258
rect 17872 15206 17924 15258
rect 17936 15206 17988 15258
rect 18000 15206 18052 15258
rect 2320 15104 2372 15156
rect 2780 15104 2832 15156
rect 3332 15104 3384 15156
rect 6460 15104 6512 15156
rect 11336 15147 11388 15156
rect 11336 15113 11345 15147
rect 11345 15113 11379 15147
rect 11379 15113 11388 15147
rect 11336 15104 11388 15113
rect 11612 15104 11664 15156
rect 13176 15147 13228 15156
rect 13176 15113 13185 15147
rect 13185 15113 13219 15147
rect 13219 15113 13228 15147
rect 13176 15104 13228 15113
rect 1768 15011 1820 15020
rect 1768 14977 1777 15011
rect 1777 14977 1811 15011
rect 1811 14977 1820 15011
rect 1768 14968 1820 14977
rect 2596 14968 2648 15020
rect 4712 14968 4764 15020
rect 1584 14900 1636 14952
rect 2320 14943 2372 14952
rect 2320 14909 2329 14943
rect 2329 14909 2363 14943
rect 2363 14909 2372 14943
rect 2320 14900 2372 14909
rect 3516 14943 3568 14952
rect 2688 14832 2740 14884
rect 3148 14764 3200 14816
rect 3516 14909 3525 14943
rect 3525 14909 3559 14943
rect 3559 14909 3568 14943
rect 3516 14900 3568 14909
rect 4528 14943 4580 14952
rect 4528 14909 4537 14943
rect 4537 14909 4571 14943
rect 4571 14909 4580 14943
rect 4528 14900 4580 14909
rect 3424 14832 3476 14884
rect 6276 14968 6328 15020
rect 8668 15036 8720 15088
rect 10508 15036 10560 15088
rect 14280 15079 14332 15088
rect 14280 15045 14298 15079
rect 14298 15045 14332 15079
rect 14280 15036 14332 15045
rect 6460 14968 6512 15020
rect 14556 15011 14608 15020
rect 14556 14977 14565 15011
rect 14565 14977 14599 15011
rect 14599 14977 14608 15011
rect 18420 15104 18472 15156
rect 18604 15104 18656 15156
rect 19800 15147 19852 15156
rect 19800 15113 19809 15147
rect 19809 15113 19843 15147
rect 19843 15113 19852 15147
rect 19800 15104 19852 15113
rect 21272 15104 21324 15156
rect 21456 15147 21508 15156
rect 21456 15113 21465 15147
rect 21465 15113 21499 15147
rect 21499 15113 21508 15147
rect 21456 15104 21508 15113
rect 21732 15104 21784 15156
rect 21824 15104 21876 15156
rect 14556 14968 14608 14977
rect 22928 15036 22980 15088
rect 6000 14764 6052 14816
rect 6184 14764 6236 14816
rect 9864 14900 9916 14952
rect 18420 15011 18472 15020
rect 18420 14977 18429 15011
rect 18429 14977 18463 15011
rect 18463 14977 18472 15011
rect 18420 14968 18472 14977
rect 16580 14900 16632 14952
rect 21088 15011 21140 15020
rect 21088 14977 21097 15011
rect 21097 14977 21131 15011
rect 21131 14977 21140 15011
rect 21088 14968 21140 14977
rect 21456 14968 21508 15020
rect 10968 14832 11020 14884
rect 20812 14943 20864 14952
rect 20812 14909 20821 14943
rect 20821 14909 20855 14943
rect 20855 14909 20864 14943
rect 20812 14900 20864 14909
rect 20996 14943 21048 14952
rect 20996 14909 21005 14943
rect 21005 14909 21039 14943
rect 21039 14909 21048 14943
rect 20996 14900 21048 14909
rect 22468 14900 22520 14952
rect 23388 14832 23440 14884
rect 9772 14764 9824 14816
rect 18144 14764 18196 14816
rect 21732 14764 21784 14816
rect 23112 14807 23164 14816
rect 23112 14773 23121 14807
rect 23121 14773 23155 14807
rect 23155 14773 23164 14807
rect 23112 14764 23164 14773
rect 3749 14662 3801 14714
rect 3813 14662 3865 14714
rect 3877 14662 3929 14714
rect 3941 14662 3993 14714
rect 4005 14662 4057 14714
rect 9347 14662 9399 14714
rect 9411 14662 9463 14714
rect 9475 14662 9527 14714
rect 9539 14662 9591 14714
rect 9603 14662 9655 14714
rect 14945 14662 14997 14714
rect 15009 14662 15061 14714
rect 15073 14662 15125 14714
rect 15137 14662 15189 14714
rect 15201 14662 15253 14714
rect 20543 14662 20595 14714
rect 20607 14662 20659 14714
rect 20671 14662 20723 14714
rect 20735 14662 20787 14714
rect 20799 14662 20851 14714
rect 2320 14560 2372 14612
rect 2412 14560 2464 14612
rect 2964 14492 3016 14544
rect 1400 14424 1452 14476
rect 2688 14424 2740 14476
rect 2320 14356 2372 14408
rect 2872 14356 2924 14408
rect 3424 14492 3476 14544
rect 3516 14467 3568 14476
rect 3516 14433 3525 14467
rect 3525 14433 3559 14467
rect 3559 14433 3568 14467
rect 3516 14424 3568 14433
rect 4068 14356 4120 14408
rect 8484 14560 8536 14612
rect 12532 14560 12584 14612
rect 16580 14560 16632 14612
rect 4620 14492 4672 14544
rect 6368 14535 6420 14544
rect 6368 14501 6377 14535
rect 6377 14501 6411 14535
rect 6411 14501 6420 14535
rect 6368 14492 6420 14501
rect 4712 14424 4764 14476
rect 6184 14399 6236 14408
rect 6184 14365 6193 14399
rect 6193 14365 6227 14399
rect 6227 14365 6236 14399
rect 6184 14356 6236 14365
rect 5816 14288 5868 14340
rect 5908 14331 5960 14340
rect 5908 14297 5948 14331
rect 5948 14297 5960 14331
rect 5908 14288 5960 14297
rect 3884 14220 3936 14272
rect 6368 14220 6420 14272
rect 7472 14331 7524 14340
rect 7472 14297 7490 14331
rect 7490 14297 7524 14331
rect 16948 14467 17000 14476
rect 16948 14433 16957 14467
rect 16957 14433 16991 14467
rect 16991 14433 17000 14467
rect 18420 14560 18472 14612
rect 18880 14492 18932 14544
rect 19432 14560 19484 14612
rect 21456 14603 21508 14612
rect 21456 14569 21465 14603
rect 21465 14569 21499 14603
rect 21499 14569 21508 14603
rect 21456 14560 21508 14569
rect 21548 14560 21600 14612
rect 21916 14560 21968 14612
rect 22744 14560 22796 14612
rect 23480 14492 23532 14544
rect 19248 14467 19300 14476
rect 16948 14424 17000 14433
rect 19248 14433 19257 14467
rect 19257 14433 19291 14467
rect 19291 14433 19300 14467
rect 19248 14424 19300 14433
rect 20812 14424 20864 14476
rect 7472 14288 7524 14297
rect 9956 14288 10008 14340
rect 9680 14220 9732 14272
rect 9864 14220 9916 14272
rect 13360 14399 13412 14408
rect 13360 14365 13378 14399
rect 13378 14365 13412 14399
rect 13360 14356 13412 14365
rect 13544 14356 13596 14408
rect 14096 14399 14148 14408
rect 14096 14365 14105 14399
rect 14105 14365 14139 14399
rect 14139 14365 14148 14399
rect 14096 14356 14148 14365
rect 13268 14288 13320 14340
rect 17224 14356 17276 14408
rect 19156 14356 19208 14408
rect 20720 14356 20772 14408
rect 21640 14399 21692 14408
rect 21640 14365 21649 14399
rect 21649 14365 21683 14399
rect 21683 14365 21692 14399
rect 21640 14356 21692 14365
rect 21732 14356 21784 14408
rect 22192 14356 22244 14408
rect 22928 14356 22980 14408
rect 14740 14288 14792 14340
rect 16672 14331 16724 14340
rect 16672 14297 16690 14331
rect 16690 14297 16724 14331
rect 16672 14288 16724 14297
rect 19432 14288 19484 14340
rect 19616 14288 19668 14340
rect 10968 14263 11020 14272
rect 10968 14229 10977 14263
rect 10977 14229 11011 14263
rect 11011 14229 11020 14263
rect 10968 14220 11020 14229
rect 15752 14220 15804 14272
rect 20260 14220 20312 14272
rect 20536 14220 20588 14272
rect 21732 14220 21784 14272
rect 6548 14118 6600 14170
rect 6612 14118 6664 14170
rect 6676 14118 6728 14170
rect 6740 14118 6792 14170
rect 6804 14118 6856 14170
rect 12146 14118 12198 14170
rect 12210 14118 12262 14170
rect 12274 14118 12326 14170
rect 12338 14118 12390 14170
rect 12402 14118 12454 14170
rect 17744 14118 17796 14170
rect 17808 14118 17860 14170
rect 17872 14118 17924 14170
rect 17936 14118 17988 14170
rect 18000 14118 18052 14170
rect 2320 14059 2372 14068
rect 2320 14025 2329 14059
rect 2329 14025 2363 14059
rect 2363 14025 2372 14059
rect 2320 14016 2372 14025
rect 3884 14016 3936 14068
rect 4160 14016 4212 14068
rect 5172 14016 5224 14068
rect 5816 14016 5868 14068
rect 8484 14059 8536 14068
rect 5632 13880 5684 13932
rect 6368 13880 6420 13932
rect 6552 13948 6604 14000
rect 8484 14025 8493 14059
rect 8493 14025 8527 14059
rect 8527 14025 8536 14059
rect 8484 14016 8536 14025
rect 9956 14059 10008 14068
rect 7472 13880 7524 13932
rect 7840 13923 7892 13932
rect 7840 13889 7858 13923
rect 7858 13889 7892 13923
rect 7840 13880 7892 13889
rect 9772 13948 9824 14000
rect 9956 14025 9965 14059
rect 9965 14025 9999 14059
rect 9999 14025 10008 14059
rect 9956 14016 10008 14025
rect 11244 14016 11296 14068
rect 14740 14059 14792 14068
rect 14740 14025 14749 14059
rect 14749 14025 14783 14059
rect 14783 14025 14792 14059
rect 14740 14016 14792 14025
rect 10968 13948 11020 14000
rect 13268 13948 13320 14000
rect 2688 13812 2740 13864
rect 4436 13855 4488 13864
rect 4436 13821 4445 13855
rect 4445 13821 4479 13855
rect 4479 13821 4488 13855
rect 4436 13812 4488 13821
rect 4712 13812 4764 13864
rect 6184 13855 6236 13864
rect 6184 13821 6193 13855
rect 6193 13821 6227 13855
rect 6227 13821 6236 13855
rect 6184 13812 6236 13821
rect 6460 13812 6512 13864
rect 9864 13855 9916 13864
rect 6184 13676 6236 13728
rect 9864 13821 9873 13855
rect 9873 13821 9907 13855
rect 9907 13821 9916 13855
rect 9864 13812 9916 13821
rect 13084 13923 13136 13932
rect 13084 13889 13093 13923
rect 13093 13889 13127 13923
rect 13127 13889 13136 13923
rect 14096 13948 14148 14000
rect 16948 14016 17000 14068
rect 18144 14016 18196 14068
rect 18880 14016 18932 14068
rect 19248 14016 19300 14068
rect 21548 14059 21600 14068
rect 13084 13880 13136 13889
rect 14188 13880 14240 13932
rect 15384 13923 15436 13932
rect 15384 13889 15418 13923
rect 15418 13889 15436 13923
rect 15384 13880 15436 13889
rect 16672 13880 16724 13932
rect 19340 13948 19392 14000
rect 19248 13880 19300 13932
rect 20536 13880 20588 13932
rect 21548 14025 21557 14059
rect 21557 14025 21591 14059
rect 21591 14025 21600 14059
rect 21548 14016 21600 14025
rect 22928 14059 22980 14068
rect 22928 14025 22937 14059
rect 22937 14025 22971 14059
rect 22971 14025 22980 14059
rect 22928 14016 22980 14025
rect 20720 13948 20772 14000
rect 22560 13948 22612 14000
rect 21916 13880 21968 13932
rect 19616 13812 19668 13864
rect 20812 13855 20864 13864
rect 20812 13821 20821 13855
rect 20821 13821 20855 13855
rect 20855 13821 20864 13855
rect 20812 13812 20864 13821
rect 20996 13855 21048 13864
rect 20996 13821 21005 13855
rect 21005 13821 21039 13855
rect 21039 13821 21048 13855
rect 20996 13812 21048 13821
rect 8392 13676 8444 13728
rect 21088 13744 21140 13796
rect 21824 13812 21876 13864
rect 23112 13923 23164 13932
rect 23112 13889 23121 13923
rect 23121 13889 23155 13923
rect 23155 13889 23164 13923
rect 23112 13880 23164 13889
rect 15752 13676 15804 13728
rect 21272 13676 21324 13728
rect 21364 13676 21416 13728
rect 21824 13676 21876 13728
rect 22652 13676 22704 13728
rect 22836 13719 22888 13728
rect 22836 13685 22845 13719
rect 22845 13685 22879 13719
rect 22879 13685 22888 13719
rect 22836 13676 22888 13685
rect 3749 13574 3801 13626
rect 3813 13574 3865 13626
rect 3877 13574 3929 13626
rect 3941 13574 3993 13626
rect 4005 13574 4057 13626
rect 9347 13574 9399 13626
rect 9411 13574 9463 13626
rect 9475 13574 9527 13626
rect 9539 13574 9591 13626
rect 9603 13574 9655 13626
rect 14945 13574 14997 13626
rect 15009 13574 15061 13626
rect 15073 13574 15125 13626
rect 15137 13574 15189 13626
rect 15201 13574 15253 13626
rect 20543 13574 20595 13626
rect 20607 13574 20659 13626
rect 20671 13574 20723 13626
rect 20735 13574 20787 13626
rect 20799 13574 20851 13626
rect 1676 13472 1728 13524
rect 2228 13472 2280 13524
rect 6276 13515 6328 13524
rect 6276 13481 6285 13515
rect 6285 13481 6319 13515
rect 6319 13481 6328 13515
rect 6276 13472 6328 13481
rect 3240 13404 3292 13456
rect 4896 13404 4948 13456
rect 6000 13404 6052 13456
rect 7840 13472 7892 13524
rect 9680 13472 9732 13524
rect 10968 13472 11020 13524
rect 3148 13379 3200 13388
rect 3148 13345 3157 13379
rect 3157 13345 3191 13379
rect 3191 13345 3200 13379
rect 3148 13336 3200 13345
rect 19156 13472 19208 13524
rect 14096 13447 14148 13456
rect 14096 13413 14105 13447
rect 14105 13413 14139 13447
rect 14139 13413 14148 13447
rect 14096 13404 14148 13413
rect 18144 13404 18196 13456
rect 20904 13472 20956 13524
rect 21548 13515 21600 13524
rect 21548 13481 21557 13515
rect 21557 13481 21591 13515
rect 21591 13481 21600 13515
rect 21548 13472 21600 13481
rect 22284 13472 22336 13524
rect 22928 13472 22980 13524
rect 18604 13379 18656 13388
rect 18604 13345 18613 13379
rect 18613 13345 18647 13379
rect 18647 13345 18656 13379
rect 18604 13336 18656 13345
rect 19248 13336 19300 13388
rect 21088 13336 21140 13388
rect 22192 13336 22244 13388
rect 2964 13311 3016 13320
rect 2964 13277 2973 13311
rect 2973 13277 3007 13311
rect 3007 13277 3016 13311
rect 2964 13268 3016 13277
rect 4712 13311 4764 13320
rect 4712 13277 4721 13311
rect 4721 13277 4755 13311
rect 4755 13277 4764 13311
rect 4712 13268 4764 13277
rect 5172 13311 5224 13320
rect 5172 13277 5206 13311
rect 5206 13277 5224 13311
rect 2688 13200 2740 13252
rect 3424 13200 3476 13252
rect 2136 13175 2188 13184
rect 2136 13141 2145 13175
rect 2145 13141 2179 13175
rect 2179 13141 2188 13175
rect 2136 13132 2188 13141
rect 3056 13175 3108 13184
rect 3056 13141 3065 13175
rect 3065 13141 3099 13175
rect 3099 13141 3108 13175
rect 3056 13132 3108 13141
rect 4804 13132 4856 13184
rect 5172 13268 5224 13277
rect 17040 13311 17092 13320
rect 6092 13200 6144 13252
rect 6184 13132 6236 13184
rect 17040 13277 17049 13311
rect 17049 13277 17083 13311
rect 17083 13277 17092 13311
rect 17040 13268 17092 13277
rect 18512 13268 18564 13320
rect 20996 13268 21048 13320
rect 21272 13268 21324 13320
rect 22560 13404 22612 13456
rect 22652 13336 22704 13388
rect 8484 13200 8536 13252
rect 11520 13200 11572 13252
rect 15660 13200 15712 13252
rect 16120 13200 16172 13252
rect 10324 13175 10376 13184
rect 10324 13141 10333 13175
rect 10333 13141 10367 13175
rect 10367 13141 10376 13175
rect 10324 13132 10376 13141
rect 19616 13200 19668 13252
rect 19064 13175 19116 13184
rect 19064 13141 19073 13175
rect 19073 13141 19107 13175
rect 19107 13141 19116 13175
rect 19064 13132 19116 13141
rect 19248 13132 19300 13184
rect 20720 13132 20772 13184
rect 22192 13200 22244 13252
rect 22008 13175 22060 13184
rect 22008 13141 22017 13175
rect 22017 13141 22051 13175
rect 22051 13141 22060 13175
rect 22008 13132 22060 13141
rect 22652 13132 22704 13184
rect 6548 13030 6600 13082
rect 6612 13030 6664 13082
rect 6676 13030 6728 13082
rect 6740 13030 6792 13082
rect 6804 13030 6856 13082
rect 12146 13030 12198 13082
rect 12210 13030 12262 13082
rect 12274 13030 12326 13082
rect 12338 13030 12390 13082
rect 12402 13030 12454 13082
rect 17744 13030 17796 13082
rect 17808 13030 17860 13082
rect 17872 13030 17924 13082
rect 17936 13030 17988 13082
rect 18000 13030 18052 13082
rect 2228 12928 2280 12980
rect 6184 12928 6236 12980
rect 6368 12971 6420 12980
rect 6368 12937 6377 12971
rect 6377 12937 6411 12971
rect 6411 12937 6420 12971
rect 6368 12928 6420 12937
rect 8392 12971 8444 12980
rect 8392 12937 8401 12971
rect 8401 12937 8435 12971
rect 8435 12937 8444 12971
rect 8392 12928 8444 12937
rect 13084 12971 13136 12980
rect 13084 12937 13093 12971
rect 13093 12937 13127 12971
rect 13127 12937 13136 12971
rect 13084 12928 13136 12937
rect 16212 12928 16264 12980
rect 17040 12928 17092 12980
rect 3608 12860 3660 12912
rect 6276 12860 6328 12912
rect 9864 12860 9916 12912
rect 2872 12835 2924 12844
rect 2872 12801 2881 12835
rect 2881 12801 2915 12835
rect 2915 12801 2924 12835
rect 2872 12792 2924 12801
rect 4252 12792 4304 12844
rect 2964 12767 3016 12776
rect 2964 12733 2973 12767
rect 2973 12733 3007 12767
rect 3007 12733 3016 12767
rect 2964 12724 3016 12733
rect 2688 12656 2740 12708
rect 3240 12724 3292 12776
rect 3424 12724 3476 12776
rect 4804 12767 4856 12776
rect 2780 12588 2832 12640
rect 4804 12733 4813 12767
rect 4813 12733 4847 12767
rect 4847 12733 4856 12767
rect 4804 12724 4856 12733
rect 6368 12792 6420 12844
rect 10324 12792 10376 12844
rect 11060 12835 11112 12844
rect 11060 12801 11089 12835
rect 11089 12801 11112 12835
rect 11060 12792 11112 12801
rect 9864 12767 9916 12776
rect 9864 12733 9873 12767
rect 9873 12733 9907 12767
rect 9907 12733 9916 12767
rect 9864 12724 9916 12733
rect 12900 12792 12952 12844
rect 13912 12792 13964 12844
rect 18144 12860 18196 12912
rect 16580 12792 16632 12844
rect 18604 12928 18656 12980
rect 20996 12928 21048 12980
rect 22100 12971 22152 12980
rect 22100 12937 22109 12971
rect 22109 12937 22143 12971
rect 22143 12937 22152 12971
rect 22100 12928 22152 12937
rect 22376 12928 22428 12980
rect 23112 12971 23164 12980
rect 23112 12937 23121 12971
rect 23121 12937 23155 12971
rect 23155 12937 23164 12971
rect 23112 12928 23164 12937
rect 19156 12860 19208 12912
rect 18420 12792 18472 12844
rect 18880 12792 18932 12844
rect 20260 12860 20312 12912
rect 20444 12792 20496 12844
rect 21088 12860 21140 12912
rect 23204 12860 23256 12912
rect 23480 12792 23532 12844
rect 4528 12656 4580 12708
rect 8484 12699 8536 12708
rect 8484 12665 8493 12699
rect 8493 12665 8527 12699
rect 8527 12665 8536 12699
rect 8484 12656 8536 12665
rect 21640 12724 21692 12776
rect 22468 12724 22520 12776
rect 23204 12724 23256 12776
rect 23388 12724 23440 12776
rect 16120 12699 16172 12708
rect 16120 12665 16129 12699
rect 16129 12665 16163 12699
rect 16163 12665 16172 12699
rect 16120 12656 16172 12665
rect 9680 12588 9732 12640
rect 16580 12588 16632 12640
rect 19248 12588 19300 12640
rect 21088 12588 21140 12640
rect 22100 12588 22152 12640
rect 3749 12486 3801 12538
rect 3813 12486 3865 12538
rect 3877 12486 3929 12538
rect 3941 12486 3993 12538
rect 4005 12486 4057 12538
rect 9347 12486 9399 12538
rect 9411 12486 9463 12538
rect 9475 12486 9527 12538
rect 9539 12486 9591 12538
rect 9603 12486 9655 12538
rect 14945 12486 14997 12538
rect 15009 12486 15061 12538
rect 15073 12486 15125 12538
rect 15137 12486 15189 12538
rect 15201 12486 15253 12538
rect 20543 12486 20595 12538
rect 20607 12486 20659 12538
rect 20671 12486 20723 12538
rect 20735 12486 20787 12538
rect 20799 12486 20851 12538
rect 1768 12384 1820 12436
rect 2872 12384 2924 12436
rect 2688 12291 2740 12300
rect 2688 12257 2697 12291
rect 2697 12257 2731 12291
rect 2731 12257 2740 12291
rect 2688 12248 2740 12257
rect 3608 12248 3660 12300
rect 3516 12180 3568 12232
rect 5908 12384 5960 12436
rect 16580 12384 16632 12436
rect 18512 12427 18564 12436
rect 18512 12393 18521 12427
rect 18521 12393 18555 12427
rect 18555 12393 18564 12427
rect 18512 12384 18564 12393
rect 20720 12384 20772 12436
rect 20812 12384 20864 12436
rect 18788 12359 18840 12368
rect 4804 12248 4856 12300
rect 9680 12248 9732 12300
rect 2872 12112 2924 12164
rect 6368 12223 6420 12232
rect 6368 12189 6377 12223
rect 6377 12189 6411 12223
rect 6411 12189 6420 12223
rect 6368 12180 6420 12189
rect 9864 12180 9916 12232
rect 5264 12112 5316 12164
rect 6184 12112 6236 12164
rect 2504 12087 2556 12096
rect 2504 12053 2513 12087
rect 2513 12053 2547 12087
rect 2547 12053 2556 12087
rect 2504 12044 2556 12053
rect 3332 12044 3384 12096
rect 3608 12087 3660 12096
rect 3608 12053 3617 12087
rect 3617 12053 3651 12087
rect 3651 12053 3660 12087
rect 3608 12044 3660 12053
rect 4068 12087 4120 12096
rect 4068 12053 4077 12087
rect 4077 12053 4111 12087
rect 4111 12053 4120 12087
rect 4068 12044 4120 12053
rect 6276 12087 6328 12096
rect 6276 12053 6285 12087
rect 6285 12053 6319 12087
rect 6319 12053 6328 12087
rect 6276 12044 6328 12053
rect 6460 12044 6512 12096
rect 9312 12112 9364 12164
rect 7840 12087 7892 12096
rect 7840 12053 7849 12087
rect 7849 12053 7883 12087
rect 7883 12053 7892 12087
rect 7840 12044 7892 12053
rect 10324 12155 10376 12164
rect 10324 12121 10358 12155
rect 10358 12121 10376 12155
rect 10324 12112 10376 12121
rect 13084 12180 13136 12232
rect 16212 12248 16264 12300
rect 18788 12325 18797 12359
rect 18797 12325 18831 12359
rect 18831 12325 18840 12359
rect 18788 12316 18840 12325
rect 19064 12359 19116 12368
rect 19064 12325 19073 12359
rect 19073 12325 19107 12359
rect 19107 12325 19116 12359
rect 19064 12316 19116 12325
rect 16580 12223 16632 12232
rect 16580 12189 16614 12223
rect 16614 12189 16632 12223
rect 16580 12180 16632 12189
rect 18880 12223 18932 12232
rect 14096 12112 14148 12164
rect 18512 12112 18564 12164
rect 18880 12189 18889 12223
rect 18889 12189 18923 12223
rect 18923 12189 18932 12223
rect 18880 12180 18932 12189
rect 19156 12248 19208 12300
rect 20812 12291 20864 12300
rect 20812 12257 20821 12291
rect 20821 12257 20855 12291
rect 20855 12257 20864 12291
rect 20812 12248 20864 12257
rect 20904 12180 20956 12232
rect 21364 12316 21416 12368
rect 21640 12291 21692 12300
rect 21640 12257 21649 12291
rect 21649 12257 21683 12291
rect 21683 12257 21692 12291
rect 21640 12248 21692 12257
rect 22836 12291 22888 12300
rect 22836 12257 22845 12291
rect 22845 12257 22879 12291
rect 22879 12257 22888 12291
rect 22836 12248 22888 12257
rect 22652 12180 22704 12232
rect 19340 12112 19392 12164
rect 19616 12112 19668 12164
rect 11336 12044 11388 12096
rect 13912 12087 13964 12096
rect 13912 12053 13921 12087
rect 13921 12053 13955 12087
rect 13955 12053 13964 12087
rect 13912 12044 13964 12053
rect 19708 12044 19760 12096
rect 20628 12087 20680 12096
rect 20628 12053 20637 12087
rect 20637 12053 20671 12087
rect 20671 12053 20680 12087
rect 20628 12044 20680 12053
rect 20720 12044 20772 12096
rect 21456 12087 21508 12096
rect 21456 12053 21465 12087
rect 21465 12053 21499 12087
rect 21499 12053 21508 12087
rect 21456 12044 21508 12053
rect 22284 12087 22336 12096
rect 22284 12053 22293 12087
rect 22293 12053 22327 12087
rect 22327 12053 22336 12087
rect 22284 12044 22336 12053
rect 23480 12044 23532 12096
rect 6548 11942 6600 11994
rect 6612 11942 6664 11994
rect 6676 11942 6728 11994
rect 6740 11942 6792 11994
rect 6804 11942 6856 11994
rect 12146 11942 12198 11994
rect 12210 11942 12262 11994
rect 12274 11942 12326 11994
rect 12338 11942 12390 11994
rect 12402 11942 12454 11994
rect 17744 11942 17796 11994
rect 17808 11942 17860 11994
rect 17872 11942 17924 11994
rect 17936 11942 17988 11994
rect 18000 11942 18052 11994
rect 2596 11883 2648 11892
rect 2596 11849 2605 11883
rect 2605 11849 2639 11883
rect 2639 11849 2648 11883
rect 2596 11840 2648 11849
rect 3056 11840 3108 11892
rect 6368 11883 6420 11892
rect 6368 11849 6377 11883
rect 6377 11849 6411 11883
rect 6411 11849 6420 11883
rect 6368 11840 6420 11849
rect 4068 11772 4120 11824
rect 2780 11747 2832 11756
rect 2780 11713 2789 11747
rect 2789 11713 2823 11747
rect 2823 11713 2832 11747
rect 2780 11704 2832 11713
rect 3332 11704 3384 11756
rect 4712 11704 4764 11756
rect 5908 11747 5960 11756
rect 5908 11713 5926 11747
rect 5926 11713 5960 11747
rect 5908 11704 5960 11713
rect 3424 11636 3476 11688
rect 4804 11636 4856 11688
rect 11520 11840 11572 11892
rect 12440 11840 12492 11892
rect 12716 11840 12768 11892
rect 18880 11840 18932 11892
rect 20444 11883 20496 11892
rect 20444 11849 20453 11883
rect 20453 11849 20487 11883
rect 20487 11849 20496 11883
rect 20444 11840 20496 11849
rect 21456 11840 21508 11892
rect 7840 11704 7892 11756
rect 9036 11704 9088 11756
rect 9312 11704 9364 11756
rect 6828 11636 6880 11688
rect 11612 11772 11664 11824
rect 10784 11704 10836 11756
rect 12624 11704 12676 11756
rect 15752 11747 15804 11756
rect 15752 11713 15770 11747
rect 15770 11713 15804 11747
rect 15752 11704 15804 11713
rect 18236 11747 18288 11756
rect 20628 11772 20680 11824
rect 21916 11772 21968 11824
rect 18236 11713 18254 11747
rect 18254 11713 18288 11747
rect 18236 11704 18288 11713
rect 19616 11704 19668 11756
rect 19708 11704 19760 11756
rect 22468 11772 22520 11824
rect 22192 11704 22244 11756
rect 22928 11704 22980 11756
rect 23204 11704 23256 11756
rect 10508 11636 10560 11688
rect 18512 11679 18564 11688
rect 18512 11645 18521 11679
rect 18521 11645 18555 11679
rect 18555 11645 18564 11679
rect 18512 11636 18564 11645
rect 16396 11568 16448 11620
rect 5816 11500 5868 11552
rect 10416 11500 10468 11552
rect 10784 11500 10836 11552
rect 13084 11543 13136 11552
rect 13084 11509 13093 11543
rect 13093 11509 13127 11543
rect 13127 11509 13136 11543
rect 13084 11500 13136 11509
rect 15292 11500 15344 11552
rect 16120 11543 16172 11552
rect 16120 11509 16129 11543
rect 16129 11509 16163 11543
rect 16163 11509 16172 11543
rect 16120 11500 16172 11509
rect 16488 11543 16540 11552
rect 16488 11509 16497 11543
rect 16497 11509 16531 11543
rect 16531 11509 16540 11543
rect 16488 11500 16540 11509
rect 17132 11543 17184 11552
rect 17132 11509 17141 11543
rect 17141 11509 17175 11543
rect 17175 11509 17184 11543
rect 17132 11500 17184 11509
rect 20812 11636 20864 11688
rect 22376 11679 22428 11688
rect 22376 11645 22385 11679
rect 22385 11645 22419 11679
rect 22419 11645 22428 11679
rect 22376 11636 22428 11645
rect 21364 11611 21416 11620
rect 21364 11577 21373 11611
rect 21373 11577 21407 11611
rect 21407 11577 21416 11611
rect 21364 11568 21416 11577
rect 22468 11568 22520 11620
rect 18328 11500 18380 11552
rect 18880 11500 18932 11552
rect 20996 11500 21048 11552
rect 21272 11543 21324 11552
rect 21272 11509 21281 11543
rect 21281 11509 21315 11543
rect 21315 11509 21324 11543
rect 21272 11500 21324 11509
rect 21824 11543 21876 11552
rect 21824 11509 21833 11543
rect 21833 11509 21867 11543
rect 21867 11509 21876 11543
rect 21824 11500 21876 11509
rect 22652 11543 22704 11552
rect 22652 11509 22661 11543
rect 22661 11509 22695 11543
rect 22695 11509 22704 11543
rect 22652 11500 22704 11509
rect 3749 11398 3801 11450
rect 3813 11398 3865 11450
rect 3877 11398 3929 11450
rect 3941 11398 3993 11450
rect 4005 11398 4057 11450
rect 9347 11398 9399 11450
rect 9411 11398 9463 11450
rect 9475 11398 9527 11450
rect 9539 11398 9591 11450
rect 9603 11398 9655 11450
rect 14945 11398 14997 11450
rect 15009 11398 15061 11450
rect 15073 11398 15125 11450
rect 15137 11398 15189 11450
rect 15201 11398 15253 11450
rect 20543 11398 20595 11450
rect 20607 11398 20659 11450
rect 20671 11398 20723 11450
rect 20735 11398 20787 11450
rect 20799 11398 20851 11450
rect 3516 11296 3568 11348
rect 4252 11339 4304 11348
rect 4252 11305 4261 11339
rect 4261 11305 4295 11339
rect 4295 11305 4304 11339
rect 4252 11296 4304 11305
rect 5264 11339 5316 11348
rect 5264 11305 5273 11339
rect 5273 11305 5307 11339
rect 5307 11305 5316 11339
rect 5264 11296 5316 11305
rect 9036 11339 9088 11348
rect 9036 11305 9045 11339
rect 9045 11305 9079 11339
rect 9079 11305 9088 11339
rect 9036 11296 9088 11305
rect 10048 11296 10100 11348
rect 12532 11296 12584 11348
rect 16396 11296 16448 11348
rect 16488 11296 16540 11348
rect 3424 11228 3476 11280
rect 4988 11228 5040 11280
rect 4804 11203 4856 11212
rect 4804 11169 4813 11203
rect 4813 11169 4847 11203
rect 4847 11169 4856 11203
rect 4804 11160 4856 11169
rect 18512 11228 18564 11280
rect 19432 11296 19484 11348
rect 22744 11296 22796 11348
rect 20352 11228 20404 11280
rect 3608 11092 3660 11144
rect 5908 11092 5960 11144
rect 6828 11092 6880 11144
rect 3148 10999 3200 11008
rect 3148 10965 3157 10999
rect 3157 10965 3191 10999
rect 3191 10965 3200 10999
rect 3148 10956 3200 10965
rect 5540 11024 5592 11076
rect 8024 11024 8076 11076
rect 9956 11024 10008 11076
rect 13084 11092 13136 11144
rect 15016 11135 15068 11144
rect 15016 11101 15025 11135
rect 15025 11101 15059 11135
rect 15059 11101 15068 11135
rect 15016 11092 15068 11101
rect 16120 11092 16172 11144
rect 12440 11024 12492 11076
rect 12624 11024 12676 11076
rect 18696 11092 18748 11144
rect 19340 11092 19392 11144
rect 20904 11228 20956 11280
rect 22928 11271 22980 11280
rect 22928 11237 22937 11271
rect 22937 11237 22971 11271
rect 22971 11237 22980 11271
rect 22928 11228 22980 11237
rect 22376 11203 22428 11212
rect 22376 11169 22385 11203
rect 22385 11169 22419 11203
rect 22419 11169 22428 11203
rect 22376 11160 22428 11169
rect 21272 11092 21324 11144
rect 8392 10956 8444 11008
rect 10508 10999 10560 11008
rect 10508 10965 10517 10999
rect 10517 10965 10551 10999
rect 10551 10965 10560 10999
rect 10508 10956 10560 10965
rect 16396 10999 16448 11008
rect 16396 10965 16405 10999
rect 16405 10965 16439 10999
rect 16439 10965 16448 10999
rect 16396 10956 16448 10965
rect 17040 10956 17092 11008
rect 21088 11024 21140 11076
rect 21456 11024 21508 11076
rect 22284 11024 22336 11076
rect 18880 10956 18932 11008
rect 6548 10854 6600 10906
rect 6612 10854 6664 10906
rect 6676 10854 6728 10906
rect 6740 10854 6792 10906
rect 6804 10854 6856 10906
rect 12146 10854 12198 10906
rect 12210 10854 12262 10906
rect 12274 10854 12326 10906
rect 12338 10854 12390 10906
rect 12402 10854 12454 10906
rect 17744 10854 17796 10906
rect 17808 10854 17860 10906
rect 17872 10854 17924 10906
rect 17936 10854 17988 10906
rect 18000 10854 18052 10906
rect 2872 10752 2924 10804
rect 3148 10752 3200 10804
rect 5540 10752 5592 10804
rect 6184 10795 6236 10804
rect 6184 10761 6193 10795
rect 6193 10761 6227 10795
rect 6227 10761 6236 10795
rect 6184 10752 6236 10761
rect 6368 10752 6420 10804
rect 13544 10795 13596 10804
rect 13544 10761 13553 10795
rect 13553 10761 13587 10795
rect 13587 10761 13596 10795
rect 13544 10752 13596 10761
rect 6460 10684 6512 10736
rect 8484 10684 8536 10736
rect 11152 10684 11204 10736
rect 12532 10684 12584 10736
rect 2780 10616 2832 10668
rect 5448 10616 5500 10668
rect 8852 10616 8904 10668
rect 4528 10591 4580 10600
rect 4528 10557 4537 10591
rect 4537 10557 4571 10591
rect 4571 10557 4580 10591
rect 4528 10548 4580 10557
rect 4712 10548 4764 10600
rect 8392 10591 8444 10600
rect 8392 10557 8401 10591
rect 8401 10557 8435 10591
rect 8435 10557 8444 10591
rect 8392 10548 8444 10557
rect 10508 10616 10560 10668
rect 15016 10659 15068 10668
rect 15016 10625 15025 10659
rect 15025 10625 15059 10659
rect 15059 10625 15068 10659
rect 15016 10616 15068 10625
rect 6460 10412 6512 10464
rect 8024 10412 8076 10464
rect 9956 10455 10008 10464
rect 9956 10421 9965 10455
rect 9965 10421 9999 10455
rect 9999 10421 10008 10455
rect 9956 10412 10008 10421
rect 11520 10455 11572 10464
rect 11520 10421 11529 10455
rect 11529 10421 11563 10455
rect 11563 10421 11572 10455
rect 11520 10412 11572 10421
rect 13636 10455 13688 10464
rect 13636 10421 13645 10455
rect 13645 10421 13679 10455
rect 13679 10421 13688 10455
rect 13636 10412 13688 10421
rect 16120 10684 16172 10736
rect 17040 10684 17092 10736
rect 22100 10752 22152 10804
rect 22468 10795 22520 10804
rect 22468 10761 22477 10795
rect 22477 10761 22511 10795
rect 22511 10761 22520 10795
rect 22468 10752 22520 10761
rect 22652 10752 22704 10804
rect 16764 10616 16816 10668
rect 18328 10659 18380 10668
rect 18328 10625 18337 10659
rect 18337 10625 18371 10659
rect 18371 10625 18380 10659
rect 18328 10616 18380 10625
rect 18788 10591 18840 10600
rect 16580 10412 16632 10464
rect 18788 10557 18797 10591
rect 18797 10557 18831 10591
rect 18831 10557 18840 10591
rect 18788 10548 18840 10557
rect 18880 10591 18932 10600
rect 18880 10557 18889 10591
rect 18889 10557 18923 10591
rect 18923 10557 18932 10591
rect 18880 10548 18932 10557
rect 19892 10480 19944 10532
rect 22284 10684 22336 10736
rect 21824 10659 21876 10668
rect 21824 10625 21833 10659
rect 21833 10625 21867 10659
rect 21867 10625 21876 10659
rect 21824 10616 21876 10625
rect 23296 10616 23348 10668
rect 21364 10591 21416 10600
rect 21364 10557 21373 10591
rect 21373 10557 21407 10591
rect 21407 10557 21416 10591
rect 21364 10548 21416 10557
rect 21456 10591 21508 10600
rect 21456 10557 21465 10591
rect 21465 10557 21499 10591
rect 21499 10557 21508 10591
rect 21456 10548 21508 10557
rect 22192 10548 22244 10600
rect 21824 10480 21876 10532
rect 17408 10412 17460 10464
rect 19248 10412 19300 10464
rect 20260 10455 20312 10464
rect 20260 10421 20269 10455
rect 20269 10421 20303 10455
rect 20303 10421 20312 10455
rect 20260 10412 20312 10421
rect 21180 10412 21232 10464
rect 22008 10455 22060 10464
rect 22008 10421 22017 10455
rect 22017 10421 22051 10455
rect 22051 10421 22060 10455
rect 22008 10412 22060 10421
rect 22100 10455 22152 10464
rect 22100 10421 22109 10455
rect 22109 10421 22143 10455
rect 22143 10421 22152 10455
rect 22100 10412 22152 10421
rect 22376 10412 22428 10464
rect 3749 10310 3801 10362
rect 3813 10310 3865 10362
rect 3877 10310 3929 10362
rect 3941 10310 3993 10362
rect 4005 10310 4057 10362
rect 9347 10310 9399 10362
rect 9411 10310 9463 10362
rect 9475 10310 9527 10362
rect 9539 10310 9591 10362
rect 9603 10310 9655 10362
rect 14945 10310 14997 10362
rect 15009 10310 15061 10362
rect 15073 10310 15125 10362
rect 15137 10310 15189 10362
rect 15201 10310 15253 10362
rect 20543 10310 20595 10362
rect 20607 10310 20659 10362
rect 20671 10310 20723 10362
rect 20735 10310 20787 10362
rect 20799 10310 20851 10362
rect 2504 10251 2556 10260
rect 2504 10217 2513 10251
rect 2513 10217 2547 10251
rect 2547 10217 2556 10251
rect 2504 10208 2556 10217
rect 2964 10208 3016 10260
rect 6368 10208 6420 10260
rect 2320 10047 2372 10056
rect 2320 10013 2329 10047
rect 2329 10013 2363 10047
rect 2363 10013 2372 10047
rect 2320 10004 2372 10013
rect 4712 10140 4764 10192
rect 3056 10072 3108 10124
rect 3424 10115 3476 10124
rect 3424 10081 3433 10115
rect 3433 10081 3467 10115
rect 3467 10081 3476 10115
rect 3424 10072 3476 10081
rect 4528 10072 4580 10124
rect 8852 10208 8904 10260
rect 18880 10208 18932 10260
rect 17040 10183 17092 10192
rect 17040 10149 17049 10183
rect 17049 10149 17083 10183
rect 17083 10149 17092 10183
rect 17040 10140 17092 10149
rect 19616 10140 19668 10192
rect 4712 10004 4764 10056
rect 4896 10004 4948 10056
rect 2872 9868 2924 9920
rect 4712 9911 4764 9920
rect 4712 9877 4721 9911
rect 4721 9877 4755 9911
rect 4755 9877 4764 9911
rect 4712 9868 4764 9877
rect 5816 9936 5868 9988
rect 7104 9979 7156 9988
rect 7104 9945 7138 9979
rect 7138 9945 7156 9979
rect 7104 9936 7156 9945
rect 6552 9868 6604 9920
rect 11520 10047 11572 10056
rect 11520 10013 11529 10047
rect 11529 10013 11563 10047
rect 11563 10013 11572 10047
rect 11520 10004 11572 10013
rect 12900 10004 12952 10056
rect 17592 10004 17644 10056
rect 18236 10072 18288 10124
rect 8392 9911 8444 9920
rect 8392 9877 8401 9911
rect 8401 9877 8435 9911
rect 8435 9877 8444 9911
rect 10232 9936 10284 9988
rect 16396 9936 16448 9988
rect 18144 9936 18196 9988
rect 8392 9868 8444 9877
rect 8576 9868 8628 9920
rect 11336 9868 11388 9920
rect 12992 9911 13044 9920
rect 12992 9877 13001 9911
rect 13001 9877 13035 9911
rect 13035 9877 13044 9911
rect 12992 9868 13044 9877
rect 14188 9911 14240 9920
rect 14188 9877 14197 9911
rect 14197 9877 14231 9911
rect 14231 9877 14240 9911
rect 14188 9868 14240 9877
rect 17316 9868 17368 9920
rect 18052 9868 18104 9920
rect 18972 10072 19024 10124
rect 20812 10208 20864 10260
rect 21916 10208 21968 10260
rect 21732 10140 21784 10192
rect 21272 10115 21324 10124
rect 21272 10081 21281 10115
rect 21281 10081 21315 10115
rect 21315 10081 21324 10115
rect 21272 10072 21324 10081
rect 21548 10072 21600 10124
rect 22192 10115 22244 10124
rect 22192 10081 22201 10115
rect 22201 10081 22235 10115
rect 22235 10081 22244 10115
rect 22192 10072 22244 10081
rect 22376 10115 22428 10124
rect 22376 10081 22385 10115
rect 22385 10081 22419 10115
rect 22419 10081 22428 10115
rect 22376 10072 22428 10081
rect 19156 10004 19208 10056
rect 21088 10004 21140 10056
rect 22008 10004 22060 10056
rect 18604 9868 18656 9920
rect 18696 9868 18748 9920
rect 20076 9868 20128 9920
rect 20996 9936 21048 9988
rect 21640 9936 21692 9988
rect 20720 9911 20772 9920
rect 20720 9877 20729 9911
rect 20729 9877 20763 9911
rect 20763 9877 20772 9911
rect 20720 9868 20772 9877
rect 20812 9868 20864 9920
rect 21456 9868 21508 9920
rect 22836 9911 22888 9920
rect 22836 9877 22845 9911
rect 22845 9877 22879 9911
rect 22879 9877 22888 9911
rect 22836 9868 22888 9877
rect 22928 9911 22980 9920
rect 22928 9877 22937 9911
rect 22937 9877 22971 9911
rect 22971 9877 22980 9911
rect 22928 9868 22980 9877
rect 6548 9766 6600 9818
rect 6612 9766 6664 9818
rect 6676 9766 6728 9818
rect 6740 9766 6792 9818
rect 6804 9766 6856 9818
rect 12146 9766 12198 9818
rect 12210 9766 12262 9818
rect 12274 9766 12326 9818
rect 12338 9766 12390 9818
rect 12402 9766 12454 9818
rect 17744 9766 17796 9818
rect 17808 9766 17860 9818
rect 17872 9766 17924 9818
rect 17936 9766 17988 9818
rect 18000 9766 18052 9818
rect 4528 9664 4580 9716
rect 6368 9707 6420 9716
rect 1400 9571 1452 9580
rect 1400 9537 1409 9571
rect 1409 9537 1443 9571
rect 1443 9537 1452 9571
rect 1400 9528 1452 9537
rect 6368 9673 6377 9707
rect 6377 9673 6411 9707
rect 6411 9673 6420 9707
rect 6644 9707 6696 9716
rect 6368 9664 6420 9673
rect 6644 9673 6653 9707
rect 6653 9673 6687 9707
rect 6687 9673 6696 9707
rect 6644 9664 6696 9673
rect 3148 9528 3200 9580
rect 3884 9528 3936 9580
rect 3240 9460 3292 9512
rect 3148 9392 3200 9444
rect 2412 9324 2464 9376
rect 4436 9324 4488 9376
rect 6644 9528 6696 9580
rect 8852 9528 8904 9580
rect 10140 9528 10192 9580
rect 11244 9664 11296 9716
rect 12624 9664 12676 9716
rect 13636 9664 13688 9716
rect 6920 9503 6972 9512
rect 6920 9469 6929 9503
rect 6929 9469 6963 9503
rect 6963 9469 6972 9503
rect 6920 9460 6972 9469
rect 9036 9503 9088 9512
rect 9036 9469 9045 9503
rect 9045 9469 9079 9503
rect 9079 9469 9088 9503
rect 9036 9460 9088 9469
rect 7104 9324 7156 9376
rect 7472 9367 7524 9376
rect 7472 9333 7481 9367
rect 7481 9333 7515 9367
rect 7515 9333 7524 9367
rect 7472 9324 7524 9333
rect 9220 9324 9272 9376
rect 10232 9324 10284 9376
rect 10692 9367 10744 9376
rect 10692 9333 10701 9367
rect 10701 9333 10735 9367
rect 10735 9333 10744 9367
rect 10692 9324 10744 9333
rect 10784 9324 10836 9376
rect 12808 9596 12860 9648
rect 17500 9664 17552 9716
rect 18052 9664 18104 9716
rect 18696 9664 18748 9716
rect 20996 9664 21048 9716
rect 21364 9707 21416 9716
rect 21364 9673 21373 9707
rect 21373 9673 21407 9707
rect 21407 9673 21416 9707
rect 21364 9664 21416 9673
rect 22192 9664 22244 9716
rect 22836 9664 22888 9716
rect 12624 9571 12676 9580
rect 12624 9537 12642 9571
rect 12642 9537 12676 9571
rect 12900 9571 12952 9580
rect 12624 9528 12676 9537
rect 12900 9537 12909 9571
rect 12909 9537 12943 9571
rect 12943 9537 12952 9571
rect 12900 9528 12952 9537
rect 12992 9528 13044 9580
rect 15384 9571 15436 9580
rect 15384 9537 15418 9571
rect 15418 9537 15436 9571
rect 15384 9528 15436 9537
rect 18236 9528 18288 9580
rect 18512 9571 18564 9580
rect 18512 9537 18530 9571
rect 18530 9537 18564 9571
rect 18512 9528 18564 9537
rect 18972 9528 19024 9580
rect 19432 9528 19484 9580
rect 18788 9503 18840 9512
rect 18788 9469 18797 9503
rect 18797 9469 18831 9503
rect 18831 9469 18840 9503
rect 18788 9460 18840 9469
rect 16304 9392 16356 9444
rect 20720 9528 20772 9580
rect 21732 9460 21784 9512
rect 22100 9528 22152 9580
rect 12624 9324 12676 9376
rect 12716 9324 12768 9376
rect 16580 9324 16632 9376
rect 17408 9367 17460 9376
rect 17408 9333 17417 9367
rect 17417 9333 17451 9367
rect 17451 9333 17460 9367
rect 17408 9324 17460 9333
rect 20076 9324 20128 9376
rect 20168 9324 20220 9376
rect 20444 9367 20496 9376
rect 20444 9333 20453 9367
rect 20453 9333 20487 9367
rect 20487 9333 20496 9367
rect 20444 9324 20496 9333
rect 21272 9367 21324 9376
rect 21272 9333 21281 9367
rect 21281 9333 21315 9367
rect 21315 9333 21324 9367
rect 21272 9324 21324 9333
rect 23020 9528 23072 9580
rect 22928 9460 22980 9512
rect 23204 9392 23256 9444
rect 22192 9324 22244 9376
rect 22284 9324 22336 9376
rect 3749 9222 3801 9274
rect 3813 9222 3865 9274
rect 3877 9222 3929 9274
rect 3941 9222 3993 9274
rect 4005 9222 4057 9274
rect 9347 9222 9399 9274
rect 9411 9222 9463 9274
rect 9475 9222 9527 9274
rect 9539 9222 9591 9274
rect 9603 9222 9655 9274
rect 14945 9222 14997 9274
rect 15009 9222 15061 9274
rect 15073 9222 15125 9274
rect 15137 9222 15189 9274
rect 15201 9222 15253 9274
rect 20543 9222 20595 9274
rect 20607 9222 20659 9274
rect 20671 9222 20723 9274
rect 20735 9222 20787 9274
rect 20799 9222 20851 9274
rect 2780 9163 2832 9172
rect 2780 9129 2789 9163
rect 2789 9129 2823 9163
rect 2823 9129 2832 9163
rect 2780 9120 2832 9129
rect 2872 9095 2924 9104
rect 2872 9061 2881 9095
rect 2881 9061 2915 9095
rect 2915 9061 2924 9095
rect 2872 9052 2924 9061
rect 3148 9052 3200 9104
rect 3516 9052 3568 9104
rect 3056 8984 3108 9036
rect 3240 8984 3292 9036
rect 4712 9120 4764 9172
rect 5448 9163 5500 9172
rect 5448 9129 5457 9163
rect 5457 9129 5491 9163
rect 5491 9129 5500 9163
rect 5448 9120 5500 9129
rect 6644 9120 6696 9172
rect 8392 9120 8444 9172
rect 9036 9163 9088 9172
rect 9036 9129 9045 9163
rect 9045 9129 9079 9163
rect 9079 9129 9088 9163
rect 9036 9120 9088 9129
rect 12900 9120 12952 9172
rect 17592 9120 17644 9172
rect 18328 9120 18380 9172
rect 19248 9120 19300 9172
rect 21456 9163 21508 9172
rect 18880 9052 18932 9104
rect 18972 9052 19024 9104
rect 21456 9129 21465 9163
rect 21465 9129 21499 9163
rect 21499 9129 21508 9163
rect 21456 9120 21508 9129
rect 21640 9120 21692 9172
rect 23572 9120 23624 9172
rect 23848 9120 23900 9172
rect 22192 9052 22244 9104
rect 23664 9052 23716 9104
rect 18788 8984 18840 9036
rect 19156 8984 19208 9036
rect 20996 8984 21048 9036
rect 2412 8959 2464 8968
rect 2412 8925 2421 8959
rect 2421 8925 2455 8959
rect 2455 8925 2464 8959
rect 2412 8916 2464 8925
rect 7472 8916 7524 8968
rect 9772 8916 9824 8968
rect 16304 8959 16356 8968
rect 16304 8925 16313 8959
rect 16313 8925 16347 8959
rect 16347 8925 16356 8959
rect 16304 8916 16356 8925
rect 16396 8916 16448 8968
rect 2872 8848 2924 8900
rect 4344 8891 4396 8900
rect 4344 8857 4378 8891
rect 4378 8857 4396 8891
rect 4344 8848 4396 8857
rect 4436 8848 4488 8900
rect 6460 8848 6512 8900
rect 12716 8848 12768 8900
rect 15936 8848 15988 8900
rect 17500 8891 17552 8900
rect 5540 8823 5592 8832
rect 5540 8789 5549 8823
rect 5549 8789 5583 8823
rect 5583 8789 5592 8823
rect 5540 8780 5592 8789
rect 8852 8780 8904 8832
rect 11152 8780 11204 8832
rect 11520 8823 11572 8832
rect 11520 8789 11529 8823
rect 11529 8789 11563 8823
rect 11563 8789 11572 8823
rect 11520 8780 11572 8789
rect 12624 8780 12676 8832
rect 15384 8780 15436 8832
rect 16396 8823 16448 8832
rect 16396 8789 16405 8823
rect 16405 8789 16439 8823
rect 16439 8789 16448 8823
rect 16396 8780 16448 8789
rect 17500 8857 17518 8891
rect 17518 8857 17552 8891
rect 17500 8848 17552 8857
rect 18236 8916 18288 8968
rect 18604 8916 18656 8968
rect 19340 8916 19392 8968
rect 19616 8916 19668 8968
rect 20536 8916 20588 8968
rect 21088 8959 21140 8968
rect 21088 8925 21097 8959
rect 21097 8925 21131 8959
rect 21131 8925 21140 8959
rect 21088 8916 21140 8925
rect 18788 8780 18840 8832
rect 19984 8780 20036 8832
rect 20352 8891 20404 8900
rect 20352 8857 20370 8891
rect 20370 8857 20404 8891
rect 21824 8984 21876 9036
rect 21456 8916 21508 8968
rect 22744 8959 22796 8968
rect 22744 8925 22753 8959
rect 22753 8925 22787 8959
rect 22787 8925 22796 8959
rect 22744 8916 22796 8925
rect 20352 8848 20404 8857
rect 22192 8848 22244 8900
rect 21640 8780 21692 8832
rect 6548 8678 6600 8730
rect 6612 8678 6664 8730
rect 6676 8678 6728 8730
rect 6740 8678 6792 8730
rect 6804 8678 6856 8730
rect 12146 8678 12198 8730
rect 12210 8678 12262 8730
rect 12274 8678 12326 8730
rect 12338 8678 12390 8730
rect 12402 8678 12454 8730
rect 17744 8678 17796 8730
rect 17808 8678 17860 8730
rect 17872 8678 17924 8730
rect 17936 8678 17988 8730
rect 18000 8678 18052 8730
rect 3332 8619 3384 8628
rect 3332 8585 3341 8619
rect 3341 8585 3375 8619
rect 3375 8585 3384 8619
rect 3332 8576 3384 8585
rect 6184 8619 6236 8628
rect 2964 8551 3016 8560
rect 2964 8517 2973 8551
rect 2973 8517 3007 8551
rect 3007 8517 3016 8551
rect 2964 8508 3016 8517
rect 2044 8483 2096 8492
rect 2044 8449 2053 8483
rect 2053 8449 2087 8483
rect 2087 8449 2096 8483
rect 2044 8440 2096 8449
rect 6184 8585 6193 8619
rect 6193 8585 6227 8619
rect 6227 8585 6236 8619
rect 6184 8576 6236 8585
rect 15752 8576 15804 8628
rect 16212 8576 16264 8628
rect 18236 8576 18288 8628
rect 4804 8508 4856 8560
rect 8300 8508 8352 8560
rect 8576 8508 8628 8560
rect 11520 8551 11572 8560
rect 4896 8440 4948 8492
rect 5816 8440 5868 8492
rect 3056 8372 3108 8424
rect 3240 8372 3292 8424
rect 2320 8304 2372 8356
rect 4436 8236 4488 8288
rect 6000 8304 6052 8356
rect 9128 8440 9180 8492
rect 11520 8517 11529 8551
rect 11529 8517 11563 8551
rect 11563 8517 11572 8551
rect 11520 8508 11572 8517
rect 10692 8440 10744 8492
rect 12532 8440 12584 8492
rect 18144 8508 18196 8560
rect 19524 8551 19576 8560
rect 19524 8517 19558 8551
rect 19558 8517 19576 8551
rect 19524 8508 19576 8517
rect 20536 8576 20588 8628
rect 21732 8576 21784 8628
rect 22468 8508 22520 8560
rect 16488 8440 16540 8492
rect 16580 8440 16632 8492
rect 18328 8440 18380 8492
rect 19064 8440 19116 8492
rect 20444 8440 20496 8492
rect 20904 8440 20956 8492
rect 21088 8483 21140 8492
rect 21088 8449 21097 8483
rect 21097 8449 21131 8483
rect 21131 8449 21140 8483
rect 21088 8440 21140 8449
rect 21180 8483 21232 8492
rect 21180 8449 21189 8483
rect 21189 8449 21223 8483
rect 21223 8449 21232 8483
rect 21180 8440 21232 8449
rect 21732 8440 21784 8492
rect 22652 8483 22704 8492
rect 8392 8415 8444 8424
rect 8392 8381 8401 8415
rect 8401 8381 8435 8415
rect 8435 8381 8444 8415
rect 8392 8372 8444 8381
rect 12072 8304 12124 8356
rect 19156 8415 19208 8424
rect 19156 8381 19165 8415
rect 19165 8381 19199 8415
rect 19199 8381 19208 8415
rect 19156 8372 19208 8381
rect 16028 8347 16080 8356
rect 16028 8313 16037 8347
rect 16037 8313 16071 8347
rect 16071 8313 16080 8347
rect 16304 8347 16356 8356
rect 16028 8304 16080 8313
rect 16304 8313 16313 8347
rect 16313 8313 16347 8347
rect 16347 8313 16356 8347
rect 16304 8304 16356 8313
rect 7012 8279 7064 8288
rect 7012 8245 7021 8279
rect 7021 8245 7055 8279
rect 7055 8245 7064 8279
rect 7012 8236 7064 8245
rect 8668 8236 8720 8288
rect 11520 8236 11572 8288
rect 11888 8236 11940 8288
rect 16396 8236 16448 8288
rect 17592 8236 17644 8288
rect 20812 8372 20864 8424
rect 22652 8449 22661 8483
rect 22661 8449 22695 8483
rect 22695 8449 22704 8483
rect 22652 8440 22704 8449
rect 22560 8372 22612 8424
rect 20996 8304 21048 8356
rect 22468 8304 22520 8356
rect 19616 8236 19668 8288
rect 20444 8236 20496 8288
rect 20812 8236 20864 8288
rect 22560 8236 22612 8288
rect 3749 8134 3801 8186
rect 3813 8134 3865 8186
rect 3877 8134 3929 8186
rect 3941 8134 3993 8186
rect 4005 8134 4057 8186
rect 9347 8134 9399 8186
rect 9411 8134 9463 8186
rect 9475 8134 9527 8186
rect 9539 8134 9591 8186
rect 9603 8134 9655 8186
rect 14945 8134 14997 8186
rect 15009 8134 15061 8186
rect 15073 8134 15125 8186
rect 15137 8134 15189 8186
rect 15201 8134 15253 8186
rect 20543 8134 20595 8186
rect 20607 8134 20659 8186
rect 20671 8134 20723 8186
rect 20735 8134 20787 8186
rect 20799 8134 20851 8186
rect 2044 8075 2096 8084
rect 2044 8041 2053 8075
rect 2053 8041 2087 8075
rect 2087 8041 2096 8075
rect 2044 8032 2096 8041
rect 2872 8075 2924 8084
rect 2872 8041 2881 8075
rect 2881 8041 2915 8075
rect 2915 8041 2924 8075
rect 2872 8032 2924 8041
rect 5816 8075 5868 8084
rect 5816 8041 5825 8075
rect 5825 8041 5859 8075
rect 5859 8041 5868 8075
rect 5816 8032 5868 8041
rect 6920 8032 6972 8084
rect 7472 8032 7524 8084
rect 11244 8032 11296 8084
rect 3240 7896 3292 7948
rect 3148 7828 3200 7880
rect 3332 7828 3384 7880
rect 4436 7871 4488 7880
rect 4436 7837 4445 7871
rect 4445 7837 4479 7871
rect 4479 7837 4488 7871
rect 4436 7828 4488 7837
rect 6000 7828 6052 7880
rect 10692 7828 10744 7880
rect 16304 7828 16356 7880
rect 22836 8032 22888 8084
rect 22192 7964 22244 8016
rect 23296 7964 23348 8016
rect 21272 7896 21324 7948
rect 21916 7896 21968 7948
rect 18420 7828 18472 7880
rect 19892 7828 19944 7880
rect 20628 7871 20680 7880
rect 20628 7837 20637 7871
rect 20637 7837 20671 7871
rect 20671 7837 20680 7871
rect 20628 7828 20680 7837
rect 21548 7828 21600 7880
rect 21824 7828 21876 7880
rect 23020 7871 23072 7880
rect 23020 7837 23029 7871
rect 23029 7837 23063 7871
rect 23063 7837 23072 7871
rect 23020 7828 23072 7837
rect 3424 7760 3476 7812
rect 3516 7760 3568 7812
rect 7196 7760 7248 7812
rect 2412 7735 2464 7744
rect 2412 7701 2421 7735
rect 2421 7701 2455 7735
rect 2455 7701 2464 7735
rect 2412 7692 2464 7701
rect 4804 7692 4856 7744
rect 7564 7760 7616 7812
rect 8392 7760 8444 7812
rect 11060 7692 11112 7744
rect 11520 7760 11572 7812
rect 11612 7760 11664 7812
rect 13360 7760 13412 7812
rect 11888 7692 11940 7744
rect 12532 7692 12584 7744
rect 13820 7735 13872 7744
rect 13820 7701 13829 7735
rect 13829 7701 13863 7735
rect 13863 7701 13872 7735
rect 13820 7692 13872 7701
rect 14740 7692 14792 7744
rect 16672 7692 16724 7744
rect 17408 7760 17460 7812
rect 20168 7760 20220 7812
rect 20260 7760 20312 7812
rect 19524 7692 19576 7744
rect 21180 7735 21232 7744
rect 21180 7701 21195 7735
rect 21195 7701 21229 7735
rect 21229 7701 21232 7735
rect 21180 7692 21232 7701
rect 22652 7735 22704 7744
rect 22652 7701 22661 7735
rect 22661 7701 22695 7735
rect 22695 7701 22704 7735
rect 22652 7692 22704 7701
rect 23572 7692 23624 7744
rect 6548 7590 6600 7642
rect 6612 7590 6664 7642
rect 6676 7590 6728 7642
rect 6740 7590 6792 7642
rect 6804 7590 6856 7642
rect 12146 7590 12198 7642
rect 12210 7590 12262 7642
rect 12274 7590 12326 7642
rect 12338 7590 12390 7642
rect 12402 7590 12454 7642
rect 17744 7590 17796 7642
rect 17808 7590 17860 7642
rect 17872 7590 17924 7642
rect 17936 7590 17988 7642
rect 18000 7590 18052 7642
rect 4344 7488 4396 7540
rect 9220 7488 9272 7540
rect 10048 7488 10100 7540
rect 10692 7531 10744 7540
rect 10692 7497 10701 7531
rect 10701 7497 10735 7531
rect 10735 7497 10744 7531
rect 10692 7488 10744 7497
rect 13360 7531 13412 7540
rect 3148 7420 3200 7472
rect 3332 7395 3384 7404
rect 3332 7361 3341 7395
rect 3341 7361 3375 7395
rect 3375 7361 3384 7395
rect 3332 7352 3384 7361
rect 5540 7420 5592 7472
rect 10416 7420 10468 7472
rect 11060 7420 11112 7472
rect 11612 7420 11664 7472
rect 5080 7352 5132 7404
rect 6092 7352 6144 7404
rect 6644 7352 6696 7404
rect 7012 7352 7064 7404
rect 7656 7352 7708 7404
rect 8392 7395 8444 7404
rect 8392 7361 8401 7395
rect 8401 7361 8435 7395
rect 8435 7361 8444 7395
rect 8392 7352 8444 7361
rect 8668 7395 8720 7404
rect 8668 7361 8702 7395
rect 8702 7361 8720 7395
rect 8668 7352 8720 7361
rect 13360 7497 13369 7531
rect 13369 7497 13403 7531
rect 13403 7497 13412 7531
rect 13360 7488 13412 7497
rect 16028 7531 16080 7540
rect 16028 7497 16037 7531
rect 16037 7497 16071 7531
rect 16071 7497 16080 7531
rect 16028 7488 16080 7497
rect 12072 7420 12124 7472
rect 13728 7352 13780 7404
rect 19524 7488 19576 7540
rect 21088 7531 21140 7540
rect 18696 7420 18748 7472
rect 19984 7420 20036 7472
rect 21088 7497 21097 7531
rect 21097 7497 21131 7531
rect 21131 7497 21140 7531
rect 21088 7488 21140 7497
rect 23020 7531 23072 7540
rect 23020 7497 23029 7531
rect 23029 7497 23063 7531
rect 23063 7497 23072 7531
rect 23020 7488 23072 7497
rect 14740 7395 14792 7404
rect 14740 7361 14774 7395
rect 14774 7361 14792 7395
rect 14740 7352 14792 7361
rect 16304 7395 16356 7404
rect 16304 7361 16313 7395
rect 16313 7361 16347 7395
rect 16347 7361 16356 7395
rect 16304 7352 16356 7361
rect 10416 7327 10468 7336
rect 10416 7293 10425 7327
rect 10425 7293 10459 7327
rect 10459 7293 10468 7327
rect 10416 7284 10468 7293
rect 16028 7284 16080 7336
rect 20444 7352 20496 7404
rect 21456 7420 21508 7472
rect 21548 7395 21600 7404
rect 19616 7327 19668 7336
rect 9772 7259 9824 7268
rect 2412 7148 2464 7200
rect 9772 7225 9781 7259
rect 9781 7225 9815 7259
rect 9815 7225 9824 7259
rect 9772 7216 9824 7225
rect 5908 7148 5960 7200
rect 8576 7148 8628 7200
rect 10048 7148 10100 7200
rect 13452 7148 13504 7200
rect 13544 7191 13596 7200
rect 13544 7157 13553 7191
rect 13553 7157 13587 7191
rect 13587 7157 13596 7191
rect 13544 7148 13596 7157
rect 13728 7148 13780 7200
rect 15844 7191 15896 7200
rect 15844 7157 15853 7191
rect 15853 7157 15887 7191
rect 15887 7157 15896 7191
rect 15844 7148 15896 7157
rect 19616 7293 19625 7327
rect 19625 7293 19659 7327
rect 19659 7293 19668 7327
rect 19616 7284 19668 7293
rect 21548 7361 21557 7395
rect 21557 7361 21591 7395
rect 21591 7361 21600 7395
rect 21548 7352 21600 7361
rect 22192 7395 22244 7404
rect 22192 7361 22201 7395
rect 22201 7361 22235 7395
rect 22235 7361 22244 7395
rect 22192 7352 22244 7361
rect 22928 7352 22980 7404
rect 22100 7327 22152 7336
rect 22100 7293 22109 7327
rect 22109 7293 22143 7327
rect 22143 7293 22152 7327
rect 22100 7284 22152 7293
rect 17960 7148 18012 7200
rect 18144 7148 18196 7200
rect 19432 7148 19484 7200
rect 21272 7216 21324 7268
rect 22560 7259 22612 7268
rect 22560 7225 22569 7259
rect 22569 7225 22603 7259
rect 22603 7225 22612 7259
rect 22560 7216 22612 7225
rect 20352 7148 20404 7200
rect 20628 7148 20680 7200
rect 21088 7148 21140 7200
rect 22652 7191 22704 7200
rect 22652 7157 22661 7191
rect 22661 7157 22695 7191
rect 22695 7157 22704 7191
rect 22652 7148 22704 7157
rect 3749 7046 3801 7098
rect 3813 7046 3865 7098
rect 3877 7046 3929 7098
rect 3941 7046 3993 7098
rect 4005 7046 4057 7098
rect 9347 7046 9399 7098
rect 9411 7046 9463 7098
rect 9475 7046 9527 7098
rect 9539 7046 9591 7098
rect 9603 7046 9655 7098
rect 14945 7046 14997 7098
rect 15009 7046 15061 7098
rect 15073 7046 15125 7098
rect 15137 7046 15189 7098
rect 15201 7046 15253 7098
rect 20543 7046 20595 7098
rect 20607 7046 20659 7098
rect 20671 7046 20723 7098
rect 20735 7046 20787 7098
rect 20799 7046 20851 7098
rect 3332 6944 3384 6996
rect 5080 6987 5132 6996
rect 5080 6953 5089 6987
rect 5089 6953 5123 6987
rect 5123 6953 5132 6987
rect 5080 6944 5132 6953
rect 6644 6987 6696 6996
rect 6644 6953 6653 6987
rect 6653 6953 6687 6987
rect 6687 6953 6696 6987
rect 6644 6944 6696 6953
rect 7196 6944 7248 6996
rect 8392 6944 8444 6996
rect 6460 6851 6512 6860
rect 6460 6817 6469 6851
rect 6469 6817 6503 6851
rect 6503 6817 6512 6851
rect 13452 6944 13504 6996
rect 22468 6944 22520 6996
rect 6460 6808 6512 6817
rect 6184 6783 6236 6792
rect 6184 6749 6202 6783
rect 6202 6749 6236 6783
rect 6184 6740 6236 6749
rect 2136 6672 2188 6724
rect 8208 6672 8260 6724
rect 8576 6672 8628 6724
rect 8760 6672 8812 6724
rect 10416 6808 10468 6860
rect 11244 6851 11296 6860
rect 11244 6817 11253 6851
rect 11253 6817 11287 6851
rect 11287 6817 11296 6851
rect 11244 6808 11296 6817
rect 12532 6808 12584 6860
rect 17960 6876 18012 6928
rect 18236 6876 18288 6928
rect 20812 6876 20864 6928
rect 21272 6876 21324 6928
rect 13360 6808 13412 6860
rect 13728 6851 13780 6860
rect 13728 6817 13737 6851
rect 13737 6817 13771 6851
rect 13771 6817 13780 6851
rect 13728 6808 13780 6817
rect 16028 6808 16080 6860
rect 9956 6740 10008 6792
rect 11152 6740 11204 6792
rect 12072 6740 12124 6792
rect 9312 6647 9364 6656
rect 9312 6613 9321 6647
rect 9321 6613 9355 6647
rect 9355 6613 9364 6647
rect 9312 6604 9364 6613
rect 9680 6604 9732 6656
rect 10232 6672 10284 6724
rect 11796 6672 11848 6724
rect 10140 6604 10192 6656
rect 10416 6647 10468 6656
rect 10416 6613 10425 6647
rect 10425 6613 10459 6647
rect 10459 6613 10468 6647
rect 10416 6604 10468 6613
rect 12072 6604 12124 6656
rect 13176 6647 13228 6656
rect 13176 6613 13185 6647
rect 13185 6613 13219 6647
rect 13219 6613 13228 6647
rect 13176 6604 13228 6613
rect 14740 6672 14792 6724
rect 15752 6672 15804 6724
rect 16396 6715 16448 6724
rect 16396 6681 16430 6715
rect 16430 6681 16448 6715
rect 16396 6672 16448 6681
rect 16488 6672 16540 6724
rect 19248 6808 19300 6860
rect 20628 6851 20680 6860
rect 20628 6817 20637 6851
rect 20637 6817 20671 6851
rect 20671 6817 20680 6851
rect 20628 6808 20680 6817
rect 20904 6851 20956 6860
rect 20904 6817 20913 6851
rect 20913 6817 20947 6851
rect 20947 6817 20956 6851
rect 20904 6808 20956 6817
rect 22100 6808 22152 6860
rect 19892 6740 19944 6792
rect 17592 6672 17644 6724
rect 15936 6604 15988 6656
rect 17500 6647 17552 6656
rect 17500 6613 17509 6647
rect 17509 6613 17543 6647
rect 17543 6613 17552 6647
rect 17500 6604 17552 6613
rect 18880 6672 18932 6724
rect 19156 6672 19208 6724
rect 20720 6740 20772 6792
rect 22468 6783 22520 6792
rect 20536 6672 20588 6724
rect 18420 6647 18472 6656
rect 18420 6613 18429 6647
rect 18429 6613 18463 6647
rect 18463 6613 18472 6647
rect 18696 6647 18748 6656
rect 18420 6604 18472 6613
rect 18696 6613 18705 6647
rect 18705 6613 18739 6647
rect 18739 6613 18748 6647
rect 18696 6604 18748 6613
rect 19064 6604 19116 6656
rect 22468 6749 22477 6783
rect 22477 6749 22511 6783
rect 22511 6749 22520 6783
rect 22468 6740 22520 6749
rect 22836 6783 22888 6792
rect 22836 6749 22845 6783
rect 22845 6749 22879 6783
rect 22879 6749 22888 6783
rect 22836 6740 22888 6749
rect 20904 6672 20956 6724
rect 21456 6672 21508 6724
rect 20996 6647 21048 6656
rect 20996 6613 21005 6647
rect 21005 6613 21039 6647
rect 21039 6613 21048 6647
rect 20996 6604 21048 6613
rect 21272 6604 21324 6656
rect 22008 6647 22060 6656
rect 22008 6613 22017 6647
rect 22017 6613 22051 6647
rect 22051 6613 22060 6647
rect 22008 6604 22060 6613
rect 22836 6604 22888 6656
rect 23020 6647 23072 6656
rect 23020 6613 23029 6647
rect 23029 6613 23063 6647
rect 23063 6613 23072 6647
rect 23020 6604 23072 6613
rect 6548 6502 6600 6554
rect 6612 6502 6664 6554
rect 6676 6502 6728 6554
rect 6740 6502 6792 6554
rect 6804 6502 6856 6554
rect 12146 6502 12198 6554
rect 12210 6502 12262 6554
rect 12274 6502 12326 6554
rect 12338 6502 12390 6554
rect 12402 6502 12454 6554
rect 17744 6502 17796 6554
rect 17808 6502 17860 6554
rect 17872 6502 17924 6554
rect 17936 6502 17988 6554
rect 18000 6502 18052 6554
rect 4804 6443 4856 6452
rect 4804 6409 4813 6443
rect 4813 6409 4847 6443
rect 4847 6409 4856 6443
rect 4804 6400 4856 6409
rect 6460 6443 6512 6452
rect 6460 6409 6469 6443
rect 6469 6409 6503 6443
rect 6503 6409 6512 6443
rect 6460 6400 6512 6409
rect 7564 6443 7616 6452
rect 7564 6409 7573 6443
rect 7573 6409 7607 6443
rect 7607 6409 7616 6443
rect 7564 6400 7616 6409
rect 7656 6400 7708 6452
rect 9220 6400 9272 6452
rect 10324 6400 10376 6452
rect 12716 6443 12768 6452
rect 12716 6409 12725 6443
rect 12725 6409 12759 6443
rect 12759 6409 12768 6443
rect 12716 6400 12768 6409
rect 12992 6400 13044 6452
rect 5908 6375 5960 6384
rect 5908 6341 5926 6375
rect 5926 6341 5960 6375
rect 5908 6332 5960 6341
rect 8300 6332 8352 6384
rect 7472 6264 7524 6316
rect 10416 6332 10468 6384
rect 7380 6239 7432 6248
rect 7380 6205 7389 6239
rect 7389 6205 7423 6239
rect 7423 6205 7432 6239
rect 8760 6239 8812 6248
rect 7380 6196 7432 6205
rect 8760 6205 8769 6239
rect 8769 6205 8803 6239
rect 8803 6205 8812 6239
rect 8760 6196 8812 6205
rect 11336 6332 11388 6384
rect 11428 6332 11480 6384
rect 15752 6400 15804 6452
rect 15936 6400 15988 6452
rect 16488 6400 16540 6452
rect 19432 6400 19484 6452
rect 20536 6400 20588 6452
rect 20720 6400 20772 6452
rect 21456 6443 21508 6452
rect 21456 6409 21465 6443
rect 21465 6409 21499 6443
rect 21499 6409 21508 6443
rect 21456 6400 21508 6409
rect 21640 6400 21692 6452
rect 15384 6332 15436 6384
rect 16764 6332 16816 6384
rect 10968 6307 11020 6316
rect 10968 6273 10977 6307
rect 10977 6273 11011 6307
rect 11011 6273 11020 6307
rect 10968 6264 11020 6273
rect 11888 6307 11940 6316
rect 11888 6273 11897 6307
rect 11897 6273 11931 6307
rect 11931 6273 11940 6307
rect 11888 6264 11940 6273
rect 15660 6264 15712 6316
rect 15844 6264 15896 6316
rect 18512 6264 18564 6316
rect 19156 6264 19208 6316
rect 19616 6332 19668 6384
rect 19800 6264 19852 6316
rect 19892 6264 19944 6316
rect 20904 6264 20956 6316
rect 21272 6264 21324 6316
rect 22468 6264 22520 6316
rect 23388 6264 23440 6316
rect 8484 6128 8536 6180
rect 9312 6196 9364 6248
rect 9956 6239 10008 6248
rect 9956 6205 9965 6239
rect 9965 6205 9999 6239
rect 9999 6205 10008 6239
rect 9956 6196 10008 6205
rect 11152 6196 11204 6248
rect 11612 6239 11664 6248
rect 11612 6205 11621 6239
rect 11621 6205 11655 6239
rect 11655 6205 11664 6239
rect 11612 6196 11664 6205
rect 12716 6196 12768 6248
rect 13544 6196 13596 6248
rect 13820 6239 13872 6248
rect 13820 6205 13829 6239
rect 13829 6205 13863 6239
rect 13863 6205 13872 6239
rect 13820 6196 13872 6205
rect 10048 6128 10100 6180
rect 14372 6171 14424 6180
rect 14372 6137 14381 6171
rect 14381 6137 14415 6171
rect 14415 6137 14424 6171
rect 14372 6128 14424 6137
rect 15292 6128 15344 6180
rect 16304 6196 16356 6248
rect 16672 6196 16724 6248
rect 16948 6239 17000 6248
rect 16948 6205 16957 6239
rect 16957 6205 16991 6239
rect 16991 6205 17000 6239
rect 16948 6196 17000 6205
rect 17776 6196 17828 6248
rect 17408 6128 17460 6180
rect 18972 6239 19024 6248
rect 18972 6205 18981 6239
rect 18981 6205 19015 6239
rect 19015 6205 19024 6239
rect 18972 6196 19024 6205
rect 17960 6128 18012 6180
rect 18788 6128 18840 6180
rect 8392 6060 8444 6112
rect 10416 6060 10468 6112
rect 11244 6060 11296 6112
rect 11336 6103 11388 6112
rect 11336 6069 11345 6103
rect 11345 6069 11379 6103
rect 11379 6069 11388 6103
rect 11336 6060 11388 6069
rect 14648 6060 14700 6112
rect 17040 6060 17092 6112
rect 17684 6060 17736 6112
rect 20536 6196 20588 6248
rect 22284 6239 22336 6248
rect 22284 6205 22293 6239
rect 22293 6205 22327 6239
rect 22327 6205 22336 6239
rect 22284 6196 22336 6205
rect 22376 6239 22428 6248
rect 22376 6205 22385 6239
rect 22385 6205 22419 6239
rect 22419 6205 22428 6239
rect 22376 6196 22428 6205
rect 22652 6171 22704 6180
rect 22652 6137 22661 6171
rect 22661 6137 22695 6171
rect 22695 6137 22704 6171
rect 22652 6128 22704 6137
rect 20352 6060 20404 6112
rect 20628 6060 20680 6112
rect 21916 6060 21968 6112
rect 22836 6060 22888 6112
rect 23020 6103 23072 6112
rect 23020 6069 23029 6103
rect 23029 6069 23063 6103
rect 23063 6069 23072 6103
rect 23020 6060 23072 6069
rect 3749 5958 3801 6010
rect 3813 5958 3865 6010
rect 3877 5958 3929 6010
rect 3941 5958 3993 6010
rect 4005 5958 4057 6010
rect 9347 5958 9399 6010
rect 9411 5958 9463 6010
rect 9475 5958 9527 6010
rect 9539 5958 9591 6010
rect 9603 5958 9655 6010
rect 14945 5958 14997 6010
rect 15009 5958 15061 6010
rect 15073 5958 15125 6010
rect 15137 5958 15189 6010
rect 15201 5958 15253 6010
rect 20543 5958 20595 6010
rect 20607 5958 20659 6010
rect 20671 5958 20723 6010
rect 20735 5958 20787 6010
rect 20799 5958 20851 6010
rect 8300 5788 8352 5840
rect 7380 5763 7432 5772
rect 7380 5729 7389 5763
rect 7389 5729 7423 5763
rect 7423 5729 7432 5763
rect 7380 5720 7432 5729
rect 10048 5899 10100 5908
rect 10048 5865 10057 5899
rect 10057 5865 10091 5899
rect 10091 5865 10100 5899
rect 10048 5856 10100 5865
rect 10968 5856 11020 5908
rect 8668 5720 8720 5772
rect 9496 5763 9548 5772
rect 9496 5729 9505 5763
rect 9505 5729 9539 5763
rect 9539 5729 9548 5763
rect 9496 5720 9548 5729
rect 7196 5652 7248 5704
rect 8392 5695 8444 5704
rect 8392 5661 8401 5695
rect 8401 5661 8435 5695
rect 8435 5661 8444 5695
rect 8392 5652 8444 5661
rect 9772 5652 9824 5704
rect 8576 5584 8628 5636
rect 9588 5584 9640 5636
rect 9956 5788 10008 5840
rect 10692 5763 10744 5772
rect 10692 5729 10701 5763
rect 10701 5729 10735 5763
rect 10735 5729 10744 5763
rect 10692 5720 10744 5729
rect 11152 5720 11204 5772
rect 12716 5763 12768 5772
rect 12716 5729 12725 5763
rect 12725 5729 12759 5763
rect 12759 5729 12768 5763
rect 12716 5720 12768 5729
rect 14648 5720 14700 5772
rect 10876 5652 10928 5704
rect 11244 5652 11296 5704
rect 15108 5652 15160 5704
rect 8944 5559 8996 5568
rect 8944 5525 8953 5559
rect 8953 5525 8987 5559
rect 8987 5525 8996 5559
rect 8944 5516 8996 5525
rect 11612 5516 11664 5568
rect 12624 5584 12676 5636
rect 16120 5763 16172 5772
rect 16120 5729 16129 5763
rect 16129 5729 16163 5763
rect 16163 5729 16172 5763
rect 17592 5856 17644 5908
rect 17776 5856 17828 5908
rect 21548 5856 21600 5908
rect 22652 5899 22704 5908
rect 22652 5865 22661 5899
rect 22661 5865 22695 5899
rect 22695 5865 22704 5899
rect 22652 5856 22704 5865
rect 20812 5788 20864 5840
rect 22100 5788 22152 5840
rect 16120 5720 16172 5729
rect 16580 5720 16632 5772
rect 18236 5763 18288 5772
rect 18236 5729 18245 5763
rect 18245 5729 18279 5763
rect 18279 5729 18288 5763
rect 18236 5720 18288 5729
rect 18512 5763 18564 5772
rect 18512 5729 18521 5763
rect 18521 5729 18555 5763
rect 18555 5729 18564 5763
rect 18512 5720 18564 5729
rect 19800 5763 19852 5772
rect 19800 5729 19809 5763
rect 19809 5729 19843 5763
rect 19843 5729 19852 5763
rect 19800 5720 19852 5729
rect 20076 5720 20128 5772
rect 21456 5763 21508 5772
rect 21456 5729 21465 5763
rect 21465 5729 21499 5763
rect 21499 5729 21508 5763
rect 23480 5788 23532 5840
rect 21456 5720 21508 5729
rect 16396 5695 16448 5704
rect 16396 5661 16405 5695
rect 16405 5661 16439 5695
rect 16439 5661 16448 5695
rect 16396 5652 16448 5661
rect 18420 5652 18472 5704
rect 19340 5652 19392 5704
rect 17316 5584 17368 5636
rect 18328 5584 18380 5636
rect 23204 5720 23256 5772
rect 22560 5652 22612 5704
rect 23112 5584 23164 5636
rect 11980 5559 12032 5568
rect 11980 5525 11989 5559
rect 11989 5525 12023 5559
rect 12023 5525 12032 5559
rect 11980 5516 12032 5525
rect 13820 5516 13872 5568
rect 14556 5559 14608 5568
rect 14556 5525 14571 5559
rect 14571 5525 14605 5559
rect 14605 5525 14608 5559
rect 14556 5516 14608 5525
rect 16672 5516 16724 5568
rect 17132 5559 17184 5568
rect 17132 5525 17141 5559
rect 17141 5525 17175 5559
rect 17175 5525 17184 5559
rect 17132 5516 17184 5525
rect 17224 5516 17276 5568
rect 17960 5516 18012 5568
rect 18236 5516 18288 5568
rect 19708 5559 19760 5568
rect 19708 5525 19717 5559
rect 19717 5525 19751 5559
rect 19751 5525 19760 5559
rect 19708 5516 19760 5525
rect 20444 5559 20496 5568
rect 20444 5525 20453 5559
rect 20453 5525 20487 5559
rect 20487 5525 20496 5559
rect 20444 5516 20496 5525
rect 21732 5516 21784 5568
rect 22652 5516 22704 5568
rect 23020 5559 23072 5568
rect 23020 5525 23029 5559
rect 23029 5525 23063 5559
rect 23063 5525 23072 5559
rect 23020 5516 23072 5525
rect 6548 5414 6600 5466
rect 6612 5414 6664 5466
rect 6676 5414 6728 5466
rect 6740 5414 6792 5466
rect 6804 5414 6856 5466
rect 12146 5414 12198 5466
rect 12210 5414 12262 5466
rect 12274 5414 12326 5466
rect 12338 5414 12390 5466
rect 12402 5414 12454 5466
rect 17744 5414 17796 5466
rect 17808 5414 17860 5466
rect 17872 5414 17924 5466
rect 17936 5414 17988 5466
rect 18000 5414 18052 5466
rect 9128 5355 9180 5364
rect 9128 5321 9137 5355
rect 9137 5321 9171 5355
rect 9171 5321 9180 5355
rect 9128 5312 9180 5321
rect 10048 5312 10100 5364
rect 12072 5312 12124 5364
rect 13176 5312 13228 5364
rect 15384 5355 15436 5364
rect 8944 5244 8996 5296
rect 14556 5287 14608 5296
rect 14556 5253 14565 5287
rect 14565 5253 14599 5287
rect 14599 5253 14608 5287
rect 14556 5244 14608 5253
rect 15384 5321 15393 5355
rect 15393 5321 15427 5355
rect 15427 5321 15436 5355
rect 15384 5312 15436 5321
rect 15660 5355 15712 5364
rect 15660 5321 15669 5355
rect 15669 5321 15703 5355
rect 15703 5321 15712 5355
rect 15660 5312 15712 5321
rect 16948 5312 17000 5364
rect 17132 5312 17184 5364
rect 17592 5312 17644 5364
rect 19340 5312 19392 5364
rect 19708 5312 19760 5364
rect 16396 5244 16448 5296
rect 16580 5244 16632 5296
rect 17500 5244 17552 5296
rect 18696 5244 18748 5296
rect 19064 5244 19116 5296
rect 22744 5355 22796 5364
rect 22744 5321 22753 5355
rect 22753 5321 22787 5355
rect 22787 5321 22796 5355
rect 22744 5312 22796 5321
rect 20260 5244 20312 5296
rect 8852 5176 8904 5228
rect 14832 5219 14884 5228
rect 14832 5185 14841 5219
rect 14841 5185 14875 5219
rect 14875 5185 14884 5219
rect 14832 5176 14884 5185
rect 8116 5151 8168 5160
rect 8116 5117 8125 5151
rect 8125 5117 8159 5151
rect 8159 5117 8168 5151
rect 8116 5108 8168 5117
rect 9312 5151 9364 5160
rect 9312 5117 9321 5151
rect 9321 5117 9355 5151
rect 9355 5117 9364 5151
rect 9312 5108 9364 5117
rect 11152 5108 11204 5160
rect 11796 5108 11848 5160
rect 15200 5176 15252 5228
rect 16028 5219 16080 5228
rect 16028 5185 16037 5219
rect 16037 5185 16071 5219
rect 16071 5185 16080 5219
rect 16028 5176 16080 5185
rect 18236 5176 18288 5228
rect 18788 5219 18840 5228
rect 18788 5185 18797 5219
rect 18797 5185 18831 5219
rect 18831 5185 18840 5219
rect 18788 5176 18840 5185
rect 18972 5176 19024 5228
rect 19892 5176 19944 5228
rect 16212 5151 16264 5160
rect 16212 5117 16221 5151
rect 16221 5117 16255 5151
rect 16255 5117 16264 5151
rect 16212 5108 16264 5117
rect 16580 5108 16632 5160
rect 16856 5108 16908 5160
rect 17408 5108 17460 5160
rect 18604 5151 18656 5160
rect 18604 5117 18613 5151
rect 18613 5117 18647 5151
rect 18647 5117 18656 5151
rect 18604 5108 18656 5117
rect 19432 5151 19484 5160
rect 14188 4972 14240 5024
rect 17132 5040 17184 5092
rect 19432 5117 19441 5151
rect 19441 5117 19475 5151
rect 19475 5117 19484 5151
rect 19432 5108 19484 5117
rect 19524 5151 19576 5160
rect 19524 5117 19533 5151
rect 19533 5117 19567 5151
rect 19567 5117 19576 5151
rect 20812 5244 20864 5296
rect 21272 5219 21324 5228
rect 21272 5185 21281 5219
rect 21281 5185 21315 5219
rect 21315 5185 21324 5219
rect 21272 5176 21324 5185
rect 22836 5219 22888 5228
rect 22836 5185 22845 5219
rect 22845 5185 22879 5219
rect 22879 5185 22888 5219
rect 22836 5176 22888 5185
rect 19524 5108 19576 5117
rect 15660 4972 15712 5024
rect 16028 4972 16080 5024
rect 17500 5015 17552 5024
rect 17500 4981 17509 5015
rect 17509 4981 17543 5015
rect 17543 4981 17552 5015
rect 17500 4972 17552 4981
rect 19340 5040 19392 5092
rect 20904 5108 20956 5160
rect 19984 5015 20036 5024
rect 19984 4981 19993 5015
rect 19993 4981 20027 5015
rect 20027 4981 20036 5015
rect 19984 4972 20036 4981
rect 20260 5040 20312 5092
rect 22376 5151 22428 5160
rect 22376 5117 22385 5151
rect 22385 5117 22419 5151
rect 22419 5117 22428 5151
rect 22376 5108 22428 5117
rect 21640 5083 21692 5092
rect 21640 5049 21649 5083
rect 21649 5049 21683 5083
rect 21683 5049 21692 5083
rect 21640 5040 21692 5049
rect 22560 5040 22612 5092
rect 21456 4972 21508 5024
rect 21824 5015 21876 5024
rect 21824 4981 21833 5015
rect 21833 4981 21867 5015
rect 21867 4981 21876 5015
rect 21824 4972 21876 4981
rect 23020 5015 23072 5024
rect 23020 4981 23029 5015
rect 23029 4981 23063 5015
rect 23063 4981 23072 5015
rect 23020 4972 23072 4981
rect 3749 4870 3801 4922
rect 3813 4870 3865 4922
rect 3877 4870 3929 4922
rect 3941 4870 3993 4922
rect 4005 4870 4057 4922
rect 9347 4870 9399 4922
rect 9411 4870 9463 4922
rect 9475 4870 9527 4922
rect 9539 4870 9591 4922
rect 9603 4870 9655 4922
rect 14945 4870 14997 4922
rect 15009 4870 15061 4922
rect 15073 4870 15125 4922
rect 15137 4870 15189 4922
rect 15201 4870 15253 4922
rect 20543 4870 20595 4922
rect 20607 4870 20659 4922
rect 20671 4870 20723 4922
rect 20735 4870 20787 4922
rect 20799 4870 20851 4922
rect 14832 4768 14884 4820
rect 19524 4768 19576 4820
rect 20260 4768 20312 4820
rect 22376 4768 22428 4820
rect 10048 4700 10100 4752
rect 18788 4700 18840 4752
rect 8116 4675 8168 4684
rect 8116 4641 8125 4675
rect 8125 4641 8159 4675
rect 8159 4641 8168 4675
rect 8300 4675 8352 4684
rect 8116 4632 8168 4641
rect 8300 4641 8309 4675
rect 8309 4641 8343 4675
rect 8343 4641 8352 4675
rect 8300 4632 8352 4641
rect 10416 4632 10468 4684
rect 8484 4564 8536 4616
rect 8208 4496 8260 4548
rect 13820 4564 13872 4616
rect 16672 4632 16724 4684
rect 17040 4675 17092 4684
rect 16764 4607 16816 4616
rect 16764 4573 16773 4607
rect 16773 4573 16807 4607
rect 16807 4573 16816 4607
rect 16764 4564 16816 4573
rect 17040 4641 17046 4675
rect 17046 4641 17080 4675
rect 17080 4641 17092 4675
rect 17040 4632 17092 4641
rect 17316 4632 17368 4684
rect 18144 4632 18196 4684
rect 18972 4632 19024 4684
rect 20076 4632 20128 4684
rect 20444 4632 20496 4684
rect 23296 4632 23348 4684
rect 17408 4564 17460 4616
rect 18236 4564 18288 4616
rect 19064 4564 19116 4616
rect 19616 4564 19668 4616
rect 20812 4607 20864 4616
rect 13728 4496 13780 4548
rect 20812 4573 20821 4607
rect 20821 4573 20855 4607
rect 20855 4573 20864 4607
rect 20812 4564 20864 4573
rect 21364 4564 21416 4616
rect 21640 4564 21692 4616
rect 15568 4471 15620 4480
rect 15568 4437 15577 4471
rect 15577 4437 15611 4471
rect 15611 4437 15620 4471
rect 15568 4428 15620 4437
rect 16856 4428 16908 4480
rect 17132 4428 17184 4480
rect 18788 4428 18840 4480
rect 19156 4428 19208 4480
rect 19616 4471 19668 4480
rect 19616 4437 19625 4471
rect 19625 4437 19659 4471
rect 19659 4437 19668 4471
rect 19616 4428 19668 4437
rect 20352 4471 20404 4480
rect 20352 4437 20361 4471
rect 20361 4437 20395 4471
rect 20395 4437 20404 4471
rect 20352 4428 20404 4437
rect 20812 4428 20864 4480
rect 21088 4428 21140 4480
rect 21180 4428 21232 4480
rect 21456 4428 21508 4480
rect 23020 4471 23072 4480
rect 23020 4437 23029 4471
rect 23029 4437 23063 4471
rect 23063 4437 23072 4471
rect 23020 4428 23072 4437
rect 6548 4326 6600 4378
rect 6612 4326 6664 4378
rect 6676 4326 6728 4378
rect 6740 4326 6792 4378
rect 6804 4326 6856 4378
rect 12146 4326 12198 4378
rect 12210 4326 12262 4378
rect 12274 4326 12326 4378
rect 12338 4326 12390 4378
rect 12402 4326 12454 4378
rect 17744 4326 17796 4378
rect 17808 4326 17860 4378
rect 17872 4326 17924 4378
rect 17936 4326 17988 4378
rect 18000 4326 18052 4378
rect 15568 4224 15620 4276
rect 18972 4224 19024 4276
rect 21272 4267 21324 4276
rect 21272 4233 21281 4267
rect 21281 4233 21315 4267
rect 21315 4233 21324 4267
rect 21272 4224 21324 4233
rect 22008 4267 22060 4276
rect 22008 4233 22017 4267
rect 22017 4233 22051 4267
rect 22051 4233 22060 4267
rect 22008 4224 22060 4233
rect 22376 4224 22428 4276
rect 15660 4199 15712 4208
rect 15660 4165 15669 4199
rect 15669 4165 15703 4199
rect 15703 4165 15712 4199
rect 15660 4156 15712 4165
rect 11888 4088 11940 4140
rect 16948 4088 17000 4140
rect 17500 4088 17552 4140
rect 17684 4088 17736 4140
rect 15568 4063 15620 4072
rect 15568 4029 15577 4063
rect 15577 4029 15611 4063
rect 15611 4029 15620 4063
rect 15568 4020 15620 4029
rect 16120 4020 16172 4072
rect 18420 4088 18472 4140
rect 17960 4020 18012 4072
rect 18144 4020 18196 4072
rect 18512 4063 18564 4072
rect 18512 4029 18521 4063
rect 18521 4029 18555 4063
rect 18555 4029 18564 4063
rect 18512 4020 18564 4029
rect 14188 3952 14240 4004
rect 16672 3927 16724 3936
rect 16672 3893 16681 3927
rect 16681 3893 16715 3927
rect 16715 3893 16724 3927
rect 16672 3884 16724 3893
rect 19432 4156 19484 4208
rect 23756 4224 23808 4276
rect 18880 4131 18932 4140
rect 18880 4097 18889 4131
rect 18889 4097 18923 4131
rect 18923 4097 18932 4131
rect 18880 4088 18932 4097
rect 19156 4131 19208 4140
rect 19156 4097 19165 4131
rect 19165 4097 19199 4131
rect 19199 4097 19208 4131
rect 19156 4088 19208 4097
rect 19524 4020 19576 4072
rect 21824 4088 21876 4140
rect 21916 4131 21968 4140
rect 21916 4097 21925 4131
rect 21925 4097 21959 4131
rect 21959 4097 21968 4131
rect 22560 4156 22612 4208
rect 21916 4088 21968 4097
rect 19340 3927 19392 3936
rect 19340 3893 19349 3927
rect 19349 3893 19383 3927
rect 19383 3893 19392 3927
rect 19340 3884 19392 3893
rect 19524 3884 19576 3936
rect 22284 3952 22336 4004
rect 20168 3927 20220 3936
rect 20168 3893 20177 3927
rect 20177 3893 20211 3927
rect 20211 3893 20220 3927
rect 20168 3884 20220 3893
rect 20444 3884 20496 3936
rect 20536 3884 20588 3936
rect 23020 3927 23072 3936
rect 23020 3893 23029 3927
rect 23029 3893 23063 3927
rect 23063 3893 23072 3927
rect 23020 3884 23072 3893
rect 3749 3782 3801 3834
rect 3813 3782 3865 3834
rect 3877 3782 3929 3834
rect 3941 3782 3993 3834
rect 4005 3782 4057 3834
rect 9347 3782 9399 3834
rect 9411 3782 9463 3834
rect 9475 3782 9527 3834
rect 9539 3782 9591 3834
rect 9603 3782 9655 3834
rect 14945 3782 14997 3834
rect 15009 3782 15061 3834
rect 15073 3782 15125 3834
rect 15137 3782 15189 3834
rect 15201 3782 15253 3834
rect 20543 3782 20595 3834
rect 20607 3782 20659 3834
rect 20671 3782 20723 3834
rect 20735 3782 20787 3834
rect 20799 3782 20851 3834
rect 17316 3680 17368 3732
rect 19432 3723 19484 3732
rect 19432 3689 19441 3723
rect 19441 3689 19475 3723
rect 19475 3689 19484 3723
rect 19432 3680 19484 3689
rect 20352 3680 20404 3732
rect 18144 3612 18196 3664
rect 18972 3612 19024 3664
rect 16856 3587 16908 3596
rect 16856 3553 16865 3587
rect 16865 3553 16899 3587
rect 16899 3553 16908 3587
rect 16856 3544 16908 3553
rect 17040 3544 17092 3596
rect 17224 3544 17276 3596
rect 16212 3476 16264 3528
rect 16580 3476 16632 3528
rect 17316 3476 17368 3528
rect 18328 3544 18380 3596
rect 19156 3612 19208 3664
rect 20260 3612 20312 3664
rect 18696 3476 18748 3528
rect 19524 3544 19576 3596
rect 20444 3587 20496 3596
rect 19156 3476 19208 3528
rect 20444 3553 20453 3587
rect 20453 3553 20487 3587
rect 20487 3553 20496 3587
rect 20444 3544 20496 3553
rect 22468 3680 22520 3732
rect 22560 3655 22612 3664
rect 22560 3621 22569 3655
rect 22569 3621 22603 3655
rect 22603 3621 22612 3655
rect 22560 3612 22612 3621
rect 21364 3544 21416 3596
rect 22192 3587 22244 3596
rect 22192 3553 22201 3587
rect 22201 3553 22235 3587
rect 22235 3553 22244 3587
rect 22192 3544 22244 3553
rect 20904 3476 20956 3528
rect 21456 3476 21508 3528
rect 23572 3680 23624 3732
rect 23664 3612 23716 3664
rect 23112 3476 23164 3528
rect 20168 3408 20220 3460
rect 1400 3383 1452 3392
rect 1400 3349 1409 3383
rect 1409 3349 1443 3383
rect 1443 3349 1452 3383
rect 1400 3340 1452 3349
rect 15752 3383 15804 3392
rect 15752 3349 15761 3383
rect 15761 3349 15795 3383
rect 15795 3349 15804 3383
rect 15752 3340 15804 3349
rect 17132 3383 17184 3392
rect 17132 3349 17134 3383
rect 17134 3349 17168 3383
rect 17168 3349 17184 3383
rect 17132 3340 17184 3349
rect 17224 3340 17276 3392
rect 19616 3340 19668 3392
rect 19892 3383 19944 3392
rect 19892 3349 19901 3383
rect 19901 3349 19935 3383
rect 19935 3349 19944 3383
rect 19892 3340 19944 3349
rect 19984 3340 20036 3392
rect 21640 3383 21692 3392
rect 21640 3349 21649 3383
rect 21649 3349 21683 3383
rect 21683 3349 21692 3383
rect 21640 3340 21692 3349
rect 22928 3408 22980 3460
rect 23020 3383 23072 3392
rect 23020 3349 23029 3383
rect 23029 3349 23063 3383
rect 23063 3349 23072 3383
rect 23020 3340 23072 3349
rect 6548 3238 6600 3290
rect 6612 3238 6664 3290
rect 6676 3238 6728 3290
rect 6740 3238 6792 3290
rect 6804 3238 6856 3290
rect 12146 3238 12198 3290
rect 12210 3238 12262 3290
rect 12274 3238 12326 3290
rect 12338 3238 12390 3290
rect 12402 3238 12454 3290
rect 17744 3238 17796 3290
rect 17808 3238 17860 3290
rect 17872 3238 17924 3290
rect 17936 3238 17988 3290
rect 18000 3238 18052 3290
rect 11336 3136 11388 3188
rect 18972 3136 19024 3188
rect 19064 3136 19116 3188
rect 21180 3136 21232 3188
rect 16212 3111 16264 3120
rect 16212 3077 16221 3111
rect 16221 3077 16255 3111
rect 16255 3077 16264 3111
rect 16212 3068 16264 3077
rect 8392 2839 8444 2848
rect 8392 2805 8401 2839
rect 8401 2805 8435 2839
rect 8435 2805 8444 2839
rect 8392 2796 8444 2805
rect 16764 3000 16816 3052
rect 19248 3000 19300 3052
rect 19708 3043 19760 3052
rect 19708 3009 19717 3043
rect 19717 3009 19751 3043
rect 19751 3009 19760 3043
rect 19708 3000 19760 3009
rect 16580 2932 16632 2984
rect 17040 2932 17092 2984
rect 17224 2932 17276 2984
rect 17408 2975 17460 2984
rect 17408 2941 17417 2975
rect 17417 2941 17451 2975
rect 17451 2941 17460 2975
rect 17408 2932 17460 2941
rect 10784 2796 10836 2848
rect 11980 2796 12032 2848
rect 18328 2796 18380 2848
rect 18420 2796 18472 2848
rect 18788 2932 18840 2984
rect 21548 3000 21600 3052
rect 22744 3136 22796 3188
rect 22652 3068 22704 3120
rect 18696 2796 18748 2848
rect 21088 2932 21140 2984
rect 22652 2932 22704 2984
rect 23388 2932 23440 2984
rect 23020 2839 23072 2848
rect 23020 2805 23029 2839
rect 23029 2805 23063 2839
rect 23063 2805 23072 2839
rect 23020 2796 23072 2805
rect 23112 2796 23164 2848
rect 23848 2796 23900 2848
rect 3749 2694 3801 2746
rect 3813 2694 3865 2746
rect 3877 2694 3929 2746
rect 3941 2694 3993 2746
rect 4005 2694 4057 2746
rect 9347 2694 9399 2746
rect 9411 2694 9463 2746
rect 9475 2694 9527 2746
rect 9539 2694 9591 2746
rect 9603 2694 9655 2746
rect 14945 2694 14997 2746
rect 15009 2694 15061 2746
rect 15073 2694 15125 2746
rect 15137 2694 15189 2746
rect 15201 2694 15253 2746
rect 20543 2694 20595 2746
rect 20607 2694 20659 2746
rect 20671 2694 20723 2746
rect 20735 2694 20787 2746
rect 20799 2694 20851 2746
rect 10784 2635 10836 2644
rect 10784 2601 10793 2635
rect 10793 2601 10827 2635
rect 10827 2601 10836 2635
rect 10784 2592 10836 2601
rect 15752 2592 15804 2644
rect 16764 2635 16816 2644
rect 16764 2601 16773 2635
rect 16773 2601 16807 2635
rect 16807 2601 16816 2635
rect 16764 2592 16816 2601
rect 23112 2592 23164 2644
rect 8392 2456 8444 2508
rect 6184 2388 6236 2440
rect 22652 2431 22704 2440
rect 22652 2397 22661 2431
rect 22661 2397 22695 2431
rect 22695 2397 22704 2431
rect 22652 2388 22704 2397
rect 2136 2252 2188 2304
rect 10232 2252 10284 2304
rect 22376 2252 22428 2304
rect 6548 2150 6600 2202
rect 6612 2150 6664 2202
rect 6676 2150 6728 2202
rect 6740 2150 6792 2202
rect 6804 2150 6856 2202
rect 12146 2150 12198 2202
rect 12210 2150 12262 2202
rect 12274 2150 12326 2202
rect 12338 2150 12390 2202
rect 12402 2150 12454 2202
rect 17744 2150 17796 2202
rect 17808 2150 17860 2202
rect 17872 2150 17924 2202
rect 17936 2150 17988 2202
rect 18000 2150 18052 2202
<< metal2 >>
rect 294 23800 350 24600
rect 938 23800 994 24600
rect 1582 23800 1638 24600
rect 2226 23800 2282 24600
rect 2870 23800 2926 24600
rect 3514 23800 3570 24600
rect 4158 23800 4214 24600
rect 4802 23800 4858 24600
rect 5446 23800 5502 24600
rect 6090 23800 6146 24600
rect 6734 23800 6790 24600
rect 7378 23800 7434 24600
rect 8022 23800 8078 24600
rect 8666 23800 8722 24600
rect 9310 23800 9366 24600
rect 9954 23800 10010 24600
rect 10598 23800 10654 24600
rect 11242 23800 11298 24600
rect 11886 23800 11942 24600
rect 12530 23800 12586 24600
rect 13174 23800 13230 24600
rect 13818 23800 13874 24600
rect 14462 23800 14518 24600
rect 14844 23854 15056 23882
rect 308 21690 336 23800
rect 296 21684 348 21690
rect 296 21626 348 21632
rect 952 21418 980 23800
rect 1596 21894 1624 23800
rect 2240 21894 2268 23800
rect 2412 22024 2464 22030
rect 2412 21966 2464 21972
rect 1584 21888 1636 21894
rect 1584 21830 1636 21836
rect 2228 21888 2280 21894
rect 2228 21830 2280 21836
rect 2424 21690 2452 21966
rect 2884 21894 2912 23800
rect 2964 22024 3016 22030
rect 2964 21966 3016 21972
rect 3240 22024 3292 22030
rect 3240 21966 3292 21972
rect 2872 21888 2924 21894
rect 2872 21830 2924 21836
rect 2976 21690 3004 21966
rect 3252 21690 3280 21966
rect 3528 21894 3556 23800
rect 3749 22332 4057 22341
rect 3749 22330 3755 22332
rect 3811 22330 3835 22332
rect 3891 22330 3915 22332
rect 3971 22330 3995 22332
rect 4051 22330 4057 22332
rect 3811 22278 3813 22330
rect 3993 22278 3995 22330
rect 3749 22276 3755 22278
rect 3811 22276 3835 22278
rect 3891 22276 3915 22278
rect 3971 22276 3995 22278
rect 4051 22276 4057 22278
rect 3749 22267 4057 22276
rect 4172 22114 4200 23800
rect 4172 22086 4292 22114
rect 4160 22024 4212 22030
rect 4160 21966 4212 21972
rect 3700 21956 3752 21962
rect 3700 21898 3752 21904
rect 3516 21888 3568 21894
rect 3516 21830 3568 21836
rect 3712 21690 3740 21898
rect 2412 21684 2464 21690
rect 2412 21626 2464 21632
rect 2964 21684 3016 21690
rect 2964 21626 3016 21632
rect 3240 21684 3292 21690
rect 3240 21626 3292 21632
rect 3700 21684 3752 21690
rect 3700 21626 3752 21632
rect 3974 21584 4030 21593
rect 2780 21548 2832 21554
rect 2780 21490 2832 21496
rect 2964 21548 3016 21554
rect 2964 21490 3016 21496
rect 3148 21548 3200 21554
rect 3148 21490 3200 21496
rect 3424 21548 3476 21554
rect 3424 21490 3476 21496
rect 3608 21548 3660 21554
rect 3974 21519 3976 21528
rect 3608 21490 3660 21496
rect 4028 21519 4030 21528
rect 3976 21490 4028 21496
rect 940 21412 992 21418
rect 940 21354 992 21360
rect 1400 21344 1452 21350
rect 1400 21286 1452 21292
rect 1412 14482 1440 21286
rect 2792 21078 2820 21490
rect 2976 21078 3004 21490
rect 2780 21072 2832 21078
rect 2778 21040 2780 21049
rect 2964 21072 3016 21078
rect 2832 21040 2834 21049
rect 2964 21014 3016 21020
rect 2778 20975 2834 20984
rect 3160 20874 3188 21490
rect 3240 21480 3292 21486
rect 3240 21422 3292 21428
rect 3148 20868 3200 20874
rect 3148 20810 3200 20816
rect 1584 20324 1636 20330
rect 1584 20266 1636 20272
rect 1492 16448 1544 16454
rect 1492 16390 1544 16396
rect 1504 16114 1532 16390
rect 1492 16108 1544 16114
rect 1492 16050 1544 16056
rect 1492 15360 1544 15366
rect 1490 15328 1492 15337
rect 1544 15328 1546 15337
rect 1490 15263 1546 15272
rect 1596 14958 1624 20266
rect 2136 20256 2188 20262
rect 2136 20198 2188 20204
rect 2044 19372 2096 19378
rect 2044 19314 2096 19320
rect 1952 19168 2004 19174
rect 1952 19110 2004 19116
rect 1964 18834 1992 19110
rect 1952 18828 2004 18834
rect 1952 18770 2004 18776
rect 1952 18692 2004 18698
rect 1952 18634 2004 18640
rect 1676 18624 1728 18630
rect 1676 18566 1728 18572
rect 1688 16250 1716 18566
rect 1860 18284 1912 18290
rect 1860 18226 1912 18232
rect 1872 17338 1900 18226
rect 1964 17882 1992 18634
rect 1952 17876 2004 17882
rect 1952 17818 2004 17824
rect 1860 17332 1912 17338
rect 1860 17274 1912 17280
rect 1860 17128 1912 17134
rect 1860 17070 1912 17076
rect 1768 16992 1820 16998
rect 1768 16934 1820 16940
rect 1676 16244 1728 16250
rect 1676 16186 1728 16192
rect 1780 16114 1808 16934
rect 1768 16108 1820 16114
rect 1768 16050 1820 16056
rect 1676 15496 1728 15502
rect 1676 15438 1728 15444
rect 1584 14952 1636 14958
rect 1584 14894 1636 14900
rect 1400 14476 1452 14482
rect 1400 14418 1452 14424
rect 1688 13530 1716 15438
rect 1872 15042 1900 17070
rect 1952 16720 2004 16726
rect 1952 16662 2004 16668
rect 1964 16250 1992 16662
rect 1952 16244 2004 16250
rect 1952 16186 2004 16192
rect 2056 15706 2084 19314
rect 2148 17746 2176 20198
rect 3148 19984 3200 19990
rect 3148 19926 3200 19932
rect 2228 19848 2280 19854
rect 2228 19790 2280 19796
rect 2136 17740 2188 17746
rect 2136 17682 2188 17688
rect 2240 17678 2268 19790
rect 2504 19712 2556 19718
rect 2504 19654 2556 19660
rect 2412 19508 2464 19514
rect 2412 19450 2464 19456
rect 2320 18624 2372 18630
rect 2320 18566 2372 18572
rect 2332 18426 2360 18566
rect 2320 18420 2372 18426
rect 2320 18362 2372 18368
rect 2424 18290 2452 19450
rect 2412 18284 2464 18290
rect 2412 18226 2464 18232
rect 2228 17672 2280 17678
rect 2228 17614 2280 17620
rect 2136 17332 2188 17338
rect 2136 17274 2188 17280
rect 2044 15700 2096 15706
rect 2044 15642 2096 15648
rect 1780 15026 1900 15042
rect 1768 15020 1900 15026
rect 1820 15014 1900 15020
rect 1768 14962 1820 14968
rect 1676 13524 1728 13530
rect 1676 13466 1728 13472
rect 1780 12442 1808 14962
rect 2148 13410 2176 17274
rect 2240 13530 2268 17614
rect 2516 17134 2544 19654
rect 2596 19440 2648 19446
rect 2596 19382 2648 19388
rect 2686 19408 2742 19417
rect 2608 17338 2636 19382
rect 2686 19343 2688 19352
rect 2740 19343 2742 19352
rect 2688 19314 2740 19320
rect 2780 19304 2832 19310
rect 2780 19246 2832 19252
rect 2686 18728 2742 18737
rect 2686 18663 2742 18672
rect 2700 18630 2728 18663
rect 2688 18624 2740 18630
rect 2688 18566 2740 18572
rect 2688 17536 2740 17542
rect 2688 17478 2740 17484
rect 2596 17332 2648 17338
rect 2596 17274 2648 17280
rect 2504 17128 2556 17134
rect 2504 17070 2556 17076
rect 2596 17128 2648 17134
rect 2700 17116 2728 17478
rect 2648 17088 2728 17116
rect 2596 17070 2648 17076
rect 2320 16584 2372 16590
rect 2320 16526 2372 16532
rect 2332 15162 2360 16526
rect 2410 16416 2466 16425
rect 2410 16351 2466 16360
rect 2424 16250 2452 16351
rect 2412 16244 2464 16250
rect 2412 16186 2464 16192
rect 2608 15450 2636 17070
rect 2792 17066 2820 19246
rect 2964 18080 3016 18086
rect 2964 18022 3016 18028
rect 2872 17196 2924 17202
rect 2872 17138 2924 17144
rect 2780 17060 2832 17066
rect 2780 17002 2832 17008
rect 2792 16674 2820 17002
rect 2884 16794 2912 17138
rect 2872 16788 2924 16794
rect 2872 16730 2924 16736
rect 2700 16658 2820 16674
rect 2976 16658 3004 18022
rect 3160 17610 3188 19926
rect 3252 19310 3280 21422
rect 3436 20942 3464 21490
rect 3424 20936 3476 20942
rect 3424 20878 3476 20884
rect 3620 20806 3648 21490
rect 3749 21244 4057 21253
rect 3749 21242 3755 21244
rect 3811 21242 3835 21244
rect 3891 21242 3915 21244
rect 3971 21242 3995 21244
rect 4051 21242 4057 21244
rect 3811 21190 3813 21242
rect 3993 21190 3995 21242
rect 3749 21188 3755 21190
rect 3811 21188 3835 21190
rect 3891 21188 3915 21190
rect 3971 21188 3995 21190
rect 4051 21188 4057 21190
rect 3749 21179 4057 21188
rect 4172 21162 4200 21966
rect 4264 21894 4292 22086
rect 4816 21894 4844 23800
rect 5172 22636 5224 22642
rect 5172 22578 5224 22584
rect 4988 22024 5040 22030
rect 4988 21966 5040 21972
rect 4252 21888 4304 21894
rect 4252 21830 4304 21836
rect 4620 21888 4672 21894
rect 4620 21830 4672 21836
rect 4804 21888 4856 21894
rect 4804 21830 4856 21836
rect 4252 21616 4304 21622
rect 4252 21558 4304 21564
rect 4264 21321 4292 21558
rect 4342 21448 4398 21457
rect 4342 21383 4398 21392
rect 4250 21312 4306 21321
rect 4250 21247 4306 21256
rect 4080 21146 4200 21162
rect 4356 21146 4384 21383
rect 4528 21344 4580 21350
rect 4528 21286 4580 21292
rect 4068 21140 4200 21146
rect 4120 21134 4200 21140
rect 4344 21140 4396 21146
rect 4068 21082 4120 21088
rect 4344 21082 4396 21088
rect 4356 20942 4384 21082
rect 3700 20936 3752 20942
rect 3698 20904 3700 20913
rect 4344 20936 4396 20942
rect 3752 20904 3754 20913
rect 4344 20878 4396 20884
rect 3698 20839 3754 20848
rect 3608 20800 3660 20806
rect 3608 20742 3660 20748
rect 3884 20800 3936 20806
rect 3884 20742 3936 20748
rect 4344 20800 4396 20806
rect 4344 20742 4396 20748
rect 3896 20505 3924 20742
rect 3882 20496 3938 20505
rect 3882 20431 3938 20440
rect 3749 20156 4057 20165
rect 3749 20154 3755 20156
rect 3811 20154 3835 20156
rect 3891 20154 3915 20156
rect 3971 20154 3995 20156
rect 4051 20154 4057 20156
rect 3811 20102 3813 20154
rect 3993 20102 3995 20154
rect 3749 20100 3755 20102
rect 3811 20100 3835 20102
rect 3891 20100 3915 20102
rect 3971 20100 3995 20102
rect 4051 20100 4057 20102
rect 3749 20091 4057 20100
rect 3516 19848 3568 19854
rect 3516 19790 3568 19796
rect 3424 19440 3476 19446
rect 3424 19382 3476 19388
rect 3332 19372 3384 19378
rect 3332 19314 3384 19320
rect 3240 19304 3292 19310
rect 3240 19246 3292 19252
rect 3240 18624 3292 18630
rect 3240 18566 3292 18572
rect 3148 17604 3200 17610
rect 3148 17546 3200 17552
rect 3160 17202 3188 17546
rect 3252 17338 3280 18566
rect 3344 17882 3372 19314
rect 3436 17882 3464 19382
rect 3528 18970 3556 19790
rect 3976 19712 4028 19718
rect 3976 19654 4028 19660
rect 3988 19514 4016 19654
rect 3976 19508 4028 19514
rect 3976 19450 4028 19456
rect 3608 19236 3660 19242
rect 3608 19178 3660 19184
rect 3516 18964 3568 18970
rect 3516 18906 3568 18912
rect 3516 18216 3568 18222
rect 3516 18158 3568 18164
rect 3332 17876 3384 17882
rect 3332 17818 3384 17824
rect 3424 17876 3476 17882
rect 3424 17818 3476 17824
rect 3528 17746 3556 18158
rect 3516 17740 3568 17746
rect 3516 17682 3568 17688
rect 3240 17332 3292 17338
rect 3240 17274 3292 17280
rect 3148 17196 3200 17202
rect 3148 17138 3200 17144
rect 3528 17134 3556 17682
rect 3516 17128 3568 17134
rect 3516 17070 3568 17076
rect 2700 16652 2832 16658
rect 2700 16646 2780 16652
rect 2700 15570 2728 16646
rect 2780 16594 2832 16600
rect 2964 16652 3016 16658
rect 2964 16594 3016 16600
rect 3528 16590 3556 17070
rect 3516 16584 3568 16590
rect 3516 16526 3568 16532
rect 2872 16448 2924 16454
rect 2872 16390 2924 16396
rect 2884 16250 2912 16390
rect 3528 16250 3556 16526
rect 3620 16454 3648 19178
rect 3749 19068 4057 19077
rect 3749 19066 3755 19068
rect 3811 19066 3835 19068
rect 3891 19066 3915 19068
rect 3971 19066 3995 19068
rect 4051 19066 4057 19068
rect 3811 19014 3813 19066
rect 3993 19014 3995 19066
rect 3749 19012 3755 19014
rect 3811 19012 3835 19014
rect 3891 19012 3915 19014
rect 3971 19012 3995 19014
rect 4051 19012 4057 19014
rect 3749 19003 4057 19012
rect 4356 18902 4384 20742
rect 4434 19816 4490 19825
rect 4434 19751 4490 19760
rect 4448 19514 4476 19751
rect 4436 19508 4488 19514
rect 4436 19450 4488 19456
rect 4436 19372 4488 19378
rect 4436 19314 4488 19320
rect 4344 18896 4396 18902
rect 4344 18838 4396 18844
rect 4252 18760 4304 18766
rect 4448 18714 4476 19314
rect 4252 18702 4304 18708
rect 4160 18692 4212 18698
rect 4160 18634 4212 18640
rect 4172 18290 4200 18634
rect 4068 18284 4120 18290
rect 4068 18226 4120 18232
rect 4160 18284 4212 18290
rect 4160 18226 4212 18232
rect 4080 18170 4108 18226
rect 4080 18142 4200 18170
rect 3749 17980 4057 17989
rect 3749 17978 3755 17980
rect 3811 17978 3835 17980
rect 3891 17978 3915 17980
rect 3971 17978 3995 17980
rect 4051 17978 4057 17980
rect 3811 17926 3813 17978
rect 3993 17926 3995 17978
rect 3749 17924 3755 17926
rect 3811 17924 3835 17926
rect 3891 17924 3915 17926
rect 3971 17924 3995 17926
rect 4051 17924 4057 17926
rect 3749 17915 4057 17924
rect 4172 17814 4200 18142
rect 4160 17808 4212 17814
rect 4160 17750 4212 17756
rect 4264 17746 4292 18702
rect 4356 18686 4476 18714
rect 4252 17740 4304 17746
rect 4252 17682 4304 17688
rect 4356 17678 4384 18686
rect 4436 18624 4488 18630
rect 4436 18566 4488 18572
rect 4344 17672 4396 17678
rect 4344 17614 4396 17620
rect 4448 17542 4476 18566
rect 4540 17746 4568 21286
rect 4632 20330 4660 21830
rect 5000 21690 5028 21966
rect 4988 21684 5040 21690
rect 4988 21626 5040 21632
rect 5184 21554 5212 22578
rect 5460 22098 5488 23800
rect 5724 22228 5776 22234
rect 5724 22170 5776 22176
rect 5448 22092 5500 22098
rect 5448 22034 5500 22040
rect 5632 21684 5684 21690
rect 5632 21626 5684 21632
rect 5448 21616 5500 21622
rect 5644 21570 5672 21626
rect 5500 21564 5672 21570
rect 5448 21558 5672 21564
rect 5172 21548 5224 21554
rect 5460 21542 5672 21558
rect 5736 21554 5764 22170
rect 6104 22098 6132 23800
rect 6748 22114 6776 23800
rect 6472 22098 6868 22114
rect 7392 22098 7420 23800
rect 7472 22704 7524 22710
rect 7472 22646 7524 22652
rect 6092 22092 6144 22098
rect 6092 22034 6144 22040
rect 6460 22092 6868 22098
rect 6512 22086 6868 22092
rect 6460 22034 6512 22040
rect 6472 22003 6500 22034
rect 6840 22030 6868 22086
rect 7380 22092 7432 22098
rect 7380 22034 7432 22040
rect 6828 22024 6880 22030
rect 6828 21966 6880 21972
rect 5816 21888 5868 21894
rect 5816 21830 5868 21836
rect 6368 21888 6420 21894
rect 6368 21830 6420 21836
rect 6460 21888 6512 21894
rect 6460 21830 6512 21836
rect 6920 21888 6972 21894
rect 6920 21830 6972 21836
rect 7102 21856 7158 21865
rect 5724 21548 5776 21554
rect 5172 21490 5224 21496
rect 5724 21490 5776 21496
rect 4804 21480 4856 21486
rect 4856 21440 4936 21468
rect 4804 21422 4856 21428
rect 4712 20460 4764 20466
rect 4712 20402 4764 20408
rect 4620 20324 4672 20330
rect 4620 20266 4672 20272
rect 4724 19514 4752 20402
rect 4804 20256 4856 20262
rect 4804 20198 4856 20204
rect 4712 19508 4764 19514
rect 4712 19450 4764 19456
rect 4816 18766 4844 20198
rect 4804 18760 4856 18766
rect 4804 18702 4856 18708
rect 4620 18284 4672 18290
rect 4620 18226 4672 18232
rect 4528 17740 4580 17746
rect 4528 17682 4580 17688
rect 4436 17536 4488 17542
rect 4436 17478 4488 17484
rect 4528 17264 4580 17270
rect 4528 17206 4580 17212
rect 4344 17196 4396 17202
rect 4344 17138 4396 17144
rect 4252 16992 4304 16998
rect 4252 16934 4304 16940
rect 3749 16892 4057 16901
rect 3749 16890 3755 16892
rect 3811 16890 3835 16892
rect 3891 16890 3915 16892
rect 3971 16890 3995 16892
rect 4051 16890 4057 16892
rect 3811 16838 3813 16890
rect 3993 16838 3995 16890
rect 3749 16836 3755 16838
rect 3811 16836 3835 16838
rect 3891 16836 3915 16838
rect 3971 16836 3995 16838
rect 4051 16836 4057 16838
rect 3749 16827 4057 16836
rect 3976 16720 4028 16726
rect 3976 16662 4028 16668
rect 3700 16516 3752 16522
rect 3700 16458 3752 16464
rect 3608 16448 3660 16454
rect 3608 16390 3660 16396
rect 3712 16250 3740 16458
rect 2872 16244 2924 16250
rect 2872 16186 2924 16192
rect 3516 16244 3568 16250
rect 3516 16186 3568 16192
rect 3700 16244 3752 16250
rect 3700 16186 3752 16192
rect 3988 16046 4016 16662
rect 4264 16658 4292 16934
rect 4252 16652 4304 16658
rect 4252 16594 4304 16600
rect 4160 16448 4212 16454
rect 4160 16390 4212 16396
rect 3332 16040 3384 16046
rect 3332 15982 3384 15988
rect 3516 16040 3568 16046
rect 3516 15982 3568 15988
rect 3976 16040 4028 16046
rect 3976 15982 4028 15988
rect 2688 15564 2740 15570
rect 2688 15506 2740 15512
rect 3240 15496 3292 15502
rect 3238 15464 3240 15473
rect 3292 15464 3294 15473
rect 2608 15422 2728 15450
rect 2412 15360 2464 15366
rect 2412 15302 2464 15308
rect 2320 15156 2372 15162
rect 2320 15098 2372 15104
rect 2320 14952 2372 14958
rect 2320 14894 2372 14900
rect 2332 14618 2360 14894
rect 2424 14618 2452 15302
rect 2596 15020 2648 15026
rect 2596 14962 2648 14968
rect 2320 14612 2372 14618
rect 2320 14554 2372 14560
rect 2412 14612 2464 14618
rect 2412 14554 2464 14560
rect 2320 14408 2372 14414
rect 2320 14350 2372 14356
rect 2332 14074 2360 14350
rect 2320 14068 2372 14074
rect 2320 14010 2372 14016
rect 2228 13524 2280 13530
rect 2228 13466 2280 13472
rect 2148 13382 2268 13410
rect 2136 13184 2188 13190
rect 2136 13126 2188 13132
rect 1768 12436 1820 12442
rect 1768 12378 1820 12384
rect 1400 9580 1452 9586
rect 1400 9522 1452 9528
rect 1412 9217 1440 9522
rect 1398 9208 1454 9217
rect 1398 9143 1454 9152
rect 2044 8492 2096 8498
rect 2044 8434 2096 8440
rect 2056 8090 2084 8434
rect 2044 8084 2096 8090
rect 2044 8026 2096 8032
rect 2148 6730 2176 13126
rect 2240 12986 2268 13382
rect 2228 12980 2280 12986
rect 2228 12922 2280 12928
rect 2504 12096 2556 12102
rect 2504 12038 2556 12044
rect 2516 10266 2544 12038
rect 2608 11898 2636 14962
rect 2700 14890 2728 15422
rect 2780 15428 2832 15434
rect 3238 15399 3294 15408
rect 2780 15370 2832 15376
rect 2792 15162 2820 15370
rect 2872 15360 2924 15366
rect 2872 15302 2924 15308
rect 2780 15156 2832 15162
rect 2780 15098 2832 15104
rect 2688 14884 2740 14890
rect 2688 14826 2740 14832
rect 2688 14476 2740 14482
rect 2688 14418 2740 14424
rect 2700 13870 2728 14418
rect 2884 14414 2912 15302
rect 3344 15162 3372 15982
rect 3332 15156 3384 15162
rect 3332 15098 3384 15104
rect 3528 14958 3556 15982
rect 4172 15978 4200 16390
rect 4356 16114 4384 17138
rect 4436 17060 4488 17066
rect 4436 17002 4488 17008
rect 4448 16658 4476 17002
rect 4436 16652 4488 16658
rect 4436 16594 4488 16600
rect 4344 16108 4396 16114
rect 4344 16050 4396 16056
rect 4160 15972 4212 15978
rect 4160 15914 4212 15920
rect 3749 15804 4057 15813
rect 3749 15802 3755 15804
rect 3811 15802 3835 15804
rect 3891 15802 3915 15804
rect 3971 15802 3995 15804
rect 4051 15802 4057 15804
rect 3811 15750 3813 15802
rect 3993 15750 3995 15802
rect 3749 15748 3755 15750
rect 3811 15748 3835 15750
rect 3891 15748 3915 15750
rect 3971 15748 3995 15750
rect 4051 15748 4057 15750
rect 3749 15739 4057 15748
rect 4356 15706 4384 16050
rect 4344 15700 4396 15706
rect 4344 15642 4396 15648
rect 4068 15564 4120 15570
rect 4540 15552 4568 17206
rect 4120 15524 4568 15552
rect 4068 15506 4120 15512
rect 3608 15360 3660 15366
rect 3608 15302 3660 15308
rect 3516 14952 3568 14958
rect 3516 14894 3568 14900
rect 3424 14884 3476 14890
rect 3424 14826 3476 14832
rect 3148 14816 3200 14822
rect 3148 14758 3200 14764
rect 2964 14544 3016 14550
rect 2964 14486 3016 14492
rect 2872 14408 2924 14414
rect 2872 14350 2924 14356
rect 2688 13864 2740 13870
rect 2688 13806 2740 13812
rect 2700 13258 2728 13806
rect 2976 13326 3004 14486
rect 3160 13394 3188 14758
rect 3436 14550 3464 14826
rect 3424 14544 3476 14550
rect 3424 14486 3476 14492
rect 3528 14482 3556 14894
rect 3516 14476 3568 14482
rect 3516 14418 3568 14424
rect 3240 13456 3292 13462
rect 3240 13398 3292 13404
rect 3148 13388 3200 13394
rect 3148 13330 3200 13336
rect 2964 13320 3016 13326
rect 2964 13262 3016 13268
rect 2688 13252 2740 13258
rect 2688 13194 2740 13200
rect 3056 13184 3108 13190
rect 3056 13126 3108 13132
rect 2872 12844 2924 12850
rect 2872 12786 2924 12792
rect 2688 12708 2740 12714
rect 2688 12650 2740 12656
rect 2700 12306 2728 12650
rect 2780 12640 2832 12646
rect 2780 12582 2832 12588
rect 2688 12300 2740 12306
rect 2688 12242 2740 12248
rect 2596 11892 2648 11898
rect 2596 11834 2648 11840
rect 2792 11762 2820 12582
rect 2884 12442 2912 12786
rect 2964 12776 3016 12782
rect 2964 12718 3016 12724
rect 2872 12436 2924 12442
rect 2872 12378 2924 12384
rect 2872 12164 2924 12170
rect 2872 12106 2924 12112
rect 2780 11756 2832 11762
rect 2780 11698 2832 11704
rect 2884 10810 2912 12106
rect 2872 10804 2924 10810
rect 2872 10746 2924 10752
rect 2780 10668 2832 10674
rect 2780 10610 2832 10616
rect 2504 10260 2556 10266
rect 2504 10202 2556 10208
rect 2320 10056 2372 10062
rect 2320 9998 2372 10004
rect 2332 8362 2360 9998
rect 2412 9376 2464 9382
rect 2412 9318 2464 9324
rect 2424 8974 2452 9318
rect 2792 9178 2820 10610
rect 2976 10266 3004 12718
rect 3068 11898 3096 13126
rect 3252 12782 3280 13398
rect 3424 13252 3476 13258
rect 3424 13194 3476 13200
rect 3436 12782 3464 13194
rect 3620 12918 3648 15302
rect 4540 14958 4568 15524
rect 4528 14952 4580 14958
rect 4528 14894 4580 14900
rect 3749 14716 4057 14725
rect 3749 14714 3755 14716
rect 3811 14714 3835 14716
rect 3891 14714 3915 14716
rect 3971 14714 3995 14716
rect 4051 14714 4057 14716
rect 3811 14662 3813 14714
rect 3993 14662 3995 14714
rect 3749 14660 3755 14662
rect 3811 14660 3835 14662
rect 3891 14660 3915 14662
rect 3971 14660 3995 14662
rect 4051 14660 4057 14662
rect 3749 14651 4057 14660
rect 4632 14550 4660 18226
rect 4804 16244 4856 16250
rect 4804 16186 4856 16192
rect 4816 15502 4844 16186
rect 4804 15496 4856 15502
rect 4804 15438 4856 15444
rect 4712 15020 4764 15026
rect 4712 14962 4764 14968
rect 4620 14544 4672 14550
rect 4620 14486 4672 14492
rect 4724 14482 4752 14962
rect 4712 14476 4764 14482
rect 4712 14418 4764 14424
rect 4068 14408 4120 14414
rect 4120 14368 4200 14396
rect 4068 14350 4120 14356
rect 3884 14272 3936 14278
rect 3884 14214 3936 14220
rect 3896 14074 3924 14214
rect 4172 14074 4200 14368
rect 3884 14068 3936 14074
rect 3884 14010 3936 14016
rect 4160 14068 4212 14074
rect 4160 14010 4212 14016
rect 4724 13870 4752 14418
rect 4436 13864 4488 13870
rect 4434 13832 4436 13841
rect 4712 13864 4764 13870
rect 4488 13832 4490 13841
rect 4712 13806 4764 13812
rect 4434 13767 4490 13776
rect 3749 13628 4057 13637
rect 3749 13626 3755 13628
rect 3811 13626 3835 13628
rect 3891 13626 3915 13628
rect 3971 13626 3995 13628
rect 4051 13626 4057 13628
rect 3811 13574 3813 13626
rect 3993 13574 3995 13626
rect 3749 13572 3755 13574
rect 3811 13572 3835 13574
rect 3891 13572 3915 13574
rect 3971 13572 3995 13574
rect 4051 13572 4057 13574
rect 3749 13563 4057 13572
rect 4724 13326 4752 13806
rect 4908 13462 4936 21440
rect 5724 21344 5776 21350
rect 5724 21286 5776 21292
rect 5448 21004 5500 21010
rect 5448 20946 5500 20952
rect 5460 20806 5488 20946
rect 4988 20800 5040 20806
rect 4988 20742 5040 20748
rect 5356 20800 5408 20806
rect 5356 20742 5408 20748
rect 5448 20800 5500 20806
rect 5448 20742 5500 20748
rect 5000 20602 5028 20742
rect 5368 20602 5396 20742
rect 4988 20596 5040 20602
rect 4988 20538 5040 20544
rect 5356 20596 5408 20602
rect 5356 20538 5408 20544
rect 5172 19780 5224 19786
rect 5172 19722 5224 19728
rect 5080 19304 5132 19310
rect 5080 19246 5132 19252
rect 5092 18086 5120 19246
rect 5080 18080 5132 18086
rect 5080 18022 5132 18028
rect 5184 17338 5212 19722
rect 5356 18624 5408 18630
rect 5356 18566 5408 18572
rect 5368 18426 5396 18566
rect 5460 18426 5488 20742
rect 5632 19712 5684 19718
rect 5632 19654 5684 19660
rect 5540 19372 5592 19378
rect 5540 19314 5592 19320
rect 5356 18420 5408 18426
rect 5356 18362 5408 18368
rect 5448 18420 5500 18426
rect 5448 18362 5500 18368
rect 5552 17882 5580 19314
rect 5644 18970 5672 19654
rect 5632 18964 5684 18970
rect 5632 18906 5684 18912
rect 5540 17876 5592 17882
rect 5540 17818 5592 17824
rect 5172 17332 5224 17338
rect 5172 17274 5224 17280
rect 5172 16992 5224 16998
rect 5552 16980 5580 17818
rect 5224 16952 5580 16980
rect 5172 16934 5224 16940
rect 5736 16794 5764 21286
rect 4988 16788 5040 16794
rect 4988 16730 5040 16736
rect 5724 16788 5776 16794
rect 5724 16730 5776 16736
rect 4896 13456 4948 13462
rect 4896 13398 4948 13404
rect 4712 13320 4764 13326
rect 4712 13262 4764 13268
rect 4804 13184 4856 13190
rect 4804 13126 4856 13132
rect 3608 12912 3660 12918
rect 3608 12854 3660 12860
rect 3240 12776 3292 12782
rect 3240 12718 3292 12724
rect 3424 12776 3476 12782
rect 3424 12718 3476 12724
rect 3332 12096 3384 12102
rect 3332 12038 3384 12044
rect 3056 11892 3108 11898
rect 3056 11834 3108 11840
rect 3344 11762 3372 12038
rect 3332 11756 3384 11762
rect 3332 11698 3384 11704
rect 3436 11694 3464 12718
rect 3620 12306 3648 12854
rect 4252 12844 4304 12850
rect 4252 12786 4304 12792
rect 3749 12540 4057 12549
rect 3749 12538 3755 12540
rect 3811 12538 3835 12540
rect 3891 12538 3915 12540
rect 3971 12538 3995 12540
rect 4051 12538 4057 12540
rect 3811 12486 3813 12538
rect 3993 12486 3995 12538
rect 3749 12484 3755 12486
rect 3811 12484 3835 12486
rect 3891 12484 3915 12486
rect 3971 12484 3995 12486
rect 4051 12484 4057 12486
rect 3749 12475 4057 12484
rect 3608 12300 3660 12306
rect 3608 12242 3660 12248
rect 3516 12232 3568 12238
rect 3516 12174 3568 12180
rect 3424 11688 3476 11694
rect 3424 11630 3476 11636
rect 3528 11354 3556 12174
rect 3608 12096 3660 12102
rect 3608 12038 3660 12044
rect 4068 12096 4120 12102
rect 4068 12038 4120 12044
rect 3516 11348 3568 11354
rect 3516 11290 3568 11296
rect 3424 11280 3476 11286
rect 3424 11222 3476 11228
rect 3148 11008 3200 11014
rect 3148 10950 3200 10956
rect 3160 10810 3188 10950
rect 3148 10804 3200 10810
rect 3148 10746 3200 10752
rect 2964 10260 3016 10266
rect 2964 10202 3016 10208
rect 3436 10130 3464 11222
rect 3620 11150 3648 12038
rect 4080 11830 4108 12038
rect 4068 11824 4120 11830
rect 4068 11766 4120 11772
rect 3749 11452 4057 11461
rect 3749 11450 3755 11452
rect 3811 11450 3835 11452
rect 3891 11450 3915 11452
rect 3971 11450 3995 11452
rect 4051 11450 4057 11452
rect 3811 11398 3813 11450
rect 3993 11398 3995 11450
rect 3749 11396 3755 11398
rect 3811 11396 3835 11398
rect 3891 11396 3915 11398
rect 3971 11396 3995 11398
rect 4051 11396 4057 11398
rect 3749 11387 4057 11396
rect 4264 11354 4292 12786
rect 4816 12782 4844 13126
rect 4804 12776 4856 12782
rect 4804 12718 4856 12724
rect 4528 12708 4580 12714
rect 4528 12650 4580 12656
rect 4252 11348 4304 11354
rect 4252 11290 4304 11296
rect 3608 11144 3660 11150
rect 3608 11086 3660 11092
rect 4540 10606 4568 12650
rect 4816 12306 4844 12718
rect 4804 12300 4856 12306
rect 4804 12242 4856 12248
rect 4712 11756 4764 11762
rect 4712 11698 4764 11704
rect 4724 10606 4752 11698
rect 4816 11694 4844 12242
rect 4804 11688 4856 11694
rect 4804 11630 4856 11636
rect 4816 11218 4844 11630
rect 5000 11286 5028 16730
rect 5540 16516 5592 16522
rect 5540 16458 5592 16464
rect 5552 15910 5580 16458
rect 5724 16176 5776 16182
rect 5724 16118 5776 16124
rect 5540 15904 5592 15910
rect 5540 15846 5592 15852
rect 5736 15366 5764 16118
rect 5828 15638 5856 21830
rect 6380 21622 6408 21830
rect 6472 21690 6500 21830
rect 6548 21788 6856 21797
rect 6548 21786 6554 21788
rect 6610 21786 6634 21788
rect 6690 21786 6714 21788
rect 6770 21786 6794 21788
rect 6850 21786 6856 21788
rect 6610 21734 6612 21786
rect 6792 21734 6794 21786
rect 6548 21732 6554 21734
rect 6610 21732 6634 21734
rect 6690 21732 6714 21734
rect 6770 21732 6794 21734
rect 6850 21732 6856 21734
rect 6548 21723 6856 21732
rect 6460 21684 6512 21690
rect 6460 21626 6512 21632
rect 6368 21616 6420 21622
rect 6368 21558 6420 21564
rect 6092 21412 6144 21418
rect 6092 21354 6144 21360
rect 5908 19780 5960 19786
rect 5908 19722 5960 19728
rect 5920 18970 5948 19722
rect 6104 19174 6132 21354
rect 6276 21344 6328 21350
rect 6276 21286 6328 21292
rect 6184 20936 6236 20942
rect 6184 20878 6236 20884
rect 6196 20398 6224 20878
rect 6184 20392 6236 20398
rect 6184 20334 6236 20340
rect 6196 19854 6224 20334
rect 6184 19848 6236 19854
rect 6184 19790 6236 19796
rect 6196 19174 6224 19790
rect 6092 19168 6144 19174
rect 6092 19110 6144 19116
rect 6184 19168 6236 19174
rect 6184 19110 6236 19116
rect 5908 18964 5960 18970
rect 5908 18906 5960 18912
rect 6196 18766 6224 19110
rect 6184 18760 6236 18766
rect 6184 18702 6236 18708
rect 6196 18222 6224 18702
rect 6184 18216 6236 18222
rect 6184 18158 6236 18164
rect 6196 17678 6224 18158
rect 6184 17672 6236 17678
rect 6184 17614 6236 17620
rect 6000 17536 6052 17542
rect 6000 17478 6052 17484
rect 6012 16522 6040 17478
rect 6196 16998 6224 17614
rect 6288 17270 6316 21286
rect 6460 20868 6512 20874
rect 6460 20810 6512 20816
rect 6472 19718 6500 20810
rect 6548 20700 6856 20709
rect 6548 20698 6554 20700
rect 6610 20698 6634 20700
rect 6690 20698 6714 20700
rect 6770 20698 6794 20700
rect 6850 20698 6856 20700
rect 6610 20646 6612 20698
rect 6792 20646 6794 20698
rect 6548 20644 6554 20646
rect 6610 20644 6634 20646
rect 6690 20644 6714 20646
rect 6770 20644 6794 20646
rect 6850 20644 6856 20646
rect 6548 20635 6856 20644
rect 6828 20256 6880 20262
rect 6828 20198 6880 20204
rect 6840 19854 6868 20198
rect 6828 19848 6880 19854
rect 6828 19790 6880 19796
rect 6460 19712 6512 19718
rect 6460 19654 6512 19660
rect 6548 19612 6856 19621
rect 6548 19610 6554 19612
rect 6610 19610 6634 19612
rect 6690 19610 6714 19612
rect 6770 19610 6794 19612
rect 6850 19610 6856 19612
rect 6610 19558 6612 19610
rect 6792 19558 6794 19610
rect 6548 19556 6554 19558
rect 6610 19556 6634 19558
rect 6690 19556 6714 19558
rect 6770 19556 6794 19558
rect 6850 19556 6856 19558
rect 6548 19547 6856 19556
rect 6932 18698 6960 21830
rect 7102 21791 7158 21800
rect 7116 20466 7144 21791
rect 7380 21344 7432 21350
rect 7378 21312 7380 21321
rect 7484 21332 7512 22646
rect 7656 22160 7708 22166
rect 7656 22102 7708 22108
rect 7564 21888 7616 21894
rect 7564 21830 7616 21836
rect 7576 21622 7604 21830
rect 7564 21616 7616 21622
rect 7564 21558 7616 21564
rect 7668 21486 7696 22102
rect 8036 22030 8064 23800
rect 8680 22094 8708 23800
rect 9036 22772 9088 22778
rect 9036 22714 9088 22720
rect 9048 22094 9076 22714
rect 9324 22522 9352 23800
rect 9232 22494 9352 22522
rect 9128 22160 9180 22166
rect 9128 22102 9180 22108
rect 8496 22066 8708 22094
rect 8956 22066 9076 22094
rect 8496 22030 8524 22066
rect 8024 22024 8076 22030
rect 8024 21966 8076 21972
rect 8484 22024 8536 22030
rect 8484 21966 8536 21972
rect 7840 21888 7892 21894
rect 7840 21830 7892 21836
rect 7852 21690 7880 21830
rect 8390 21720 8446 21729
rect 7840 21684 7892 21690
rect 8496 21690 8524 21966
rect 8390 21655 8446 21664
rect 8484 21684 8536 21690
rect 7840 21626 7892 21632
rect 7656 21480 7708 21486
rect 7656 21422 7708 21428
rect 7840 21480 7892 21486
rect 8404 21434 8432 21655
rect 8484 21626 8536 21632
rect 7840 21422 7892 21428
rect 7432 21312 7512 21332
rect 7434 21304 7512 21312
rect 7378 21247 7434 21256
rect 7852 21146 7880 21422
rect 8312 21406 8432 21434
rect 8852 21480 8904 21486
rect 8852 21422 8904 21428
rect 7840 21140 7892 21146
rect 7840 21082 7892 21088
rect 8312 21010 8340 21406
rect 8392 21344 8444 21350
rect 8392 21286 8444 21292
rect 8484 21344 8536 21350
rect 8484 21286 8536 21292
rect 8404 21049 8432 21286
rect 8496 21078 8524 21286
rect 8484 21072 8536 21078
rect 8390 21040 8446 21049
rect 7288 21004 7340 21010
rect 7288 20946 7340 20952
rect 8300 21004 8352 21010
rect 8484 21014 8536 21020
rect 8668 21072 8720 21078
rect 8668 21014 8720 21020
rect 8390 20975 8446 20984
rect 8576 21004 8628 21010
rect 8300 20946 8352 20952
rect 8576 20946 8628 20952
rect 7196 20528 7248 20534
rect 7196 20470 7248 20476
rect 7104 20460 7156 20466
rect 7104 20402 7156 20408
rect 7208 19854 7236 20470
rect 7196 19848 7248 19854
rect 7196 19790 7248 19796
rect 6920 18692 6972 18698
rect 6920 18634 6972 18640
rect 6548 18524 6856 18533
rect 6548 18522 6554 18524
rect 6610 18522 6634 18524
rect 6690 18522 6714 18524
rect 6770 18522 6794 18524
rect 6850 18522 6856 18524
rect 6610 18470 6612 18522
rect 6792 18470 6794 18522
rect 6548 18468 6554 18470
rect 6610 18468 6634 18470
rect 6690 18468 6714 18470
rect 6770 18468 6794 18470
rect 6850 18468 6856 18470
rect 6548 18459 6856 18468
rect 7208 17882 7236 19790
rect 7300 19786 7328 20946
rect 7840 20936 7892 20942
rect 7840 20878 7892 20884
rect 7472 20800 7524 20806
rect 7472 20742 7524 20748
rect 7484 20602 7512 20742
rect 7472 20596 7524 20602
rect 7472 20538 7524 20544
rect 7748 20460 7800 20466
rect 7748 20402 7800 20408
rect 7288 19780 7340 19786
rect 7288 19722 7340 19728
rect 7760 19514 7788 20402
rect 7748 19508 7800 19514
rect 7748 19450 7800 19456
rect 7852 18426 7880 20878
rect 7932 20800 7984 20806
rect 7932 20742 7984 20748
rect 8300 20800 8352 20806
rect 8300 20742 8352 20748
rect 8484 20800 8536 20806
rect 8484 20742 8536 20748
rect 7944 20466 7972 20742
rect 7932 20460 7984 20466
rect 7932 20402 7984 20408
rect 8024 20392 8076 20398
rect 8312 20346 8340 20742
rect 8496 20602 8524 20742
rect 8484 20596 8536 20602
rect 8484 20538 8536 20544
rect 8024 20334 8076 20340
rect 8036 18970 8064 20334
rect 8128 20318 8340 20346
rect 8392 20392 8444 20398
rect 8392 20334 8444 20340
rect 8128 19310 8156 20318
rect 8404 19990 8432 20334
rect 8392 19984 8444 19990
rect 8392 19926 8444 19932
rect 8300 19712 8352 19718
rect 8300 19654 8352 19660
rect 8116 19304 8168 19310
rect 8116 19246 8168 19252
rect 8024 18964 8076 18970
rect 8024 18906 8076 18912
rect 8128 18630 8156 19246
rect 8312 18630 8340 19654
rect 8588 19514 8616 20946
rect 8576 19508 8628 19514
rect 8576 19450 8628 19456
rect 8680 19258 8708 21014
rect 8760 20800 8812 20806
rect 8760 20742 8812 20748
rect 8772 20262 8800 20742
rect 8864 20262 8892 21422
rect 8956 21350 8984 22066
rect 9036 21480 9088 21486
rect 9036 21422 9088 21428
rect 8944 21344 8996 21350
rect 8944 21286 8996 21292
rect 8944 20868 8996 20874
rect 8944 20810 8996 20816
rect 8956 20466 8984 20810
rect 8944 20460 8996 20466
rect 8944 20402 8996 20408
rect 8760 20256 8812 20262
rect 8760 20198 8812 20204
rect 8852 20256 8904 20262
rect 8852 20198 8904 20204
rect 8852 19848 8904 19854
rect 8852 19790 8904 19796
rect 8864 19378 8892 19790
rect 8852 19372 8904 19378
rect 8852 19314 8904 19320
rect 8680 19230 8892 19258
rect 8864 18698 8892 19230
rect 9048 18834 9076 21422
rect 9036 18828 9088 18834
rect 9036 18770 9088 18776
rect 8852 18692 8904 18698
rect 8852 18634 8904 18640
rect 8116 18624 8168 18630
rect 8116 18566 8168 18572
rect 8300 18624 8352 18630
rect 8300 18566 8352 18572
rect 7840 18420 7892 18426
rect 7840 18362 7892 18368
rect 7196 17876 7248 17882
rect 7196 17818 7248 17824
rect 6368 17604 6420 17610
rect 6368 17546 6420 17552
rect 6276 17264 6328 17270
rect 6276 17206 6328 17212
rect 6184 16992 6236 16998
rect 6184 16934 6236 16940
rect 6196 16522 6224 16934
rect 6000 16516 6052 16522
rect 6000 16458 6052 16464
rect 6184 16516 6236 16522
rect 6184 16458 6236 16464
rect 6090 16416 6146 16425
rect 6090 16351 6146 16360
rect 5816 15632 5868 15638
rect 5816 15574 5868 15580
rect 5724 15360 5776 15366
rect 5724 15302 5776 15308
rect 6000 14816 6052 14822
rect 6000 14758 6052 14764
rect 5816 14340 5868 14346
rect 5816 14282 5868 14288
rect 5908 14340 5960 14346
rect 5908 14282 5960 14288
rect 5828 14074 5856 14282
rect 5172 14068 5224 14074
rect 5172 14010 5224 14016
rect 5816 14068 5868 14074
rect 5816 14010 5868 14016
rect 5184 13326 5212 14010
rect 5630 13968 5686 13977
rect 5630 13903 5632 13912
rect 5684 13903 5686 13912
rect 5632 13874 5684 13880
rect 5172 13320 5224 13326
rect 5172 13262 5224 13268
rect 5920 12442 5948 14282
rect 6012 13462 6040 14758
rect 6000 13456 6052 13462
rect 6000 13398 6052 13404
rect 6104 13258 6132 16351
rect 6196 15910 6224 16458
rect 6276 16448 6328 16454
rect 6274 16416 6276 16425
rect 6328 16416 6330 16425
rect 6274 16351 6330 16360
rect 6184 15904 6236 15910
rect 6184 15846 6236 15852
rect 6196 15434 6224 15846
rect 6184 15428 6236 15434
rect 6184 15370 6236 15376
rect 6196 14822 6224 15370
rect 6276 15020 6328 15026
rect 6276 14962 6328 14968
rect 6184 14816 6236 14822
rect 6184 14758 6236 14764
rect 6196 14414 6224 14758
rect 6184 14408 6236 14414
rect 6184 14350 6236 14356
rect 6196 13870 6224 14350
rect 6184 13864 6236 13870
rect 6184 13806 6236 13812
rect 6196 13734 6224 13806
rect 6184 13728 6236 13734
rect 6184 13670 6236 13676
rect 6092 13252 6144 13258
rect 6092 13194 6144 13200
rect 6196 13190 6224 13670
rect 6288 13530 6316 14962
rect 6380 14550 6408 17546
rect 6548 17436 6856 17445
rect 6548 17434 6554 17436
rect 6610 17434 6634 17436
rect 6690 17434 6714 17436
rect 6770 17434 6794 17436
rect 6850 17434 6856 17436
rect 6610 17382 6612 17434
rect 6792 17382 6794 17434
rect 6548 17380 6554 17382
rect 6610 17380 6634 17382
rect 6690 17380 6714 17382
rect 6770 17380 6794 17382
rect 6850 17380 6856 17382
rect 6548 17371 6856 17380
rect 7852 16522 7880 18362
rect 8312 18290 8340 18566
rect 8300 18284 8352 18290
rect 8300 18226 8352 18232
rect 8312 17542 8340 18226
rect 8576 18080 8628 18086
rect 8576 18022 8628 18028
rect 8300 17536 8352 17542
rect 8300 17478 8352 17484
rect 8484 17536 8536 17542
rect 8484 17478 8536 17484
rect 8496 17134 8524 17478
rect 8588 17270 8616 18022
rect 8864 17338 8892 18634
rect 9048 17882 9076 18770
rect 9036 17876 9088 17882
rect 9036 17818 9088 17824
rect 8852 17332 8904 17338
rect 8852 17274 8904 17280
rect 9140 17270 9168 22102
rect 9232 22030 9260 22494
rect 9347 22332 9655 22341
rect 9347 22330 9353 22332
rect 9409 22330 9433 22332
rect 9489 22330 9513 22332
rect 9569 22330 9593 22332
rect 9649 22330 9655 22332
rect 9409 22278 9411 22330
rect 9591 22278 9593 22330
rect 9347 22276 9353 22278
rect 9409 22276 9433 22278
rect 9489 22276 9513 22278
rect 9569 22276 9593 22278
rect 9649 22276 9655 22278
rect 9347 22267 9655 22276
rect 9968 22030 9996 23800
rect 9220 22024 9272 22030
rect 9220 21966 9272 21972
rect 9956 22024 10008 22030
rect 9956 21966 10008 21972
rect 10232 22024 10284 22030
rect 10232 21966 10284 21972
rect 9220 21888 9272 21894
rect 9220 21830 9272 21836
rect 9496 21888 9548 21894
rect 9496 21830 9548 21836
rect 9772 21888 9824 21894
rect 10048 21888 10100 21894
rect 9772 21830 9824 21836
rect 10046 21856 10048 21865
rect 10100 21856 10102 21865
rect 9232 21729 9260 21830
rect 9218 21720 9274 21729
rect 9508 21690 9536 21830
rect 9218 21655 9274 21664
rect 9496 21684 9548 21690
rect 9496 21626 9548 21632
rect 9496 21548 9548 21554
rect 9548 21508 9720 21536
rect 9496 21490 9548 21496
rect 9220 21480 9272 21486
rect 9220 21422 9272 21428
rect 9232 20058 9260 21422
rect 9347 21244 9655 21253
rect 9347 21242 9353 21244
rect 9409 21242 9433 21244
rect 9489 21242 9513 21244
rect 9569 21242 9593 21244
rect 9649 21242 9655 21244
rect 9409 21190 9411 21242
rect 9591 21190 9593 21242
rect 9347 21188 9353 21190
rect 9409 21188 9433 21190
rect 9489 21188 9513 21190
rect 9569 21188 9593 21190
rect 9649 21188 9655 21190
rect 9347 21179 9655 21188
rect 9347 20156 9655 20165
rect 9347 20154 9353 20156
rect 9409 20154 9433 20156
rect 9489 20154 9513 20156
rect 9569 20154 9593 20156
rect 9649 20154 9655 20156
rect 9409 20102 9411 20154
rect 9591 20102 9593 20154
rect 9347 20100 9353 20102
rect 9409 20100 9433 20102
rect 9489 20100 9513 20102
rect 9569 20100 9593 20102
rect 9649 20100 9655 20102
rect 9347 20091 9655 20100
rect 9220 20052 9272 20058
rect 9220 19994 9272 20000
rect 9220 19916 9272 19922
rect 9220 19858 9272 19864
rect 9232 18086 9260 19858
rect 9494 19816 9550 19825
rect 9494 19751 9496 19760
rect 9548 19751 9550 19760
rect 9496 19722 9548 19728
rect 9508 19417 9536 19722
rect 9494 19408 9550 19417
rect 9494 19343 9550 19352
rect 9692 19242 9720 21508
rect 9784 21146 9812 21830
rect 10046 21791 10102 21800
rect 9864 21480 9916 21486
rect 9864 21422 9916 21428
rect 9772 21140 9824 21146
rect 9772 21082 9824 21088
rect 9876 21078 9904 21422
rect 10244 21146 10272 21966
rect 10612 21962 10640 23800
rect 11256 22094 11284 23800
rect 11900 22098 11928 23800
rect 11980 22840 12032 22846
rect 11980 22782 12032 22788
rect 11072 22066 11284 22094
rect 11888 22092 11940 22098
rect 11072 22030 11100 22066
rect 11888 22034 11940 22040
rect 11060 22024 11112 22030
rect 11520 22024 11572 22030
rect 11060 21966 11112 21972
rect 11242 21992 11298 22001
rect 10600 21956 10652 21962
rect 10600 21898 10652 21904
rect 10876 21888 10928 21894
rect 10876 21830 10928 21836
rect 10782 21720 10838 21729
rect 10782 21655 10838 21664
rect 10324 21480 10376 21486
rect 10324 21422 10376 21428
rect 10232 21140 10284 21146
rect 10232 21082 10284 21088
rect 9864 21072 9916 21078
rect 9864 21014 9916 21020
rect 10336 21010 10364 21422
rect 10508 21344 10560 21350
rect 10508 21286 10560 21292
rect 10324 21004 10376 21010
rect 10324 20946 10376 20952
rect 9956 20868 10008 20874
rect 9956 20810 10008 20816
rect 9772 20800 9824 20806
rect 9772 20742 9824 20748
rect 9784 20602 9812 20742
rect 9968 20602 9996 20810
rect 9772 20596 9824 20602
rect 9772 20538 9824 20544
rect 9956 20596 10008 20602
rect 9956 20538 10008 20544
rect 9784 19378 9812 20538
rect 10336 19718 10364 20946
rect 10520 20806 10548 21286
rect 10600 21004 10652 21010
rect 10600 20946 10652 20952
rect 10508 20800 10560 20806
rect 10508 20742 10560 20748
rect 10612 20466 10640 20946
rect 10692 20800 10744 20806
rect 10692 20742 10744 20748
rect 10704 20602 10732 20742
rect 10796 20618 10824 21655
rect 10888 21593 10916 21830
rect 10874 21584 10930 21593
rect 10874 21519 10930 21528
rect 10968 21548 11020 21554
rect 10968 21490 11020 21496
rect 10692 20596 10744 20602
rect 10796 20590 10916 20618
rect 10692 20538 10744 20544
rect 10600 20460 10652 20466
rect 10600 20402 10652 20408
rect 10612 19990 10640 20402
rect 10784 20392 10836 20398
rect 10784 20334 10836 20340
rect 10600 19984 10652 19990
rect 10600 19926 10652 19932
rect 9864 19712 9916 19718
rect 9864 19654 9916 19660
rect 10324 19712 10376 19718
rect 10324 19654 10376 19660
rect 9876 19378 9904 19654
rect 9772 19372 9824 19378
rect 9772 19314 9824 19320
rect 9864 19372 9916 19378
rect 9864 19314 9916 19320
rect 9680 19236 9732 19242
rect 9680 19178 9732 19184
rect 9347 19068 9655 19077
rect 9347 19066 9353 19068
rect 9409 19066 9433 19068
rect 9489 19066 9513 19068
rect 9569 19066 9593 19068
rect 9649 19066 9655 19068
rect 9409 19014 9411 19066
rect 9591 19014 9593 19066
rect 9347 19012 9353 19014
rect 9409 19012 9433 19014
rect 9489 19012 9513 19014
rect 9569 19012 9593 19014
rect 9649 19012 9655 19014
rect 9347 19003 9655 19012
rect 9588 18760 9640 18766
rect 9588 18702 9640 18708
rect 9600 18426 9628 18702
rect 9588 18420 9640 18426
rect 9692 18408 9720 19178
rect 9772 18420 9824 18426
rect 9692 18380 9772 18408
rect 9588 18362 9640 18368
rect 9772 18362 9824 18368
rect 9220 18080 9272 18086
rect 9220 18022 9272 18028
rect 9680 18080 9732 18086
rect 9680 18022 9732 18028
rect 9347 17980 9655 17989
rect 9347 17978 9353 17980
rect 9409 17978 9433 17980
rect 9489 17978 9513 17980
rect 9569 17978 9593 17980
rect 9649 17978 9655 17980
rect 9409 17926 9411 17978
rect 9591 17926 9593 17978
rect 9347 17924 9353 17926
rect 9409 17924 9433 17926
rect 9489 17924 9513 17926
rect 9569 17924 9593 17926
rect 9649 17924 9655 17926
rect 9347 17915 9655 17924
rect 9692 17864 9720 18022
rect 9600 17836 9720 17864
rect 8576 17264 8628 17270
rect 8576 17206 8628 17212
rect 8760 17264 8812 17270
rect 8760 17206 8812 17212
rect 9128 17264 9180 17270
rect 9128 17206 9180 17212
rect 8484 17128 8536 17134
rect 8484 17070 8536 17076
rect 8496 16658 8524 17070
rect 8772 16794 8800 17206
rect 9600 16980 9628 17836
rect 10796 17678 10824 20334
rect 10888 20058 10916 20590
rect 10876 20052 10928 20058
rect 10876 19994 10928 20000
rect 10876 19508 10928 19514
rect 10876 19450 10928 19456
rect 10888 18970 10916 19450
rect 10876 18964 10928 18970
rect 10876 18906 10928 18912
rect 10980 17882 11008 21490
rect 11072 20602 11100 21966
rect 11520 21966 11572 21972
rect 11242 21927 11298 21936
rect 11152 21888 11204 21894
rect 11152 21830 11204 21836
rect 11164 21418 11192 21830
rect 11152 21412 11204 21418
rect 11152 21354 11204 21360
rect 11150 20904 11206 20913
rect 11150 20839 11206 20848
rect 11060 20596 11112 20602
rect 11060 20538 11112 20544
rect 11164 20505 11192 20839
rect 11256 20777 11284 21927
rect 11532 21690 11560 21966
rect 11704 21888 11756 21894
rect 11704 21830 11756 21836
rect 11888 21888 11940 21894
rect 11888 21830 11940 21836
rect 11520 21684 11572 21690
rect 11520 21626 11572 21632
rect 11520 21548 11572 21554
rect 11520 21490 11572 21496
rect 11242 20768 11298 20777
rect 11242 20703 11298 20712
rect 11150 20496 11206 20505
rect 11150 20431 11206 20440
rect 11164 20058 11192 20431
rect 11152 20052 11204 20058
rect 11152 19994 11204 20000
rect 11256 19990 11284 20703
rect 11532 20262 11560 21490
rect 11716 21486 11744 21830
rect 11900 21622 11928 21830
rect 11888 21616 11940 21622
rect 11888 21558 11940 21564
rect 11796 21548 11848 21554
rect 11796 21490 11848 21496
rect 11704 21480 11756 21486
rect 11704 21422 11756 21428
rect 11808 20466 11836 21490
rect 11796 20460 11848 20466
rect 11796 20402 11848 20408
rect 11520 20256 11572 20262
rect 11520 20198 11572 20204
rect 11244 19984 11296 19990
rect 11244 19926 11296 19932
rect 11426 19816 11482 19825
rect 11426 19751 11428 19760
rect 11480 19751 11482 19760
rect 11428 19722 11480 19728
rect 11152 19712 11204 19718
rect 11152 19654 11204 19660
rect 11520 19712 11572 19718
rect 11520 19654 11572 19660
rect 11164 19174 11192 19654
rect 11532 19258 11560 19654
rect 11808 19553 11836 20402
rect 11992 20074 12020 22782
rect 12440 22094 12492 22098
rect 12544 22094 12572 23800
rect 12440 22092 12572 22094
rect 12492 22066 12572 22092
rect 12716 22092 12768 22098
rect 12440 22034 12492 22040
rect 12716 22034 12768 22040
rect 12532 22024 12584 22030
rect 12532 21966 12584 21972
rect 12072 21888 12124 21894
rect 12072 21830 12124 21836
rect 12084 21078 12112 21830
rect 12146 21788 12454 21797
rect 12146 21786 12152 21788
rect 12208 21786 12232 21788
rect 12288 21786 12312 21788
rect 12368 21786 12392 21788
rect 12448 21786 12454 21788
rect 12208 21734 12210 21786
rect 12390 21734 12392 21786
rect 12146 21732 12152 21734
rect 12208 21732 12232 21734
rect 12288 21732 12312 21734
rect 12368 21732 12392 21734
rect 12448 21732 12454 21734
rect 12146 21723 12454 21732
rect 12544 21690 12572 21966
rect 12532 21684 12584 21690
rect 12532 21626 12584 21632
rect 12728 21486 12756 22034
rect 13188 22030 13216 23800
rect 13832 22438 13860 23800
rect 14096 22500 14148 22506
rect 14096 22442 14148 22448
rect 13820 22432 13872 22438
rect 13820 22374 13872 22380
rect 13636 22160 13688 22166
rect 13636 22102 13688 22108
rect 13648 22030 13676 22102
rect 13176 22024 13228 22030
rect 13176 21966 13228 21972
rect 13636 22024 13688 22030
rect 13636 21966 13688 21972
rect 12900 21888 12952 21894
rect 12900 21830 12952 21836
rect 12992 21888 13044 21894
rect 13820 21888 13872 21894
rect 12992 21830 13044 21836
rect 13726 21856 13782 21865
rect 12716 21480 12768 21486
rect 12716 21422 12768 21428
rect 12912 21078 12940 21830
rect 12072 21072 12124 21078
rect 12072 21014 12124 21020
rect 12900 21072 12952 21078
rect 12900 21014 12952 21020
rect 12808 20936 12860 20942
rect 12808 20878 12860 20884
rect 12072 20868 12124 20874
rect 12072 20810 12124 20816
rect 11900 20046 12020 20074
rect 11900 19718 11928 20046
rect 11980 19984 12032 19990
rect 11978 19952 11980 19961
rect 12032 19952 12034 19961
rect 11978 19887 12034 19896
rect 11888 19712 11940 19718
rect 11888 19654 11940 19660
rect 11794 19544 11850 19553
rect 11612 19508 11664 19514
rect 11794 19479 11850 19488
rect 11612 19450 11664 19456
rect 11440 19230 11560 19258
rect 11152 19168 11204 19174
rect 11152 19110 11204 19116
rect 11164 18766 11192 19110
rect 11152 18760 11204 18766
rect 11152 18702 11204 18708
rect 10968 17876 11020 17882
rect 10968 17818 11020 17824
rect 10784 17672 10836 17678
rect 10784 17614 10836 17620
rect 10796 17338 10824 17614
rect 10784 17332 10836 17338
rect 10784 17274 10836 17280
rect 10980 17270 11008 17818
rect 10968 17264 11020 17270
rect 10968 17206 11020 17212
rect 11336 17264 11388 17270
rect 11336 17206 11388 17212
rect 10508 17196 10560 17202
rect 10508 17138 10560 17144
rect 9772 17128 9824 17134
rect 9772 17070 9824 17076
rect 9600 16952 9720 16980
rect 9347 16892 9655 16901
rect 9347 16890 9353 16892
rect 9409 16890 9433 16892
rect 9489 16890 9513 16892
rect 9569 16890 9593 16892
rect 9649 16890 9655 16892
rect 9409 16838 9411 16890
rect 9591 16838 9593 16890
rect 9347 16836 9353 16838
rect 9409 16836 9433 16838
rect 9489 16836 9513 16838
rect 9569 16836 9593 16838
rect 9649 16836 9655 16838
rect 9347 16827 9655 16836
rect 8760 16788 8812 16794
rect 8760 16730 8812 16736
rect 9692 16674 9720 16952
rect 8484 16652 8536 16658
rect 8484 16594 8536 16600
rect 9600 16646 9720 16674
rect 7840 16516 7892 16522
rect 7840 16458 7892 16464
rect 6548 16348 6856 16357
rect 6548 16346 6554 16348
rect 6610 16346 6634 16348
rect 6690 16346 6714 16348
rect 6770 16346 6794 16348
rect 6850 16346 6856 16348
rect 6610 16294 6612 16346
rect 6792 16294 6794 16346
rect 6548 16292 6554 16294
rect 6610 16292 6634 16294
rect 6690 16292 6714 16294
rect 6770 16292 6794 16294
rect 6850 16292 6856 16294
rect 6548 16283 6856 16292
rect 9600 16250 9628 16646
rect 9784 16590 9812 17070
rect 9772 16584 9824 16590
rect 9772 16526 9824 16532
rect 9588 16244 9640 16250
rect 9588 16186 9640 16192
rect 9784 16114 9812 16526
rect 9864 16244 9916 16250
rect 9864 16186 9916 16192
rect 9772 16108 9824 16114
rect 9772 16050 9824 16056
rect 8392 15904 8444 15910
rect 8392 15846 8444 15852
rect 8404 15434 8432 15846
rect 9347 15804 9655 15813
rect 9347 15802 9353 15804
rect 9409 15802 9433 15804
rect 9489 15802 9513 15804
rect 9569 15802 9593 15804
rect 9649 15802 9655 15804
rect 9409 15750 9411 15802
rect 9591 15750 9593 15802
rect 9347 15748 9353 15750
rect 9409 15748 9433 15750
rect 9489 15748 9513 15750
rect 9569 15748 9593 15750
rect 9649 15748 9655 15750
rect 9347 15739 9655 15748
rect 9876 15502 9904 16186
rect 10520 15706 10548 17138
rect 11060 16516 11112 16522
rect 11060 16458 11112 16464
rect 10508 15700 10560 15706
rect 10508 15642 10560 15648
rect 9864 15496 9916 15502
rect 8666 15464 8722 15473
rect 6460 15428 6512 15434
rect 6460 15370 6512 15376
rect 8392 15428 8444 15434
rect 9864 15438 9916 15444
rect 8666 15399 8722 15408
rect 8392 15370 8444 15376
rect 6472 15162 6500 15370
rect 8680 15366 8708 15399
rect 8668 15360 8720 15366
rect 8668 15302 8720 15308
rect 6548 15260 6856 15269
rect 6548 15258 6554 15260
rect 6610 15258 6634 15260
rect 6690 15258 6714 15260
rect 6770 15258 6794 15260
rect 6850 15258 6856 15260
rect 6610 15206 6612 15258
rect 6792 15206 6794 15258
rect 6548 15204 6554 15206
rect 6610 15204 6634 15206
rect 6690 15204 6714 15206
rect 6770 15204 6794 15206
rect 6850 15204 6856 15206
rect 6548 15195 6856 15204
rect 6460 15156 6512 15162
rect 6460 15098 6512 15104
rect 8680 15094 8708 15302
rect 10520 15094 10548 15642
rect 11072 15366 11100 16458
rect 11244 16448 11296 16454
rect 11244 16390 11296 16396
rect 11152 16108 11204 16114
rect 11256 16096 11284 16390
rect 11204 16068 11284 16096
rect 11152 16050 11204 16056
rect 11060 15360 11112 15366
rect 11060 15302 11112 15308
rect 11348 15162 11376 17206
rect 11336 15156 11388 15162
rect 11336 15098 11388 15104
rect 8668 15088 8720 15094
rect 8668 15030 8720 15036
rect 10508 15088 10560 15094
rect 10508 15030 10560 15036
rect 6460 15020 6512 15026
rect 6460 14962 6512 14968
rect 6368 14544 6420 14550
rect 6368 14486 6420 14492
rect 6380 14278 6408 14486
rect 6368 14272 6420 14278
rect 6368 14214 6420 14220
rect 6472 13954 6500 14962
rect 9864 14952 9916 14958
rect 9864 14894 9916 14900
rect 9772 14816 9824 14822
rect 9772 14758 9824 14764
rect 9347 14716 9655 14725
rect 9347 14714 9353 14716
rect 9409 14714 9433 14716
rect 9489 14714 9513 14716
rect 9569 14714 9593 14716
rect 9649 14714 9655 14716
rect 9409 14662 9411 14714
rect 9591 14662 9593 14714
rect 9347 14660 9353 14662
rect 9409 14660 9433 14662
rect 9489 14660 9513 14662
rect 9569 14660 9593 14662
rect 9649 14660 9655 14662
rect 9347 14651 9655 14660
rect 8484 14612 8536 14618
rect 8484 14554 8536 14560
rect 7472 14340 7524 14346
rect 7472 14282 7524 14288
rect 6548 14172 6856 14181
rect 6548 14170 6554 14172
rect 6610 14170 6634 14172
rect 6690 14170 6714 14172
rect 6770 14170 6794 14172
rect 6850 14170 6856 14172
rect 6610 14118 6612 14170
rect 6792 14118 6794 14170
rect 6548 14116 6554 14118
rect 6610 14116 6634 14118
rect 6690 14116 6714 14118
rect 6770 14116 6794 14118
rect 6850 14116 6856 14118
rect 6548 14107 6856 14116
rect 6552 14000 6604 14006
rect 6380 13938 6500 13954
rect 6368 13932 6500 13938
rect 6420 13926 6500 13932
rect 6368 13874 6420 13880
rect 6472 13870 6500 13926
rect 6550 13968 6552 13977
rect 6604 13968 6606 13977
rect 7484 13938 7512 14282
rect 8496 14074 8524 14554
rect 9680 14272 9732 14278
rect 9680 14214 9732 14220
rect 8484 14068 8536 14074
rect 8484 14010 8536 14016
rect 6550 13903 6606 13912
rect 7472 13932 7524 13938
rect 7472 13874 7524 13880
rect 7840 13932 7892 13938
rect 7840 13874 7892 13880
rect 6460 13864 6512 13870
rect 6460 13806 6512 13812
rect 7852 13530 7880 13874
rect 8390 13832 8446 13841
rect 8390 13767 8446 13776
rect 8404 13734 8432 13767
rect 8392 13728 8444 13734
rect 8392 13670 8444 13676
rect 6276 13524 6328 13530
rect 6276 13466 6328 13472
rect 7840 13524 7892 13530
rect 7840 13466 7892 13472
rect 6184 13184 6236 13190
rect 6184 13126 6236 13132
rect 6196 12986 6224 13126
rect 6548 13084 6856 13093
rect 6548 13082 6554 13084
rect 6610 13082 6634 13084
rect 6690 13082 6714 13084
rect 6770 13082 6794 13084
rect 6850 13082 6856 13084
rect 6610 13030 6612 13082
rect 6792 13030 6794 13082
rect 6548 13028 6554 13030
rect 6610 13028 6634 13030
rect 6690 13028 6714 13030
rect 6770 13028 6794 13030
rect 6850 13028 6856 13030
rect 6548 13019 6856 13028
rect 8404 12986 8432 13670
rect 8496 13258 8524 14010
rect 9347 13628 9655 13637
rect 9347 13626 9353 13628
rect 9409 13626 9433 13628
rect 9489 13626 9513 13628
rect 9569 13626 9593 13628
rect 9649 13626 9655 13628
rect 9409 13574 9411 13626
rect 9591 13574 9593 13626
rect 9347 13572 9353 13574
rect 9409 13572 9433 13574
rect 9489 13572 9513 13574
rect 9569 13572 9593 13574
rect 9649 13572 9655 13574
rect 9347 13563 9655 13572
rect 9692 13530 9720 14214
rect 9784 14006 9812 14758
rect 9876 14278 9904 14894
rect 10968 14884 11020 14890
rect 10968 14826 11020 14832
rect 9956 14340 10008 14346
rect 9956 14282 10008 14288
rect 9864 14272 9916 14278
rect 9864 14214 9916 14220
rect 9772 14000 9824 14006
rect 9772 13942 9824 13948
rect 9876 13870 9904 14214
rect 9968 14074 9996 14282
rect 10980 14278 11008 14826
rect 10968 14272 11020 14278
rect 10968 14214 11020 14220
rect 9956 14068 10008 14074
rect 9956 14010 10008 14016
rect 10980 14006 11008 14214
rect 11244 14068 11296 14074
rect 11244 14010 11296 14016
rect 10968 14000 11020 14006
rect 10968 13942 11020 13948
rect 9864 13864 9916 13870
rect 9864 13806 9916 13812
rect 9680 13524 9732 13530
rect 9680 13466 9732 13472
rect 8484 13252 8536 13258
rect 8484 13194 8536 13200
rect 6184 12980 6236 12986
rect 6184 12922 6236 12928
rect 6368 12980 6420 12986
rect 6368 12922 6420 12928
rect 8392 12980 8444 12986
rect 8392 12922 8444 12928
rect 6276 12912 6328 12918
rect 6276 12854 6328 12860
rect 5908 12436 5960 12442
rect 5908 12378 5960 12384
rect 5264 12164 5316 12170
rect 5264 12106 5316 12112
rect 6184 12164 6236 12170
rect 6184 12106 6236 12112
rect 5276 11354 5304 12106
rect 5908 11756 5960 11762
rect 5908 11698 5960 11704
rect 5816 11552 5868 11558
rect 5816 11494 5868 11500
rect 5264 11348 5316 11354
rect 5264 11290 5316 11296
rect 4988 11280 5040 11286
rect 4988 11222 5040 11228
rect 4804 11212 4856 11218
rect 4804 11154 4856 11160
rect 5540 11076 5592 11082
rect 5540 11018 5592 11024
rect 5552 10810 5580 11018
rect 5540 10804 5592 10810
rect 5540 10746 5592 10752
rect 5448 10668 5500 10674
rect 5448 10610 5500 10616
rect 4528 10600 4580 10606
rect 4528 10542 4580 10548
rect 4712 10600 4764 10606
rect 4712 10542 4764 10548
rect 3749 10364 4057 10373
rect 3749 10362 3755 10364
rect 3811 10362 3835 10364
rect 3891 10362 3915 10364
rect 3971 10362 3995 10364
rect 4051 10362 4057 10364
rect 3811 10310 3813 10362
rect 3993 10310 3995 10362
rect 3749 10308 3755 10310
rect 3811 10308 3835 10310
rect 3891 10308 3915 10310
rect 3971 10308 3995 10310
rect 4051 10308 4057 10310
rect 3749 10299 4057 10308
rect 4540 10130 4568 10542
rect 4724 10198 4752 10542
rect 4712 10192 4764 10198
rect 4712 10134 4764 10140
rect 3056 10124 3108 10130
rect 3056 10066 3108 10072
rect 3424 10124 3476 10130
rect 3424 10066 3476 10072
rect 4528 10124 4580 10130
rect 4528 10066 4580 10072
rect 2872 9920 2924 9926
rect 2872 9862 2924 9868
rect 2780 9172 2832 9178
rect 2780 9114 2832 9120
rect 2884 9110 2912 9862
rect 2872 9104 2924 9110
rect 2872 9046 2924 9052
rect 3068 9042 3096 10066
rect 4540 9722 4568 10066
rect 4712 10056 4764 10062
rect 4896 10056 4948 10062
rect 4764 10016 4896 10044
rect 4712 9998 4764 10004
rect 4896 9998 4948 10004
rect 4712 9920 4764 9926
rect 4712 9862 4764 9868
rect 4528 9716 4580 9722
rect 4528 9658 4580 9664
rect 3160 9586 3924 9602
rect 3148 9580 3936 9586
rect 3200 9574 3884 9580
rect 3148 9522 3200 9528
rect 3884 9522 3936 9528
rect 3240 9512 3292 9518
rect 3240 9454 3292 9460
rect 3148 9444 3200 9450
rect 3148 9386 3200 9392
rect 3160 9110 3188 9386
rect 3252 9194 3280 9454
rect 4436 9376 4488 9382
rect 4436 9318 4488 9324
rect 3749 9276 4057 9285
rect 3749 9274 3755 9276
rect 3811 9274 3835 9276
rect 3891 9274 3915 9276
rect 3971 9274 3995 9276
rect 4051 9274 4057 9276
rect 3811 9222 3813 9274
rect 3993 9222 3995 9274
rect 3749 9220 3755 9222
rect 3811 9220 3835 9222
rect 3891 9220 3915 9222
rect 3971 9220 3995 9222
rect 4051 9220 4057 9222
rect 3749 9211 4057 9220
rect 3252 9166 3372 9194
rect 3148 9104 3200 9110
rect 3148 9046 3200 9052
rect 3056 9036 3108 9042
rect 3056 8978 3108 8984
rect 3240 9036 3292 9042
rect 3240 8978 3292 8984
rect 2412 8968 2464 8974
rect 2412 8910 2464 8916
rect 2872 8900 2924 8906
rect 2872 8842 2924 8848
rect 2320 8356 2372 8362
rect 2320 8298 2372 8304
rect 2884 8090 2912 8842
rect 2964 8560 3016 8566
rect 2962 8528 2964 8537
rect 3016 8528 3018 8537
rect 2962 8463 3018 8472
rect 3068 8430 3096 8978
rect 3252 8430 3280 8978
rect 3344 8634 3372 9166
rect 3516 9104 3568 9110
rect 3516 9046 3568 9052
rect 3332 8628 3384 8634
rect 3332 8570 3384 8576
rect 3056 8424 3108 8430
rect 3056 8366 3108 8372
rect 3240 8424 3292 8430
rect 3240 8366 3292 8372
rect 2872 8084 2924 8090
rect 2872 8026 2924 8032
rect 3252 7954 3280 8366
rect 3344 7970 3372 8570
rect 3240 7948 3292 7954
rect 3344 7942 3464 7970
rect 3240 7890 3292 7896
rect 3148 7880 3200 7886
rect 3148 7822 3200 7828
rect 3332 7880 3384 7886
rect 3332 7822 3384 7828
rect 2412 7744 2464 7750
rect 2412 7686 2464 7692
rect 2424 7206 2452 7686
rect 3160 7478 3188 7822
rect 3148 7472 3200 7478
rect 3148 7414 3200 7420
rect 3344 7410 3372 7822
rect 3436 7818 3464 7942
rect 3528 7818 3556 9046
rect 4448 8906 4476 9318
rect 4724 9178 4752 9862
rect 5460 9178 5488 10610
rect 5828 9994 5856 11494
rect 5920 11150 5948 11698
rect 5908 11144 5960 11150
rect 5908 11086 5960 11092
rect 6196 10810 6224 12106
rect 6288 12102 6316 12854
rect 6380 12850 6408 12922
rect 9876 12918 9904 13806
rect 10980 13530 11008 13942
rect 10968 13524 11020 13530
rect 10968 13466 11020 13472
rect 10324 13184 10376 13190
rect 10324 13126 10376 13132
rect 9864 12912 9916 12918
rect 9864 12854 9916 12860
rect 6368 12844 6420 12850
rect 6368 12786 6420 12792
rect 6380 12238 6408 12786
rect 9876 12782 9904 12854
rect 10336 12850 10364 13126
rect 10324 12844 10376 12850
rect 10324 12786 10376 12792
rect 11060 12844 11112 12850
rect 11060 12786 11112 12792
rect 9864 12776 9916 12782
rect 9864 12718 9916 12724
rect 8484 12708 8536 12714
rect 8484 12650 8536 12656
rect 6368 12232 6420 12238
rect 6368 12174 6420 12180
rect 6276 12096 6328 12102
rect 6276 12038 6328 12044
rect 6380 11898 6408 12174
rect 6460 12096 6512 12102
rect 6460 12038 6512 12044
rect 7840 12096 7892 12102
rect 7840 12038 7892 12044
rect 6368 11892 6420 11898
rect 6368 11834 6420 11840
rect 6380 10810 6408 11834
rect 6184 10804 6236 10810
rect 6184 10746 6236 10752
rect 6368 10804 6420 10810
rect 6368 10746 6420 10752
rect 6380 10266 6408 10746
rect 6472 10742 6500 12038
rect 6548 11996 6856 12005
rect 6548 11994 6554 11996
rect 6610 11994 6634 11996
rect 6690 11994 6714 11996
rect 6770 11994 6794 11996
rect 6850 11994 6856 11996
rect 6610 11942 6612 11994
rect 6792 11942 6794 11994
rect 6548 11940 6554 11942
rect 6610 11940 6634 11942
rect 6690 11940 6714 11942
rect 6770 11940 6794 11942
rect 6850 11940 6856 11942
rect 6548 11931 6856 11940
rect 7852 11762 7880 12038
rect 7840 11756 7892 11762
rect 7840 11698 7892 11704
rect 6828 11688 6880 11694
rect 6828 11630 6880 11636
rect 6840 11150 6868 11630
rect 6828 11144 6880 11150
rect 6828 11086 6880 11092
rect 8024 11076 8076 11082
rect 8024 11018 8076 11024
rect 6548 10908 6856 10917
rect 6548 10906 6554 10908
rect 6610 10906 6634 10908
rect 6690 10906 6714 10908
rect 6770 10906 6794 10908
rect 6850 10906 6856 10908
rect 6610 10854 6612 10906
rect 6792 10854 6794 10906
rect 6548 10852 6554 10854
rect 6610 10852 6634 10854
rect 6690 10852 6714 10854
rect 6770 10852 6794 10854
rect 6850 10852 6856 10854
rect 6548 10843 6856 10852
rect 6460 10736 6512 10742
rect 6460 10678 6512 10684
rect 8036 10470 8064 11018
rect 8392 11008 8444 11014
rect 8392 10950 8444 10956
rect 8404 10606 8432 10950
rect 8496 10742 8524 12650
rect 9680 12640 9732 12646
rect 9680 12582 9732 12588
rect 9347 12540 9655 12549
rect 9347 12538 9353 12540
rect 9409 12538 9433 12540
rect 9489 12538 9513 12540
rect 9569 12538 9593 12540
rect 9649 12538 9655 12540
rect 9409 12486 9411 12538
rect 9591 12486 9593 12538
rect 9347 12484 9353 12486
rect 9409 12484 9433 12486
rect 9489 12484 9513 12486
rect 9569 12484 9593 12486
rect 9649 12484 9655 12486
rect 9347 12475 9655 12484
rect 9692 12306 9720 12582
rect 9680 12300 9732 12306
rect 9680 12242 9732 12248
rect 9876 12238 9904 12718
rect 9864 12232 9916 12238
rect 9864 12174 9916 12180
rect 9312 12164 9364 12170
rect 9312 12106 9364 12112
rect 10324 12164 10376 12170
rect 10324 12106 10376 12112
rect 9324 11762 9352 12106
rect 9036 11756 9088 11762
rect 9036 11698 9088 11704
rect 9312 11756 9364 11762
rect 9312 11698 9364 11704
rect 9048 11354 9076 11698
rect 9347 11452 9655 11461
rect 9347 11450 9353 11452
rect 9409 11450 9433 11452
rect 9489 11450 9513 11452
rect 9569 11450 9593 11452
rect 9649 11450 9655 11452
rect 9409 11398 9411 11450
rect 9591 11398 9593 11450
rect 9347 11396 9353 11398
rect 9409 11396 9433 11398
rect 9489 11396 9513 11398
rect 9569 11396 9593 11398
rect 9649 11396 9655 11398
rect 9347 11387 9655 11396
rect 9036 11348 9088 11354
rect 9036 11290 9088 11296
rect 10048 11348 10100 11354
rect 10048 11290 10100 11296
rect 9956 11076 10008 11082
rect 9956 11018 10008 11024
rect 8484 10736 8536 10742
rect 8484 10678 8536 10684
rect 8852 10668 8904 10674
rect 8852 10610 8904 10616
rect 8392 10600 8444 10606
rect 8392 10542 8444 10548
rect 6460 10464 6512 10470
rect 6460 10406 6512 10412
rect 8024 10464 8076 10470
rect 8024 10406 8076 10412
rect 6368 10260 6420 10266
rect 6368 10202 6420 10208
rect 5816 9988 5868 9994
rect 5816 9930 5868 9936
rect 6380 9722 6408 10202
rect 6472 10010 6500 10406
rect 6472 9982 6592 10010
rect 6368 9716 6420 9722
rect 6368 9658 6420 9664
rect 4712 9172 4764 9178
rect 4712 9114 4764 9120
rect 5448 9172 5500 9178
rect 5448 9114 5500 9120
rect 6472 8906 6500 9982
rect 6564 9926 6592 9982
rect 7104 9988 7156 9994
rect 7104 9930 7156 9936
rect 6552 9920 6604 9926
rect 6552 9862 6604 9868
rect 6548 9820 6856 9829
rect 6548 9818 6554 9820
rect 6610 9818 6634 9820
rect 6690 9818 6714 9820
rect 6770 9818 6794 9820
rect 6850 9818 6856 9820
rect 6610 9766 6612 9818
rect 6792 9766 6794 9818
rect 6548 9764 6554 9766
rect 6610 9764 6634 9766
rect 6690 9764 6714 9766
rect 6770 9764 6794 9766
rect 6850 9764 6856 9766
rect 6548 9755 6856 9764
rect 6644 9716 6696 9722
rect 6644 9658 6696 9664
rect 6656 9586 6684 9658
rect 6644 9580 6696 9586
rect 6644 9522 6696 9528
rect 6656 9178 6684 9522
rect 6920 9512 6972 9518
rect 6920 9454 6972 9460
rect 6644 9172 6696 9178
rect 6644 9114 6696 9120
rect 4344 8900 4396 8906
rect 4344 8842 4396 8848
rect 4436 8900 4488 8906
rect 4436 8842 4488 8848
rect 6460 8900 6512 8906
rect 6460 8842 6512 8848
rect 3749 8188 4057 8197
rect 3749 8186 3755 8188
rect 3811 8186 3835 8188
rect 3891 8186 3915 8188
rect 3971 8186 3995 8188
rect 4051 8186 4057 8188
rect 3811 8134 3813 8186
rect 3993 8134 3995 8186
rect 3749 8132 3755 8134
rect 3811 8132 3835 8134
rect 3891 8132 3915 8134
rect 3971 8132 3995 8134
rect 4051 8132 4057 8134
rect 3749 8123 4057 8132
rect 3424 7812 3476 7818
rect 3424 7754 3476 7760
rect 3516 7812 3568 7818
rect 3516 7754 3568 7760
rect 4356 7546 4384 8842
rect 4448 8294 4476 8842
rect 5540 8832 5592 8838
rect 5540 8774 5592 8780
rect 4804 8560 4856 8566
rect 4804 8502 4856 8508
rect 4894 8528 4950 8537
rect 4436 8288 4488 8294
rect 4436 8230 4488 8236
rect 4448 7886 4476 8230
rect 4436 7880 4488 7886
rect 4436 7822 4488 7828
rect 4816 7750 4844 8502
rect 4894 8463 4896 8472
rect 4948 8463 4950 8472
rect 4896 8434 4948 8440
rect 4804 7744 4856 7750
rect 4804 7686 4856 7692
rect 4344 7540 4396 7546
rect 4344 7482 4396 7488
rect 3332 7404 3384 7410
rect 3332 7346 3384 7352
rect 2412 7200 2464 7206
rect 2412 7142 2464 7148
rect 3344 7002 3372 7346
rect 3749 7100 4057 7109
rect 3749 7098 3755 7100
rect 3811 7098 3835 7100
rect 3891 7098 3915 7100
rect 3971 7098 3995 7100
rect 4051 7098 4057 7100
rect 3811 7046 3813 7098
rect 3993 7046 3995 7098
rect 3749 7044 3755 7046
rect 3811 7044 3835 7046
rect 3891 7044 3915 7046
rect 3971 7044 3995 7046
rect 4051 7044 4057 7046
rect 3749 7035 4057 7044
rect 3332 6996 3384 7002
rect 3332 6938 3384 6944
rect 2136 6724 2188 6730
rect 2136 6666 2188 6672
rect 4816 6458 4844 7686
rect 5552 7478 5580 8774
rect 6548 8732 6856 8741
rect 6548 8730 6554 8732
rect 6610 8730 6634 8732
rect 6690 8730 6714 8732
rect 6770 8730 6794 8732
rect 6850 8730 6856 8732
rect 6610 8678 6612 8730
rect 6792 8678 6794 8730
rect 6548 8676 6554 8678
rect 6610 8676 6634 8678
rect 6690 8676 6714 8678
rect 6770 8676 6794 8678
rect 6850 8676 6856 8678
rect 6548 8667 6856 8676
rect 6184 8628 6236 8634
rect 6184 8570 6236 8576
rect 5816 8492 5868 8498
rect 5816 8434 5868 8440
rect 5828 8090 5856 8434
rect 6000 8356 6052 8362
rect 6000 8298 6052 8304
rect 5816 8084 5868 8090
rect 5816 8026 5868 8032
rect 6012 7886 6040 8298
rect 6000 7880 6052 7886
rect 6000 7822 6052 7828
rect 5540 7472 5592 7478
rect 5540 7414 5592 7420
rect 6012 7426 6040 7822
rect 6012 7410 6132 7426
rect 5080 7404 5132 7410
rect 6012 7404 6144 7410
rect 6012 7398 6092 7404
rect 5080 7346 5132 7352
rect 6092 7346 6144 7352
rect 5092 7002 5120 7346
rect 5908 7200 5960 7206
rect 5908 7142 5960 7148
rect 5080 6996 5132 7002
rect 5080 6938 5132 6944
rect 4804 6452 4856 6458
rect 4804 6394 4856 6400
rect 5920 6390 5948 7142
rect 6196 6798 6224 8570
rect 6932 8090 6960 9454
rect 7116 9382 7144 9930
rect 8404 9926 8432 10542
rect 8864 10266 8892 10610
rect 9968 10470 9996 11018
rect 9956 10464 10008 10470
rect 9956 10406 10008 10412
rect 9347 10364 9655 10373
rect 9347 10362 9353 10364
rect 9409 10362 9433 10364
rect 9489 10362 9513 10364
rect 9569 10362 9593 10364
rect 9649 10362 9655 10364
rect 9409 10310 9411 10362
rect 9591 10310 9593 10362
rect 9347 10308 9353 10310
rect 9409 10308 9433 10310
rect 9489 10308 9513 10310
rect 9569 10308 9593 10310
rect 9649 10308 9655 10310
rect 9347 10299 9655 10308
rect 8852 10260 8904 10266
rect 8852 10202 8904 10208
rect 8392 9920 8444 9926
rect 8392 9862 8444 9868
rect 8576 9920 8628 9926
rect 8576 9862 8628 9868
rect 7104 9376 7156 9382
rect 7104 9318 7156 9324
rect 7472 9376 7524 9382
rect 7472 9318 7524 9324
rect 7484 8974 7512 9318
rect 8404 9178 8432 9862
rect 8392 9172 8444 9178
rect 8392 9114 8444 9120
rect 7472 8968 7524 8974
rect 7472 8910 7524 8916
rect 8300 8560 8352 8566
rect 8300 8502 8352 8508
rect 7012 8288 7064 8294
rect 7012 8230 7064 8236
rect 6920 8084 6972 8090
rect 6920 8026 6972 8032
rect 6548 7644 6856 7653
rect 6548 7642 6554 7644
rect 6610 7642 6634 7644
rect 6690 7642 6714 7644
rect 6770 7642 6794 7644
rect 6850 7642 6856 7644
rect 6610 7590 6612 7642
rect 6792 7590 6794 7642
rect 6548 7588 6554 7590
rect 6610 7588 6634 7590
rect 6690 7588 6714 7590
rect 6770 7588 6794 7590
rect 6850 7588 6856 7590
rect 6548 7579 6856 7588
rect 7024 7410 7052 8230
rect 7472 8084 7524 8090
rect 7472 8026 7524 8032
rect 7196 7812 7248 7818
rect 7196 7754 7248 7760
rect 6644 7404 6696 7410
rect 6644 7346 6696 7352
rect 7012 7404 7064 7410
rect 7012 7346 7064 7352
rect 6656 7002 6684 7346
rect 7208 7002 7236 7754
rect 6644 6996 6696 7002
rect 6644 6938 6696 6944
rect 7196 6996 7248 7002
rect 7196 6938 7248 6944
rect 6460 6860 6512 6866
rect 6460 6802 6512 6808
rect 6184 6792 6236 6798
rect 6184 6734 6236 6740
rect 6472 6458 6500 6802
rect 6548 6556 6856 6565
rect 6548 6554 6554 6556
rect 6610 6554 6634 6556
rect 6690 6554 6714 6556
rect 6770 6554 6794 6556
rect 6850 6554 6856 6556
rect 6610 6502 6612 6554
rect 6792 6502 6794 6554
rect 6548 6500 6554 6502
rect 6610 6500 6634 6502
rect 6690 6500 6714 6502
rect 6770 6500 6794 6502
rect 6850 6500 6856 6502
rect 6548 6491 6856 6500
rect 6460 6452 6512 6458
rect 6460 6394 6512 6400
rect 5908 6384 5960 6390
rect 5908 6326 5960 6332
rect 3749 6012 4057 6021
rect 3749 6010 3755 6012
rect 3811 6010 3835 6012
rect 3891 6010 3915 6012
rect 3971 6010 3995 6012
rect 4051 6010 4057 6012
rect 3811 5958 3813 6010
rect 3993 5958 3995 6010
rect 3749 5956 3755 5958
rect 3811 5956 3835 5958
rect 3891 5956 3915 5958
rect 3971 5956 3995 5958
rect 4051 5956 4057 5958
rect 3749 5947 4057 5956
rect 7208 5710 7236 6938
rect 7484 6322 7512 8026
rect 7564 7812 7616 7818
rect 7564 7754 7616 7760
rect 7576 6458 7604 7754
rect 7656 7404 7708 7410
rect 7656 7346 7708 7352
rect 7668 6458 7696 7346
rect 8208 6724 8260 6730
rect 8208 6666 8260 6672
rect 7564 6452 7616 6458
rect 7564 6394 7616 6400
rect 7656 6452 7708 6458
rect 7656 6394 7708 6400
rect 7472 6316 7524 6322
rect 7472 6258 7524 6264
rect 7380 6248 7432 6254
rect 7380 6190 7432 6196
rect 7392 5778 7420 6190
rect 7380 5772 7432 5778
rect 7380 5714 7432 5720
rect 7196 5704 7248 5710
rect 7196 5646 7248 5652
rect 6548 5468 6856 5477
rect 6548 5466 6554 5468
rect 6610 5466 6634 5468
rect 6690 5466 6714 5468
rect 6770 5466 6794 5468
rect 6850 5466 6856 5468
rect 6610 5414 6612 5466
rect 6792 5414 6794 5466
rect 6548 5412 6554 5414
rect 6610 5412 6634 5414
rect 6690 5412 6714 5414
rect 6770 5412 6794 5414
rect 6850 5412 6856 5414
rect 6548 5403 6856 5412
rect 8116 5160 8168 5166
rect 8116 5102 8168 5108
rect 3749 4924 4057 4933
rect 3749 4922 3755 4924
rect 3811 4922 3835 4924
rect 3891 4922 3915 4924
rect 3971 4922 3995 4924
rect 4051 4922 4057 4924
rect 3811 4870 3813 4922
rect 3993 4870 3995 4922
rect 3749 4868 3755 4870
rect 3811 4868 3835 4870
rect 3891 4868 3915 4870
rect 3971 4868 3995 4870
rect 4051 4868 4057 4870
rect 3749 4859 4057 4868
rect 8128 4690 8156 5102
rect 8116 4684 8168 4690
rect 8116 4626 8168 4632
rect 8220 4554 8248 6666
rect 8312 6390 8340 8502
rect 8404 8430 8432 9114
rect 8588 8566 8616 9862
rect 8852 9580 8904 9586
rect 8852 9522 8904 9528
rect 8864 8838 8892 9522
rect 9036 9512 9088 9518
rect 9036 9454 9088 9460
rect 9048 9178 9076 9454
rect 9220 9376 9272 9382
rect 9140 9336 9220 9364
rect 9036 9172 9088 9178
rect 9036 9114 9088 9120
rect 8852 8832 8904 8838
rect 8852 8774 8904 8780
rect 8576 8560 8628 8566
rect 8576 8502 8628 8508
rect 8392 8424 8444 8430
rect 8392 8366 8444 8372
rect 8404 7818 8432 8366
rect 8668 8288 8720 8294
rect 8668 8230 8720 8236
rect 8392 7812 8444 7818
rect 8392 7754 8444 7760
rect 8404 7410 8432 7754
rect 8680 7410 8708 8230
rect 8392 7404 8444 7410
rect 8392 7346 8444 7352
rect 8668 7404 8720 7410
rect 8668 7346 8720 7352
rect 8404 7002 8432 7346
rect 8576 7200 8628 7206
rect 8576 7142 8628 7148
rect 8392 6996 8444 7002
rect 8392 6938 8444 6944
rect 8588 6730 8616 7142
rect 8576 6724 8628 6730
rect 8576 6666 8628 6672
rect 8300 6384 8352 6390
rect 8300 6326 8352 6332
rect 8484 6180 8536 6186
rect 8484 6122 8536 6128
rect 8392 6112 8444 6118
rect 8392 6054 8444 6060
rect 8300 5840 8352 5846
rect 8300 5782 8352 5788
rect 8312 4690 8340 5782
rect 8404 5710 8432 6054
rect 8392 5704 8444 5710
rect 8392 5646 8444 5652
rect 8300 4684 8352 4690
rect 8300 4626 8352 4632
rect 8496 4622 8524 6122
rect 8588 5642 8616 6666
rect 8680 5778 8708 7346
rect 8760 6724 8812 6730
rect 8760 6666 8812 6672
rect 8772 6254 8800 6666
rect 8760 6248 8812 6254
rect 8760 6190 8812 6196
rect 8668 5772 8720 5778
rect 8668 5714 8720 5720
rect 8576 5636 8628 5642
rect 8576 5578 8628 5584
rect 8864 5234 8892 8774
rect 9140 8498 9168 9336
rect 9220 9318 9272 9324
rect 9347 9276 9655 9285
rect 9347 9274 9353 9276
rect 9409 9274 9433 9276
rect 9489 9274 9513 9276
rect 9569 9274 9593 9276
rect 9649 9274 9655 9276
rect 9409 9222 9411 9274
rect 9591 9222 9593 9274
rect 9347 9220 9353 9222
rect 9409 9220 9433 9222
rect 9489 9220 9513 9222
rect 9569 9220 9593 9222
rect 9649 9220 9655 9222
rect 9347 9211 9655 9220
rect 9772 8968 9824 8974
rect 9772 8910 9824 8916
rect 9128 8492 9180 8498
rect 9128 8434 9180 8440
rect 8944 5568 8996 5574
rect 8944 5510 8996 5516
rect 8956 5302 8984 5510
rect 9140 5370 9168 8434
rect 9347 8188 9655 8197
rect 9347 8186 9353 8188
rect 9409 8186 9433 8188
rect 9489 8186 9513 8188
rect 9569 8186 9593 8188
rect 9649 8186 9655 8188
rect 9409 8134 9411 8186
rect 9591 8134 9593 8186
rect 9347 8132 9353 8134
rect 9409 8132 9433 8134
rect 9489 8132 9513 8134
rect 9569 8132 9593 8134
rect 9649 8132 9655 8134
rect 9347 8123 9655 8132
rect 9220 7540 9272 7546
rect 9220 7482 9272 7488
rect 9232 6458 9260 7482
rect 9784 7274 9812 8910
rect 9772 7268 9824 7274
rect 9772 7210 9824 7216
rect 9347 7100 9655 7109
rect 9347 7098 9353 7100
rect 9409 7098 9433 7100
rect 9489 7098 9513 7100
rect 9569 7098 9593 7100
rect 9649 7098 9655 7100
rect 9409 7046 9411 7098
rect 9591 7046 9593 7098
rect 9347 7044 9353 7046
rect 9409 7044 9433 7046
rect 9489 7044 9513 7046
rect 9569 7044 9593 7046
rect 9649 7044 9655 7046
rect 9347 7035 9655 7044
rect 9312 6656 9364 6662
rect 9312 6598 9364 6604
rect 9680 6656 9732 6662
rect 9680 6598 9732 6604
rect 9220 6452 9272 6458
rect 9220 6394 9272 6400
rect 9324 6254 9352 6598
rect 9312 6248 9364 6254
rect 9232 6196 9312 6202
rect 9232 6190 9364 6196
rect 9232 6174 9352 6190
rect 9232 5794 9260 6174
rect 9324 6125 9352 6174
rect 9347 6012 9655 6021
rect 9347 6010 9353 6012
rect 9409 6010 9433 6012
rect 9489 6010 9513 6012
rect 9569 6010 9593 6012
rect 9649 6010 9655 6012
rect 9409 5958 9411 6010
rect 9591 5958 9593 6010
rect 9347 5956 9353 5958
rect 9409 5956 9433 5958
rect 9489 5956 9513 5958
rect 9569 5956 9593 5958
rect 9649 5956 9655 5958
rect 9347 5947 9655 5956
rect 9232 5778 9536 5794
rect 9232 5772 9548 5778
rect 9232 5766 9496 5772
rect 9128 5364 9180 5370
rect 9128 5306 9180 5312
rect 8944 5296 8996 5302
rect 8944 5238 8996 5244
rect 8852 5228 8904 5234
rect 8852 5170 8904 5176
rect 9324 5166 9352 5766
rect 9496 5714 9548 5720
rect 9588 5636 9640 5642
rect 9692 5624 9720 6598
rect 9784 5710 9812 7210
rect 9968 6798 9996 10406
rect 10060 7546 10088 11290
rect 10232 9988 10284 9994
rect 10232 9930 10284 9936
rect 10140 9580 10192 9586
rect 10140 9522 10192 9528
rect 10048 7540 10100 7546
rect 10048 7482 10100 7488
rect 10048 7200 10100 7206
rect 10048 7142 10100 7148
rect 9956 6792 10008 6798
rect 9956 6734 10008 6740
rect 9956 6248 10008 6254
rect 9956 6190 10008 6196
rect 9968 5846 9996 6190
rect 10060 6186 10088 7142
rect 10152 6662 10180 9522
rect 10244 9382 10272 9930
rect 10232 9376 10284 9382
rect 10232 9318 10284 9324
rect 10244 6730 10272 9318
rect 10232 6724 10284 6730
rect 10232 6666 10284 6672
rect 10140 6656 10192 6662
rect 10140 6598 10192 6604
rect 10336 6458 10364 12106
rect 10784 11756 10836 11762
rect 10784 11698 10836 11704
rect 10508 11688 10560 11694
rect 10508 11630 10560 11636
rect 10416 11552 10468 11558
rect 10416 11494 10468 11500
rect 10428 7478 10456 11494
rect 10520 11014 10548 11630
rect 10796 11558 10824 11698
rect 10784 11552 10836 11558
rect 10784 11494 10836 11500
rect 10508 11008 10560 11014
rect 10508 10950 10560 10956
rect 10520 10674 10548 10950
rect 10508 10668 10560 10674
rect 10508 10610 10560 10616
rect 11072 9704 11100 12786
rect 11152 10736 11204 10742
rect 11152 10678 11204 10684
rect 10888 9676 11100 9704
rect 10692 9376 10744 9382
rect 10692 9318 10744 9324
rect 10784 9376 10836 9382
rect 10784 9318 10836 9324
rect 10704 8498 10732 9318
rect 10692 8492 10744 8498
rect 10692 8434 10744 8440
rect 10692 7880 10744 7886
rect 10692 7822 10744 7828
rect 10704 7546 10732 7822
rect 10692 7540 10744 7546
rect 10692 7482 10744 7488
rect 10416 7472 10468 7478
rect 10796 7426 10824 9318
rect 10416 7414 10468 7420
rect 10704 7398 10824 7426
rect 10416 7336 10468 7342
rect 10416 7278 10468 7284
rect 10428 6866 10456 7278
rect 10416 6860 10468 6866
rect 10416 6802 10468 6808
rect 10416 6656 10468 6662
rect 10416 6598 10468 6604
rect 10324 6452 10376 6458
rect 10324 6394 10376 6400
rect 10428 6390 10456 6598
rect 10416 6384 10468 6390
rect 10416 6326 10468 6332
rect 10048 6180 10100 6186
rect 10048 6122 10100 6128
rect 10060 5914 10088 6122
rect 10416 6112 10468 6118
rect 10416 6054 10468 6060
rect 10048 5908 10100 5914
rect 10048 5850 10100 5856
rect 9956 5840 10008 5846
rect 9956 5782 10008 5788
rect 9772 5704 9824 5710
rect 9772 5646 9824 5652
rect 9640 5596 9720 5624
rect 9588 5578 9640 5584
rect 10060 5370 10088 5850
rect 10048 5364 10100 5370
rect 10048 5306 10100 5312
rect 9312 5160 9364 5166
rect 9312 5102 9364 5108
rect 9347 4924 9655 4933
rect 9347 4922 9353 4924
rect 9409 4922 9433 4924
rect 9489 4922 9513 4924
rect 9569 4922 9593 4924
rect 9649 4922 9655 4924
rect 9409 4870 9411 4922
rect 9591 4870 9593 4922
rect 9347 4868 9353 4870
rect 9409 4868 9433 4870
rect 9489 4868 9513 4870
rect 9569 4868 9593 4870
rect 9649 4868 9655 4870
rect 9347 4859 9655 4868
rect 10060 4758 10088 5306
rect 10048 4752 10100 4758
rect 10048 4694 10100 4700
rect 10428 4690 10456 6054
rect 10704 5778 10732 7398
rect 10692 5772 10744 5778
rect 10692 5714 10744 5720
rect 10888 5710 10916 9676
rect 11164 8838 11192 10678
rect 11256 9722 11284 14010
rect 11336 12096 11388 12102
rect 11336 12038 11388 12044
rect 11348 9926 11376 12038
rect 11336 9920 11388 9926
rect 11336 9862 11388 9868
rect 11244 9716 11296 9722
rect 11244 9658 11296 9664
rect 11152 8832 11204 8838
rect 11152 8774 11204 8780
rect 11060 7744 11112 7750
rect 11060 7686 11112 7692
rect 11072 7478 11100 7686
rect 11060 7472 11112 7478
rect 11060 7414 11112 7420
rect 11164 6798 11192 8774
rect 11244 8084 11296 8090
rect 11244 8026 11296 8032
rect 11256 6866 11284 8026
rect 11244 6860 11296 6866
rect 11244 6802 11296 6808
rect 11152 6792 11204 6798
rect 11152 6734 11204 6740
rect 11348 6390 11376 9862
rect 11440 6390 11468 19230
rect 11624 15502 11652 19450
rect 12084 17338 12112 20810
rect 12532 20800 12584 20806
rect 12532 20742 12584 20748
rect 12146 20700 12454 20709
rect 12146 20698 12152 20700
rect 12208 20698 12232 20700
rect 12288 20698 12312 20700
rect 12368 20698 12392 20700
rect 12448 20698 12454 20700
rect 12208 20646 12210 20698
rect 12390 20646 12392 20698
rect 12146 20644 12152 20646
rect 12208 20644 12232 20646
rect 12288 20644 12312 20646
rect 12368 20644 12392 20646
rect 12448 20644 12454 20646
rect 12146 20635 12454 20644
rect 12544 20602 12572 20742
rect 12532 20596 12584 20602
rect 12532 20538 12584 20544
rect 12162 20496 12218 20505
rect 12162 20431 12218 20440
rect 12440 20460 12492 20466
rect 12176 19990 12204 20431
rect 12492 20420 12572 20448
rect 12440 20402 12492 20408
rect 12256 20392 12308 20398
rect 12256 20334 12308 20340
rect 12268 20058 12296 20334
rect 12256 20052 12308 20058
rect 12256 19994 12308 20000
rect 12164 19984 12216 19990
rect 12164 19926 12216 19932
rect 12146 19612 12454 19621
rect 12146 19610 12152 19612
rect 12208 19610 12232 19612
rect 12288 19610 12312 19612
rect 12368 19610 12392 19612
rect 12448 19610 12454 19612
rect 12208 19558 12210 19610
rect 12390 19558 12392 19610
rect 12146 19556 12152 19558
rect 12208 19556 12232 19558
rect 12288 19556 12312 19558
rect 12368 19556 12392 19558
rect 12448 19556 12454 19558
rect 12146 19547 12454 19556
rect 12146 18524 12454 18533
rect 12146 18522 12152 18524
rect 12208 18522 12232 18524
rect 12288 18522 12312 18524
rect 12368 18522 12392 18524
rect 12448 18522 12454 18524
rect 12208 18470 12210 18522
rect 12390 18470 12392 18522
rect 12146 18468 12152 18470
rect 12208 18468 12232 18470
rect 12288 18468 12312 18470
rect 12368 18468 12392 18470
rect 12448 18468 12454 18470
rect 12146 18459 12454 18468
rect 12544 17882 12572 20420
rect 12622 20360 12678 20369
rect 12622 20295 12678 20304
rect 12636 19922 12664 20295
rect 12624 19916 12676 19922
rect 12624 19858 12676 19864
rect 12624 19712 12676 19718
rect 12624 19654 12676 19660
rect 12716 19712 12768 19718
rect 12716 19654 12768 19660
rect 12532 17876 12584 17882
rect 12532 17818 12584 17824
rect 12532 17536 12584 17542
rect 12532 17478 12584 17484
rect 12146 17436 12454 17445
rect 12146 17434 12152 17436
rect 12208 17434 12232 17436
rect 12288 17434 12312 17436
rect 12368 17434 12392 17436
rect 12448 17434 12454 17436
rect 12208 17382 12210 17434
rect 12390 17382 12392 17434
rect 12146 17380 12152 17382
rect 12208 17380 12232 17382
rect 12288 17380 12312 17382
rect 12368 17380 12392 17382
rect 12448 17380 12454 17382
rect 12146 17371 12454 17380
rect 12544 17338 12572 17478
rect 12072 17332 12124 17338
rect 12072 17274 12124 17280
rect 12532 17332 12584 17338
rect 12532 17274 12584 17280
rect 11796 17128 11848 17134
rect 11796 17070 11848 17076
rect 11808 16658 11836 17070
rect 11796 16652 11848 16658
rect 11796 16594 11848 16600
rect 11796 16448 11848 16454
rect 11796 16390 11848 16396
rect 11808 16250 11836 16390
rect 12146 16348 12454 16357
rect 12146 16346 12152 16348
rect 12208 16346 12232 16348
rect 12288 16346 12312 16348
rect 12368 16346 12392 16348
rect 12448 16346 12454 16348
rect 12208 16294 12210 16346
rect 12390 16294 12392 16346
rect 12146 16292 12152 16294
rect 12208 16292 12232 16294
rect 12288 16292 12312 16294
rect 12368 16292 12392 16294
rect 12448 16292 12454 16294
rect 12146 16283 12454 16292
rect 11796 16244 11848 16250
rect 11796 16186 11848 16192
rect 11980 16108 12032 16114
rect 11980 16050 12032 16056
rect 11992 15706 12020 16050
rect 11980 15700 12032 15706
rect 11980 15642 12032 15648
rect 11612 15496 11664 15502
rect 11612 15438 11664 15444
rect 12532 15428 12584 15434
rect 12532 15370 12584 15376
rect 12146 15260 12454 15269
rect 12146 15258 12152 15260
rect 12208 15258 12232 15260
rect 12288 15258 12312 15260
rect 12368 15258 12392 15260
rect 12448 15258 12454 15260
rect 12208 15206 12210 15258
rect 12390 15206 12392 15258
rect 12146 15204 12152 15206
rect 12208 15204 12232 15206
rect 12288 15204 12312 15206
rect 12368 15204 12392 15206
rect 12448 15204 12454 15206
rect 12146 15195 12454 15204
rect 11612 15156 11664 15162
rect 11612 15098 11664 15104
rect 11520 13252 11572 13258
rect 11520 13194 11572 13200
rect 11532 11898 11560 13194
rect 11520 11892 11572 11898
rect 11520 11834 11572 11840
rect 11624 11830 11652 15098
rect 12544 14618 12572 15370
rect 12532 14612 12584 14618
rect 12532 14554 12584 14560
rect 12146 14172 12454 14181
rect 12146 14170 12152 14172
rect 12208 14170 12232 14172
rect 12288 14170 12312 14172
rect 12368 14170 12392 14172
rect 12448 14170 12454 14172
rect 12208 14118 12210 14170
rect 12390 14118 12392 14170
rect 12146 14116 12152 14118
rect 12208 14116 12232 14118
rect 12288 14116 12312 14118
rect 12368 14116 12392 14118
rect 12448 14116 12454 14118
rect 12146 14107 12454 14116
rect 12146 13084 12454 13093
rect 12146 13082 12152 13084
rect 12208 13082 12232 13084
rect 12288 13082 12312 13084
rect 12368 13082 12392 13084
rect 12448 13082 12454 13084
rect 12208 13030 12210 13082
rect 12390 13030 12392 13082
rect 12146 13028 12152 13030
rect 12208 13028 12232 13030
rect 12288 13028 12312 13030
rect 12368 13028 12392 13030
rect 12448 13028 12454 13030
rect 12146 13019 12454 13028
rect 12636 12434 12664 19654
rect 12544 12406 12664 12434
rect 12146 11996 12454 12005
rect 12146 11994 12152 11996
rect 12208 11994 12232 11996
rect 12288 11994 12312 11996
rect 12368 11994 12392 11996
rect 12448 11994 12454 11996
rect 12208 11942 12210 11994
rect 12390 11942 12392 11994
rect 12146 11940 12152 11942
rect 12208 11940 12232 11942
rect 12288 11940 12312 11942
rect 12368 11940 12392 11942
rect 12448 11940 12454 11942
rect 12146 11931 12454 11940
rect 12440 11892 12492 11898
rect 12440 11834 12492 11840
rect 11612 11824 11664 11830
rect 11612 11766 11664 11772
rect 12452 11082 12480 11834
rect 12544 11354 12572 12406
rect 12728 11898 12756 19654
rect 12820 16998 12848 20878
rect 12900 20800 12952 20806
rect 12900 20742 12952 20748
rect 12912 20534 12940 20742
rect 12900 20528 12952 20534
rect 12900 20470 12952 20476
rect 13004 20262 13032 21830
rect 13820 21830 13872 21836
rect 13726 21791 13782 21800
rect 13740 21690 13768 21791
rect 13360 21684 13412 21690
rect 13728 21684 13780 21690
rect 13412 21644 13676 21672
rect 13360 21626 13412 21632
rect 13648 21536 13676 21644
rect 13728 21626 13780 21632
rect 13648 21508 13768 21536
rect 13176 21480 13228 21486
rect 13228 21428 13308 21434
rect 13176 21422 13308 21428
rect 13188 21406 13308 21422
rect 13084 20460 13136 20466
rect 13084 20402 13136 20408
rect 12992 20256 13044 20262
rect 12992 20198 13044 20204
rect 12900 19916 12952 19922
rect 12900 19858 12952 19864
rect 12912 19446 12940 19858
rect 12900 19440 12952 19446
rect 12900 19382 12952 19388
rect 12992 19372 13044 19378
rect 12992 19314 13044 19320
rect 12900 19304 12952 19310
rect 12900 19246 12952 19252
rect 12912 18766 12940 19246
rect 13004 18970 13032 19314
rect 13096 19174 13124 20402
rect 13176 20392 13228 20398
rect 13176 20334 13228 20340
rect 13084 19168 13136 19174
rect 13084 19110 13136 19116
rect 12992 18964 13044 18970
rect 12992 18906 13044 18912
rect 13084 18896 13136 18902
rect 12990 18864 13046 18873
rect 13084 18838 13136 18844
rect 12990 18799 13046 18808
rect 12900 18760 12952 18766
rect 12900 18702 12952 18708
rect 12808 16992 12860 16998
rect 12808 16934 12860 16940
rect 12820 16114 12848 16934
rect 13004 16454 13032 18799
rect 13096 18358 13124 18838
rect 13084 18352 13136 18358
rect 13084 18294 13136 18300
rect 13188 18154 13216 20334
rect 13280 19836 13308 21406
rect 13636 21412 13688 21418
rect 13636 21354 13688 21360
rect 13544 21140 13596 21146
rect 13544 21082 13596 21088
rect 13452 20800 13504 20806
rect 13452 20742 13504 20748
rect 13360 19848 13412 19854
rect 13280 19808 13360 19836
rect 13360 19790 13412 19796
rect 13268 19372 13320 19378
rect 13268 19314 13320 19320
rect 13176 18148 13228 18154
rect 13176 18090 13228 18096
rect 13084 17536 13136 17542
rect 13084 17478 13136 17484
rect 12992 16448 13044 16454
rect 12992 16390 13044 16396
rect 12808 16108 12860 16114
rect 12808 16050 12860 16056
rect 13096 15434 13124 17478
rect 13176 17264 13228 17270
rect 13176 17206 13228 17212
rect 13084 15428 13136 15434
rect 13084 15370 13136 15376
rect 13188 15162 13216 17206
rect 13280 15366 13308 19314
rect 13372 18737 13400 19790
rect 13464 18873 13492 20742
rect 13556 19854 13584 21082
rect 13648 21010 13676 21354
rect 13740 21146 13768 21508
rect 13728 21140 13780 21146
rect 13728 21082 13780 21088
rect 13636 21004 13688 21010
rect 13636 20946 13688 20952
rect 13648 20330 13676 20946
rect 13636 20324 13688 20330
rect 13636 20266 13688 20272
rect 13728 19984 13780 19990
rect 13726 19952 13728 19961
rect 13780 19952 13782 19961
rect 13726 19887 13782 19896
rect 13544 19848 13596 19854
rect 13544 19790 13596 19796
rect 13636 19712 13688 19718
rect 13636 19654 13688 19660
rect 13544 19304 13596 19310
rect 13544 19246 13596 19252
rect 13450 18864 13506 18873
rect 13450 18799 13506 18808
rect 13452 18760 13504 18766
rect 13358 18728 13414 18737
rect 13452 18702 13504 18708
rect 13358 18663 13414 18672
rect 13464 17746 13492 18702
rect 13452 17740 13504 17746
rect 13452 17682 13504 17688
rect 13360 17536 13412 17542
rect 13360 17478 13412 17484
rect 13268 15360 13320 15366
rect 13268 15302 13320 15308
rect 13176 15156 13228 15162
rect 13176 15098 13228 15104
rect 13372 14414 13400 17478
rect 13556 16658 13584 19246
rect 13648 19174 13676 19654
rect 13636 19168 13688 19174
rect 13636 19110 13688 19116
rect 13636 18964 13688 18970
rect 13636 18906 13688 18912
rect 13648 18358 13676 18906
rect 13832 18834 13860 21830
rect 14004 21344 14056 21350
rect 14004 21286 14056 21292
rect 13912 20936 13964 20942
rect 13912 20878 13964 20884
rect 13924 20602 13952 20878
rect 13912 20596 13964 20602
rect 13912 20538 13964 20544
rect 13912 20256 13964 20262
rect 13912 20198 13964 20204
rect 13820 18828 13872 18834
rect 13820 18770 13872 18776
rect 13728 18692 13780 18698
rect 13728 18634 13780 18640
rect 13636 18352 13688 18358
rect 13636 18294 13688 18300
rect 13740 18222 13768 18634
rect 13832 18222 13860 18770
rect 13728 18216 13780 18222
rect 13728 18158 13780 18164
rect 13820 18216 13872 18222
rect 13820 18158 13872 18164
rect 13636 18148 13688 18154
rect 13636 18090 13688 18096
rect 13648 17270 13676 18090
rect 13636 17264 13688 17270
rect 13636 17206 13688 17212
rect 13740 17066 13768 18158
rect 13924 18086 13952 20198
rect 14016 20058 14044 21286
rect 14004 20052 14056 20058
rect 14004 19994 14056 20000
rect 14108 19990 14136 22442
rect 14476 22234 14504 23800
rect 14556 22568 14608 22574
rect 14556 22510 14608 22516
rect 14464 22228 14516 22234
rect 14464 22170 14516 22176
rect 14372 21956 14424 21962
rect 14372 21898 14424 21904
rect 14384 21486 14412 21898
rect 14372 21480 14424 21486
rect 14372 21422 14424 21428
rect 14188 21412 14240 21418
rect 14188 21354 14240 21360
rect 14096 19984 14148 19990
rect 14096 19926 14148 19932
rect 13912 18080 13964 18086
rect 13912 18022 13964 18028
rect 13910 17912 13966 17921
rect 14200 17898 14228 21354
rect 14280 20936 14332 20942
rect 14280 20878 14332 20884
rect 14292 20534 14320 20878
rect 14280 20528 14332 20534
rect 14280 20470 14332 20476
rect 14372 20460 14424 20466
rect 14372 20402 14424 20408
rect 14384 20058 14412 20402
rect 14464 20256 14516 20262
rect 14464 20198 14516 20204
rect 14372 20052 14424 20058
rect 14372 19994 14424 20000
rect 14476 19854 14504 20198
rect 14568 19990 14596 22510
rect 14844 22166 14872 23854
rect 15028 23746 15056 23854
rect 15106 23800 15162 24600
rect 15750 23800 15806 24600
rect 15856 23854 16344 23882
rect 15120 23746 15148 23800
rect 15028 23718 15148 23746
rect 15764 23746 15792 23800
rect 15856 23746 15884 23854
rect 15764 23718 15884 23746
rect 16316 22658 16344 23854
rect 16394 23800 16450 24600
rect 17038 23800 17094 24600
rect 17682 23800 17738 24600
rect 18326 23800 18382 24600
rect 18970 23800 19026 24600
rect 19614 23800 19670 24600
rect 20258 23800 20314 24600
rect 20902 23800 20958 24600
rect 21546 23800 21602 24600
rect 22190 23800 22246 24600
rect 22834 23800 22890 24600
rect 23478 23800 23534 24600
rect 24122 23800 24178 24600
rect 16316 22630 16436 22658
rect 16304 22568 16356 22574
rect 16304 22510 16356 22516
rect 15568 22432 15620 22438
rect 15568 22374 15620 22380
rect 14945 22332 15253 22341
rect 14945 22330 14951 22332
rect 15007 22330 15031 22332
rect 15087 22330 15111 22332
rect 15167 22330 15191 22332
rect 15247 22330 15253 22332
rect 15007 22278 15009 22330
rect 15189 22278 15191 22330
rect 14945 22276 14951 22278
rect 15007 22276 15031 22278
rect 15087 22276 15111 22278
rect 15167 22276 15191 22278
rect 15247 22276 15253 22278
rect 14945 22267 15253 22276
rect 14832 22160 14884 22166
rect 14832 22102 14884 22108
rect 14740 21888 14792 21894
rect 14740 21830 14792 21836
rect 14646 21448 14702 21457
rect 14646 21383 14702 21392
rect 14660 20777 14688 21383
rect 14752 21049 14780 21830
rect 14844 21146 14872 22102
rect 15476 22024 15528 22030
rect 15580 22012 15608 22374
rect 16316 22234 16344 22510
rect 16028 22228 16080 22234
rect 16028 22170 16080 22176
rect 16304 22228 16356 22234
rect 16304 22170 16356 22176
rect 16040 22030 16068 22170
rect 16120 22160 16172 22166
rect 16120 22102 16172 22108
rect 16408 22114 16436 22630
rect 16488 22160 16540 22166
rect 16408 22108 16488 22114
rect 16408 22102 16540 22108
rect 16132 22030 16160 22102
rect 16408 22086 16528 22102
rect 16948 22092 17000 22098
rect 15752 22024 15804 22030
rect 15580 21984 15752 22012
rect 15476 21966 15528 21972
rect 15752 21966 15804 21972
rect 16028 22024 16080 22030
rect 16028 21966 16080 21972
rect 16120 22024 16172 22030
rect 16120 21966 16172 21972
rect 15016 21956 15068 21962
rect 15016 21898 15068 21904
rect 15028 21729 15056 21898
rect 15200 21888 15252 21894
rect 15384 21888 15436 21894
rect 15200 21830 15252 21836
rect 15304 21848 15384 21876
rect 15014 21720 15070 21729
rect 15014 21655 15070 21664
rect 15028 21486 15056 21655
rect 15108 21548 15160 21554
rect 15212 21536 15240 21830
rect 15304 21690 15332 21848
rect 15384 21830 15436 21836
rect 15292 21684 15344 21690
rect 15292 21626 15344 21632
rect 15160 21508 15240 21536
rect 15108 21490 15160 21496
rect 15016 21480 15068 21486
rect 15016 21422 15068 21428
rect 15212 21350 15240 21508
rect 15292 21480 15344 21486
rect 15292 21422 15344 21428
rect 15200 21344 15252 21350
rect 15200 21286 15252 21292
rect 14945 21244 15253 21253
rect 14945 21242 14951 21244
rect 15007 21242 15031 21244
rect 15087 21242 15111 21244
rect 15167 21242 15191 21244
rect 15247 21242 15253 21244
rect 15007 21190 15009 21242
rect 15189 21190 15191 21242
rect 14945 21188 14951 21190
rect 15007 21188 15031 21190
rect 15087 21188 15111 21190
rect 15167 21188 15191 21190
rect 15247 21188 15253 21190
rect 14945 21179 15253 21188
rect 14832 21140 14884 21146
rect 14832 21082 14884 21088
rect 14924 21140 14976 21146
rect 14924 21082 14976 21088
rect 14738 21040 14794 21049
rect 14936 21010 14964 21082
rect 14738 20975 14794 20984
rect 14924 21004 14976 21010
rect 14752 20890 14780 20975
rect 14924 20946 14976 20952
rect 14752 20862 14872 20890
rect 14844 20806 14872 20862
rect 14832 20800 14884 20806
rect 14646 20768 14702 20777
rect 14832 20742 14884 20748
rect 14646 20703 14702 20712
rect 15304 20602 15332 21422
rect 15488 21321 15516 21966
rect 15658 21720 15714 21729
rect 15658 21655 15660 21664
rect 15712 21655 15714 21664
rect 15660 21626 15712 21632
rect 15474 21312 15530 21321
rect 15474 21247 15530 21256
rect 15488 21146 15516 21247
rect 15658 21176 15714 21185
rect 15476 21140 15528 21146
rect 15764 21146 15792 21966
rect 15936 21956 15988 21962
rect 15936 21898 15988 21904
rect 15948 21865 15976 21898
rect 15934 21856 15990 21865
rect 15934 21791 15990 21800
rect 15936 21684 15988 21690
rect 15936 21626 15988 21632
rect 15658 21111 15714 21120
rect 15752 21140 15804 21146
rect 15476 21082 15528 21088
rect 15384 20936 15436 20942
rect 15384 20878 15436 20884
rect 15396 20806 15424 20878
rect 15384 20800 15436 20806
rect 15672 20777 15700 21111
rect 15752 21082 15804 21088
rect 15384 20742 15436 20748
rect 15658 20768 15714 20777
rect 15658 20703 15714 20712
rect 15672 20602 15700 20703
rect 14648 20596 14700 20602
rect 14648 20538 14700 20544
rect 15292 20596 15344 20602
rect 15660 20596 15712 20602
rect 15292 20538 15344 20544
rect 15580 20556 15660 20584
rect 14556 19984 14608 19990
rect 14556 19926 14608 19932
rect 14464 19848 14516 19854
rect 14464 19790 14516 19796
rect 14556 19848 14608 19854
rect 14556 19790 14608 19796
rect 14280 19168 14332 19174
rect 14280 19110 14332 19116
rect 14372 19168 14424 19174
rect 14372 19110 14424 19116
rect 14292 18766 14320 19110
rect 14280 18760 14332 18766
rect 14280 18702 14332 18708
rect 14292 18426 14320 18702
rect 14280 18420 14332 18426
rect 14280 18362 14332 18368
rect 14384 18170 14412 19110
rect 14292 18142 14412 18170
rect 14292 18086 14320 18142
rect 14280 18080 14332 18086
rect 14280 18022 14332 18028
rect 14372 18080 14424 18086
rect 14372 18022 14424 18028
rect 14200 17870 14320 17898
rect 13910 17847 13912 17856
rect 13964 17847 13966 17856
rect 13912 17818 13964 17824
rect 14188 17672 14240 17678
rect 14188 17614 14240 17620
rect 14004 17604 14056 17610
rect 14004 17546 14056 17552
rect 13728 17060 13780 17066
rect 13728 17002 13780 17008
rect 14016 16998 14044 17546
rect 14200 17338 14228 17614
rect 14292 17542 14320 17870
rect 14280 17536 14332 17542
rect 14280 17478 14332 17484
rect 14188 17332 14240 17338
rect 14188 17274 14240 17280
rect 14004 16992 14056 16998
rect 14004 16934 14056 16940
rect 13544 16652 13596 16658
rect 13544 16594 13596 16600
rect 14280 15904 14332 15910
rect 14280 15846 14332 15852
rect 14292 15094 14320 15846
rect 14384 15434 14412 18022
rect 14372 15428 14424 15434
rect 14372 15370 14424 15376
rect 14280 15088 14332 15094
rect 14280 15030 14332 15036
rect 13360 14408 13412 14414
rect 13360 14350 13412 14356
rect 13544 14408 13596 14414
rect 13544 14350 13596 14356
rect 14096 14408 14148 14414
rect 14096 14350 14148 14356
rect 13268 14340 13320 14346
rect 13268 14282 13320 14288
rect 13280 14006 13308 14282
rect 13268 14000 13320 14006
rect 13268 13942 13320 13948
rect 13084 13932 13136 13938
rect 13084 13874 13136 13880
rect 13096 12986 13124 13874
rect 13084 12980 13136 12986
rect 13084 12922 13136 12928
rect 12900 12844 12952 12850
rect 12900 12786 12952 12792
rect 12912 12434 12940 12786
rect 12820 12406 12940 12434
rect 12716 11892 12768 11898
rect 12716 11834 12768 11840
rect 12624 11756 12676 11762
rect 12624 11698 12676 11704
rect 12532 11348 12584 11354
rect 12532 11290 12584 11296
rect 12440 11076 12492 11082
rect 12440 11018 12492 11024
rect 12146 10908 12454 10917
rect 12146 10906 12152 10908
rect 12208 10906 12232 10908
rect 12288 10906 12312 10908
rect 12368 10906 12392 10908
rect 12448 10906 12454 10908
rect 12208 10854 12210 10906
rect 12390 10854 12392 10906
rect 12146 10852 12152 10854
rect 12208 10852 12232 10854
rect 12288 10852 12312 10854
rect 12368 10852 12392 10854
rect 12448 10852 12454 10854
rect 12146 10843 12454 10852
rect 12544 10742 12572 11290
rect 12636 11082 12664 11698
rect 12624 11076 12676 11082
rect 12624 11018 12676 11024
rect 12532 10736 12584 10742
rect 12532 10678 12584 10684
rect 11520 10464 11572 10470
rect 11520 10406 11572 10412
rect 11532 10062 11560 10406
rect 11520 10056 11572 10062
rect 11520 9998 11572 10004
rect 12146 9820 12454 9829
rect 12146 9818 12152 9820
rect 12208 9818 12232 9820
rect 12288 9818 12312 9820
rect 12368 9818 12392 9820
rect 12448 9818 12454 9820
rect 12208 9766 12210 9818
rect 12390 9766 12392 9818
rect 12146 9764 12152 9766
rect 12208 9764 12232 9766
rect 12288 9764 12312 9766
rect 12368 9764 12392 9766
rect 12448 9764 12454 9766
rect 12146 9755 12454 9764
rect 12624 9716 12676 9722
rect 12624 9658 12676 9664
rect 12636 9586 12664 9658
rect 12820 9654 12848 12406
rect 13096 12238 13124 12922
rect 13084 12232 13136 12238
rect 13084 12174 13136 12180
rect 13084 11552 13136 11558
rect 13084 11494 13136 11500
rect 13096 11150 13124 11494
rect 13084 11144 13136 11150
rect 13084 11086 13136 11092
rect 13556 10810 13584 14350
rect 14108 14006 14136 14350
rect 14096 14000 14148 14006
rect 14096 13942 14148 13948
rect 14188 13932 14240 13938
rect 14188 13874 14240 13880
rect 14096 13456 14148 13462
rect 14094 13424 14096 13433
rect 14148 13424 14150 13433
rect 14094 13359 14150 13368
rect 13912 12844 13964 12850
rect 13912 12786 13964 12792
rect 13924 12102 13952 12786
rect 14108 12170 14136 13359
rect 14096 12164 14148 12170
rect 14096 12106 14148 12112
rect 13912 12096 13964 12102
rect 13912 12038 13964 12044
rect 13544 10804 13596 10810
rect 13544 10746 13596 10752
rect 13636 10464 13688 10470
rect 13636 10406 13688 10412
rect 12900 10056 12952 10062
rect 12900 9998 12952 10004
rect 12808 9648 12860 9654
rect 12808 9590 12860 9596
rect 12912 9586 12940 9998
rect 12992 9920 13044 9926
rect 12992 9862 13044 9868
rect 13004 9586 13032 9862
rect 13648 9722 13676 10406
rect 14200 9926 14228 13874
rect 14188 9920 14240 9926
rect 14188 9862 14240 9868
rect 13636 9716 13688 9722
rect 13636 9658 13688 9664
rect 12624 9580 12676 9586
rect 12624 9522 12676 9528
rect 12900 9580 12952 9586
rect 12900 9522 12952 9528
rect 12992 9580 13044 9586
rect 12992 9522 13044 9528
rect 12624 9376 12676 9382
rect 12624 9318 12676 9324
rect 12716 9376 12768 9382
rect 12716 9318 12768 9324
rect 12636 8838 12664 9318
rect 12728 8906 12756 9318
rect 12912 9178 12940 9522
rect 12900 9172 12952 9178
rect 12900 9114 12952 9120
rect 12716 8900 12768 8906
rect 12716 8842 12768 8848
rect 11520 8832 11572 8838
rect 11520 8774 11572 8780
rect 12624 8832 12676 8838
rect 12624 8774 12676 8780
rect 11532 8566 11560 8774
rect 12146 8732 12454 8741
rect 12146 8730 12152 8732
rect 12208 8730 12232 8732
rect 12288 8730 12312 8732
rect 12368 8730 12392 8732
rect 12448 8730 12454 8732
rect 12208 8678 12210 8730
rect 12390 8678 12392 8730
rect 12146 8676 12152 8678
rect 12208 8676 12232 8678
rect 12288 8676 12312 8678
rect 12368 8676 12392 8678
rect 12448 8676 12454 8678
rect 12146 8667 12454 8676
rect 11520 8560 11572 8566
rect 11520 8502 11572 8508
rect 12532 8492 12584 8498
rect 12532 8434 12584 8440
rect 12072 8356 12124 8362
rect 12072 8298 12124 8304
rect 11520 8288 11572 8294
rect 11520 8230 11572 8236
rect 11888 8288 11940 8294
rect 11888 8230 11940 8236
rect 11532 7818 11560 8230
rect 11520 7812 11572 7818
rect 11520 7754 11572 7760
rect 11612 7812 11664 7818
rect 11612 7754 11664 7760
rect 11336 6384 11388 6390
rect 11336 6326 11388 6332
rect 11428 6384 11480 6390
rect 11428 6326 11480 6332
rect 10968 6316 11020 6322
rect 10968 6258 11020 6264
rect 10980 5914 11008 6258
rect 11152 6248 11204 6254
rect 11152 6190 11204 6196
rect 10968 5908 11020 5914
rect 10968 5850 11020 5856
rect 11164 5778 11192 6190
rect 11244 6112 11296 6118
rect 11244 6054 11296 6060
rect 11336 6112 11388 6118
rect 11336 6054 11388 6060
rect 11532 6066 11560 7754
rect 11624 7478 11652 7754
rect 11900 7750 11928 8230
rect 11888 7744 11940 7750
rect 11888 7686 11940 7692
rect 12084 7478 12112 8298
rect 12544 7750 12572 8434
rect 12532 7744 12584 7750
rect 12532 7686 12584 7692
rect 12146 7644 12454 7653
rect 12146 7642 12152 7644
rect 12208 7642 12232 7644
rect 12288 7642 12312 7644
rect 12368 7642 12392 7644
rect 12448 7642 12454 7644
rect 12208 7590 12210 7642
rect 12390 7590 12392 7642
rect 12146 7588 12152 7590
rect 12208 7588 12232 7590
rect 12288 7588 12312 7590
rect 12368 7588 12392 7590
rect 12448 7588 12454 7590
rect 12146 7579 12454 7588
rect 11612 7472 11664 7478
rect 11612 7414 11664 7420
rect 12072 7472 12124 7478
rect 12072 7414 12124 7420
rect 11624 6254 11652 7414
rect 12084 6798 12112 7414
rect 12544 6866 12572 7686
rect 12532 6860 12584 6866
rect 12532 6802 12584 6808
rect 12072 6792 12124 6798
rect 12072 6734 12124 6740
rect 11796 6724 11848 6730
rect 11796 6666 11848 6672
rect 11612 6248 11664 6254
rect 11612 6190 11664 6196
rect 11152 5772 11204 5778
rect 11152 5714 11204 5720
rect 10876 5704 10928 5710
rect 10876 5646 10928 5652
rect 11164 5166 11192 5714
rect 11256 5710 11284 6054
rect 11244 5704 11296 5710
rect 11244 5646 11296 5652
rect 11152 5160 11204 5166
rect 11152 5102 11204 5108
rect 10416 4684 10468 4690
rect 10416 4626 10468 4632
rect 8484 4616 8536 4622
rect 8484 4558 8536 4564
rect 8208 4548 8260 4554
rect 8208 4490 8260 4496
rect 6548 4380 6856 4389
rect 6548 4378 6554 4380
rect 6610 4378 6634 4380
rect 6690 4378 6714 4380
rect 6770 4378 6794 4380
rect 6850 4378 6856 4380
rect 6610 4326 6612 4378
rect 6792 4326 6794 4378
rect 6548 4324 6554 4326
rect 6610 4324 6634 4326
rect 6690 4324 6714 4326
rect 6770 4324 6794 4326
rect 6850 4324 6856 4326
rect 6548 4315 6856 4324
rect 3749 3836 4057 3845
rect 3749 3834 3755 3836
rect 3811 3834 3835 3836
rect 3891 3834 3915 3836
rect 3971 3834 3995 3836
rect 4051 3834 4057 3836
rect 3811 3782 3813 3834
rect 3993 3782 3995 3834
rect 3749 3780 3755 3782
rect 3811 3780 3835 3782
rect 3891 3780 3915 3782
rect 3971 3780 3995 3782
rect 4051 3780 4057 3782
rect 3749 3771 4057 3780
rect 9347 3836 9655 3845
rect 9347 3834 9353 3836
rect 9409 3834 9433 3836
rect 9489 3834 9513 3836
rect 9569 3834 9593 3836
rect 9649 3834 9655 3836
rect 9409 3782 9411 3834
rect 9591 3782 9593 3834
rect 9347 3780 9353 3782
rect 9409 3780 9433 3782
rect 9489 3780 9513 3782
rect 9569 3780 9593 3782
rect 9649 3780 9655 3782
rect 9347 3771 9655 3780
rect 1400 3392 1452 3398
rect 1400 3334 1452 3340
rect 1412 3097 1440 3334
rect 6548 3292 6856 3301
rect 6548 3290 6554 3292
rect 6610 3290 6634 3292
rect 6690 3290 6714 3292
rect 6770 3290 6794 3292
rect 6850 3290 6856 3292
rect 6610 3238 6612 3290
rect 6792 3238 6794 3290
rect 6548 3236 6554 3238
rect 6610 3236 6634 3238
rect 6690 3236 6714 3238
rect 6770 3236 6794 3238
rect 6850 3236 6856 3238
rect 6548 3227 6856 3236
rect 11348 3194 11376 6054
rect 11532 6038 11652 6066
rect 11624 5574 11652 6038
rect 11612 5568 11664 5574
rect 11612 5510 11664 5516
rect 11808 5166 11836 6666
rect 12072 6656 12124 6662
rect 12072 6598 12124 6604
rect 11888 6316 11940 6322
rect 11888 6258 11940 6264
rect 11796 5160 11848 5166
rect 11796 5102 11848 5108
rect 11900 4146 11928 6258
rect 11980 5568 12032 5574
rect 11980 5510 12032 5516
rect 11888 4140 11940 4146
rect 11888 4082 11940 4088
rect 11336 3188 11388 3194
rect 11336 3130 11388 3136
rect 1398 3088 1454 3097
rect 1398 3023 1454 3032
rect 11992 2854 12020 5510
rect 12084 5370 12112 6598
rect 12146 6556 12454 6565
rect 12146 6554 12152 6556
rect 12208 6554 12232 6556
rect 12288 6554 12312 6556
rect 12368 6554 12392 6556
rect 12448 6554 12454 6556
rect 12208 6502 12210 6554
rect 12390 6502 12392 6554
rect 12146 6500 12152 6502
rect 12208 6500 12232 6502
rect 12288 6500 12312 6502
rect 12368 6500 12392 6502
rect 12448 6500 12454 6502
rect 12146 6491 12454 6500
rect 12636 5642 12664 8774
rect 12728 6458 12756 8842
rect 13004 6458 13032 9522
rect 13360 7812 13412 7818
rect 13360 7754 13412 7760
rect 13372 7546 13400 7754
rect 13820 7744 13872 7750
rect 13820 7686 13872 7692
rect 13360 7540 13412 7546
rect 13360 7482 13412 7488
rect 13372 6866 13400 7482
rect 13728 7404 13780 7410
rect 13728 7346 13780 7352
rect 13740 7206 13768 7346
rect 13452 7200 13504 7206
rect 13452 7142 13504 7148
rect 13544 7200 13596 7206
rect 13544 7142 13596 7148
rect 13728 7200 13780 7206
rect 13728 7142 13780 7148
rect 13464 7002 13492 7142
rect 13452 6996 13504 7002
rect 13452 6938 13504 6944
rect 13360 6860 13412 6866
rect 13360 6802 13412 6808
rect 13176 6656 13228 6662
rect 13176 6598 13228 6604
rect 12716 6452 12768 6458
rect 12716 6394 12768 6400
rect 12992 6452 13044 6458
rect 12992 6394 13044 6400
rect 12716 6248 12768 6254
rect 12716 6190 12768 6196
rect 12728 5778 12756 6190
rect 12716 5772 12768 5778
rect 12716 5714 12768 5720
rect 12624 5636 12676 5642
rect 12624 5578 12676 5584
rect 12146 5468 12454 5477
rect 12146 5466 12152 5468
rect 12208 5466 12232 5468
rect 12288 5466 12312 5468
rect 12368 5466 12392 5468
rect 12448 5466 12454 5468
rect 12208 5414 12210 5466
rect 12390 5414 12392 5466
rect 12146 5412 12152 5414
rect 12208 5412 12232 5414
rect 12288 5412 12312 5414
rect 12368 5412 12392 5414
rect 12448 5412 12454 5414
rect 12146 5403 12454 5412
rect 13188 5370 13216 6598
rect 13556 6254 13584 7142
rect 13740 6866 13768 7142
rect 13728 6860 13780 6866
rect 13728 6802 13780 6808
rect 13832 6254 13860 7686
rect 14476 7449 14504 19790
rect 14568 19378 14596 19790
rect 14556 19372 14608 19378
rect 14556 19314 14608 19320
rect 14568 18630 14596 19314
rect 14556 18624 14608 18630
rect 14556 18566 14608 18572
rect 14568 18306 14596 18566
rect 14660 18426 14688 20538
rect 15200 20392 15252 20398
rect 15384 20392 15436 20398
rect 15252 20352 15332 20380
rect 15200 20334 15252 20340
rect 14945 20156 15253 20165
rect 14945 20154 14951 20156
rect 15007 20154 15031 20156
rect 15087 20154 15111 20156
rect 15167 20154 15191 20156
rect 15247 20154 15253 20156
rect 15007 20102 15009 20154
rect 15189 20102 15191 20154
rect 14945 20100 14951 20102
rect 15007 20100 15031 20102
rect 15087 20100 15111 20102
rect 15167 20100 15191 20102
rect 15247 20100 15253 20102
rect 14945 20091 15253 20100
rect 15304 20058 15332 20352
rect 15384 20334 15436 20340
rect 15292 20052 15344 20058
rect 15292 19994 15344 20000
rect 15292 19916 15344 19922
rect 15292 19858 15344 19864
rect 14740 19712 14792 19718
rect 14740 19654 14792 19660
rect 14832 19712 14884 19718
rect 14832 19654 14884 19660
rect 14752 19514 14780 19654
rect 14740 19508 14792 19514
rect 14740 19450 14792 19456
rect 14648 18420 14700 18426
rect 14648 18362 14700 18368
rect 14752 18358 14780 19450
rect 14844 19446 14872 19654
rect 14832 19440 14884 19446
rect 14832 19382 14884 19388
rect 14740 18352 14792 18358
rect 14568 18290 14688 18306
rect 14740 18294 14792 18300
rect 14568 18284 14700 18290
rect 14568 18278 14648 18284
rect 14648 18226 14700 18232
rect 14648 17536 14700 17542
rect 14648 17478 14700 17484
rect 14556 15428 14608 15434
rect 14556 15370 14608 15376
rect 14568 15026 14596 15370
rect 14556 15020 14608 15026
rect 14556 14962 14608 14968
rect 14660 12434 14688 17478
rect 14844 16250 14872 19382
rect 14945 19068 15253 19077
rect 14945 19066 14951 19068
rect 15007 19066 15031 19068
rect 15087 19066 15111 19068
rect 15167 19066 15191 19068
rect 15247 19066 15253 19068
rect 15007 19014 15009 19066
rect 15189 19014 15191 19066
rect 14945 19012 14951 19014
rect 15007 19012 15031 19014
rect 15087 19012 15111 19014
rect 15167 19012 15191 19014
rect 15247 19012 15253 19014
rect 14945 19003 15253 19012
rect 15304 18970 15332 19858
rect 15292 18964 15344 18970
rect 15292 18906 15344 18912
rect 15292 18284 15344 18290
rect 15292 18226 15344 18232
rect 14945 17980 15253 17989
rect 14945 17978 14951 17980
rect 15007 17978 15031 17980
rect 15087 17978 15111 17980
rect 15167 17978 15191 17980
rect 15247 17978 15253 17980
rect 15007 17926 15009 17978
rect 15189 17926 15191 17978
rect 14945 17924 14951 17926
rect 15007 17924 15031 17926
rect 15087 17924 15111 17926
rect 15167 17924 15191 17926
rect 15247 17924 15253 17926
rect 14945 17915 15253 17924
rect 15200 17876 15252 17882
rect 15200 17818 15252 17824
rect 15212 17542 15240 17818
rect 15200 17536 15252 17542
rect 15200 17478 15252 17484
rect 14945 16892 15253 16901
rect 14945 16890 14951 16892
rect 15007 16890 15031 16892
rect 15087 16890 15111 16892
rect 15167 16890 15191 16892
rect 15247 16890 15253 16892
rect 15007 16838 15009 16890
rect 15189 16838 15191 16890
rect 14945 16836 14951 16838
rect 15007 16836 15031 16838
rect 15087 16836 15111 16838
rect 15167 16836 15191 16838
rect 15247 16836 15253 16838
rect 14945 16827 15253 16836
rect 14832 16244 14884 16250
rect 14832 16186 14884 16192
rect 15304 16114 15332 18226
rect 15396 17610 15424 20334
rect 15476 19984 15528 19990
rect 15476 19926 15528 19932
rect 15488 17882 15516 19926
rect 15476 17876 15528 17882
rect 15476 17818 15528 17824
rect 15384 17604 15436 17610
rect 15384 17546 15436 17552
rect 15488 16590 15516 17818
rect 15580 17542 15608 20556
rect 15660 20538 15712 20544
rect 15844 20460 15896 20466
rect 15844 20402 15896 20408
rect 15660 19712 15712 19718
rect 15660 19654 15712 19660
rect 15672 19417 15700 19654
rect 15856 19514 15884 20402
rect 15844 19508 15896 19514
rect 15844 19450 15896 19456
rect 15658 19408 15714 19417
rect 15658 19343 15714 19352
rect 15752 19372 15804 19378
rect 15752 19314 15804 19320
rect 15764 18834 15792 19314
rect 15844 18964 15896 18970
rect 15844 18906 15896 18912
rect 15752 18828 15804 18834
rect 15752 18770 15804 18776
rect 15764 18426 15792 18770
rect 15752 18420 15804 18426
rect 15752 18362 15804 18368
rect 15764 17882 15792 18362
rect 15752 17876 15804 17882
rect 15752 17818 15804 17824
rect 15856 17678 15884 18906
rect 15948 18698 15976 21626
rect 16040 21350 16068 21966
rect 16120 21888 16172 21894
rect 16120 21830 16172 21836
rect 16304 21888 16356 21894
rect 16304 21830 16356 21836
rect 16132 21622 16160 21830
rect 16316 21729 16344 21830
rect 16302 21720 16358 21729
rect 16302 21655 16358 21664
rect 16120 21616 16172 21622
rect 16120 21558 16172 21564
rect 16120 21480 16172 21486
rect 16120 21422 16172 21428
rect 16028 21344 16080 21350
rect 16028 21286 16080 21292
rect 16132 20874 16160 21422
rect 16304 21004 16356 21010
rect 16304 20946 16356 20952
rect 16120 20868 16172 20874
rect 16120 20810 16172 20816
rect 16028 20800 16080 20806
rect 16028 20742 16080 20748
rect 16212 20800 16264 20806
rect 16212 20742 16264 20748
rect 16040 19718 16068 20742
rect 16224 20534 16252 20742
rect 16212 20528 16264 20534
rect 16212 20470 16264 20476
rect 16120 19916 16172 19922
rect 16120 19858 16172 19864
rect 16028 19712 16080 19718
rect 16028 19654 16080 19660
rect 15936 18692 15988 18698
rect 15936 18634 15988 18640
rect 15948 18086 15976 18634
rect 15936 18080 15988 18086
rect 15936 18022 15988 18028
rect 15844 17672 15896 17678
rect 15844 17614 15896 17620
rect 16028 17604 16080 17610
rect 16028 17546 16080 17552
rect 15568 17536 15620 17542
rect 15568 17478 15620 17484
rect 16040 17338 16068 17546
rect 16028 17332 16080 17338
rect 16028 17274 16080 17280
rect 15476 16584 15528 16590
rect 15476 16526 15528 16532
rect 15292 16108 15344 16114
rect 15292 16050 15344 16056
rect 14945 15804 15253 15813
rect 14945 15802 14951 15804
rect 15007 15802 15031 15804
rect 15087 15802 15111 15804
rect 15167 15802 15191 15804
rect 15247 15802 15253 15804
rect 15007 15750 15009 15802
rect 15189 15750 15191 15802
rect 14945 15748 14951 15750
rect 15007 15748 15031 15750
rect 15087 15748 15111 15750
rect 15167 15748 15191 15750
rect 15247 15748 15253 15750
rect 14945 15739 15253 15748
rect 15304 15706 15332 16050
rect 16132 15910 16160 19858
rect 16224 19530 16252 20470
rect 16316 20330 16344 20946
rect 16408 20369 16436 22086
rect 16948 22034 17000 22040
rect 16486 21720 16542 21729
rect 16960 21690 16988 22034
rect 16486 21655 16542 21664
rect 16948 21684 17000 21690
rect 16500 21185 16528 21655
rect 16948 21626 17000 21632
rect 16764 21480 16816 21486
rect 16764 21422 16816 21428
rect 16776 21321 16804 21422
rect 16762 21312 16818 21321
rect 16762 21247 16818 21256
rect 16486 21176 16542 21185
rect 16486 21111 16542 21120
rect 16948 21072 17000 21078
rect 16948 21014 17000 21020
rect 16856 21004 16908 21010
rect 16856 20946 16908 20952
rect 16488 20800 16540 20806
rect 16488 20742 16540 20748
rect 16764 20800 16816 20806
rect 16764 20742 16816 20748
rect 16394 20360 16450 20369
rect 16304 20324 16356 20330
rect 16394 20295 16450 20304
rect 16304 20266 16356 20272
rect 16396 20256 16448 20262
rect 16396 20198 16448 20204
rect 16224 19502 16344 19530
rect 16408 19514 16436 20198
rect 16500 19854 16528 20742
rect 16776 20602 16804 20742
rect 16764 20596 16816 20602
rect 16764 20538 16816 20544
rect 16868 20482 16896 20946
rect 16580 20460 16632 20466
rect 16580 20402 16632 20408
rect 16776 20454 16896 20482
rect 16488 19848 16540 19854
rect 16488 19790 16540 19796
rect 16592 19514 16620 20402
rect 16672 20392 16724 20398
rect 16672 20334 16724 20340
rect 16684 19514 16712 20334
rect 16316 19446 16344 19502
rect 16396 19508 16448 19514
rect 16396 19450 16448 19456
rect 16580 19508 16632 19514
rect 16580 19450 16632 19456
rect 16672 19508 16724 19514
rect 16672 19450 16724 19456
rect 16304 19440 16356 19446
rect 16304 19382 16356 19388
rect 16776 17082 16804 20454
rect 16856 20392 16908 20398
rect 16856 20334 16908 20340
rect 16868 20058 16896 20334
rect 16856 20052 16908 20058
rect 16856 19994 16908 20000
rect 16960 18698 16988 21014
rect 17052 20505 17080 23800
rect 17316 22160 17368 22166
rect 17316 22102 17368 22108
rect 17406 22128 17462 22137
rect 17132 21888 17184 21894
rect 17132 21830 17184 21836
rect 17222 21856 17278 21865
rect 17144 21185 17172 21830
rect 17222 21791 17278 21800
rect 17236 21321 17264 21791
rect 17222 21312 17278 21321
rect 17222 21247 17278 21256
rect 17130 21176 17186 21185
rect 17130 21111 17186 21120
rect 17236 21078 17264 21247
rect 17224 21072 17276 21078
rect 17224 21014 17276 21020
rect 17038 20496 17094 20505
rect 17038 20431 17094 20440
rect 17224 20392 17276 20398
rect 17144 20352 17224 20380
rect 17040 19780 17092 19786
rect 17040 19722 17092 19728
rect 17052 19514 17080 19722
rect 17040 19508 17092 19514
rect 17040 19450 17092 19456
rect 16948 18692 17000 18698
rect 16948 18634 17000 18640
rect 16960 17882 16988 18634
rect 16948 17876 17000 17882
rect 16948 17818 17000 17824
rect 17040 17876 17092 17882
rect 17040 17818 17092 17824
rect 16948 17196 17000 17202
rect 16948 17138 17000 17144
rect 16684 17054 16804 17082
rect 16684 16522 16712 17054
rect 16764 16992 16816 16998
rect 16960 16980 16988 17138
rect 17052 16998 17080 17818
rect 17144 17338 17172 20352
rect 17224 20334 17276 20340
rect 17328 18970 17356 22102
rect 17406 22063 17462 22072
rect 17696 22094 17724 23800
rect 18340 22094 18368 23800
rect 18602 22128 18658 22137
rect 17696 22066 18000 22094
rect 18340 22066 18552 22094
rect 17420 21554 17448 22063
rect 17972 22030 18000 22066
rect 17960 22024 18012 22030
rect 17960 21966 18012 21972
rect 17592 21956 17644 21962
rect 17592 21898 17644 21904
rect 18144 21956 18196 21962
rect 18144 21898 18196 21904
rect 17500 21888 17552 21894
rect 17500 21830 17552 21836
rect 17408 21548 17460 21554
rect 17408 21490 17460 21496
rect 17408 21412 17460 21418
rect 17408 21354 17460 21360
rect 17420 20398 17448 21354
rect 17512 20942 17540 21830
rect 17604 21690 17632 21898
rect 17744 21788 18052 21797
rect 17744 21786 17750 21788
rect 17806 21786 17830 21788
rect 17886 21786 17910 21788
rect 17966 21786 17990 21788
rect 18046 21786 18052 21788
rect 17806 21734 17808 21786
rect 17988 21734 17990 21786
rect 17744 21732 17750 21734
rect 17806 21732 17830 21734
rect 17886 21732 17910 21734
rect 17966 21732 17990 21734
rect 18046 21732 18052 21734
rect 17744 21723 18052 21732
rect 17592 21684 17644 21690
rect 17592 21626 17644 21632
rect 17868 21344 17920 21350
rect 17866 21312 17868 21321
rect 17920 21312 17922 21321
rect 17866 21247 17922 21256
rect 18156 21146 18184 21898
rect 18236 21888 18288 21894
rect 18236 21830 18288 21836
rect 18328 21888 18380 21894
rect 18328 21830 18380 21836
rect 18248 21622 18276 21830
rect 18236 21616 18288 21622
rect 18236 21558 18288 21564
rect 18144 21140 18196 21146
rect 18144 21082 18196 21088
rect 18340 21078 18368 21830
rect 18418 21176 18474 21185
rect 18418 21111 18474 21120
rect 18328 21072 18380 21078
rect 18142 21040 18198 21049
rect 17592 21004 17644 21010
rect 17868 21004 17920 21010
rect 17644 20964 17868 20992
rect 17592 20946 17644 20952
rect 18328 21014 18380 21020
rect 18142 20975 18198 20984
rect 17868 20946 17920 20952
rect 17500 20936 17552 20942
rect 17500 20878 17552 20884
rect 17500 20800 17552 20806
rect 17684 20800 17736 20806
rect 17500 20742 17552 20748
rect 17604 20760 17684 20788
rect 17512 20602 17540 20742
rect 17500 20596 17552 20602
rect 17500 20538 17552 20544
rect 17408 20392 17460 20398
rect 17408 20334 17460 20340
rect 17604 20058 17632 20760
rect 17684 20742 17736 20748
rect 17744 20700 18052 20709
rect 17744 20698 17750 20700
rect 17806 20698 17830 20700
rect 17886 20698 17910 20700
rect 17966 20698 17990 20700
rect 18046 20698 18052 20700
rect 17806 20646 17808 20698
rect 17988 20646 17990 20698
rect 17744 20644 17750 20646
rect 17806 20644 17830 20646
rect 17886 20644 17910 20646
rect 17966 20644 17990 20646
rect 18046 20644 18052 20646
rect 17744 20635 18052 20644
rect 18156 20602 18184 20975
rect 18144 20596 18196 20602
rect 18144 20538 18196 20544
rect 18328 20392 18380 20398
rect 18328 20334 18380 20340
rect 18144 20256 18196 20262
rect 18144 20198 18196 20204
rect 17592 20052 17644 20058
rect 17592 19994 17644 20000
rect 18050 19952 18106 19961
rect 17500 19916 17552 19922
rect 18156 19922 18184 20198
rect 18050 19887 18106 19896
rect 18144 19916 18196 19922
rect 17500 19858 17552 19864
rect 17408 19372 17460 19378
rect 17408 19314 17460 19320
rect 17316 18964 17368 18970
rect 17316 18906 17368 18912
rect 17420 18850 17448 19314
rect 17328 18822 17448 18850
rect 17224 18624 17276 18630
rect 17224 18566 17276 18572
rect 17236 18290 17264 18566
rect 17224 18284 17276 18290
rect 17224 18226 17276 18232
rect 17328 18170 17356 18822
rect 17408 18624 17460 18630
rect 17408 18566 17460 18572
rect 17236 18142 17356 18170
rect 17236 17542 17264 18142
rect 17314 17640 17370 17649
rect 17314 17575 17370 17584
rect 17224 17536 17276 17542
rect 17224 17478 17276 17484
rect 17132 17332 17184 17338
rect 17132 17274 17184 17280
rect 16816 16952 16988 16980
rect 17040 16992 17092 16998
rect 16764 16934 16816 16940
rect 17040 16934 17092 16940
rect 16672 16516 16724 16522
rect 16672 16458 16724 16464
rect 16304 16448 16356 16454
rect 16304 16390 16356 16396
rect 16316 16250 16344 16390
rect 16304 16244 16356 16250
rect 16304 16186 16356 16192
rect 16120 15904 16172 15910
rect 16120 15846 16172 15852
rect 15292 15700 15344 15706
rect 15292 15642 15344 15648
rect 16684 15434 16712 16458
rect 16672 15428 16724 15434
rect 16672 15370 16724 15376
rect 16592 14958 16620 14989
rect 16580 14952 16632 14958
rect 16578 14920 16580 14929
rect 16632 14920 16634 14929
rect 16578 14855 16634 14864
rect 14945 14716 15253 14725
rect 14945 14714 14951 14716
rect 15007 14714 15031 14716
rect 15087 14714 15111 14716
rect 15167 14714 15191 14716
rect 15247 14714 15253 14716
rect 15007 14662 15009 14714
rect 15189 14662 15191 14714
rect 14945 14660 14951 14662
rect 15007 14660 15031 14662
rect 15087 14660 15111 14662
rect 15167 14660 15191 14662
rect 15247 14660 15253 14662
rect 14945 14651 15253 14660
rect 16592 14618 16620 14855
rect 16580 14612 16632 14618
rect 16580 14554 16632 14560
rect 14738 14376 14794 14385
rect 14738 14311 14740 14320
rect 14792 14311 14794 14320
rect 16672 14340 16724 14346
rect 14740 14282 14792 14288
rect 16672 14282 16724 14288
rect 14752 14074 14780 14282
rect 15752 14272 15804 14278
rect 15752 14214 15804 14220
rect 14740 14068 14792 14074
rect 14740 14010 14792 14016
rect 15384 13932 15436 13938
rect 15384 13874 15436 13880
rect 14945 13628 15253 13637
rect 14945 13626 14951 13628
rect 15007 13626 15031 13628
rect 15087 13626 15111 13628
rect 15167 13626 15191 13628
rect 15247 13626 15253 13628
rect 15007 13574 15009 13626
rect 15189 13574 15191 13626
rect 14945 13572 14951 13574
rect 15007 13572 15031 13574
rect 15087 13572 15111 13574
rect 15167 13572 15191 13574
rect 15247 13572 15253 13574
rect 14945 13563 15253 13572
rect 14945 12540 15253 12549
rect 14945 12538 14951 12540
rect 15007 12538 15031 12540
rect 15087 12538 15111 12540
rect 15167 12538 15191 12540
rect 15247 12538 15253 12540
rect 15007 12486 15009 12538
rect 15189 12486 15191 12538
rect 14945 12484 14951 12486
rect 15007 12484 15031 12486
rect 15087 12484 15111 12486
rect 15167 12484 15191 12486
rect 15247 12484 15253 12486
rect 14945 12475 15253 12484
rect 15396 12434 15424 13874
rect 15764 13734 15792 14214
rect 16684 13938 16712 14282
rect 16672 13932 16724 13938
rect 16672 13874 16724 13880
rect 15752 13728 15804 13734
rect 15752 13670 15804 13676
rect 15660 13252 15712 13258
rect 15764 13240 15792 13670
rect 16578 13288 16634 13297
rect 15712 13212 15792 13240
rect 16120 13252 16172 13258
rect 15660 13194 15712 13200
rect 16578 13223 16634 13232
rect 16120 13194 16172 13200
rect 16132 12714 16160 13194
rect 16212 12980 16264 12986
rect 16212 12922 16264 12928
rect 16120 12708 16172 12714
rect 16120 12650 16172 12656
rect 14568 12406 14688 12434
rect 15304 12406 15424 12434
rect 14462 7440 14518 7449
rect 14462 7375 14518 7384
rect 13544 6248 13596 6254
rect 13544 6190 13596 6196
rect 13820 6248 13872 6254
rect 13820 6190 13872 6196
rect 14370 6216 14426 6225
rect 14370 6151 14372 6160
rect 14424 6151 14426 6160
rect 14372 6122 14424 6128
rect 14568 5574 14596 12406
rect 15304 11558 15332 12406
rect 16224 12306 16252 12922
rect 16592 12850 16620 13223
rect 16580 12844 16632 12850
rect 16580 12786 16632 12792
rect 16580 12640 16632 12646
rect 16580 12582 16632 12588
rect 16592 12442 16620 12582
rect 16580 12436 16632 12442
rect 16776 12434 16804 16934
rect 17144 16794 17172 17274
rect 17132 16788 17184 16794
rect 17132 16730 17184 16736
rect 16948 14476 17000 14482
rect 16948 14418 17000 14424
rect 16960 14074 16988 14418
rect 17236 14414 17264 17478
rect 17328 17338 17356 17575
rect 17420 17338 17448 18566
rect 17316 17332 17368 17338
rect 17316 17274 17368 17280
rect 17408 17332 17460 17338
rect 17408 17274 17460 17280
rect 17408 17060 17460 17066
rect 17408 17002 17460 17008
rect 17224 14408 17276 14414
rect 17224 14350 17276 14356
rect 16948 14068 17000 14074
rect 16948 14010 17000 14016
rect 17040 13320 17092 13326
rect 17040 13262 17092 13268
rect 17052 12986 17080 13262
rect 17040 12980 17092 12986
rect 17040 12922 17092 12928
rect 17420 12434 17448 17002
rect 17512 16590 17540 19858
rect 18064 19854 18092 19887
rect 18144 19858 18196 19864
rect 18340 19854 18368 20334
rect 18432 19854 18460 21111
rect 18524 21026 18552 22066
rect 18602 22063 18658 22072
rect 18616 21146 18644 22063
rect 18880 22024 18932 22030
rect 18880 21966 18932 21972
rect 18696 21888 18748 21894
rect 18696 21830 18748 21836
rect 18604 21140 18656 21146
rect 18604 21082 18656 21088
rect 18524 20998 18644 21026
rect 18616 20942 18644 20998
rect 18512 20936 18564 20942
rect 18512 20878 18564 20884
rect 18604 20936 18656 20942
rect 18604 20878 18656 20884
rect 18524 20505 18552 20878
rect 18510 20496 18566 20505
rect 18510 20431 18566 20440
rect 18512 20392 18564 20398
rect 18512 20334 18564 20340
rect 18052 19848 18104 19854
rect 18052 19790 18104 19796
rect 18328 19848 18380 19854
rect 18328 19790 18380 19796
rect 18420 19848 18472 19854
rect 18420 19790 18472 19796
rect 17744 19612 18052 19621
rect 17744 19610 17750 19612
rect 17806 19610 17830 19612
rect 17886 19610 17910 19612
rect 17966 19610 17990 19612
rect 18046 19610 18052 19612
rect 17806 19558 17808 19610
rect 17988 19558 17990 19610
rect 17744 19556 17750 19558
rect 17806 19556 17830 19558
rect 17886 19556 17910 19558
rect 17966 19556 17990 19558
rect 18046 19556 18052 19558
rect 17744 19547 18052 19556
rect 18524 19514 18552 20334
rect 18616 19825 18644 20878
rect 18602 19816 18658 19825
rect 18708 19786 18736 21830
rect 18892 21690 18920 21966
rect 18880 21684 18932 21690
rect 18880 21626 18932 21632
rect 18984 21146 19012 23800
rect 19064 22840 19116 22846
rect 19064 22782 19116 22788
rect 19076 21554 19104 22782
rect 19340 22636 19392 22642
rect 19340 22578 19392 22584
rect 19156 22160 19208 22166
rect 19156 22102 19208 22108
rect 19064 21548 19116 21554
rect 19064 21490 19116 21496
rect 18972 21140 19024 21146
rect 18972 21082 19024 21088
rect 18880 20936 18932 20942
rect 18880 20878 18932 20884
rect 18788 20052 18840 20058
rect 18892 20040 18920 20878
rect 18840 20012 18920 20040
rect 18788 19994 18840 20000
rect 19168 19802 19196 22102
rect 19352 22030 19380 22578
rect 19340 22024 19392 22030
rect 19340 21966 19392 21972
rect 19352 21690 19380 21966
rect 19628 21894 19656 23800
rect 20168 22772 20220 22778
rect 20168 22714 20220 22720
rect 19708 22704 19760 22710
rect 19708 22646 19760 22652
rect 19720 22030 19748 22646
rect 20180 22030 20208 22714
rect 19708 22024 19760 22030
rect 19708 21966 19760 21972
rect 20168 22024 20220 22030
rect 20168 21966 20220 21972
rect 20272 21894 20300 23800
rect 20543 22332 20851 22341
rect 20543 22330 20549 22332
rect 20605 22330 20629 22332
rect 20685 22330 20709 22332
rect 20765 22330 20789 22332
rect 20845 22330 20851 22332
rect 20605 22278 20607 22330
rect 20787 22278 20789 22330
rect 20543 22276 20549 22278
rect 20605 22276 20629 22278
rect 20685 22276 20709 22278
rect 20765 22276 20789 22278
rect 20845 22276 20851 22278
rect 20543 22267 20851 22276
rect 20534 22128 20590 22137
rect 20534 22063 20590 22072
rect 19616 21888 19668 21894
rect 19616 21830 19668 21836
rect 20260 21888 20312 21894
rect 20260 21830 20312 21836
rect 20548 21690 20576 22063
rect 20916 21894 20944 23800
rect 20996 22500 21048 22506
rect 20996 22442 21048 22448
rect 21008 22030 21036 22442
rect 20996 22024 21048 22030
rect 20996 21966 21048 21972
rect 21088 22024 21140 22030
rect 21456 22024 21508 22030
rect 21088 21966 21140 21972
rect 21376 21984 21456 22012
rect 20812 21888 20864 21894
rect 20812 21830 20864 21836
rect 20904 21888 20956 21894
rect 20904 21830 20956 21836
rect 19340 21684 19392 21690
rect 19340 21626 19392 21632
rect 20536 21684 20588 21690
rect 20536 21626 20588 21632
rect 20628 21684 20680 21690
rect 20628 21626 20680 21632
rect 19892 21548 19944 21554
rect 19892 21490 19944 21496
rect 20352 21548 20404 21554
rect 20352 21490 20404 21496
rect 19524 21480 19576 21486
rect 19524 21422 19576 21428
rect 18602 19751 18658 19760
rect 18696 19780 18748 19786
rect 18696 19722 18748 19728
rect 19076 19774 19196 19802
rect 19248 19848 19300 19854
rect 19248 19790 19300 19796
rect 18144 19508 18196 19514
rect 18144 19450 18196 19456
rect 18512 19508 18564 19514
rect 18512 19450 18564 19456
rect 17592 18692 17644 18698
rect 17592 18634 17644 18640
rect 17604 18426 17632 18634
rect 17744 18524 18052 18533
rect 17744 18522 17750 18524
rect 17806 18522 17830 18524
rect 17886 18522 17910 18524
rect 17966 18522 17990 18524
rect 18046 18522 18052 18524
rect 17806 18470 17808 18522
rect 17988 18470 17990 18522
rect 17744 18468 17750 18470
rect 17806 18468 17830 18470
rect 17886 18468 17910 18470
rect 17966 18468 17990 18470
rect 18046 18468 18052 18470
rect 17744 18459 18052 18468
rect 17592 18420 17644 18426
rect 17592 18362 17644 18368
rect 18156 17678 18184 19450
rect 19076 19378 19104 19774
rect 19156 19712 19208 19718
rect 19156 19654 19208 19660
rect 19064 19372 19116 19378
rect 19064 19314 19116 19320
rect 18878 19272 18934 19281
rect 18878 19207 18934 19216
rect 18512 19168 18564 19174
rect 18512 19110 18564 19116
rect 18524 18358 18552 19110
rect 18892 18766 18920 19207
rect 18880 18760 18932 18766
rect 18880 18702 18932 18708
rect 18602 18592 18658 18601
rect 18602 18527 18658 18536
rect 18512 18352 18564 18358
rect 18512 18294 18564 18300
rect 18420 17740 18472 17746
rect 18420 17682 18472 17688
rect 18144 17672 18196 17678
rect 18144 17614 18196 17620
rect 17744 17436 18052 17445
rect 17744 17434 17750 17436
rect 17806 17434 17830 17436
rect 17886 17434 17910 17436
rect 17966 17434 17990 17436
rect 18046 17434 18052 17436
rect 17806 17382 17808 17434
rect 17988 17382 17990 17434
rect 17744 17380 17750 17382
rect 17806 17380 17830 17382
rect 17886 17380 17910 17382
rect 17966 17380 17990 17382
rect 18046 17380 18052 17382
rect 17744 17371 18052 17380
rect 17960 17332 18012 17338
rect 17960 17274 18012 17280
rect 17592 17196 17644 17202
rect 17592 17138 17644 17144
rect 17868 17196 17920 17202
rect 17972 17184 18000 17274
rect 18432 17270 18460 17682
rect 18512 17604 18564 17610
rect 18512 17546 18564 17552
rect 18524 17513 18552 17546
rect 18510 17504 18566 17513
rect 18510 17439 18566 17448
rect 18512 17332 18564 17338
rect 18512 17274 18564 17280
rect 18420 17264 18472 17270
rect 18420 17206 18472 17212
rect 17920 17156 18000 17184
rect 17868 17138 17920 17144
rect 17500 16584 17552 16590
rect 17500 16526 17552 16532
rect 17512 15638 17540 16526
rect 17500 15632 17552 15638
rect 17500 15574 17552 15580
rect 17604 12434 17632 17138
rect 18432 16794 18460 17206
rect 18420 16788 18472 16794
rect 18420 16730 18472 16736
rect 18144 16584 18196 16590
rect 18144 16526 18196 16532
rect 17744 16348 18052 16357
rect 17744 16346 17750 16348
rect 17806 16346 17830 16348
rect 17886 16346 17910 16348
rect 17966 16346 17990 16348
rect 18046 16346 18052 16348
rect 17806 16294 17808 16346
rect 17988 16294 17990 16346
rect 17744 16292 17750 16294
rect 17806 16292 17830 16294
rect 17886 16292 17910 16294
rect 17966 16292 17990 16294
rect 18046 16292 18052 16294
rect 17744 16283 18052 16292
rect 18156 16182 18184 16526
rect 18432 16250 18460 16730
rect 18524 16697 18552 17274
rect 18510 16688 18566 16697
rect 18510 16623 18566 16632
rect 18420 16244 18472 16250
rect 18420 16186 18472 16192
rect 18144 16176 18196 16182
rect 18144 16118 18196 16124
rect 18524 16046 18552 16623
rect 18616 16454 18644 18527
rect 18892 18193 18920 18702
rect 18972 18352 19024 18358
rect 18972 18294 19024 18300
rect 18878 18184 18934 18193
rect 18878 18119 18934 18128
rect 18880 17672 18932 17678
rect 18880 17614 18932 17620
rect 18604 16448 18656 16454
rect 18604 16390 18656 16396
rect 18604 16244 18656 16250
rect 18604 16186 18656 16192
rect 18512 16040 18564 16046
rect 18512 15982 18564 15988
rect 18420 15904 18472 15910
rect 18420 15846 18472 15852
rect 18236 15700 18288 15706
rect 18236 15642 18288 15648
rect 17744 15260 18052 15269
rect 17744 15258 17750 15260
rect 17806 15258 17830 15260
rect 17886 15258 17910 15260
rect 17966 15258 17990 15260
rect 18046 15258 18052 15260
rect 17806 15206 17808 15258
rect 17988 15206 17990 15258
rect 17744 15204 17750 15206
rect 17806 15204 17830 15206
rect 17886 15204 17910 15206
rect 17966 15204 17990 15206
rect 18046 15204 18052 15206
rect 17744 15195 18052 15204
rect 18144 14816 18196 14822
rect 18144 14758 18196 14764
rect 17744 14172 18052 14181
rect 17744 14170 17750 14172
rect 17806 14170 17830 14172
rect 17886 14170 17910 14172
rect 17966 14170 17990 14172
rect 18046 14170 18052 14172
rect 17806 14118 17808 14170
rect 17988 14118 17990 14170
rect 17744 14116 17750 14118
rect 17806 14116 17830 14118
rect 17886 14116 17910 14118
rect 17966 14116 17990 14118
rect 18046 14116 18052 14118
rect 17744 14107 18052 14116
rect 18156 14074 18184 14758
rect 18144 14068 18196 14074
rect 18144 14010 18196 14016
rect 18144 13456 18196 13462
rect 18144 13398 18196 13404
rect 17744 13084 18052 13093
rect 17744 13082 17750 13084
rect 17806 13082 17830 13084
rect 17886 13082 17910 13084
rect 17966 13082 17990 13084
rect 18046 13082 18052 13084
rect 17806 13030 17808 13082
rect 17988 13030 17990 13082
rect 17744 13028 17750 13030
rect 17806 13028 17830 13030
rect 17886 13028 17910 13030
rect 17966 13028 17990 13030
rect 18046 13028 18052 13030
rect 17744 13019 18052 13028
rect 18156 12918 18184 13398
rect 18144 12912 18196 12918
rect 18144 12854 18196 12860
rect 16776 12406 16896 12434
rect 16580 12378 16632 12384
rect 16212 12300 16264 12306
rect 16212 12242 16264 12248
rect 16592 12238 16620 12378
rect 16580 12232 16632 12238
rect 16580 12174 16632 12180
rect 15752 11756 15804 11762
rect 15752 11698 15804 11704
rect 15292 11552 15344 11558
rect 15292 11494 15344 11500
rect 14945 11452 15253 11461
rect 14945 11450 14951 11452
rect 15007 11450 15031 11452
rect 15087 11450 15111 11452
rect 15167 11450 15191 11452
rect 15247 11450 15253 11452
rect 15007 11398 15009 11450
rect 15189 11398 15191 11450
rect 14945 11396 14951 11398
rect 15007 11396 15031 11398
rect 15087 11396 15111 11398
rect 15167 11396 15191 11398
rect 15247 11396 15253 11398
rect 14945 11387 15253 11396
rect 15016 11144 15068 11150
rect 15016 11086 15068 11092
rect 15028 10674 15056 11086
rect 15016 10668 15068 10674
rect 15016 10610 15068 10616
rect 14945 10364 15253 10373
rect 14945 10362 14951 10364
rect 15007 10362 15031 10364
rect 15087 10362 15111 10364
rect 15167 10362 15191 10364
rect 15247 10362 15253 10364
rect 15007 10310 15009 10362
rect 15189 10310 15191 10362
rect 14945 10308 14951 10310
rect 15007 10308 15031 10310
rect 15087 10308 15111 10310
rect 15167 10308 15191 10310
rect 15247 10308 15253 10310
rect 14945 10299 15253 10308
rect 14945 9276 15253 9285
rect 14945 9274 14951 9276
rect 15007 9274 15031 9276
rect 15087 9274 15111 9276
rect 15167 9274 15191 9276
rect 15247 9274 15253 9276
rect 15007 9222 15009 9274
rect 15189 9222 15191 9274
rect 14945 9220 14951 9222
rect 15007 9220 15031 9222
rect 15087 9220 15111 9222
rect 15167 9220 15191 9222
rect 15247 9220 15253 9222
rect 14945 9211 15253 9220
rect 14945 8188 15253 8197
rect 14945 8186 14951 8188
rect 15007 8186 15031 8188
rect 15087 8186 15111 8188
rect 15167 8186 15191 8188
rect 15247 8186 15253 8188
rect 15007 8134 15009 8186
rect 15189 8134 15191 8186
rect 14945 8132 14951 8134
rect 15007 8132 15031 8134
rect 15087 8132 15111 8134
rect 15167 8132 15191 8134
rect 15247 8132 15253 8134
rect 14945 8123 15253 8132
rect 14740 7744 14792 7750
rect 14740 7686 14792 7692
rect 14752 7410 14780 7686
rect 14740 7404 14792 7410
rect 14740 7346 14792 7352
rect 14752 6730 14780 7346
rect 14945 7100 15253 7109
rect 14945 7098 14951 7100
rect 15007 7098 15031 7100
rect 15087 7098 15111 7100
rect 15167 7098 15191 7100
rect 15247 7098 15253 7100
rect 15007 7046 15009 7098
rect 15189 7046 15191 7098
rect 14945 7044 14951 7046
rect 15007 7044 15031 7046
rect 15087 7044 15111 7046
rect 15167 7044 15191 7046
rect 15247 7044 15253 7046
rect 14945 7035 15253 7044
rect 14740 6724 14792 6730
rect 14740 6666 14792 6672
rect 15304 6186 15332 11494
rect 15384 9580 15436 9586
rect 15384 9522 15436 9528
rect 15396 8838 15424 9522
rect 15384 8832 15436 8838
rect 15384 8774 15436 8780
rect 15764 8634 15792 11698
rect 16396 11620 16448 11626
rect 16396 11562 16448 11568
rect 16120 11552 16172 11558
rect 16120 11494 16172 11500
rect 16132 11150 16160 11494
rect 16408 11354 16436 11562
rect 16488 11552 16540 11558
rect 16488 11494 16540 11500
rect 16500 11354 16528 11494
rect 16396 11348 16448 11354
rect 16396 11290 16448 11296
rect 16488 11348 16540 11354
rect 16488 11290 16540 11296
rect 16120 11144 16172 11150
rect 16120 11086 16172 11092
rect 16132 10742 16160 11086
rect 16396 11008 16448 11014
rect 16396 10950 16448 10956
rect 16120 10736 16172 10742
rect 16120 10678 16172 10684
rect 16408 9994 16436 10950
rect 16764 10668 16816 10674
rect 16764 10610 16816 10616
rect 16580 10464 16632 10470
rect 16580 10406 16632 10412
rect 16592 10169 16620 10406
rect 16578 10160 16634 10169
rect 16578 10095 16634 10104
rect 16776 10010 16804 10610
rect 16396 9988 16448 9994
rect 16396 9930 16448 9936
rect 16592 9982 16804 10010
rect 16868 10010 16896 12406
rect 17236 12406 17448 12434
rect 17512 12406 17632 12434
rect 17132 11552 17184 11558
rect 17132 11494 17184 11500
rect 17040 11008 17092 11014
rect 17040 10950 17092 10956
rect 17052 10742 17080 10950
rect 17040 10736 17092 10742
rect 17040 10678 17092 10684
rect 17052 10198 17080 10678
rect 17040 10192 17092 10198
rect 17040 10134 17092 10140
rect 16868 9982 17080 10010
rect 16304 9444 16356 9450
rect 16304 9386 16356 9392
rect 16316 8974 16344 9386
rect 16408 8974 16436 9930
rect 16592 9382 16620 9982
rect 16580 9376 16632 9382
rect 16580 9318 16632 9324
rect 16304 8968 16356 8974
rect 16304 8910 16356 8916
rect 16396 8968 16448 8974
rect 16396 8910 16448 8916
rect 15936 8900 15988 8906
rect 15936 8842 15988 8848
rect 15752 8628 15804 8634
rect 15752 8570 15804 8576
rect 15844 7200 15896 7206
rect 15844 7142 15896 7148
rect 15856 6746 15884 7142
rect 15764 6730 15884 6746
rect 15752 6724 15884 6730
rect 15804 6718 15884 6724
rect 15752 6666 15804 6672
rect 15752 6452 15804 6458
rect 15752 6394 15804 6400
rect 15384 6384 15436 6390
rect 15384 6326 15436 6332
rect 15292 6180 15344 6186
rect 15292 6122 15344 6128
rect 14648 6112 14700 6118
rect 14648 6054 14700 6060
rect 14660 5778 14688 6054
rect 14945 6012 15253 6021
rect 14945 6010 14951 6012
rect 15007 6010 15031 6012
rect 15087 6010 15111 6012
rect 15167 6010 15191 6012
rect 15247 6010 15253 6012
rect 15007 5958 15009 6010
rect 15189 5958 15191 6010
rect 14945 5956 14951 5958
rect 15007 5956 15031 5958
rect 15087 5956 15111 5958
rect 15167 5956 15191 5958
rect 15247 5956 15253 5958
rect 14945 5947 15253 5956
rect 14648 5772 14700 5778
rect 14648 5714 14700 5720
rect 15108 5704 15160 5710
rect 15108 5646 15160 5652
rect 13820 5568 13872 5574
rect 13820 5510 13872 5516
rect 14556 5568 14608 5574
rect 14556 5510 14608 5516
rect 12072 5364 12124 5370
rect 12072 5306 12124 5312
rect 13176 5364 13228 5370
rect 13176 5306 13228 5312
rect 13832 4622 13860 5510
rect 14568 5302 14596 5510
rect 14556 5296 14608 5302
rect 14556 5238 14608 5244
rect 15120 5250 15148 5646
rect 15396 5370 15424 6326
rect 15660 6316 15712 6322
rect 15660 6258 15712 6264
rect 15672 5370 15700 6258
rect 15384 5364 15436 5370
rect 15384 5306 15436 5312
rect 15660 5364 15712 5370
rect 15660 5306 15712 5312
rect 15120 5234 15240 5250
rect 14832 5228 14884 5234
rect 15120 5228 15252 5234
rect 15120 5222 15200 5228
rect 14832 5170 14884 5176
rect 15200 5170 15252 5176
rect 14188 5024 14240 5030
rect 14188 4966 14240 4972
rect 13820 4616 13872 4622
rect 13820 4558 13872 4564
rect 13728 4548 13780 4554
rect 13728 4490 13780 4496
rect 12146 4380 12454 4389
rect 12146 4378 12152 4380
rect 12208 4378 12232 4380
rect 12288 4378 12312 4380
rect 12368 4378 12392 4380
rect 12448 4378 12454 4380
rect 12208 4326 12210 4378
rect 12390 4326 12392 4378
rect 12146 4324 12152 4326
rect 12208 4324 12232 4326
rect 12288 4324 12312 4326
rect 12368 4324 12392 4326
rect 12448 4324 12454 4326
rect 12146 4315 12454 4324
rect 13740 4185 13768 4490
rect 13726 4176 13782 4185
rect 13726 4111 13782 4120
rect 14200 4010 14228 4966
rect 14844 4826 14872 5170
rect 15660 5024 15712 5030
rect 15660 4966 15712 4972
rect 14945 4924 15253 4933
rect 14945 4922 14951 4924
rect 15007 4922 15031 4924
rect 15087 4922 15111 4924
rect 15167 4922 15191 4924
rect 15247 4922 15253 4924
rect 15007 4870 15009 4922
rect 15189 4870 15191 4922
rect 14945 4868 14951 4870
rect 15007 4868 15031 4870
rect 15087 4868 15111 4870
rect 15167 4868 15191 4870
rect 15247 4868 15253 4870
rect 14945 4859 15253 4868
rect 14832 4820 14884 4826
rect 14832 4762 14884 4768
rect 15568 4480 15620 4486
rect 15568 4422 15620 4428
rect 15580 4282 15608 4422
rect 15568 4276 15620 4282
rect 15568 4218 15620 4224
rect 15672 4214 15700 4966
rect 15660 4208 15712 4214
rect 15660 4150 15712 4156
rect 15568 4072 15620 4078
rect 15568 4014 15620 4020
rect 14188 4004 14240 4010
rect 14188 3946 14240 3952
rect 14945 3836 15253 3845
rect 14945 3834 14951 3836
rect 15007 3834 15031 3836
rect 15087 3834 15111 3836
rect 15167 3834 15191 3836
rect 15247 3834 15253 3836
rect 15007 3782 15009 3834
rect 15189 3782 15191 3834
rect 14945 3780 14951 3782
rect 15007 3780 15031 3782
rect 15087 3780 15111 3782
rect 15167 3780 15191 3782
rect 15247 3780 15253 3782
rect 14945 3771 15253 3780
rect 15580 3641 15608 4014
rect 15566 3632 15622 3641
rect 15566 3567 15622 3576
rect 15764 3398 15792 6394
rect 15856 6322 15884 6718
rect 15948 6662 15976 8842
rect 16212 8628 16264 8634
rect 16212 8570 16264 8576
rect 16028 8356 16080 8362
rect 16028 8298 16080 8304
rect 16040 7546 16068 8298
rect 16028 7540 16080 7546
rect 16028 7482 16080 7488
rect 16040 7342 16068 7482
rect 16028 7336 16080 7342
rect 16028 7278 16080 7284
rect 16040 6866 16068 7278
rect 16028 6860 16080 6866
rect 16028 6802 16080 6808
rect 15936 6656 15988 6662
rect 15936 6598 15988 6604
rect 15948 6458 15976 6598
rect 15936 6452 15988 6458
rect 15936 6394 15988 6400
rect 15844 6316 15896 6322
rect 15844 6258 15896 6264
rect 16120 5772 16172 5778
rect 16120 5714 16172 5720
rect 16028 5228 16080 5234
rect 16028 5170 16080 5176
rect 16040 5030 16068 5170
rect 16028 5024 16080 5030
rect 16028 4966 16080 4972
rect 16132 4078 16160 5714
rect 16224 5166 16252 8570
rect 16316 8362 16344 8910
rect 16396 8832 16448 8838
rect 16396 8774 16448 8780
rect 16304 8356 16356 8362
rect 16304 8298 16356 8304
rect 16316 7886 16344 8298
rect 16408 8294 16436 8774
rect 16592 8498 16620 9318
rect 16488 8492 16540 8498
rect 16488 8434 16540 8440
rect 16580 8492 16632 8498
rect 16580 8434 16632 8440
rect 16500 8401 16528 8434
rect 16486 8392 16542 8401
rect 16486 8327 16542 8336
rect 16396 8288 16448 8294
rect 16448 8248 16620 8276
rect 16396 8230 16448 8236
rect 16408 8165 16436 8230
rect 16304 7880 16356 7886
rect 16304 7822 16356 7828
rect 16304 7404 16356 7410
rect 16304 7346 16356 7352
rect 16316 6254 16344 7346
rect 16396 6724 16448 6730
rect 16396 6666 16448 6672
rect 16488 6724 16540 6730
rect 16488 6666 16540 6672
rect 16408 6361 16436 6666
rect 16500 6458 16528 6666
rect 16488 6452 16540 6458
rect 16488 6394 16540 6400
rect 16394 6352 16450 6361
rect 16394 6287 16450 6296
rect 16304 6248 16356 6254
rect 16304 6190 16356 6196
rect 16212 5160 16264 5166
rect 16212 5102 16264 5108
rect 16120 4072 16172 4078
rect 16120 4014 16172 4020
rect 16212 3528 16264 3534
rect 16316 3505 16344 6190
rect 16592 5778 16620 8248
rect 16672 7744 16724 7750
rect 16672 7686 16724 7692
rect 16684 6254 16712 7686
rect 16946 7304 17002 7313
rect 16946 7239 17002 7248
rect 16764 6384 16816 6390
rect 16960 6338 16988 7239
rect 16764 6326 16816 6332
rect 16672 6248 16724 6254
rect 16672 6190 16724 6196
rect 16580 5772 16632 5778
rect 16580 5714 16632 5720
rect 16396 5704 16448 5710
rect 16396 5646 16448 5652
rect 16408 5302 16436 5646
rect 16672 5568 16724 5574
rect 16672 5510 16724 5516
rect 16396 5296 16448 5302
rect 16396 5238 16448 5244
rect 16580 5296 16632 5302
rect 16580 5238 16632 5244
rect 16592 5166 16620 5238
rect 16580 5160 16632 5166
rect 16580 5102 16632 5108
rect 16684 4690 16712 5510
rect 16672 4684 16724 4690
rect 16672 4626 16724 4632
rect 16776 4622 16804 6326
rect 16868 6310 16988 6338
rect 16868 5250 16896 6310
rect 16948 6248 17000 6254
rect 17052 6225 17080 9982
rect 17144 6361 17172 11494
rect 17236 6769 17264 12406
rect 17408 10464 17460 10470
rect 17408 10406 17460 10412
rect 17316 9920 17368 9926
rect 17316 9862 17368 9868
rect 17222 6760 17278 6769
rect 17222 6695 17278 6704
rect 17130 6352 17186 6361
rect 17130 6287 17186 6296
rect 16948 6190 17000 6196
rect 17038 6216 17094 6225
rect 16960 5370 16988 6190
rect 17038 6151 17094 6160
rect 17040 6112 17092 6118
rect 17040 6054 17092 6060
rect 16948 5364 17000 5370
rect 16948 5306 17000 5312
rect 16868 5222 16988 5250
rect 16856 5160 16908 5166
rect 16856 5102 16908 5108
rect 16764 4616 16816 4622
rect 16764 4558 16816 4564
rect 16868 4486 16896 5102
rect 16856 4480 16908 4486
rect 16856 4422 16908 4428
rect 16672 3936 16724 3942
rect 16672 3878 16724 3884
rect 16580 3528 16632 3534
rect 16212 3470 16264 3476
rect 16302 3496 16358 3505
rect 15752 3392 15804 3398
rect 15752 3334 15804 3340
rect 12146 3292 12454 3301
rect 12146 3290 12152 3292
rect 12208 3290 12232 3292
rect 12288 3290 12312 3292
rect 12368 3290 12392 3292
rect 12448 3290 12454 3292
rect 12208 3238 12210 3290
rect 12390 3238 12392 3290
rect 12146 3236 12152 3238
rect 12208 3236 12232 3238
rect 12288 3236 12312 3238
rect 12368 3236 12392 3238
rect 12448 3236 12454 3238
rect 12146 3227 12454 3236
rect 8392 2848 8444 2854
rect 8392 2790 8444 2796
rect 10784 2848 10836 2854
rect 10784 2790 10836 2796
rect 11980 2848 12032 2854
rect 11980 2790 12032 2796
rect 3749 2748 4057 2757
rect 3749 2746 3755 2748
rect 3811 2746 3835 2748
rect 3891 2746 3915 2748
rect 3971 2746 3995 2748
rect 4051 2746 4057 2748
rect 3811 2694 3813 2746
rect 3993 2694 3995 2746
rect 3749 2692 3755 2694
rect 3811 2692 3835 2694
rect 3891 2692 3915 2694
rect 3971 2692 3995 2694
rect 4051 2692 4057 2694
rect 3749 2683 4057 2692
rect 8404 2514 8432 2790
rect 9347 2748 9655 2757
rect 9347 2746 9353 2748
rect 9409 2746 9433 2748
rect 9489 2746 9513 2748
rect 9569 2746 9593 2748
rect 9649 2746 9655 2748
rect 9409 2694 9411 2746
rect 9591 2694 9593 2746
rect 9347 2692 9353 2694
rect 9409 2692 9433 2694
rect 9489 2692 9513 2694
rect 9569 2692 9593 2694
rect 9649 2692 9655 2694
rect 9347 2683 9655 2692
rect 10796 2650 10824 2790
rect 14945 2748 15253 2757
rect 14945 2746 14951 2748
rect 15007 2746 15031 2748
rect 15087 2746 15111 2748
rect 15167 2746 15191 2748
rect 15247 2746 15253 2748
rect 15007 2694 15009 2746
rect 15189 2694 15191 2746
rect 14945 2692 14951 2694
rect 15007 2692 15031 2694
rect 15087 2692 15111 2694
rect 15167 2692 15191 2694
rect 15247 2692 15253 2694
rect 14945 2683 15253 2692
rect 15764 2650 15792 3334
rect 16224 3126 16252 3470
rect 16580 3470 16632 3476
rect 16302 3431 16358 3440
rect 16212 3120 16264 3126
rect 16212 3062 16264 3068
rect 16592 2990 16620 3470
rect 16684 3097 16712 3878
rect 16868 3602 16896 4422
rect 16960 4146 16988 5222
rect 17052 4690 17080 6054
rect 17236 5574 17264 6695
rect 17328 6066 17356 9862
rect 17420 9382 17448 10406
rect 17512 9722 17540 12406
rect 18248 12209 18276 15642
rect 18432 15502 18460 15846
rect 18616 15706 18644 16186
rect 18604 15700 18656 15706
rect 18604 15642 18656 15648
rect 18420 15496 18472 15502
rect 18420 15438 18472 15444
rect 18616 15162 18644 15642
rect 18892 15609 18920 17614
rect 18878 15600 18934 15609
rect 18878 15535 18934 15544
rect 18880 15496 18932 15502
rect 18880 15438 18932 15444
rect 18420 15156 18472 15162
rect 18420 15098 18472 15104
rect 18604 15156 18656 15162
rect 18604 15098 18656 15104
rect 18432 15026 18460 15098
rect 18420 15020 18472 15026
rect 18420 14962 18472 14968
rect 18432 14618 18460 14962
rect 18420 14612 18472 14618
rect 18420 14554 18472 14560
rect 18892 14550 18920 15438
rect 18880 14544 18932 14550
rect 18880 14486 18932 14492
rect 18880 14068 18932 14074
rect 18880 14010 18932 14016
rect 18604 13388 18656 13394
rect 18604 13330 18656 13336
rect 18512 13320 18564 13326
rect 18512 13262 18564 13268
rect 18420 12844 18472 12850
rect 18420 12786 18472 12792
rect 18234 12200 18290 12209
rect 18432 12186 18460 12786
rect 18524 12753 18552 13262
rect 18616 12986 18644 13330
rect 18604 12980 18656 12986
rect 18604 12922 18656 12928
rect 18892 12850 18920 14010
rect 18880 12844 18932 12850
rect 18880 12786 18932 12792
rect 18510 12744 18566 12753
rect 18510 12679 18566 12688
rect 18524 12442 18552 12679
rect 18512 12436 18564 12442
rect 18512 12378 18564 12384
rect 18788 12368 18840 12374
rect 18788 12310 18840 12316
rect 18878 12336 18934 12345
rect 18432 12170 18552 12186
rect 18432 12164 18564 12170
rect 18432 12158 18512 12164
rect 18234 12135 18290 12144
rect 17744 11996 18052 12005
rect 17744 11994 17750 11996
rect 17806 11994 17830 11996
rect 17886 11994 17910 11996
rect 17966 11994 17990 11996
rect 18046 11994 18052 11996
rect 17806 11942 17808 11994
rect 17988 11942 17990 11994
rect 17744 11940 17750 11942
rect 17806 11940 17830 11942
rect 17886 11940 17910 11942
rect 17966 11940 17990 11942
rect 18046 11940 18052 11942
rect 17744 11931 18052 11940
rect 18248 11762 18276 12135
rect 18512 12106 18564 12112
rect 18236 11756 18288 11762
rect 18236 11698 18288 11704
rect 18524 11694 18552 12106
rect 18512 11688 18564 11694
rect 18800 11665 18828 12310
rect 18878 12271 18934 12280
rect 18892 12238 18920 12271
rect 18880 12232 18932 12238
rect 18880 12174 18932 12180
rect 18892 11898 18920 12174
rect 18880 11892 18932 11898
rect 18880 11834 18932 11840
rect 18512 11630 18564 11636
rect 18786 11656 18842 11665
rect 18786 11591 18842 11600
rect 18328 11552 18380 11558
rect 18328 11494 18380 11500
rect 18880 11552 18932 11558
rect 18880 11494 18932 11500
rect 17744 10908 18052 10917
rect 17744 10906 17750 10908
rect 17806 10906 17830 10908
rect 17886 10906 17910 10908
rect 17966 10906 17990 10908
rect 18046 10906 18052 10908
rect 17806 10854 17808 10906
rect 17988 10854 17990 10906
rect 17744 10852 17750 10854
rect 17806 10852 17830 10854
rect 17886 10852 17910 10854
rect 17966 10852 17990 10854
rect 18046 10852 18052 10854
rect 17744 10843 18052 10852
rect 18340 10792 18368 11494
rect 18512 11280 18564 11286
rect 18512 11222 18564 11228
rect 18340 10764 18460 10792
rect 18328 10668 18380 10674
rect 18328 10610 18380 10616
rect 18236 10124 18288 10130
rect 18236 10066 18288 10072
rect 17592 10056 17644 10062
rect 17592 9998 17644 10004
rect 18050 10024 18106 10033
rect 17500 9716 17552 9722
rect 17500 9658 17552 9664
rect 17408 9376 17460 9382
rect 17408 9318 17460 9324
rect 17604 9178 17632 9998
rect 18050 9959 18106 9968
rect 18144 9988 18196 9994
rect 18064 9926 18092 9959
rect 18144 9930 18196 9936
rect 18052 9920 18104 9926
rect 18052 9862 18104 9868
rect 17744 9820 18052 9829
rect 17744 9818 17750 9820
rect 17806 9818 17830 9820
rect 17886 9818 17910 9820
rect 17966 9818 17990 9820
rect 18046 9818 18052 9820
rect 17806 9766 17808 9818
rect 17988 9766 17990 9818
rect 17744 9764 17750 9766
rect 17806 9764 17830 9766
rect 17886 9764 17910 9766
rect 17966 9764 17990 9766
rect 18046 9764 18052 9766
rect 17744 9755 18052 9764
rect 18052 9716 18104 9722
rect 18052 9658 18104 9664
rect 17592 9172 17644 9178
rect 17592 9114 17644 9120
rect 17500 8900 17552 8906
rect 17500 8842 17552 8848
rect 17408 7812 17460 7818
rect 17408 7754 17460 7760
rect 17420 6186 17448 7754
rect 17512 6662 17540 8842
rect 17604 8294 17632 9114
rect 18064 8945 18092 9658
rect 18050 8936 18106 8945
rect 18050 8871 18106 8880
rect 17744 8732 18052 8741
rect 17744 8730 17750 8732
rect 17806 8730 17830 8732
rect 17886 8730 17910 8732
rect 17966 8730 17990 8732
rect 18046 8730 18052 8732
rect 17806 8678 17808 8730
rect 17988 8678 17990 8730
rect 17744 8676 17750 8678
rect 17806 8676 17830 8678
rect 17886 8676 17910 8678
rect 17966 8676 17990 8678
rect 18046 8676 18052 8678
rect 17744 8667 18052 8676
rect 18156 8566 18184 9930
rect 18248 9586 18276 10066
rect 18236 9580 18288 9586
rect 18236 9522 18288 9528
rect 18340 9178 18368 10610
rect 18432 10033 18460 10764
rect 18418 10024 18474 10033
rect 18418 9959 18474 9968
rect 18418 9888 18474 9897
rect 18418 9823 18474 9832
rect 18328 9172 18380 9178
rect 18328 9114 18380 9120
rect 18236 8968 18288 8974
rect 18236 8910 18288 8916
rect 18248 8634 18276 8910
rect 18236 8628 18288 8634
rect 18236 8570 18288 8576
rect 18144 8560 18196 8566
rect 18144 8502 18196 8508
rect 18328 8492 18380 8498
rect 18328 8434 18380 8440
rect 17592 8288 17644 8294
rect 17592 8230 17644 8236
rect 17744 7644 18052 7653
rect 17744 7642 17750 7644
rect 17806 7642 17830 7644
rect 17886 7642 17910 7644
rect 17966 7642 17990 7644
rect 18046 7642 18052 7644
rect 17806 7590 17808 7642
rect 17988 7590 17990 7642
rect 17744 7588 17750 7590
rect 17806 7588 17830 7590
rect 17886 7588 17910 7590
rect 17966 7588 17990 7590
rect 18046 7588 18052 7590
rect 17744 7579 18052 7588
rect 17960 7200 18012 7206
rect 17960 7142 18012 7148
rect 18144 7200 18196 7206
rect 18144 7142 18196 7148
rect 17972 6934 18000 7142
rect 17960 6928 18012 6934
rect 17960 6870 18012 6876
rect 17592 6724 17644 6730
rect 17592 6666 17644 6672
rect 17500 6656 17552 6662
rect 17500 6598 17552 6604
rect 17408 6180 17460 6186
rect 17408 6122 17460 6128
rect 17328 6038 17448 6066
rect 17316 5636 17368 5642
rect 17316 5578 17368 5584
rect 17132 5568 17184 5574
rect 17132 5510 17184 5516
rect 17224 5568 17276 5574
rect 17224 5510 17276 5516
rect 17144 5370 17172 5510
rect 17132 5364 17184 5370
rect 17132 5306 17184 5312
rect 17132 5092 17184 5098
rect 17132 5034 17184 5040
rect 17040 4684 17092 4690
rect 17040 4626 17092 4632
rect 17144 4486 17172 5034
rect 17328 4690 17356 5578
rect 17420 5166 17448 6038
rect 17512 5302 17540 6598
rect 17604 5914 17632 6666
rect 17744 6556 18052 6565
rect 17744 6554 17750 6556
rect 17806 6554 17830 6556
rect 17886 6554 17910 6556
rect 17966 6554 17990 6556
rect 18046 6554 18052 6556
rect 17806 6502 17808 6554
rect 17988 6502 17990 6554
rect 17744 6500 17750 6502
rect 17806 6500 17830 6502
rect 17886 6500 17910 6502
rect 17966 6500 17990 6502
rect 18046 6500 18052 6502
rect 17744 6491 18052 6500
rect 17776 6248 17828 6254
rect 17776 6190 17828 6196
rect 17684 6112 17736 6118
rect 17684 6054 17736 6060
rect 17592 5908 17644 5914
rect 17592 5850 17644 5856
rect 17696 5556 17724 6054
rect 17788 5914 17816 6190
rect 17960 6180 18012 6186
rect 17960 6122 18012 6128
rect 17776 5908 17828 5914
rect 17776 5850 17828 5856
rect 17972 5574 18000 6122
rect 17604 5528 17724 5556
rect 17960 5568 18012 5574
rect 17604 5370 17632 5528
rect 17960 5510 18012 5516
rect 17744 5468 18052 5477
rect 17744 5466 17750 5468
rect 17806 5466 17830 5468
rect 17886 5466 17910 5468
rect 17966 5466 17990 5468
rect 18046 5466 18052 5468
rect 17806 5414 17808 5466
rect 17988 5414 17990 5466
rect 17744 5412 17750 5414
rect 17806 5412 17830 5414
rect 17886 5412 17910 5414
rect 17966 5412 17990 5414
rect 18046 5412 18052 5414
rect 17744 5403 18052 5412
rect 17592 5364 17644 5370
rect 17592 5306 17644 5312
rect 17500 5296 17552 5302
rect 17500 5238 17552 5244
rect 17408 5160 17460 5166
rect 17408 5102 17460 5108
rect 17500 5024 17552 5030
rect 17500 4966 17552 4972
rect 17316 4684 17368 4690
rect 17316 4626 17368 4632
rect 17132 4480 17184 4486
rect 17132 4422 17184 4428
rect 16948 4140 17000 4146
rect 16948 4082 17000 4088
rect 16960 3618 16988 4082
rect 16960 3602 17080 3618
rect 16856 3596 16908 3602
rect 16960 3596 17092 3602
rect 16960 3590 17040 3596
rect 16856 3538 16908 3544
rect 17040 3538 17092 3544
rect 17144 3584 17172 4422
rect 17328 3738 17356 4626
rect 17408 4616 17460 4622
rect 17408 4558 17460 4564
rect 17316 3732 17368 3738
rect 17316 3674 17368 3680
rect 17224 3596 17276 3602
rect 17144 3556 17224 3584
rect 17144 3398 17172 3556
rect 17224 3538 17276 3544
rect 17328 3534 17356 3674
rect 17316 3528 17368 3534
rect 17316 3470 17368 3476
rect 17132 3392 17184 3398
rect 17132 3334 17184 3340
rect 17224 3392 17276 3398
rect 17224 3334 17276 3340
rect 16670 3088 16726 3097
rect 17144 3074 17172 3334
rect 16670 3023 16726 3032
rect 16764 3052 16816 3058
rect 16764 2994 16816 3000
rect 17052 3046 17172 3074
rect 16580 2984 16632 2990
rect 16580 2926 16632 2932
rect 16776 2650 16804 2994
rect 17052 2990 17080 3046
rect 17236 2990 17264 3334
rect 17420 2990 17448 4558
rect 17512 4146 17540 4966
rect 18156 4690 18184 7142
rect 18236 6928 18288 6934
rect 18236 6870 18288 6876
rect 18248 5778 18276 6870
rect 18236 5772 18288 5778
rect 18236 5714 18288 5720
rect 18340 5642 18368 8434
rect 18432 7886 18460 9823
rect 18524 9586 18552 11222
rect 18696 11144 18748 11150
rect 18696 11086 18748 11092
rect 18708 10112 18736 11086
rect 18892 11014 18920 11494
rect 18880 11008 18932 11014
rect 18880 10950 18932 10956
rect 18892 10606 18920 10950
rect 18788 10600 18840 10606
rect 18788 10542 18840 10548
rect 18880 10600 18932 10606
rect 18880 10542 18932 10548
rect 18699 10084 18736 10112
rect 18800 10112 18828 10542
rect 18892 10266 18920 10542
rect 18880 10260 18932 10266
rect 18880 10202 18932 10208
rect 18984 10130 19012 18294
rect 19064 17808 19116 17814
rect 19062 17776 19064 17785
rect 19116 17776 19118 17785
rect 19062 17711 19118 17720
rect 19168 16017 19196 19654
rect 19260 19310 19288 19790
rect 19432 19712 19484 19718
rect 19432 19654 19484 19660
rect 19340 19508 19392 19514
rect 19340 19450 19392 19456
rect 19248 19304 19300 19310
rect 19248 19246 19300 19252
rect 19248 18760 19300 18766
rect 19248 18702 19300 18708
rect 19260 18290 19288 18702
rect 19248 18284 19300 18290
rect 19248 18226 19300 18232
rect 19260 17746 19288 18226
rect 19248 17740 19300 17746
rect 19248 17682 19300 17688
rect 19352 17610 19380 19450
rect 19444 18902 19472 19654
rect 19432 18896 19484 18902
rect 19432 18838 19484 18844
rect 19536 18442 19564 21422
rect 19708 21412 19760 21418
rect 19708 21354 19760 21360
rect 19800 21412 19852 21418
rect 19800 21354 19852 21360
rect 19720 20874 19748 21354
rect 19708 20868 19760 20874
rect 19708 20810 19760 20816
rect 19812 18698 19840 21354
rect 19904 20602 19932 21490
rect 20168 21480 20220 21486
rect 20168 21422 20220 21428
rect 19892 20596 19944 20602
rect 19892 20538 19944 20544
rect 19984 20460 20036 20466
rect 19984 20402 20036 20408
rect 19996 19417 20024 20402
rect 20180 19786 20208 21422
rect 20260 20936 20312 20942
rect 20260 20878 20312 20884
rect 20168 19780 20220 19786
rect 20168 19722 20220 19728
rect 19982 19408 20038 19417
rect 19982 19343 20038 19352
rect 20076 19372 20128 19378
rect 19800 18692 19852 18698
rect 19800 18634 19852 18640
rect 19708 18624 19760 18630
rect 19708 18566 19760 18572
rect 19444 18426 19564 18442
rect 19432 18420 19564 18426
rect 19484 18414 19564 18420
rect 19616 18420 19668 18426
rect 19432 18362 19484 18368
rect 19616 18362 19668 18368
rect 19340 17604 19392 17610
rect 19340 17546 19392 17552
rect 19340 16992 19392 16998
rect 19340 16934 19392 16940
rect 19352 16794 19380 16934
rect 19340 16788 19392 16794
rect 19340 16730 19392 16736
rect 19154 16008 19210 16017
rect 19154 15943 19210 15952
rect 19154 15600 19210 15609
rect 19154 15535 19210 15544
rect 19168 15502 19196 15535
rect 19352 15502 19380 16730
rect 19432 16652 19484 16658
rect 19432 16594 19484 16600
rect 19444 16153 19472 16594
rect 19430 16144 19486 16153
rect 19628 16114 19656 18362
rect 19720 18290 19748 18566
rect 19708 18284 19760 18290
rect 19708 18226 19760 18232
rect 19706 18184 19762 18193
rect 19706 18119 19762 18128
rect 19430 16079 19486 16088
rect 19616 16108 19668 16114
rect 19616 16050 19668 16056
rect 19156 15496 19208 15502
rect 19156 15438 19208 15444
rect 19340 15496 19392 15502
rect 19340 15438 19392 15444
rect 19432 14612 19484 14618
rect 19432 14554 19484 14560
rect 19248 14476 19300 14482
rect 19248 14418 19300 14424
rect 19156 14408 19208 14414
rect 19156 14350 19208 14356
rect 19168 13530 19196 14350
rect 19260 14074 19288 14418
rect 19444 14346 19472 14554
rect 19432 14340 19484 14346
rect 19432 14282 19484 14288
rect 19616 14340 19668 14346
rect 19616 14282 19668 14288
rect 19248 14068 19300 14074
rect 19248 14010 19300 14016
rect 19260 13938 19288 14010
rect 19340 14000 19392 14006
rect 19340 13942 19392 13948
rect 19248 13932 19300 13938
rect 19248 13874 19300 13880
rect 19156 13524 19208 13530
rect 19156 13466 19208 13472
rect 19260 13394 19288 13874
rect 19248 13388 19300 13394
rect 19248 13330 19300 13336
rect 19064 13184 19116 13190
rect 19064 13126 19116 13132
rect 19248 13184 19300 13190
rect 19352 13161 19380 13942
rect 19628 13870 19656 14282
rect 19616 13864 19668 13870
rect 19616 13806 19668 13812
rect 19616 13252 19668 13258
rect 19616 13194 19668 13200
rect 19248 13126 19300 13132
rect 19338 13152 19394 13161
rect 19076 12889 19104 13126
rect 19156 12912 19208 12918
rect 19062 12880 19118 12889
rect 19156 12854 19208 12860
rect 19062 12815 19118 12824
rect 19064 12368 19116 12374
rect 19064 12310 19116 12316
rect 18972 10124 19024 10130
rect 18800 10084 18920 10112
rect 18699 9926 18727 10084
rect 18892 9976 18920 10084
rect 18972 10066 19024 10072
rect 18800 9948 18920 9976
rect 18970 10024 19026 10033
rect 18970 9959 19026 9968
rect 18604 9920 18656 9926
rect 18604 9862 18656 9868
rect 18696 9920 18748 9926
rect 18696 9862 18748 9868
rect 18512 9580 18564 9586
rect 18512 9522 18564 9528
rect 18524 8786 18552 9522
rect 18616 8974 18644 9862
rect 18708 9722 18736 9862
rect 18800 9761 18828 9948
rect 18878 9888 18934 9897
rect 18878 9823 18934 9832
rect 18786 9752 18842 9761
rect 18696 9716 18748 9722
rect 18786 9687 18842 9696
rect 18696 9658 18748 9664
rect 18892 9602 18920 9823
rect 18708 9574 18920 9602
rect 18984 9586 19012 9959
rect 18972 9580 19024 9586
rect 18604 8968 18656 8974
rect 18604 8910 18656 8916
rect 18524 8758 18644 8786
rect 18420 7880 18472 7886
rect 18420 7822 18472 7828
rect 18420 6656 18472 6662
rect 18420 6598 18472 6604
rect 18432 5710 18460 6598
rect 18512 6316 18564 6322
rect 18512 6258 18564 6264
rect 18524 5778 18552 6258
rect 18512 5772 18564 5778
rect 18512 5714 18564 5720
rect 18420 5704 18472 5710
rect 18420 5646 18472 5652
rect 18328 5636 18380 5642
rect 18328 5578 18380 5584
rect 18236 5568 18288 5574
rect 18236 5510 18288 5516
rect 18248 5234 18276 5510
rect 18236 5228 18288 5234
rect 18236 5170 18288 5176
rect 18144 4684 18196 4690
rect 18144 4626 18196 4632
rect 18248 4622 18276 5170
rect 18616 5166 18644 8758
rect 18708 7478 18736 9574
rect 18972 9522 19024 9528
rect 18788 9512 18840 9518
rect 18788 9454 18840 9460
rect 18800 9042 18828 9454
rect 18984 9110 19012 9522
rect 19076 9489 19104 12310
rect 19168 12306 19196 12854
rect 19260 12646 19288 13126
rect 19338 13087 19394 13096
rect 19248 12640 19300 12646
rect 19248 12582 19300 12588
rect 19156 12300 19208 12306
rect 19156 12242 19208 12248
rect 19628 12170 19656 13194
rect 19720 12434 19748 18119
rect 19800 17604 19852 17610
rect 19800 17546 19852 17552
rect 19812 15162 19840 17546
rect 19892 16448 19944 16454
rect 19892 16390 19944 16396
rect 19904 16114 19932 16390
rect 19892 16108 19944 16114
rect 19892 16050 19944 16056
rect 19904 15502 19932 16050
rect 19892 15496 19944 15502
rect 19892 15438 19944 15444
rect 19996 15434 20024 19343
rect 20076 19314 20128 19320
rect 20088 18873 20116 19314
rect 20074 18864 20130 18873
rect 20074 18799 20130 18808
rect 20272 18358 20300 20878
rect 20260 18352 20312 18358
rect 20260 18294 20312 18300
rect 20364 17882 20392 21490
rect 20640 21350 20668 21626
rect 20824 21400 20852 21830
rect 21100 21706 21128 21966
rect 21272 21888 21324 21894
rect 21272 21830 21324 21836
rect 21008 21678 21128 21706
rect 21008 21457 21036 21678
rect 21088 21548 21140 21554
rect 21088 21490 21140 21496
rect 20994 21448 21050 21457
rect 20824 21372 20944 21400
rect 20994 21383 21050 21392
rect 20628 21344 20680 21350
rect 20628 21286 20680 21292
rect 20543 21244 20851 21253
rect 20543 21242 20549 21244
rect 20605 21242 20629 21244
rect 20685 21242 20709 21244
rect 20765 21242 20789 21244
rect 20845 21242 20851 21244
rect 20605 21190 20607 21242
rect 20787 21190 20789 21242
rect 20543 21188 20549 21190
rect 20605 21188 20629 21190
rect 20685 21188 20709 21190
rect 20765 21188 20789 21190
rect 20845 21188 20851 21190
rect 20543 21179 20851 21188
rect 20444 21140 20496 21146
rect 20444 21082 20496 21088
rect 20456 20058 20484 21082
rect 20810 21040 20866 21049
rect 20810 20975 20866 20984
rect 20824 20806 20852 20975
rect 20720 20800 20772 20806
rect 20720 20742 20772 20748
rect 20812 20800 20864 20806
rect 20812 20742 20864 20748
rect 20732 20602 20760 20742
rect 20916 20602 20944 21372
rect 21100 21010 21128 21490
rect 21180 21480 21232 21486
rect 21180 21422 21232 21428
rect 21088 21004 21140 21010
rect 21088 20946 21140 20952
rect 20996 20936 21048 20942
rect 20996 20878 21048 20884
rect 20720 20596 20772 20602
rect 20720 20538 20772 20544
rect 20904 20596 20956 20602
rect 20904 20538 20956 20544
rect 20543 20156 20851 20165
rect 20543 20154 20549 20156
rect 20605 20154 20629 20156
rect 20685 20154 20709 20156
rect 20765 20154 20789 20156
rect 20845 20154 20851 20156
rect 20605 20102 20607 20154
rect 20787 20102 20789 20154
rect 20543 20100 20549 20102
rect 20605 20100 20629 20102
rect 20685 20100 20709 20102
rect 20765 20100 20789 20102
rect 20845 20100 20851 20102
rect 20543 20091 20851 20100
rect 20444 20052 20496 20058
rect 20444 19994 20496 20000
rect 20536 20052 20588 20058
rect 20536 19994 20588 20000
rect 20548 19854 20576 19994
rect 20536 19848 20588 19854
rect 20904 19848 20956 19854
rect 20536 19790 20588 19796
rect 20902 19816 20904 19825
rect 21008 19836 21036 20878
rect 21088 20256 21140 20262
rect 21088 20198 21140 20204
rect 20956 19816 21036 19836
rect 20958 19808 21036 19816
rect 20548 19378 20576 19790
rect 20902 19751 20958 19760
rect 20720 19712 20772 19718
rect 20720 19654 20772 19660
rect 20732 19446 20760 19654
rect 21100 19446 21128 20198
rect 21192 19530 21220 21422
rect 21284 19922 21312 21830
rect 21376 21690 21404 21984
rect 21456 21966 21508 21972
rect 21560 21876 21588 23800
rect 21824 22024 21876 22030
rect 21822 21992 21824 22001
rect 21876 21992 21878 22001
rect 21822 21927 21878 21936
rect 22204 21894 22232 23800
rect 22560 22228 22612 22234
rect 22560 22170 22612 22176
rect 22468 22024 22520 22030
rect 22468 21966 22520 21972
rect 21640 21888 21692 21894
rect 21560 21848 21640 21876
rect 21640 21830 21692 21836
rect 22192 21888 22244 21894
rect 22192 21830 22244 21836
rect 21364 21684 21416 21690
rect 21364 21626 21416 21632
rect 21824 21616 21876 21622
rect 22480 21593 22508 21966
rect 21824 21558 21876 21564
rect 22466 21584 22522 21593
rect 21732 21480 21784 21486
rect 21732 21422 21784 21428
rect 21364 21344 21416 21350
rect 21364 21286 21416 21292
rect 21376 20913 21404 21286
rect 21362 20904 21418 20913
rect 21362 20839 21418 20848
rect 21376 20466 21404 20839
rect 21548 20800 21600 20806
rect 21548 20742 21600 20748
rect 21640 20800 21692 20806
rect 21640 20742 21692 20748
rect 21364 20460 21416 20466
rect 21364 20402 21416 20408
rect 21456 20324 21508 20330
rect 21456 20266 21508 20272
rect 21468 19922 21496 20266
rect 21272 19916 21324 19922
rect 21272 19858 21324 19864
rect 21456 19916 21508 19922
rect 21456 19858 21508 19864
rect 21560 19718 21588 20742
rect 21548 19712 21600 19718
rect 21548 19654 21600 19660
rect 21652 19530 21680 20742
rect 21744 19854 21772 21422
rect 21836 20262 21864 21558
rect 22192 21548 22244 21554
rect 22466 21519 22522 21528
rect 22192 21490 22244 21496
rect 22100 21344 22152 21350
rect 22100 21286 22152 21292
rect 22112 20618 22140 21286
rect 22204 20777 22232 21490
rect 22572 20942 22600 22170
rect 22848 21894 22876 23800
rect 23204 21956 23256 21962
rect 23204 21898 23256 21904
rect 22836 21888 22888 21894
rect 22836 21830 22888 21836
rect 22650 21584 22706 21593
rect 22650 21519 22706 21528
rect 22664 21146 22692 21519
rect 23020 21344 23072 21350
rect 23020 21286 23072 21292
rect 22652 21140 22704 21146
rect 22652 21082 22704 21088
rect 23032 21049 23060 21286
rect 23216 21078 23244 21898
rect 23204 21072 23256 21078
rect 23018 21040 23074 21049
rect 23204 21014 23256 21020
rect 23018 20975 23074 20984
rect 22284 20936 22336 20942
rect 22284 20878 22336 20884
rect 22560 20936 22612 20942
rect 22560 20878 22612 20884
rect 22190 20768 22246 20777
rect 22190 20703 22246 20712
rect 22020 20602 22140 20618
rect 22008 20596 22140 20602
rect 22060 20590 22140 20596
rect 22008 20538 22060 20544
rect 21824 20256 21876 20262
rect 21824 20198 21876 20204
rect 22112 20074 22140 20590
rect 22296 20398 22324 20878
rect 23112 20868 23164 20874
rect 23112 20810 23164 20816
rect 23020 20800 23072 20806
rect 23020 20742 23072 20748
rect 23032 20505 23060 20742
rect 23018 20496 23074 20505
rect 22836 20460 22888 20466
rect 23018 20431 23074 20440
rect 22836 20402 22888 20408
rect 22284 20392 22336 20398
rect 22284 20334 22336 20340
rect 22560 20392 22612 20398
rect 22560 20334 22612 20340
rect 22020 20058 22140 20074
rect 22296 20058 22324 20334
rect 22008 20052 22140 20058
rect 22060 20046 22140 20052
rect 22284 20052 22336 20058
rect 22008 19994 22060 20000
rect 22284 19994 22336 20000
rect 21732 19848 21784 19854
rect 21732 19790 21784 19796
rect 21192 19502 21680 19530
rect 20720 19440 20772 19446
rect 20720 19382 20772 19388
rect 21088 19440 21140 19446
rect 21088 19382 21140 19388
rect 20536 19372 20588 19378
rect 20456 19332 20536 19360
rect 20456 18952 20484 19332
rect 20536 19314 20588 19320
rect 20904 19372 20956 19378
rect 20904 19314 20956 19320
rect 20543 19068 20851 19077
rect 20543 19066 20549 19068
rect 20605 19066 20629 19068
rect 20685 19066 20709 19068
rect 20765 19066 20789 19068
rect 20845 19066 20851 19068
rect 20605 19014 20607 19066
rect 20787 19014 20789 19066
rect 20543 19012 20549 19014
rect 20605 19012 20629 19014
rect 20685 19012 20709 19014
rect 20765 19012 20789 19014
rect 20845 19012 20851 19014
rect 20543 19003 20851 19012
rect 20456 18924 20760 18952
rect 20732 18766 20760 18924
rect 20812 18896 20864 18902
rect 20810 18864 20812 18873
rect 20864 18864 20866 18873
rect 20810 18799 20866 18808
rect 20720 18760 20772 18766
rect 20720 18702 20772 18708
rect 20444 18692 20496 18698
rect 20444 18634 20496 18640
rect 20456 17882 20484 18634
rect 20628 18420 20680 18426
rect 20628 18362 20680 18368
rect 20640 18170 20668 18362
rect 20640 18154 20760 18170
rect 20640 18148 20772 18154
rect 20640 18142 20720 18148
rect 20720 18090 20772 18096
rect 20543 17980 20851 17989
rect 20543 17978 20549 17980
rect 20605 17978 20629 17980
rect 20685 17978 20709 17980
rect 20765 17978 20789 17980
rect 20845 17978 20851 17980
rect 20605 17926 20607 17978
rect 20787 17926 20789 17978
rect 20543 17924 20549 17926
rect 20605 17924 20629 17926
rect 20685 17924 20709 17926
rect 20765 17924 20789 17926
rect 20845 17924 20851 17926
rect 20543 17915 20851 17924
rect 20352 17876 20404 17882
rect 20352 17818 20404 17824
rect 20444 17876 20496 17882
rect 20444 17818 20496 17824
rect 20720 17536 20772 17542
rect 20916 17513 20944 19314
rect 21180 19168 21232 19174
rect 21180 19110 21232 19116
rect 21192 18290 21220 19110
rect 21272 18352 21324 18358
rect 21272 18294 21324 18300
rect 21180 18284 21232 18290
rect 21180 18226 21232 18232
rect 20996 18080 21048 18086
rect 20996 18022 21048 18028
rect 21008 17678 21036 18022
rect 21088 17876 21140 17882
rect 21088 17818 21140 17824
rect 21100 17678 21128 17818
rect 21284 17678 21312 18294
rect 20996 17672 21048 17678
rect 20996 17614 21048 17620
rect 21088 17672 21140 17678
rect 21088 17614 21140 17620
rect 21272 17672 21324 17678
rect 21272 17614 21324 17620
rect 20720 17478 20772 17484
rect 20902 17504 20958 17513
rect 20732 17202 20760 17478
rect 20902 17439 20958 17448
rect 21008 17270 21036 17614
rect 20996 17264 21048 17270
rect 20996 17206 21048 17212
rect 20720 17196 20772 17202
rect 20720 17138 20772 17144
rect 21272 17196 21324 17202
rect 21272 17138 21324 17144
rect 20904 17128 20956 17134
rect 20904 17070 20956 17076
rect 21088 17128 21140 17134
rect 21088 17070 21140 17076
rect 20543 16892 20851 16901
rect 20543 16890 20549 16892
rect 20605 16890 20629 16892
rect 20685 16890 20709 16892
rect 20765 16890 20789 16892
rect 20845 16890 20851 16892
rect 20605 16838 20607 16890
rect 20787 16838 20789 16890
rect 20543 16836 20549 16838
rect 20605 16836 20629 16838
rect 20685 16836 20709 16838
rect 20765 16836 20789 16838
rect 20845 16836 20851 16838
rect 20543 16827 20851 16836
rect 20916 16726 20944 17070
rect 20904 16720 20956 16726
rect 20904 16662 20956 16668
rect 21100 16658 21128 17070
rect 21284 16794 21312 17138
rect 21272 16788 21324 16794
rect 21272 16730 21324 16736
rect 21088 16652 21140 16658
rect 21088 16594 21140 16600
rect 20904 16584 20956 16590
rect 20904 16526 20956 16532
rect 20352 16516 20404 16522
rect 20352 16458 20404 16464
rect 20536 16516 20588 16522
rect 20536 16458 20588 16464
rect 20168 16176 20220 16182
rect 20168 16118 20220 16124
rect 20180 15706 20208 16118
rect 20364 15706 20392 16458
rect 20548 16250 20576 16458
rect 20536 16244 20588 16250
rect 20536 16186 20588 16192
rect 20916 16114 20944 16526
rect 20904 16108 20956 16114
rect 20904 16050 20956 16056
rect 20543 15804 20851 15813
rect 20543 15802 20549 15804
rect 20605 15802 20629 15804
rect 20685 15802 20709 15804
rect 20765 15802 20789 15804
rect 20845 15802 20851 15804
rect 20605 15750 20607 15802
rect 20787 15750 20789 15802
rect 20543 15748 20549 15750
rect 20605 15748 20629 15750
rect 20685 15748 20709 15750
rect 20765 15748 20789 15750
rect 20845 15748 20851 15750
rect 20543 15739 20851 15748
rect 20168 15700 20220 15706
rect 20168 15642 20220 15648
rect 20352 15700 20404 15706
rect 20352 15642 20404 15648
rect 20812 15564 20864 15570
rect 20916 15552 20944 16050
rect 21272 15972 21324 15978
rect 21272 15914 21324 15920
rect 21088 15904 21140 15910
rect 21088 15846 21140 15852
rect 21100 15638 21128 15846
rect 21088 15632 21140 15638
rect 21088 15574 21140 15580
rect 20864 15524 20944 15552
rect 20812 15506 20864 15512
rect 19984 15428 20036 15434
rect 19984 15370 20036 15376
rect 19800 15156 19852 15162
rect 19800 15098 19852 15104
rect 20824 14958 20852 15506
rect 21284 15162 21312 15914
rect 21272 15156 21324 15162
rect 21272 15098 21324 15104
rect 21088 15020 21140 15026
rect 21088 14962 21140 14968
rect 20812 14952 20864 14958
rect 20812 14894 20864 14900
rect 20996 14952 21048 14958
rect 21100 14929 21128 14962
rect 20996 14894 21048 14900
rect 21086 14920 21142 14929
rect 20543 14716 20851 14725
rect 20543 14714 20549 14716
rect 20605 14714 20629 14716
rect 20685 14714 20709 14716
rect 20765 14714 20789 14716
rect 20845 14714 20851 14716
rect 20605 14662 20607 14714
rect 20787 14662 20789 14714
rect 20543 14660 20549 14662
rect 20605 14660 20629 14662
rect 20685 14660 20709 14662
rect 20765 14660 20789 14662
rect 20845 14660 20851 14662
rect 20543 14651 20851 14660
rect 20812 14476 20864 14482
rect 20812 14418 20864 14424
rect 20720 14408 20772 14414
rect 20720 14350 20772 14356
rect 20260 14272 20312 14278
rect 20260 14214 20312 14220
rect 20536 14272 20588 14278
rect 20536 14214 20588 14220
rect 20272 12918 20300 14214
rect 20548 13938 20576 14214
rect 20732 14006 20760 14350
rect 20720 14000 20772 14006
rect 20720 13942 20772 13948
rect 20536 13932 20588 13938
rect 20536 13874 20588 13880
rect 20824 13870 20852 14418
rect 21008 14385 21036 14894
rect 21086 14855 21142 14864
rect 20994 14376 21050 14385
rect 20994 14311 21050 14320
rect 20812 13864 20864 13870
rect 20812 13806 20864 13812
rect 20996 13864 21048 13870
rect 20996 13806 21048 13812
rect 20543 13628 20851 13637
rect 20543 13626 20549 13628
rect 20605 13626 20629 13628
rect 20685 13626 20709 13628
rect 20765 13626 20789 13628
rect 20845 13626 20851 13628
rect 20605 13574 20607 13626
rect 20787 13574 20789 13626
rect 20543 13572 20549 13574
rect 20605 13572 20629 13574
rect 20685 13572 20709 13574
rect 20765 13572 20789 13574
rect 20845 13572 20851 13574
rect 20543 13563 20851 13572
rect 20904 13524 20956 13530
rect 20904 13466 20956 13472
rect 20718 13288 20774 13297
rect 20718 13223 20774 13232
rect 20732 13190 20760 13223
rect 20720 13184 20772 13190
rect 20720 13126 20772 13132
rect 20260 12912 20312 12918
rect 20260 12854 20312 12860
rect 20444 12844 20496 12850
rect 20444 12786 20496 12792
rect 19720 12406 19840 12434
rect 19340 12164 19392 12170
rect 19340 12106 19392 12112
rect 19616 12164 19668 12170
rect 19616 12106 19668 12112
rect 19352 11801 19380 12106
rect 19708 12096 19760 12102
rect 19708 12038 19760 12044
rect 19338 11792 19394 11801
rect 19720 11762 19748 12038
rect 19338 11727 19394 11736
rect 19616 11756 19668 11762
rect 19616 11698 19668 11704
rect 19708 11756 19760 11762
rect 19708 11698 19760 11704
rect 19432 11348 19484 11354
rect 19432 11290 19484 11296
rect 19340 11144 19392 11150
rect 19340 11086 19392 11092
rect 19352 10713 19380 11086
rect 19338 10704 19394 10713
rect 19338 10639 19394 10648
rect 19248 10464 19300 10470
rect 19248 10406 19300 10412
rect 19156 10056 19208 10062
rect 19156 9998 19208 10004
rect 19168 9625 19196 9998
rect 19260 9897 19288 10406
rect 19338 10024 19394 10033
rect 19338 9959 19394 9968
rect 19246 9888 19302 9897
rect 19246 9823 19302 9832
rect 19352 9704 19380 9959
rect 19260 9676 19380 9704
rect 19154 9616 19210 9625
rect 19154 9551 19210 9560
rect 19062 9480 19118 9489
rect 19062 9415 19118 9424
rect 19260 9178 19288 9676
rect 19444 9586 19472 11290
rect 19628 11257 19656 11698
rect 19614 11248 19670 11257
rect 19614 11183 19670 11192
rect 19616 10192 19668 10198
rect 19616 10134 19668 10140
rect 19432 9580 19484 9586
rect 19432 9522 19484 9528
rect 19248 9172 19300 9178
rect 19248 9114 19300 9120
rect 18880 9104 18932 9110
rect 18880 9046 18932 9052
rect 18972 9104 19024 9110
rect 19628 9081 19656 10134
rect 18972 9046 19024 9052
rect 19614 9072 19670 9081
rect 18788 9036 18840 9042
rect 18788 8978 18840 8984
rect 18788 8832 18840 8838
rect 18788 8774 18840 8780
rect 18696 7472 18748 7478
rect 18696 7414 18748 7420
rect 18696 6656 18748 6662
rect 18696 6598 18748 6604
rect 18708 5302 18736 6598
rect 18800 6186 18828 8774
rect 18892 8106 18920 9046
rect 19156 9036 19208 9042
rect 19614 9007 19670 9016
rect 19156 8978 19208 8984
rect 19064 8492 19116 8498
rect 19064 8434 19116 8440
rect 18892 8078 19012 8106
rect 18880 6724 18932 6730
rect 18880 6666 18932 6672
rect 18788 6180 18840 6186
rect 18788 6122 18840 6128
rect 18696 5296 18748 5302
rect 18696 5238 18748 5244
rect 18788 5228 18840 5234
rect 18788 5170 18840 5176
rect 18604 5160 18656 5166
rect 18604 5102 18656 5108
rect 18800 4758 18828 5170
rect 18788 4752 18840 4758
rect 18788 4694 18840 4700
rect 18236 4616 18288 4622
rect 18236 4558 18288 4564
rect 18788 4480 18840 4486
rect 18788 4422 18840 4428
rect 17744 4380 18052 4389
rect 17744 4378 17750 4380
rect 17806 4378 17830 4380
rect 17886 4378 17910 4380
rect 17966 4378 17990 4380
rect 18046 4378 18052 4380
rect 17806 4326 17808 4378
rect 17988 4326 17990 4378
rect 17744 4324 17750 4326
rect 17806 4324 17830 4326
rect 17886 4324 17910 4326
rect 17966 4324 17990 4326
rect 18046 4324 18052 4326
rect 17744 4315 18052 4324
rect 17500 4140 17552 4146
rect 17500 4082 17552 4088
rect 17684 4140 17736 4146
rect 17684 4082 17736 4088
rect 18420 4140 18472 4146
rect 18420 4082 18472 4088
rect 17696 4026 17724 4082
rect 17960 4072 18012 4078
rect 17696 4020 17960 4026
rect 17696 4014 18012 4020
rect 18144 4072 18196 4078
rect 18144 4014 18196 4020
rect 17696 3998 18000 4014
rect 18156 3670 18184 4014
rect 18144 3664 18196 3670
rect 18144 3606 18196 3612
rect 18328 3596 18380 3602
rect 18328 3538 18380 3544
rect 17744 3292 18052 3301
rect 17744 3290 17750 3292
rect 17806 3290 17830 3292
rect 17886 3290 17910 3292
rect 17966 3290 17990 3292
rect 18046 3290 18052 3292
rect 17806 3238 17808 3290
rect 17988 3238 17990 3290
rect 17744 3236 17750 3238
rect 17806 3236 17830 3238
rect 17886 3236 17910 3238
rect 17966 3236 17990 3238
rect 18046 3236 18052 3238
rect 17744 3227 18052 3236
rect 17040 2984 17092 2990
rect 17040 2926 17092 2932
rect 17224 2984 17276 2990
rect 17224 2926 17276 2932
rect 17408 2984 17460 2990
rect 17408 2926 17460 2932
rect 18340 2854 18368 3538
rect 18432 2854 18460 4082
rect 18512 4072 18564 4078
rect 18564 4020 18736 4026
rect 18512 4014 18736 4020
rect 18524 3998 18736 4014
rect 18708 3534 18736 3998
rect 18696 3528 18748 3534
rect 18696 3470 18748 3476
rect 18708 2854 18736 3470
rect 18800 2990 18828 4422
rect 18892 4146 18920 6666
rect 18984 6254 19012 8078
rect 19076 6662 19104 8434
rect 19168 8430 19196 8978
rect 19340 8968 19392 8974
rect 19340 8910 19392 8916
rect 19616 8968 19668 8974
rect 19616 8910 19668 8916
rect 19352 8537 19380 8910
rect 19524 8560 19576 8566
rect 19338 8528 19394 8537
rect 19260 8486 19338 8514
rect 19156 8424 19208 8430
rect 19156 8366 19208 8372
rect 19260 6866 19288 8486
rect 19338 8463 19394 8472
rect 19444 8520 19524 8548
rect 19444 7206 19472 8520
rect 19524 8502 19576 8508
rect 19628 8294 19656 8910
rect 19616 8288 19668 8294
rect 19616 8230 19668 8236
rect 19524 7744 19576 7750
rect 19524 7686 19576 7692
rect 19536 7546 19564 7686
rect 19524 7540 19576 7546
rect 19524 7482 19576 7488
rect 19432 7200 19484 7206
rect 19536 7177 19564 7482
rect 19628 7342 19656 8230
rect 19812 7528 19840 12406
rect 20456 11898 20484 12786
rect 20543 12540 20851 12549
rect 20543 12538 20549 12540
rect 20605 12538 20629 12540
rect 20685 12538 20709 12540
rect 20765 12538 20789 12540
rect 20845 12538 20851 12540
rect 20605 12486 20607 12538
rect 20787 12486 20789 12538
rect 20543 12484 20549 12486
rect 20605 12484 20629 12486
rect 20685 12484 20709 12486
rect 20765 12484 20789 12486
rect 20845 12484 20851 12486
rect 20543 12475 20851 12484
rect 20720 12436 20772 12442
rect 20720 12378 20772 12384
rect 20812 12436 20864 12442
rect 20812 12378 20864 12384
rect 20732 12102 20760 12378
rect 20824 12306 20852 12378
rect 20812 12300 20864 12306
rect 20812 12242 20864 12248
rect 20628 12096 20680 12102
rect 20628 12038 20680 12044
rect 20720 12096 20772 12102
rect 20720 12038 20772 12044
rect 20444 11892 20496 11898
rect 20444 11834 20496 11840
rect 20640 11830 20668 12038
rect 20628 11824 20680 11830
rect 20628 11766 20680 11772
rect 20824 11694 20852 12242
rect 20916 12238 20944 13466
rect 21008 13326 21036 13806
rect 21088 13796 21140 13802
rect 21088 13738 21140 13744
rect 21100 13394 21128 13738
rect 21376 13734 21404 19502
rect 22100 19372 22152 19378
rect 22100 19314 22152 19320
rect 22376 19372 22428 19378
rect 22376 19314 22428 19320
rect 21732 19304 21784 19310
rect 21732 19246 21784 19252
rect 21916 19304 21968 19310
rect 21916 19246 21968 19252
rect 21456 18284 21508 18290
rect 21456 18226 21508 18232
rect 21468 16454 21496 18226
rect 21744 17882 21772 19246
rect 21928 18698 21956 19246
rect 22008 19236 22060 19242
rect 22008 19178 22060 19184
rect 22020 18970 22048 19178
rect 22112 18970 22140 19314
rect 22284 19168 22336 19174
rect 22284 19110 22336 19116
rect 22008 18964 22060 18970
rect 22008 18906 22060 18912
rect 22100 18964 22152 18970
rect 22100 18906 22152 18912
rect 22296 18748 22324 19110
rect 22388 18873 22416 19314
rect 22468 19304 22520 19310
rect 22468 19246 22520 19252
rect 22374 18864 22430 18873
rect 22480 18834 22508 19246
rect 22374 18799 22430 18808
rect 22468 18828 22520 18834
rect 22468 18770 22520 18776
rect 22376 18760 22428 18766
rect 22296 18720 22376 18748
rect 22376 18702 22428 18708
rect 21916 18692 21968 18698
rect 21916 18634 21968 18640
rect 21732 17876 21784 17882
rect 21732 17818 21784 17824
rect 21548 17740 21600 17746
rect 21548 17682 21600 17688
rect 21456 16448 21508 16454
rect 21456 16390 21508 16396
rect 21560 16182 21588 17682
rect 21640 16992 21692 16998
rect 21640 16934 21692 16940
rect 21652 16658 21680 16934
rect 21640 16652 21692 16658
rect 21640 16594 21692 16600
rect 21744 16590 21772 17818
rect 21824 16720 21876 16726
rect 21824 16662 21876 16668
rect 21732 16584 21784 16590
rect 21732 16526 21784 16532
rect 21548 16176 21600 16182
rect 21548 16118 21600 16124
rect 21456 16108 21508 16114
rect 21456 16050 21508 16056
rect 21468 15162 21496 16050
rect 21744 16046 21772 16526
rect 21732 16040 21784 16046
rect 21546 16008 21602 16017
rect 21732 15982 21784 15988
rect 21546 15943 21602 15952
rect 21560 15502 21588 15943
rect 21548 15496 21600 15502
rect 21548 15438 21600 15444
rect 21640 15360 21692 15366
rect 21836 15314 21864 16662
rect 21928 16250 21956 18634
rect 22468 18624 22520 18630
rect 22468 18566 22520 18572
rect 22192 18216 22244 18222
rect 22192 18158 22244 18164
rect 22376 18216 22428 18222
rect 22376 18158 22428 18164
rect 22204 18086 22232 18158
rect 22100 18080 22152 18086
rect 22100 18022 22152 18028
rect 22192 18080 22244 18086
rect 22192 18022 22244 18028
rect 22008 16448 22060 16454
rect 22008 16390 22060 16396
rect 21916 16244 21968 16250
rect 21916 16186 21968 16192
rect 22020 15706 22048 16390
rect 22008 15700 22060 15706
rect 22008 15642 22060 15648
rect 21640 15302 21692 15308
rect 21456 15156 21508 15162
rect 21456 15098 21508 15104
rect 21456 15020 21508 15026
rect 21456 14962 21508 14968
rect 21468 14618 21496 14962
rect 21456 14612 21508 14618
rect 21456 14554 21508 14560
rect 21548 14612 21600 14618
rect 21548 14554 21600 14560
rect 21560 14074 21588 14554
rect 21652 14414 21680 15302
rect 21744 15286 21956 15314
rect 21744 15162 21772 15286
rect 21732 15156 21784 15162
rect 21732 15098 21784 15104
rect 21824 15156 21876 15162
rect 21824 15098 21876 15104
rect 21732 14816 21784 14822
rect 21732 14758 21784 14764
rect 21744 14414 21772 14758
rect 21640 14408 21692 14414
rect 21640 14350 21692 14356
rect 21732 14408 21784 14414
rect 21732 14350 21784 14356
rect 21732 14272 21784 14278
rect 21732 14214 21784 14220
rect 21548 14068 21600 14074
rect 21548 14010 21600 14016
rect 21272 13728 21324 13734
rect 21272 13670 21324 13676
rect 21364 13728 21416 13734
rect 21364 13670 21416 13676
rect 21088 13388 21140 13394
rect 21088 13330 21140 13336
rect 20996 13320 21048 13326
rect 20996 13262 21048 13268
rect 21008 12986 21036 13262
rect 20996 12980 21048 12986
rect 20996 12922 21048 12928
rect 21100 12918 21128 13330
rect 21284 13326 21312 13670
rect 21560 13530 21588 14010
rect 21548 13524 21600 13530
rect 21548 13466 21600 13472
rect 21272 13320 21324 13326
rect 21272 13262 21324 13268
rect 21088 12912 21140 12918
rect 21088 12854 21140 12860
rect 21640 12776 21692 12782
rect 21640 12718 21692 12724
rect 21088 12640 21140 12646
rect 21088 12582 21140 12588
rect 20904 12232 20956 12238
rect 20904 12174 20956 12180
rect 20812 11688 20864 11694
rect 20812 11630 20864 11636
rect 20996 11552 21048 11558
rect 20996 11494 21048 11500
rect 20543 11452 20851 11461
rect 20543 11450 20549 11452
rect 20605 11450 20629 11452
rect 20685 11450 20709 11452
rect 20765 11450 20789 11452
rect 20845 11450 20851 11452
rect 20605 11398 20607 11450
rect 20787 11398 20789 11450
rect 20543 11396 20549 11398
rect 20605 11396 20629 11398
rect 20685 11396 20709 11398
rect 20765 11396 20789 11398
rect 20845 11396 20851 11398
rect 20543 11387 20851 11396
rect 20352 11280 20404 11286
rect 20352 11222 20404 11228
rect 20904 11280 20956 11286
rect 20904 11222 20956 11228
rect 19892 10532 19944 10538
rect 19892 10474 19944 10480
rect 19904 7886 19932 10474
rect 20260 10464 20312 10470
rect 20260 10406 20312 10412
rect 20076 9920 20128 9926
rect 20076 9862 20128 9868
rect 20088 9674 20116 9862
rect 20088 9646 20208 9674
rect 20180 9382 20208 9646
rect 20076 9376 20128 9382
rect 20076 9318 20128 9324
rect 20168 9376 20220 9382
rect 20168 9318 20220 9324
rect 19984 8832 20036 8838
rect 19984 8774 20036 8780
rect 19892 7880 19944 7886
rect 19892 7822 19944 7828
rect 19812 7500 19932 7528
rect 19616 7336 19668 7342
rect 19616 7278 19668 7284
rect 19432 7142 19484 7148
rect 19522 7168 19578 7177
rect 19444 7041 19472 7142
rect 19522 7103 19578 7112
rect 19430 7032 19486 7041
rect 19430 6967 19486 6976
rect 19798 7032 19854 7041
rect 19798 6967 19854 6976
rect 19248 6860 19300 6866
rect 19248 6802 19300 6808
rect 19156 6724 19208 6730
rect 19156 6666 19208 6672
rect 19064 6656 19116 6662
rect 19064 6598 19116 6604
rect 19168 6322 19196 6666
rect 19156 6316 19208 6322
rect 19156 6258 19208 6264
rect 18972 6248 19024 6254
rect 18972 6190 19024 6196
rect 19064 5296 19116 5302
rect 19064 5238 19116 5244
rect 18972 5228 19024 5234
rect 18972 5170 19024 5176
rect 18984 4690 19012 5170
rect 18972 4684 19024 4690
rect 18972 4626 19024 4632
rect 19076 4622 19104 5238
rect 19064 4616 19116 4622
rect 19064 4558 19116 4564
rect 19076 4298 19104 4558
rect 19168 4486 19196 6258
rect 19156 4480 19208 4486
rect 19156 4422 19208 4428
rect 18984 4282 19104 4298
rect 18972 4276 19104 4282
rect 19024 4270 19104 4276
rect 18972 4218 19024 4224
rect 18880 4140 18932 4146
rect 18880 4082 18932 4088
rect 19156 4140 19208 4146
rect 19156 4082 19208 4088
rect 19168 3670 19196 4082
rect 18972 3664 19024 3670
rect 19156 3664 19208 3670
rect 19024 3612 19104 3618
rect 18972 3606 19104 3612
rect 19156 3606 19208 3612
rect 18984 3590 19104 3606
rect 19076 3194 19104 3590
rect 19156 3528 19208 3534
rect 19156 3470 19208 3476
rect 18972 3188 19024 3194
rect 18972 3130 19024 3136
rect 19064 3188 19116 3194
rect 19064 3130 19116 3136
rect 18984 3074 19012 3130
rect 19168 3074 19196 3470
rect 18984 3046 19196 3074
rect 19260 3058 19288 6802
rect 19430 6488 19486 6497
rect 19812 6440 19840 6967
rect 19904 6882 19932 7500
rect 19996 7478 20024 8774
rect 19984 7472 20036 7478
rect 19984 7414 20036 7420
rect 19996 7041 20024 7414
rect 19982 7032 20038 7041
rect 19982 6967 20038 6976
rect 19904 6854 20024 6882
rect 19892 6792 19944 6798
rect 19892 6734 19944 6740
rect 19904 6497 19932 6734
rect 19430 6423 19432 6432
rect 19484 6423 19486 6432
rect 19432 6394 19484 6400
rect 19720 6412 19840 6440
rect 19890 6488 19946 6497
rect 19890 6423 19946 6432
rect 19616 6384 19668 6390
rect 19720 6372 19748 6412
rect 19668 6344 19748 6372
rect 19616 6326 19668 6332
rect 19800 6316 19852 6322
rect 19892 6316 19944 6322
rect 19852 6276 19892 6304
rect 19800 6258 19852 6264
rect 19892 6258 19944 6264
rect 19430 6080 19486 6089
rect 19430 6015 19486 6024
rect 19798 6080 19854 6089
rect 19798 6015 19854 6024
rect 19340 5704 19392 5710
rect 19340 5646 19392 5652
rect 19352 5370 19380 5646
rect 19340 5364 19392 5370
rect 19340 5306 19392 5312
rect 19444 5166 19472 6015
rect 19812 5778 19840 6015
rect 19800 5772 19852 5778
rect 19800 5714 19852 5720
rect 19708 5568 19760 5574
rect 19708 5510 19760 5516
rect 19720 5370 19748 5510
rect 19708 5364 19760 5370
rect 19708 5306 19760 5312
rect 19892 5228 19944 5234
rect 19892 5170 19944 5176
rect 19432 5160 19484 5166
rect 19432 5102 19484 5108
rect 19524 5160 19576 5166
rect 19524 5102 19576 5108
rect 19340 5092 19392 5098
rect 19340 5034 19392 5040
rect 19352 3942 19380 5034
rect 19536 4826 19564 5102
rect 19614 4856 19670 4865
rect 19524 4820 19576 4826
rect 19614 4791 19670 4800
rect 19524 4762 19576 4768
rect 19628 4622 19656 4791
rect 19616 4616 19668 4622
rect 19536 4576 19616 4604
rect 19432 4208 19484 4214
rect 19432 4150 19484 4156
rect 19340 3936 19392 3942
rect 19340 3878 19392 3884
rect 19444 3738 19472 4150
rect 19536 4078 19564 4576
rect 19616 4558 19668 4564
rect 19616 4480 19668 4486
rect 19616 4422 19668 4428
rect 19524 4072 19576 4078
rect 19524 4014 19576 4020
rect 19524 3936 19576 3942
rect 19524 3878 19576 3884
rect 19432 3732 19484 3738
rect 19432 3674 19484 3680
rect 19536 3602 19564 3878
rect 19524 3596 19576 3602
rect 19524 3538 19576 3544
rect 19628 3398 19656 4422
rect 19904 3398 19932 5170
rect 19996 5030 20024 6854
rect 20088 5778 20116 9318
rect 20180 8809 20208 9318
rect 20166 8800 20222 8809
rect 20166 8735 20222 8744
rect 20272 7818 20300 10406
rect 20364 8906 20392 11222
rect 20543 10364 20851 10373
rect 20543 10362 20549 10364
rect 20605 10362 20629 10364
rect 20685 10362 20709 10364
rect 20765 10362 20789 10364
rect 20845 10362 20851 10364
rect 20605 10310 20607 10362
rect 20787 10310 20789 10362
rect 20543 10308 20549 10310
rect 20605 10308 20629 10310
rect 20685 10308 20709 10310
rect 20765 10308 20789 10310
rect 20845 10308 20851 10310
rect 20543 10299 20851 10308
rect 20812 10260 20864 10266
rect 20812 10202 20864 10208
rect 20824 9926 20852 10202
rect 20720 9920 20772 9926
rect 20720 9862 20772 9868
rect 20812 9920 20864 9926
rect 20812 9862 20864 9868
rect 20732 9586 20760 9862
rect 20720 9580 20772 9586
rect 20720 9522 20772 9528
rect 20444 9376 20496 9382
rect 20444 9318 20496 9324
rect 20456 8956 20484 9318
rect 20543 9276 20851 9285
rect 20543 9274 20549 9276
rect 20605 9274 20629 9276
rect 20685 9274 20709 9276
rect 20765 9274 20789 9276
rect 20845 9274 20851 9276
rect 20605 9222 20607 9274
rect 20787 9222 20789 9274
rect 20543 9220 20549 9222
rect 20605 9220 20629 9222
rect 20685 9220 20709 9222
rect 20765 9220 20789 9222
rect 20845 9220 20851 9222
rect 20543 9211 20851 9220
rect 20916 9058 20944 11222
rect 21008 9994 21036 11494
rect 21100 11082 21128 12582
rect 21364 12368 21416 12374
rect 21364 12310 21416 12316
rect 21376 12209 21404 12310
rect 21652 12306 21680 12718
rect 21640 12300 21692 12306
rect 21640 12242 21692 12248
rect 21362 12200 21418 12209
rect 21362 12135 21418 12144
rect 21456 12096 21508 12102
rect 21456 12038 21508 12044
rect 21468 11898 21496 12038
rect 21456 11892 21508 11898
rect 21456 11834 21508 11840
rect 21364 11620 21416 11626
rect 21364 11562 21416 11568
rect 21272 11552 21324 11558
rect 21272 11494 21324 11500
rect 21284 11150 21312 11494
rect 21272 11144 21324 11150
rect 21376 11121 21404 11562
rect 21272 11086 21324 11092
rect 21362 11112 21418 11121
rect 21088 11076 21140 11082
rect 21362 11047 21418 11056
rect 21456 11076 21508 11082
rect 21088 11018 21140 11024
rect 21456 11018 21508 11024
rect 21468 10606 21496 11018
rect 21364 10600 21416 10606
rect 21364 10542 21416 10548
rect 21456 10600 21508 10606
rect 21456 10542 21508 10548
rect 21180 10464 21232 10470
rect 21180 10406 21232 10412
rect 21088 10056 21140 10062
rect 21088 9998 21140 10004
rect 20996 9988 21048 9994
rect 20996 9930 21048 9936
rect 20996 9716 21048 9722
rect 20996 9658 21048 9664
rect 20824 9030 20944 9058
rect 21008 9042 21036 9658
rect 20996 9036 21048 9042
rect 20536 8968 20588 8974
rect 20456 8928 20536 8956
rect 20536 8910 20588 8916
rect 20718 8936 20774 8945
rect 20352 8900 20404 8906
rect 20352 8842 20404 8848
rect 20364 8786 20392 8842
rect 20364 8758 20484 8786
rect 20456 8498 20484 8758
rect 20548 8634 20576 8910
rect 20718 8871 20774 8880
rect 20536 8628 20588 8634
rect 20536 8570 20588 8576
rect 20444 8492 20496 8498
rect 20444 8434 20496 8440
rect 20444 8288 20496 8294
rect 20732 8276 20760 8871
rect 20824 8430 20852 9030
rect 20996 8978 21048 8984
rect 21100 8974 21128 9998
rect 21088 8968 21140 8974
rect 21088 8910 21140 8916
rect 21192 8498 21220 10406
rect 21270 10160 21326 10169
rect 21270 10095 21272 10104
rect 21324 10095 21326 10104
rect 21272 10066 21324 10072
rect 21376 9722 21404 10542
rect 21744 10198 21772 14214
rect 21836 13870 21864 15098
rect 21928 14618 21956 15286
rect 21916 14612 21968 14618
rect 21916 14554 21968 14560
rect 22112 14226 22140 18022
rect 22388 17338 22416 18158
rect 22480 18154 22508 18566
rect 22468 18148 22520 18154
rect 22468 18090 22520 18096
rect 22572 18086 22600 20334
rect 22652 20256 22704 20262
rect 22652 20198 22704 20204
rect 22664 19281 22692 20198
rect 22650 19272 22706 19281
rect 22848 19242 22876 20402
rect 23020 20256 23072 20262
rect 23020 20198 23072 20204
rect 23032 19961 23060 20198
rect 23018 19952 23074 19961
rect 23018 19887 23074 19896
rect 22928 19848 22980 19854
rect 22928 19790 22980 19796
rect 22650 19207 22706 19216
rect 22836 19236 22888 19242
rect 22836 19178 22888 19184
rect 22744 19168 22796 19174
rect 22744 19110 22796 19116
rect 22652 18828 22704 18834
rect 22652 18770 22704 18776
rect 22560 18080 22612 18086
rect 22560 18022 22612 18028
rect 22664 17746 22692 18770
rect 22756 18426 22784 19110
rect 22744 18420 22796 18426
rect 22744 18362 22796 18368
rect 22652 17740 22704 17746
rect 22652 17682 22704 17688
rect 22652 17536 22704 17542
rect 22652 17478 22704 17484
rect 22376 17332 22428 17338
rect 22376 17274 22428 17280
rect 22192 17196 22244 17202
rect 22192 17138 22244 17144
rect 22204 16794 22232 17138
rect 22376 17128 22428 17134
rect 22376 17070 22428 17076
rect 22192 16788 22244 16794
rect 22192 16730 22244 16736
rect 22388 15978 22416 17070
rect 22560 16992 22612 16998
rect 22560 16934 22612 16940
rect 22376 15972 22428 15978
rect 22376 15914 22428 15920
rect 22468 15564 22520 15570
rect 22468 15506 22520 15512
rect 22284 15360 22336 15366
rect 22284 15302 22336 15308
rect 22376 15360 22428 15366
rect 22376 15302 22428 15308
rect 22192 14408 22244 14414
rect 22192 14350 22244 14356
rect 21928 14198 22140 14226
rect 21928 13938 21956 14198
rect 21916 13932 21968 13938
rect 21916 13874 21968 13880
rect 21824 13864 21876 13870
rect 21824 13806 21876 13812
rect 21824 13728 21876 13734
rect 21824 13670 21876 13676
rect 21836 11642 21864 13670
rect 21928 11830 21956 13874
rect 22098 13424 22154 13433
rect 22204 13394 22232 14350
rect 22296 13530 22324 15302
rect 22284 13524 22336 13530
rect 22284 13466 22336 13472
rect 22098 13359 22154 13368
rect 22192 13388 22244 13394
rect 22008 13184 22060 13190
rect 22006 13152 22008 13161
rect 22060 13152 22062 13161
rect 22006 13087 22062 13096
rect 22112 12986 22140 13359
rect 22192 13330 22244 13336
rect 22192 13252 22244 13258
rect 22192 13194 22244 13200
rect 22100 12980 22152 12986
rect 22100 12922 22152 12928
rect 22100 12640 22152 12646
rect 22100 12582 22152 12588
rect 21916 11824 21968 11830
rect 21916 11766 21968 11772
rect 21836 11614 21956 11642
rect 21824 11552 21876 11558
rect 21824 11494 21876 11500
rect 21836 10674 21864 11494
rect 21824 10668 21876 10674
rect 21824 10610 21876 10616
rect 21824 10532 21876 10538
rect 21824 10474 21876 10480
rect 21732 10192 21784 10198
rect 21732 10134 21784 10140
rect 21548 10124 21600 10130
rect 21548 10066 21600 10072
rect 21456 9920 21508 9926
rect 21456 9862 21508 9868
rect 21364 9716 21416 9722
rect 21364 9658 21416 9664
rect 21272 9376 21324 9382
rect 21272 9318 21324 9324
rect 20904 8492 20956 8498
rect 20904 8434 20956 8440
rect 21088 8492 21140 8498
rect 21088 8434 21140 8440
rect 21180 8492 21232 8498
rect 21180 8434 21232 8440
rect 20812 8424 20864 8430
rect 20812 8366 20864 8372
rect 20812 8288 20864 8294
rect 20732 8248 20812 8276
rect 20444 8230 20496 8236
rect 20812 8230 20864 8236
rect 20168 7812 20220 7818
rect 20168 7754 20220 7760
rect 20260 7812 20312 7818
rect 20260 7754 20312 7760
rect 20076 5772 20128 5778
rect 20076 5714 20128 5720
rect 20074 5672 20130 5681
rect 20074 5607 20130 5616
rect 19984 5024 20036 5030
rect 19984 4966 20036 4972
rect 19996 3398 20024 4966
rect 20088 4690 20116 5607
rect 20076 4684 20128 4690
rect 20076 4626 20128 4632
rect 20180 4026 20208 7754
rect 20272 5302 20300 7754
rect 20456 7410 20484 8230
rect 20543 8188 20851 8197
rect 20543 8186 20549 8188
rect 20605 8186 20629 8188
rect 20685 8186 20709 8188
rect 20765 8186 20789 8188
rect 20845 8186 20851 8188
rect 20605 8134 20607 8186
rect 20787 8134 20789 8186
rect 20543 8132 20549 8134
rect 20605 8132 20629 8134
rect 20685 8132 20709 8134
rect 20765 8132 20789 8134
rect 20845 8132 20851 8134
rect 20543 8123 20851 8132
rect 20628 7880 20680 7886
rect 20628 7822 20680 7828
rect 20444 7404 20496 7410
rect 20444 7346 20496 7352
rect 20352 7200 20404 7206
rect 20352 7142 20404 7148
rect 20364 6118 20392 7142
rect 20352 6112 20404 6118
rect 20352 6054 20404 6060
rect 20260 5296 20312 5302
rect 20260 5238 20312 5244
rect 20260 5092 20312 5098
rect 20260 5034 20312 5040
rect 20272 4826 20300 5034
rect 20260 4820 20312 4826
rect 20260 4762 20312 4768
rect 20364 4486 20392 6054
rect 20456 5681 20484 7346
rect 20640 7206 20668 7822
rect 20628 7200 20680 7206
rect 20628 7142 20680 7148
rect 20543 7100 20851 7109
rect 20543 7098 20549 7100
rect 20605 7098 20629 7100
rect 20685 7098 20709 7100
rect 20765 7098 20789 7100
rect 20845 7098 20851 7100
rect 20605 7046 20607 7098
rect 20787 7046 20789 7098
rect 20543 7044 20549 7046
rect 20605 7044 20629 7046
rect 20685 7044 20709 7046
rect 20765 7044 20789 7046
rect 20845 7044 20851 7046
rect 20543 7035 20851 7044
rect 20812 6928 20864 6934
rect 20812 6870 20864 6876
rect 20628 6860 20680 6866
rect 20628 6802 20680 6808
rect 20536 6724 20588 6730
rect 20536 6666 20588 6672
rect 20548 6458 20576 6666
rect 20536 6452 20588 6458
rect 20536 6394 20588 6400
rect 20548 6254 20576 6394
rect 20536 6248 20588 6254
rect 20536 6190 20588 6196
rect 20640 6118 20668 6802
rect 20720 6792 20772 6798
rect 20720 6734 20772 6740
rect 20732 6458 20760 6734
rect 20720 6452 20772 6458
rect 20720 6394 20772 6400
rect 20824 6202 20852 6870
rect 20916 6866 20944 8434
rect 20996 8356 21048 8362
rect 20996 8298 21048 8304
rect 20904 6860 20956 6866
rect 20904 6802 20956 6808
rect 21008 6746 21036 8298
rect 21100 7546 21128 8434
rect 21178 8392 21234 8401
rect 21178 8327 21234 8336
rect 21192 7834 21220 8327
rect 21284 7954 21312 9318
rect 21468 9178 21496 9862
rect 21456 9172 21508 9178
rect 21456 9114 21508 9120
rect 21468 8974 21496 9114
rect 21456 8968 21508 8974
rect 21456 8910 21508 8916
rect 21560 7970 21588 10066
rect 21640 9988 21692 9994
rect 21640 9930 21692 9936
rect 21652 9178 21680 9930
rect 21732 9512 21784 9518
rect 21732 9454 21784 9460
rect 21640 9172 21692 9178
rect 21640 9114 21692 9120
rect 21640 8832 21692 8838
rect 21640 8774 21692 8780
rect 21272 7948 21324 7954
rect 21272 7890 21324 7896
rect 21376 7942 21588 7970
rect 21192 7806 21312 7834
rect 21180 7744 21232 7750
rect 21180 7686 21232 7692
rect 21088 7540 21140 7546
rect 21088 7482 21140 7488
rect 21088 7200 21140 7206
rect 21088 7142 21140 7148
rect 20916 6730 21036 6746
rect 20904 6724 21036 6730
rect 20956 6718 21036 6724
rect 20904 6666 20956 6672
rect 20916 6322 20944 6666
rect 20996 6656 21048 6662
rect 20996 6598 21048 6604
rect 20904 6316 20956 6322
rect 20904 6258 20956 6264
rect 20824 6174 20944 6202
rect 20628 6112 20680 6118
rect 20628 6054 20680 6060
rect 20543 6012 20851 6021
rect 20543 6010 20549 6012
rect 20605 6010 20629 6012
rect 20685 6010 20709 6012
rect 20765 6010 20789 6012
rect 20845 6010 20851 6012
rect 20605 5958 20607 6010
rect 20787 5958 20789 6010
rect 20543 5956 20549 5958
rect 20605 5956 20629 5958
rect 20685 5956 20709 5958
rect 20765 5956 20789 5958
rect 20845 5956 20851 5958
rect 20543 5947 20851 5956
rect 20812 5840 20864 5846
rect 20812 5782 20864 5788
rect 20442 5672 20498 5681
rect 20442 5607 20498 5616
rect 20444 5568 20496 5574
rect 20444 5510 20496 5516
rect 20456 4690 20484 5510
rect 20824 5302 20852 5782
rect 20812 5296 20864 5302
rect 20812 5238 20864 5244
rect 20824 5012 20852 5238
rect 20916 5166 20944 6174
rect 20904 5160 20956 5166
rect 20904 5102 20956 5108
rect 20824 4984 20944 5012
rect 20543 4924 20851 4933
rect 20543 4922 20549 4924
rect 20605 4922 20629 4924
rect 20685 4922 20709 4924
rect 20765 4922 20789 4924
rect 20845 4922 20851 4924
rect 20605 4870 20607 4922
rect 20787 4870 20789 4922
rect 20543 4868 20549 4870
rect 20605 4868 20629 4870
rect 20685 4868 20709 4870
rect 20765 4868 20789 4870
rect 20845 4868 20851 4870
rect 20543 4859 20851 4868
rect 20534 4720 20590 4729
rect 20444 4684 20496 4690
rect 20534 4655 20590 4664
rect 20444 4626 20496 4632
rect 20352 4480 20404 4486
rect 20352 4422 20404 4428
rect 20180 3998 20300 4026
rect 20168 3936 20220 3942
rect 20168 3878 20220 3884
rect 20180 3466 20208 3878
rect 20272 3670 20300 3998
rect 20364 3738 20392 4422
rect 20548 3942 20576 4655
rect 20812 4616 20864 4622
rect 20812 4558 20864 4564
rect 20824 4486 20852 4558
rect 20812 4480 20864 4486
rect 20812 4422 20864 4428
rect 20444 3936 20496 3942
rect 20444 3878 20496 3884
rect 20536 3936 20588 3942
rect 20536 3878 20588 3884
rect 20352 3732 20404 3738
rect 20352 3674 20404 3680
rect 20260 3664 20312 3670
rect 20260 3606 20312 3612
rect 20456 3602 20484 3878
rect 20543 3836 20851 3845
rect 20543 3834 20549 3836
rect 20605 3834 20629 3836
rect 20685 3834 20709 3836
rect 20765 3834 20789 3836
rect 20845 3834 20851 3836
rect 20605 3782 20607 3834
rect 20787 3782 20789 3834
rect 20543 3780 20549 3782
rect 20605 3780 20629 3782
rect 20685 3780 20709 3782
rect 20765 3780 20789 3782
rect 20845 3780 20851 3782
rect 20543 3771 20851 3780
rect 20444 3596 20496 3602
rect 20444 3538 20496 3544
rect 20916 3534 20944 4984
rect 20904 3528 20956 3534
rect 20904 3470 20956 3476
rect 20168 3460 20220 3466
rect 20168 3402 20220 3408
rect 19616 3392 19668 3398
rect 19616 3334 19668 3340
rect 19892 3392 19944 3398
rect 19892 3334 19944 3340
rect 19984 3392 20036 3398
rect 19984 3334 20036 3340
rect 21008 3097 21036 6598
rect 21100 4486 21128 7142
rect 21192 4486 21220 7686
rect 21284 7274 21312 7806
rect 21272 7268 21324 7274
rect 21272 7210 21324 7216
rect 21284 6934 21312 7210
rect 21272 6928 21324 6934
rect 21272 6870 21324 6876
rect 21272 6656 21324 6662
rect 21270 6624 21272 6633
rect 21324 6624 21326 6633
rect 21270 6559 21326 6568
rect 21272 6316 21324 6322
rect 21272 6258 21324 6264
rect 21284 6089 21312 6258
rect 21270 6080 21326 6089
rect 21270 6015 21326 6024
rect 21272 5228 21324 5234
rect 21272 5170 21324 5176
rect 21088 4480 21140 4486
rect 21088 4422 21140 4428
rect 21180 4480 21232 4486
rect 21180 4422 21232 4428
rect 19706 3088 19762 3097
rect 19248 3052 19300 3058
rect 19706 3023 19708 3032
rect 19248 2994 19300 3000
rect 19760 3023 19762 3032
rect 20994 3088 21050 3097
rect 20994 3023 21050 3032
rect 19708 2994 19760 3000
rect 21100 2990 21128 4422
rect 21192 3194 21220 4422
rect 21284 4282 21312 5170
rect 21376 4622 21404 7942
rect 21548 7880 21600 7886
rect 21548 7822 21600 7828
rect 21456 7472 21508 7478
rect 21560 7449 21588 7822
rect 21456 7414 21508 7420
rect 21546 7440 21602 7449
rect 21468 6848 21496 7414
rect 21546 7375 21548 7384
rect 21600 7375 21602 7384
rect 21548 7346 21600 7352
rect 21468 6820 21588 6848
rect 21456 6724 21508 6730
rect 21456 6666 21508 6672
rect 21468 6458 21496 6666
rect 21456 6452 21508 6458
rect 21456 6394 21508 6400
rect 21454 6352 21510 6361
rect 21454 6287 21510 6296
rect 21468 5778 21496 6287
rect 21560 6202 21588 6820
rect 21652 6458 21680 8774
rect 21744 8634 21772 9454
rect 21836 9042 21864 10474
rect 21928 10266 21956 11614
rect 22112 10810 22140 12582
rect 22204 11762 22232 13194
rect 22388 12986 22416 15302
rect 22480 14958 22508 15506
rect 22468 14952 22520 14958
rect 22468 14894 22520 14900
rect 22376 12980 22428 12986
rect 22376 12922 22428 12928
rect 22480 12866 22508 14894
rect 22572 14006 22600 16934
rect 22664 16590 22692 17478
rect 22756 17134 22784 18362
rect 22836 18284 22888 18290
rect 22836 18226 22888 18232
rect 22744 17128 22796 17134
rect 22744 17070 22796 17076
rect 22756 16794 22784 17070
rect 22744 16788 22796 16794
rect 22744 16730 22796 16736
rect 22652 16584 22704 16590
rect 22652 16526 22704 16532
rect 22652 15360 22704 15366
rect 22652 15302 22704 15308
rect 22560 14000 22612 14006
rect 22560 13942 22612 13948
rect 22572 13462 22600 13942
rect 22664 13734 22692 15302
rect 22744 14612 22796 14618
rect 22744 14554 22796 14560
rect 22652 13728 22704 13734
rect 22652 13670 22704 13676
rect 22560 13456 22612 13462
rect 22560 13398 22612 13404
rect 22652 13388 22704 13394
rect 22652 13330 22704 13336
rect 22664 13274 22692 13330
rect 22388 12838 22508 12866
rect 22572 13246 22692 13274
rect 22284 12096 22336 12102
rect 22284 12038 22336 12044
rect 22192 11756 22244 11762
rect 22192 11698 22244 11704
rect 22296 11082 22324 12038
rect 22388 11694 22416 12838
rect 22468 12776 22520 12782
rect 22468 12718 22520 12724
rect 22480 11830 22508 12718
rect 22468 11824 22520 11830
rect 22468 11766 22520 11772
rect 22376 11688 22428 11694
rect 22376 11630 22428 11636
rect 22388 11218 22416 11630
rect 22468 11620 22520 11626
rect 22468 11562 22520 11568
rect 22376 11212 22428 11218
rect 22376 11154 22428 11160
rect 22284 11076 22336 11082
rect 22284 11018 22336 11024
rect 22480 10810 22508 11562
rect 22100 10804 22152 10810
rect 22100 10746 22152 10752
rect 22468 10804 22520 10810
rect 22468 10746 22520 10752
rect 22284 10736 22336 10742
rect 22284 10678 22336 10684
rect 22192 10600 22244 10606
rect 22192 10542 22244 10548
rect 22008 10464 22060 10470
rect 22008 10406 22060 10412
rect 22100 10464 22152 10470
rect 22100 10406 22152 10412
rect 21916 10260 21968 10266
rect 21916 10202 21968 10208
rect 21824 9036 21876 9042
rect 21824 8978 21876 8984
rect 21732 8628 21784 8634
rect 21732 8570 21784 8576
rect 21732 8492 21784 8498
rect 21732 8434 21784 8440
rect 21640 6452 21692 6458
rect 21640 6394 21692 6400
rect 21560 6174 21680 6202
rect 21546 6080 21602 6089
rect 21546 6015 21602 6024
rect 21560 5914 21588 6015
rect 21548 5908 21600 5914
rect 21548 5850 21600 5856
rect 21456 5772 21508 5778
rect 21456 5714 21508 5720
rect 21456 5024 21508 5030
rect 21456 4966 21508 4972
rect 21364 4616 21416 4622
rect 21364 4558 21416 4564
rect 21468 4486 21496 4966
rect 21456 4480 21508 4486
rect 21362 4448 21418 4457
rect 21456 4422 21508 4428
rect 21362 4383 21418 4392
rect 21272 4276 21324 4282
rect 21272 4218 21324 4224
rect 21376 3602 21404 4383
rect 21454 4176 21510 4185
rect 21454 4111 21510 4120
rect 21364 3596 21416 3602
rect 21364 3538 21416 3544
rect 21468 3534 21496 4111
rect 21456 3528 21508 3534
rect 21456 3470 21508 3476
rect 21180 3188 21232 3194
rect 21180 3130 21232 3136
rect 21560 3058 21588 5850
rect 21652 5098 21680 6174
rect 21744 5574 21772 8434
rect 21928 7954 21956 10202
rect 22020 10062 22048 10406
rect 22008 10056 22060 10062
rect 22008 9998 22060 10004
rect 22112 9586 22140 10406
rect 22204 10130 22232 10542
rect 22192 10124 22244 10130
rect 22192 10066 22244 10072
rect 22204 9722 22232 10066
rect 22192 9716 22244 9722
rect 22192 9658 22244 9664
rect 22100 9580 22152 9586
rect 22100 9522 22152 9528
rect 22296 9382 22324 10678
rect 22376 10464 22428 10470
rect 22376 10406 22428 10412
rect 22388 10130 22416 10406
rect 22376 10124 22428 10130
rect 22376 10066 22428 10072
rect 22466 9888 22522 9897
rect 22466 9823 22522 9832
rect 22192 9376 22244 9382
rect 22192 9318 22244 9324
rect 22284 9376 22336 9382
rect 22284 9318 22336 9324
rect 22204 9110 22232 9318
rect 22192 9104 22244 9110
rect 22192 9046 22244 9052
rect 22192 8900 22244 8906
rect 22192 8842 22244 8848
rect 22204 8022 22232 8842
rect 22374 8800 22430 8809
rect 22374 8735 22430 8744
rect 22192 8016 22244 8022
rect 22192 7958 22244 7964
rect 21916 7948 21968 7954
rect 21916 7890 21968 7896
rect 21824 7880 21876 7886
rect 21824 7822 21876 7828
rect 21732 5568 21784 5574
rect 21836 5556 21864 7822
rect 22192 7404 22244 7410
rect 22192 7346 22244 7352
rect 22100 7336 22152 7342
rect 22100 7278 22152 7284
rect 22112 6866 22140 7278
rect 22100 6860 22152 6866
rect 22100 6802 22152 6808
rect 22008 6656 22060 6662
rect 21914 6624 21970 6633
rect 22008 6598 22060 6604
rect 21914 6559 21970 6568
rect 21928 6118 21956 6559
rect 21916 6112 21968 6118
rect 21916 6054 21968 6060
rect 21836 5528 21956 5556
rect 21732 5510 21784 5516
rect 21640 5092 21692 5098
rect 21640 5034 21692 5040
rect 21824 5024 21876 5030
rect 21824 4966 21876 4972
rect 21640 4616 21692 4622
rect 21640 4558 21692 4564
rect 21652 3398 21680 4558
rect 21836 4146 21864 4966
rect 21928 4146 21956 5528
rect 22020 4282 22048 6598
rect 22098 6488 22154 6497
rect 22098 6423 22154 6432
rect 22112 5846 22140 6423
rect 22100 5840 22152 5846
rect 22100 5782 22152 5788
rect 22008 4276 22060 4282
rect 22008 4218 22060 4224
rect 21824 4140 21876 4146
rect 21824 4082 21876 4088
rect 21916 4140 21968 4146
rect 21916 4082 21968 4088
rect 22204 3602 22232 7346
rect 22388 6254 22416 8735
rect 22480 8566 22508 9823
rect 22468 8560 22520 8566
rect 22468 8502 22520 8508
rect 22572 8430 22600 13246
rect 22652 13184 22704 13190
rect 22652 13126 22704 13132
rect 22664 12238 22692 13126
rect 22652 12232 22704 12238
rect 22652 12174 22704 12180
rect 22652 11552 22704 11558
rect 22652 11494 22704 11500
rect 22664 10810 22692 11494
rect 22756 11354 22784 14554
rect 22848 13818 22876 18226
rect 22940 17921 22968 19790
rect 23020 19712 23072 19718
rect 23020 19654 23072 19660
rect 23032 19417 23060 19654
rect 23018 19408 23074 19417
rect 23018 19343 23074 19352
rect 23020 19168 23072 19174
rect 23020 19110 23072 19116
rect 23032 18873 23060 19110
rect 23018 18864 23074 18873
rect 23018 18799 23074 18808
rect 23020 18420 23072 18426
rect 23020 18362 23072 18368
rect 23032 18329 23060 18362
rect 23018 18320 23074 18329
rect 23018 18255 23074 18264
rect 22926 17912 22982 17921
rect 22926 17847 22982 17856
rect 22928 17740 22980 17746
rect 22928 17682 22980 17688
rect 22940 17338 22968 17682
rect 23124 17649 23152 20810
rect 23216 17785 23244 21014
rect 23492 20330 23520 23800
rect 24136 22098 24164 23800
rect 24124 22092 24176 22098
rect 24124 22034 24176 22040
rect 23480 20324 23532 20330
rect 23480 20266 23532 20272
rect 23202 17776 23258 17785
rect 23202 17711 23258 17720
rect 23110 17640 23166 17649
rect 23110 17575 23166 17584
rect 22928 17332 22980 17338
rect 22928 17274 22980 17280
rect 23204 16584 23256 16590
rect 23204 16526 23256 16532
rect 23020 16448 23072 16454
rect 23020 16390 23072 16396
rect 22928 15904 22980 15910
rect 22928 15846 22980 15852
rect 22940 15094 22968 15846
rect 22928 15088 22980 15094
rect 22928 15030 22980 15036
rect 22928 14408 22980 14414
rect 22928 14350 22980 14356
rect 22940 14074 22968 14350
rect 22928 14068 22980 14074
rect 22928 14010 22980 14016
rect 22848 13790 22968 13818
rect 22836 13728 22888 13734
rect 22836 13670 22888 13676
rect 22848 12306 22876 13670
rect 22940 13530 22968 13790
rect 22928 13524 22980 13530
rect 22928 13466 22980 13472
rect 22836 12300 22888 12306
rect 22836 12242 22888 12248
rect 22928 11756 22980 11762
rect 22928 11698 22980 11704
rect 22744 11348 22796 11354
rect 22744 11290 22796 11296
rect 22940 11286 22968 11698
rect 22928 11280 22980 11286
rect 22928 11222 22980 11228
rect 22652 10804 22704 10810
rect 22652 10746 22704 10752
rect 22836 9920 22888 9926
rect 22836 9862 22888 9868
rect 22928 9920 22980 9926
rect 22928 9862 22980 9868
rect 22742 9752 22798 9761
rect 22848 9722 22876 9862
rect 22742 9687 22798 9696
rect 22836 9716 22888 9722
rect 22756 8974 22784 9687
rect 22836 9658 22888 9664
rect 22940 9518 22968 9862
rect 23032 9586 23060 16390
rect 23112 16108 23164 16114
rect 23112 16050 23164 16056
rect 23124 14822 23152 16050
rect 23216 15065 23244 16526
rect 23296 15632 23348 15638
rect 23296 15574 23348 15580
rect 23202 15056 23258 15065
rect 23202 14991 23258 15000
rect 23112 14816 23164 14822
rect 23112 14758 23164 14764
rect 23124 14521 23152 14758
rect 23110 14512 23166 14521
rect 23110 14447 23166 14456
rect 23112 13932 23164 13938
rect 23112 13874 23164 13880
rect 23124 12986 23152 13874
rect 23202 13424 23258 13433
rect 23202 13359 23258 13368
rect 23112 12980 23164 12986
rect 23112 12922 23164 12928
rect 23216 12918 23244 13359
rect 23204 12912 23256 12918
rect 23204 12854 23256 12860
rect 23204 12776 23256 12782
rect 23204 12718 23256 12724
rect 23216 11762 23244 12718
rect 23204 11756 23256 11762
rect 23204 11698 23256 11704
rect 23308 10674 23336 15574
rect 23664 15564 23716 15570
rect 23664 15506 23716 15512
rect 23388 14884 23440 14890
rect 23388 14826 23440 14832
rect 23400 12782 23428 14826
rect 23480 14544 23532 14550
rect 23480 14486 23532 14492
rect 23492 13977 23520 14486
rect 23478 13968 23534 13977
rect 23478 13903 23534 13912
rect 23492 12850 23520 13903
rect 23480 12844 23532 12850
rect 23480 12786 23532 12792
rect 23388 12776 23440 12782
rect 23388 12718 23440 12724
rect 23676 12434 23704 15506
rect 23584 12406 23704 12434
rect 23480 12096 23532 12102
rect 23480 12038 23532 12044
rect 23296 10668 23348 10674
rect 23296 10610 23348 10616
rect 23020 9580 23072 9586
rect 23020 9522 23072 9528
rect 22928 9512 22980 9518
rect 22928 9454 22980 9460
rect 23110 9480 23166 9489
rect 23110 9415 23166 9424
rect 23204 9444 23256 9450
rect 22744 8968 22796 8974
rect 22744 8910 22796 8916
rect 22650 8528 22706 8537
rect 22706 8472 22784 8480
rect 22650 8463 22652 8472
rect 22704 8452 22784 8472
rect 22652 8434 22704 8440
rect 22560 8424 22612 8430
rect 22560 8366 22612 8372
rect 22468 8356 22520 8362
rect 22468 8298 22520 8304
rect 22480 7002 22508 8298
rect 22560 8288 22612 8294
rect 22560 8230 22612 8236
rect 22572 7274 22600 8230
rect 22652 7744 22704 7750
rect 22652 7686 22704 7692
rect 22560 7268 22612 7274
rect 22560 7210 22612 7216
rect 22468 6996 22520 7002
rect 22468 6938 22520 6944
rect 22468 6792 22520 6798
rect 22466 6760 22468 6769
rect 22520 6760 22522 6769
rect 22466 6695 22522 6704
rect 22468 6316 22520 6322
rect 22468 6258 22520 6264
rect 22284 6248 22336 6254
rect 22284 6190 22336 6196
rect 22376 6248 22428 6254
rect 22376 6190 22428 6196
rect 22296 4010 22324 6190
rect 22376 5160 22428 5166
rect 22376 5102 22428 5108
rect 22388 4826 22416 5102
rect 22376 4820 22428 4826
rect 22376 4762 22428 4768
rect 22376 4276 22428 4282
rect 22376 4218 22428 4224
rect 22284 4004 22336 4010
rect 22284 3946 22336 3952
rect 22192 3596 22244 3602
rect 22192 3538 22244 3544
rect 22388 3505 22416 4218
rect 22480 3738 22508 6258
rect 22572 5710 22600 7210
rect 22664 7206 22692 7686
rect 22652 7200 22704 7206
rect 22652 7142 22704 7148
rect 22664 6186 22692 7142
rect 22652 6180 22704 6186
rect 22652 6122 22704 6128
rect 22664 5914 22692 6122
rect 22652 5908 22704 5914
rect 22652 5850 22704 5856
rect 22560 5704 22612 5710
rect 22560 5646 22612 5652
rect 22652 5568 22704 5574
rect 22652 5510 22704 5516
rect 22560 5092 22612 5098
rect 22560 5034 22612 5040
rect 22572 4214 22600 5034
rect 22560 4208 22612 4214
rect 22560 4150 22612 4156
rect 22468 3732 22520 3738
rect 22468 3674 22520 3680
rect 22560 3664 22612 3670
rect 22558 3632 22560 3641
rect 22612 3632 22614 3641
rect 22558 3567 22614 3576
rect 22374 3496 22430 3505
rect 22374 3431 22430 3440
rect 21640 3392 21692 3398
rect 21640 3334 21692 3340
rect 22664 3126 22692 5510
rect 22756 5370 22784 8452
rect 22836 8084 22888 8090
rect 22836 8026 22888 8032
rect 22848 6798 22876 8026
rect 23018 7984 23074 7993
rect 23018 7919 23074 7928
rect 23032 7886 23060 7919
rect 23020 7880 23072 7886
rect 23020 7822 23072 7828
rect 23020 7540 23072 7546
rect 23020 7482 23072 7488
rect 23032 7449 23060 7482
rect 23018 7440 23074 7449
rect 22928 7404 22980 7410
rect 23018 7375 23074 7384
rect 22928 7346 22980 7352
rect 22836 6792 22888 6798
rect 22836 6734 22888 6740
rect 22836 6656 22888 6662
rect 22836 6598 22888 6604
rect 22848 6361 22876 6598
rect 22834 6352 22890 6361
rect 22834 6287 22890 6296
rect 22836 6112 22888 6118
rect 22836 6054 22888 6060
rect 22744 5364 22796 5370
rect 22744 5306 22796 5312
rect 22756 3194 22784 5306
rect 22848 5234 22876 6054
rect 22836 5228 22888 5234
rect 22836 5170 22888 5176
rect 22940 3466 22968 7346
rect 23018 6896 23074 6905
rect 23018 6831 23074 6840
rect 23032 6662 23060 6831
rect 23020 6656 23072 6662
rect 23020 6598 23072 6604
rect 23020 6112 23072 6118
rect 23020 6054 23072 6060
rect 23032 5817 23060 6054
rect 23018 5808 23074 5817
rect 23018 5743 23074 5752
rect 23124 5642 23152 9415
rect 23204 9386 23256 9392
rect 23216 5778 23244 9386
rect 23296 8016 23348 8022
rect 23296 7958 23348 7964
rect 23204 5772 23256 5778
rect 23204 5714 23256 5720
rect 23112 5636 23164 5642
rect 23112 5578 23164 5584
rect 23020 5568 23072 5574
rect 23020 5510 23072 5516
rect 23032 5273 23060 5510
rect 23018 5264 23074 5273
rect 23018 5199 23074 5208
rect 23020 5024 23072 5030
rect 23020 4966 23072 4972
rect 23032 4729 23060 4966
rect 23018 4720 23074 4729
rect 23308 4690 23336 7958
rect 23388 6316 23440 6322
rect 23388 6258 23440 6264
rect 23400 6225 23428 6258
rect 23386 6216 23442 6225
rect 23386 6151 23442 6160
rect 23018 4655 23074 4664
rect 23296 4684 23348 4690
rect 23296 4626 23348 4632
rect 23020 4480 23072 4486
rect 23020 4422 23072 4428
rect 23032 4185 23060 4422
rect 23018 4176 23074 4185
rect 23018 4111 23074 4120
rect 23020 3936 23072 3942
rect 23020 3878 23072 3884
rect 23032 3641 23060 3878
rect 23018 3632 23074 3641
rect 23018 3567 23074 3576
rect 23112 3528 23164 3534
rect 23112 3470 23164 3476
rect 22928 3460 22980 3466
rect 22928 3402 22980 3408
rect 23020 3392 23072 3398
rect 23020 3334 23072 3340
rect 22744 3188 22796 3194
rect 22744 3130 22796 3136
rect 22652 3120 22704 3126
rect 23032 3097 23060 3334
rect 22652 3062 22704 3068
rect 23018 3088 23074 3097
rect 21548 3052 21600 3058
rect 23018 3023 23074 3032
rect 21548 2994 21600 3000
rect 18788 2984 18840 2990
rect 18788 2926 18840 2932
rect 21088 2984 21140 2990
rect 21088 2926 21140 2932
rect 22652 2984 22704 2990
rect 22652 2926 22704 2932
rect 18328 2848 18380 2854
rect 18328 2790 18380 2796
rect 18420 2848 18472 2854
rect 18420 2790 18472 2796
rect 18696 2848 18748 2854
rect 18696 2790 18748 2796
rect 20543 2748 20851 2757
rect 20543 2746 20549 2748
rect 20605 2746 20629 2748
rect 20685 2746 20709 2748
rect 20765 2746 20789 2748
rect 20845 2746 20851 2748
rect 20605 2694 20607 2746
rect 20787 2694 20789 2746
rect 20543 2692 20549 2694
rect 20605 2692 20629 2694
rect 20685 2692 20709 2694
rect 20765 2692 20789 2694
rect 20845 2692 20851 2694
rect 20543 2683 20851 2692
rect 10784 2644 10836 2650
rect 10784 2586 10836 2592
rect 15752 2644 15804 2650
rect 15752 2586 15804 2592
rect 16764 2644 16816 2650
rect 16764 2586 16816 2592
rect 8392 2508 8444 2514
rect 8392 2450 8444 2456
rect 22664 2446 22692 2926
rect 23124 2854 23152 3470
rect 23400 2990 23428 6151
rect 23492 5846 23520 12038
rect 23584 9178 23612 12406
rect 23662 11656 23718 11665
rect 23718 11614 23796 11642
rect 23662 11591 23718 11600
rect 23572 9172 23624 9178
rect 23572 9114 23624 9120
rect 23664 9104 23716 9110
rect 23664 9046 23716 9052
rect 23572 7744 23624 7750
rect 23572 7686 23624 7692
rect 23480 5840 23532 5846
rect 23480 5782 23532 5788
rect 23584 3738 23612 7686
rect 23572 3732 23624 3738
rect 23572 3674 23624 3680
rect 23676 3670 23704 9046
rect 23768 4282 23796 11614
rect 23848 9172 23900 9178
rect 23848 9114 23900 9120
rect 23756 4276 23808 4282
rect 23756 4218 23808 4224
rect 23664 3664 23716 3670
rect 23664 3606 23716 3612
rect 23388 2984 23440 2990
rect 23388 2926 23440 2932
rect 23860 2854 23888 9114
rect 23020 2848 23072 2854
rect 23020 2790 23072 2796
rect 23112 2848 23164 2854
rect 23112 2790 23164 2796
rect 23848 2848 23900 2854
rect 23848 2790 23900 2796
rect 23032 2553 23060 2790
rect 23124 2650 23152 2790
rect 23112 2644 23164 2650
rect 23112 2586 23164 2592
rect 23018 2544 23074 2553
rect 23018 2479 23074 2488
rect 6184 2440 6236 2446
rect 6184 2382 6236 2388
rect 22652 2440 22704 2446
rect 22652 2382 22704 2388
rect 2136 2304 2188 2310
rect 2136 2246 2188 2252
rect 2148 800 2176 2246
rect 6196 800 6224 2382
rect 10232 2304 10284 2310
rect 10232 2246 10284 2252
rect 22376 2304 22428 2310
rect 22376 2246 22428 2252
rect 6548 2204 6856 2213
rect 6548 2202 6554 2204
rect 6610 2202 6634 2204
rect 6690 2202 6714 2204
rect 6770 2202 6794 2204
rect 6850 2202 6856 2204
rect 6610 2150 6612 2202
rect 6792 2150 6794 2202
rect 6548 2148 6554 2150
rect 6610 2148 6634 2150
rect 6690 2148 6714 2150
rect 6770 2148 6794 2150
rect 6850 2148 6856 2150
rect 6548 2139 6856 2148
rect 10244 800 10272 2246
rect 12146 2204 12454 2213
rect 12146 2202 12152 2204
rect 12208 2202 12232 2204
rect 12288 2202 12312 2204
rect 12368 2202 12392 2204
rect 12448 2202 12454 2204
rect 12208 2150 12210 2202
rect 12390 2150 12392 2202
rect 12146 2148 12152 2150
rect 12208 2148 12232 2150
rect 12288 2148 12312 2150
rect 12368 2148 12392 2150
rect 12448 2148 12454 2150
rect 12146 2139 12454 2148
rect 17744 2204 18052 2213
rect 17744 2202 17750 2204
rect 17806 2202 17830 2204
rect 17886 2202 17910 2204
rect 17966 2202 17990 2204
rect 18046 2202 18052 2204
rect 17806 2150 17808 2202
rect 17988 2150 17990 2202
rect 17744 2148 17750 2150
rect 17806 2148 17830 2150
rect 17886 2148 17910 2150
rect 17966 2148 17990 2150
rect 18046 2148 18052 2150
rect 17744 2139 18052 2148
rect 22388 800 22416 2246
rect 2134 0 2190 800
rect 6182 0 6238 800
rect 10230 0 10286 800
rect 14278 0 14334 800
rect 18326 0 18382 800
rect 22374 0 22430 800
<< via2 >>
rect 3755 22330 3811 22332
rect 3835 22330 3891 22332
rect 3915 22330 3971 22332
rect 3995 22330 4051 22332
rect 3755 22278 3801 22330
rect 3801 22278 3811 22330
rect 3835 22278 3865 22330
rect 3865 22278 3877 22330
rect 3877 22278 3891 22330
rect 3915 22278 3929 22330
rect 3929 22278 3941 22330
rect 3941 22278 3971 22330
rect 3995 22278 4005 22330
rect 4005 22278 4051 22330
rect 3755 22276 3811 22278
rect 3835 22276 3891 22278
rect 3915 22276 3971 22278
rect 3995 22276 4051 22278
rect 3974 21548 4030 21584
rect 3974 21528 3976 21548
rect 3976 21528 4028 21548
rect 4028 21528 4030 21548
rect 2778 21020 2780 21040
rect 2780 21020 2832 21040
rect 2832 21020 2834 21040
rect 2778 20984 2834 21020
rect 1490 15308 1492 15328
rect 1492 15308 1544 15328
rect 1544 15308 1546 15328
rect 1490 15272 1546 15308
rect 2686 19372 2742 19408
rect 2686 19352 2688 19372
rect 2688 19352 2740 19372
rect 2740 19352 2742 19372
rect 2686 18672 2742 18728
rect 2410 16360 2466 16416
rect 3755 21242 3811 21244
rect 3835 21242 3891 21244
rect 3915 21242 3971 21244
rect 3995 21242 4051 21244
rect 3755 21190 3801 21242
rect 3801 21190 3811 21242
rect 3835 21190 3865 21242
rect 3865 21190 3877 21242
rect 3877 21190 3891 21242
rect 3915 21190 3929 21242
rect 3929 21190 3941 21242
rect 3941 21190 3971 21242
rect 3995 21190 4005 21242
rect 4005 21190 4051 21242
rect 3755 21188 3811 21190
rect 3835 21188 3891 21190
rect 3915 21188 3971 21190
rect 3995 21188 4051 21190
rect 4342 21392 4398 21448
rect 4250 21256 4306 21312
rect 3698 20884 3700 20904
rect 3700 20884 3752 20904
rect 3752 20884 3754 20904
rect 3698 20848 3754 20884
rect 3882 20440 3938 20496
rect 3755 20154 3811 20156
rect 3835 20154 3891 20156
rect 3915 20154 3971 20156
rect 3995 20154 4051 20156
rect 3755 20102 3801 20154
rect 3801 20102 3811 20154
rect 3835 20102 3865 20154
rect 3865 20102 3877 20154
rect 3877 20102 3891 20154
rect 3915 20102 3929 20154
rect 3929 20102 3941 20154
rect 3941 20102 3971 20154
rect 3995 20102 4005 20154
rect 4005 20102 4051 20154
rect 3755 20100 3811 20102
rect 3835 20100 3891 20102
rect 3915 20100 3971 20102
rect 3995 20100 4051 20102
rect 3755 19066 3811 19068
rect 3835 19066 3891 19068
rect 3915 19066 3971 19068
rect 3995 19066 4051 19068
rect 3755 19014 3801 19066
rect 3801 19014 3811 19066
rect 3835 19014 3865 19066
rect 3865 19014 3877 19066
rect 3877 19014 3891 19066
rect 3915 19014 3929 19066
rect 3929 19014 3941 19066
rect 3941 19014 3971 19066
rect 3995 19014 4005 19066
rect 4005 19014 4051 19066
rect 3755 19012 3811 19014
rect 3835 19012 3891 19014
rect 3915 19012 3971 19014
rect 3995 19012 4051 19014
rect 4434 19760 4490 19816
rect 3755 17978 3811 17980
rect 3835 17978 3891 17980
rect 3915 17978 3971 17980
rect 3995 17978 4051 17980
rect 3755 17926 3801 17978
rect 3801 17926 3811 17978
rect 3835 17926 3865 17978
rect 3865 17926 3877 17978
rect 3877 17926 3891 17978
rect 3915 17926 3929 17978
rect 3929 17926 3941 17978
rect 3941 17926 3971 17978
rect 3995 17926 4005 17978
rect 4005 17926 4051 17978
rect 3755 17924 3811 17926
rect 3835 17924 3891 17926
rect 3915 17924 3971 17926
rect 3995 17924 4051 17926
rect 3755 16890 3811 16892
rect 3835 16890 3891 16892
rect 3915 16890 3971 16892
rect 3995 16890 4051 16892
rect 3755 16838 3801 16890
rect 3801 16838 3811 16890
rect 3835 16838 3865 16890
rect 3865 16838 3877 16890
rect 3877 16838 3891 16890
rect 3915 16838 3929 16890
rect 3929 16838 3941 16890
rect 3941 16838 3971 16890
rect 3995 16838 4005 16890
rect 4005 16838 4051 16890
rect 3755 16836 3811 16838
rect 3835 16836 3891 16838
rect 3915 16836 3971 16838
rect 3995 16836 4051 16838
rect 3238 15444 3240 15464
rect 3240 15444 3292 15464
rect 3292 15444 3294 15464
rect 1398 9152 1454 9208
rect 3238 15408 3294 15444
rect 3755 15802 3811 15804
rect 3835 15802 3891 15804
rect 3915 15802 3971 15804
rect 3995 15802 4051 15804
rect 3755 15750 3801 15802
rect 3801 15750 3811 15802
rect 3835 15750 3865 15802
rect 3865 15750 3877 15802
rect 3877 15750 3891 15802
rect 3915 15750 3929 15802
rect 3929 15750 3941 15802
rect 3941 15750 3971 15802
rect 3995 15750 4005 15802
rect 4005 15750 4051 15802
rect 3755 15748 3811 15750
rect 3835 15748 3891 15750
rect 3915 15748 3971 15750
rect 3995 15748 4051 15750
rect 3755 14714 3811 14716
rect 3835 14714 3891 14716
rect 3915 14714 3971 14716
rect 3995 14714 4051 14716
rect 3755 14662 3801 14714
rect 3801 14662 3811 14714
rect 3835 14662 3865 14714
rect 3865 14662 3877 14714
rect 3877 14662 3891 14714
rect 3915 14662 3929 14714
rect 3929 14662 3941 14714
rect 3941 14662 3971 14714
rect 3995 14662 4005 14714
rect 4005 14662 4051 14714
rect 3755 14660 3811 14662
rect 3835 14660 3891 14662
rect 3915 14660 3971 14662
rect 3995 14660 4051 14662
rect 4434 13812 4436 13832
rect 4436 13812 4488 13832
rect 4488 13812 4490 13832
rect 4434 13776 4490 13812
rect 3755 13626 3811 13628
rect 3835 13626 3891 13628
rect 3915 13626 3971 13628
rect 3995 13626 4051 13628
rect 3755 13574 3801 13626
rect 3801 13574 3811 13626
rect 3835 13574 3865 13626
rect 3865 13574 3877 13626
rect 3877 13574 3891 13626
rect 3915 13574 3929 13626
rect 3929 13574 3941 13626
rect 3941 13574 3971 13626
rect 3995 13574 4005 13626
rect 4005 13574 4051 13626
rect 3755 13572 3811 13574
rect 3835 13572 3891 13574
rect 3915 13572 3971 13574
rect 3995 13572 4051 13574
rect 3755 12538 3811 12540
rect 3835 12538 3891 12540
rect 3915 12538 3971 12540
rect 3995 12538 4051 12540
rect 3755 12486 3801 12538
rect 3801 12486 3811 12538
rect 3835 12486 3865 12538
rect 3865 12486 3877 12538
rect 3877 12486 3891 12538
rect 3915 12486 3929 12538
rect 3929 12486 3941 12538
rect 3941 12486 3971 12538
rect 3995 12486 4005 12538
rect 4005 12486 4051 12538
rect 3755 12484 3811 12486
rect 3835 12484 3891 12486
rect 3915 12484 3971 12486
rect 3995 12484 4051 12486
rect 3755 11450 3811 11452
rect 3835 11450 3891 11452
rect 3915 11450 3971 11452
rect 3995 11450 4051 11452
rect 3755 11398 3801 11450
rect 3801 11398 3811 11450
rect 3835 11398 3865 11450
rect 3865 11398 3877 11450
rect 3877 11398 3891 11450
rect 3915 11398 3929 11450
rect 3929 11398 3941 11450
rect 3941 11398 3971 11450
rect 3995 11398 4005 11450
rect 4005 11398 4051 11450
rect 3755 11396 3811 11398
rect 3835 11396 3891 11398
rect 3915 11396 3971 11398
rect 3995 11396 4051 11398
rect 6554 21786 6610 21788
rect 6634 21786 6690 21788
rect 6714 21786 6770 21788
rect 6794 21786 6850 21788
rect 6554 21734 6600 21786
rect 6600 21734 6610 21786
rect 6634 21734 6664 21786
rect 6664 21734 6676 21786
rect 6676 21734 6690 21786
rect 6714 21734 6728 21786
rect 6728 21734 6740 21786
rect 6740 21734 6770 21786
rect 6794 21734 6804 21786
rect 6804 21734 6850 21786
rect 6554 21732 6610 21734
rect 6634 21732 6690 21734
rect 6714 21732 6770 21734
rect 6794 21732 6850 21734
rect 6554 20698 6610 20700
rect 6634 20698 6690 20700
rect 6714 20698 6770 20700
rect 6794 20698 6850 20700
rect 6554 20646 6600 20698
rect 6600 20646 6610 20698
rect 6634 20646 6664 20698
rect 6664 20646 6676 20698
rect 6676 20646 6690 20698
rect 6714 20646 6728 20698
rect 6728 20646 6740 20698
rect 6740 20646 6770 20698
rect 6794 20646 6804 20698
rect 6804 20646 6850 20698
rect 6554 20644 6610 20646
rect 6634 20644 6690 20646
rect 6714 20644 6770 20646
rect 6794 20644 6850 20646
rect 6554 19610 6610 19612
rect 6634 19610 6690 19612
rect 6714 19610 6770 19612
rect 6794 19610 6850 19612
rect 6554 19558 6600 19610
rect 6600 19558 6610 19610
rect 6634 19558 6664 19610
rect 6664 19558 6676 19610
rect 6676 19558 6690 19610
rect 6714 19558 6728 19610
rect 6728 19558 6740 19610
rect 6740 19558 6770 19610
rect 6794 19558 6804 19610
rect 6804 19558 6850 19610
rect 6554 19556 6610 19558
rect 6634 19556 6690 19558
rect 6714 19556 6770 19558
rect 6794 19556 6850 19558
rect 7102 21800 7158 21856
rect 8390 21664 8446 21720
rect 7378 21292 7380 21312
rect 7380 21292 7432 21312
rect 7432 21292 7434 21312
rect 7378 21256 7434 21292
rect 8390 20984 8446 21040
rect 6554 18522 6610 18524
rect 6634 18522 6690 18524
rect 6714 18522 6770 18524
rect 6794 18522 6850 18524
rect 6554 18470 6600 18522
rect 6600 18470 6610 18522
rect 6634 18470 6664 18522
rect 6664 18470 6676 18522
rect 6676 18470 6690 18522
rect 6714 18470 6728 18522
rect 6728 18470 6740 18522
rect 6740 18470 6770 18522
rect 6794 18470 6804 18522
rect 6804 18470 6850 18522
rect 6554 18468 6610 18470
rect 6634 18468 6690 18470
rect 6714 18468 6770 18470
rect 6794 18468 6850 18470
rect 6090 16360 6146 16416
rect 5630 13932 5686 13968
rect 5630 13912 5632 13932
rect 5632 13912 5684 13932
rect 5684 13912 5686 13932
rect 6274 16396 6276 16416
rect 6276 16396 6328 16416
rect 6328 16396 6330 16416
rect 6274 16360 6330 16396
rect 6554 17434 6610 17436
rect 6634 17434 6690 17436
rect 6714 17434 6770 17436
rect 6794 17434 6850 17436
rect 6554 17382 6600 17434
rect 6600 17382 6610 17434
rect 6634 17382 6664 17434
rect 6664 17382 6676 17434
rect 6676 17382 6690 17434
rect 6714 17382 6728 17434
rect 6728 17382 6740 17434
rect 6740 17382 6770 17434
rect 6794 17382 6804 17434
rect 6804 17382 6850 17434
rect 6554 17380 6610 17382
rect 6634 17380 6690 17382
rect 6714 17380 6770 17382
rect 6794 17380 6850 17382
rect 9353 22330 9409 22332
rect 9433 22330 9489 22332
rect 9513 22330 9569 22332
rect 9593 22330 9649 22332
rect 9353 22278 9399 22330
rect 9399 22278 9409 22330
rect 9433 22278 9463 22330
rect 9463 22278 9475 22330
rect 9475 22278 9489 22330
rect 9513 22278 9527 22330
rect 9527 22278 9539 22330
rect 9539 22278 9569 22330
rect 9593 22278 9603 22330
rect 9603 22278 9649 22330
rect 9353 22276 9409 22278
rect 9433 22276 9489 22278
rect 9513 22276 9569 22278
rect 9593 22276 9649 22278
rect 10046 21836 10048 21856
rect 10048 21836 10100 21856
rect 10100 21836 10102 21856
rect 9218 21664 9274 21720
rect 9353 21242 9409 21244
rect 9433 21242 9489 21244
rect 9513 21242 9569 21244
rect 9593 21242 9649 21244
rect 9353 21190 9399 21242
rect 9399 21190 9409 21242
rect 9433 21190 9463 21242
rect 9463 21190 9475 21242
rect 9475 21190 9489 21242
rect 9513 21190 9527 21242
rect 9527 21190 9539 21242
rect 9539 21190 9569 21242
rect 9593 21190 9603 21242
rect 9603 21190 9649 21242
rect 9353 21188 9409 21190
rect 9433 21188 9489 21190
rect 9513 21188 9569 21190
rect 9593 21188 9649 21190
rect 9353 20154 9409 20156
rect 9433 20154 9489 20156
rect 9513 20154 9569 20156
rect 9593 20154 9649 20156
rect 9353 20102 9399 20154
rect 9399 20102 9409 20154
rect 9433 20102 9463 20154
rect 9463 20102 9475 20154
rect 9475 20102 9489 20154
rect 9513 20102 9527 20154
rect 9527 20102 9539 20154
rect 9539 20102 9569 20154
rect 9593 20102 9603 20154
rect 9603 20102 9649 20154
rect 9353 20100 9409 20102
rect 9433 20100 9489 20102
rect 9513 20100 9569 20102
rect 9593 20100 9649 20102
rect 9494 19780 9550 19816
rect 9494 19760 9496 19780
rect 9496 19760 9548 19780
rect 9548 19760 9550 19780
rect 9494 19352 9550 19408
rect 10046 21800 10102 21836
rect 10782 21664 10838 21720
rect 10874 21528 10930 21584
rect 9353 19066 9409 19068
rect 9433 19066 9489 19068
rect 9513 19066 9569 19068
rect 9593 19066 9649 19068
rect 9353 19014 9399 19066
rect 9399 19014 9409 19066
rect 9433 19014 9463 19066
rect 9463 19014 9475 19066
rect 9475 19014 9489 19066
rect 9513 19014 9527 19066
rect 9527 19014 9539 19066
rect 9539 19014 9569 19066
rect 9593 19014 9603 19066
rect 9603 19014 9649 19066
rect 9353 19012 9409 19014
rect 9433 19012 9489 19014
rect 9513 19012 9569 19014
rect 9593 19012 9649 19014
rect 9353 17978 9409 17980
rect 9433 17978 9489 17980
rect 9513 17978 9569 17980
rect 9593 17978 9649 17980
rect 9353 17926 9399 17978
rect 9399 17926 9409 17978
rect 9433 17926 9463 17978
rect 9463 17926 9475 17978
rect 9475 17926 9489 17978
rect 9513 17926 9527 17978
rect 9527 17926 9539 17978
rect 9539 17926 9569 17978
rect 9593 17926 9603 17978
rect 9603 17926 9649 17978
rect 9353 17924 9409 17926
rect 9433 17924 9489 17926
rect 9513 17924 9569 17926
rect 9593 17924 9649 17926
rect 11242 21936 11298 21992
rect 11150 20848 11206 20904
rect 11242 20712 11298 20768
rect 11150 20440 11206 20496
rect 11426 19780 11482 19816
rect 11426 19760 11428 19780
rect 11428 19760 11480 19780
rect 11480 19760 11482 19780
rect 12152 21786 12208 21788
rect 12232 21786 12288 21788
rect 12312 21786 12368 21788
rect 12392 21786 12448 21788
rect 12152 21734 12198 21786
rect 12198 21734 12208 21786
rect 12232 21734 12262 21786
rect 12262 21734 12274 21786
rect 12274 21734 12288 21786
rect 12312 21734 12326 21786
rect 12326 21734 12338 21786
rect 12338 21734 12368 21786
rect 12392 21734 12402 21786
rect 12402 21734 12448 21786
rect 12152 21732 12208 21734
rect 12232 21732 12288 21734
rect 12312 21732 12368 21734
rect 12392 21732 12448 21734
rect 11978 19932 11980 19952
rect 11980 19932 12032 19952
rect 12032 19932 12034 19952
rect 11978 19896 12034 19932
rect 11794 19488 11850 19544
rect 9353 16890 9409 16892
rect 9433 16890 9489 16892
rect 9513 16890 9569 16892
rect 9593 16890 9649 16892
rect 9353 16838 9399 16890
rect 9399 16838 9409 16890
rect 9433 16838 9463 16890
rect 9463 16838 9475 16890
rect 9475 16838 9489 16890
rect 9513 16838 9527 16890
rect 9527 16838 9539 16890
rect 9539 16838 9569 16890
rect 9593 16838 9603 16890
rect 9603 16838 9649 16890
rect 9353 16836 9409 16838
rect 9433 16836 9489 16838
rect 9513 16836 9569 16838
rect 9593 16836 9649 16838
rect 6554 16346 6610 16348
rect 6634 16346 6690 16348
rect 6714 16346 6770 16348
rect 6794 16346 6850 16348
rect 6554 16294 6600 16346
rect 6600 16294 6610 16346
rect 6634 16294 6664 16346
rect 6664 16294 6676 16346
rect 6676 16294 6690 16346
rect 6714 16294 6728 16346
rect 6728 16294 6740 16346
rect 6740 16294 6770 16346
rect 6794 16294 6804 16346
rect 6804 16294 6850 16346
rect 6554 16292 6610 16294
rect 6634 16292 6690 16294
rect 6714 16292 6770 16294
rect 6794 16292 6850 16294
rect 9353 15802 9409 15804
rect 9433 15802 9489 15804
rect 9513 15802 9569 15804
rect 9593 15802 9649 15804
rect 9353 15750 9399 15802
rect 9399 15750 9409 15802
rect 9433 15750 9463 15802
rect 9463 15750 9475 15802
rect 9475 15750 9489 15802
rect 9513 15750 9527 15802
rect 9527 15750 9539 15802
rect 9539 15750 9569 15802
rect 9593 15750 9603 15802
rect 9603 15750 9649 15802
rect 9353 15748 9409 15750
rect 9433 15748 9489 15750
rect 9513 15748 9569 15750
rect 9593 15748 9649 15750
rect 8666 15408 8722 15464
rect 6554 15258 6610 15260
rect 6634 15258 6690 15260
rect 6714 15258 6770 15260
rect 6794 15258 6850 15260
rect 6554 15206 6600 15258
rect 6600 15206 6610 15258
rect 6634 15206 6664 15258
rect 6664 15206 6676 15258
rect 6676 15206 6690 15258
rect 6714 15206 6728 15258
rect 6728 15206 6740 15258
rect 6740 15206 6770 15258
rect 6794 15206 6804 15258
rect 6804 15206 6850 15258
rect 6554 15204 6610 15206
rect 6634 15204 6690 15206
rect 6714 15204 6770 15206
rect 6794 15204 6850 15206
rect 9353 14714 9409 14716
rect 9433 14714 9489 14716
rect 9513 14714 9569 14716
rect 9593 14714 9649 14716
rect 9353 14662 9399 14714
rect 9399 14662 9409 14714
rect 9433 14662 9463 14714
rect 9463 14662 9475 14714
rect 9475 14662 9489 14714
rect 9513 14662 9527 14714
rect 9527 14662 9539 14714
rect 9539 14662 9569 14714
rect 9593 14662 9603 14714
rect 9603 14662 9649 14714
rect 9353 14660 9409 14662
rect 9433 14660 9489 14662
rect 9513 14660 9569 14662
rect 9593 14660 9649 14662
rect 6554 14170 6610 14172
rect 6634 14170 6690 14172
rect 6714 14170 6770 14172
rect 6794 14170 6850 14172
rect 6554 14118 6600 14170
rect 6600 14118 6610 14170
rect 6634 14118 6664 14170
rect 6664 14118 6676 14170
rect 6676 14118 6690 14170
rect 6714 14118 6728 14170
rect 6728 14118 6740 14170
rect 6740 14118 6770 14170
rect 6794 14118 6804 14170
rect 6804 14118 6850 14170
rect 6554 14116 6610 14118
rect 6634 14116 6690 14118
rect 6714 14116 6770 14118
rect 6794 14116 6850 14118
rect 6550 13948 6552 13968
rect 6552 13948 6604 13968
rect 6604 13948 6606 13968
rect 6550 13912 6606 13948
rect 8390 13776 8446 13832
rect 6554 13082 6610 13084
rect 6634 13082 6690 13084
rect 6714 13082 6770 13084
rect 6794 13082 6850 13084
rect 6554 13030 6600 13082
rect 6600 13030 6610 13082
rect 6634 13030 6664 13082
rect 6664 13030 6676 13082
rect 6676 13030 6690 13082
rect 6714 13030 6728 13082
rect 6728 13030 6740 13082
rect 6740 13030 6770 13082
rect 6794 13030 6804 13082
rect 6804 13030 6850 13082
rect 6554 13028 6610 13030
rect 6634 13028 6690 13030
rect 6714 13028 6770 13030
rect 6794 13028 6850 13030
rect 9353 13626 9409 13628
rect 9433 13626 9489 13628
rect 9513 13626 9569 13628
rect 9593 13626 9649 13628
rect 9353 13574 9399 13626
rect 9399 13574 9409 13626
rect 9433 13574 9463 13626
rect 9463 13574 9475 13626
rect 9475 13574 9489 13626
rect 9513 13574 9527 13626
rect 9527 13574 9539 13626
rect 9539 13574 9569 13626
rect 9593 13574 9603 13626
rect 9603 13574 9649 13626
rect 9353 13572 9409 13574
rect 9433 13572 9489 13574
rect 9513 13572 9569 13574
rect 9593 13572 9649 13574
rect 3755 10362 3811 10364
rect 3835 10362 3891 10364
rect 3915 10362 3971 10364
rect 3995 10362 4051 10364
rect 3755 10310 3801 10362
rect 3801 10310 3811 10362
rect 3835 10310 3865 10362
rect 3865 10310 3877 10362
rect 3877 10310 3891 10362
rect 3915 10310 3929 10362
rect 3929 10310 3941 10362
rect 3941 10310 3971 10362
rect 3995 10310 4005 10362
rect 4005 10310 4051 10362
rect 3755 10308 3811 10310
rect 3835 10308 3891 10310
rect 3915 10308 3971 10310
rect 3995 10308 4051 10310
rect 3755 9274 3811 9276
rect 3835 9274 3891 9276
rect 3915 9274 3971 9276
rect 3995 9274 4051 9276
rect 3755 9222 3801 9274
rect 3801 9222 3811 9274
rect 3835 9222 3865 9274
rect 3865 9222 3877 9274
rect 3877 9222 3891 9274
rect 3915 9222 3929 9274
rect 3929 9222 3941 9274
rect 3941 9222 3971 9274
rect 3995 9222 4005 9274
rect 4005 9222 4051 9274
rect 3755 9220 3811 9222
rect 3835 9220 3891 9222
rect 3915 9220 3971 9222
rect 3995 9220 4051 9222
rect 2962 8508 2964 8528
rect 2964 8508 3016 8528
rect 3016 8508 3018 8528
rect 2962 8472 3018 8508
rect 6554 11994 6610 11996
rect 6634 11994 6690 11996
rect 6714 11994 6770 11996
rect 6794 11994 6850 11996
rect 6554 11942 6600 11994
rect 6600 11942 6610 11994
rect 6634 11942 6664 11994
rect 6664 11942 6676 11994
rect 6676 11942 6690 11994
rect 6714 11942 6728 11994
rect 6728 11942 6740 11994
rect 6740 11942 6770 11994
rect 6794 11942 6804 11994
rect 6804 11942 6850 11994
rect 6554 11940 6610 11942
rect 6634 11940 6690 11942
rect 6714 11940 6770 11942
rect 6794 11940 6850 11942
rect 6554 10906 6610 10908
rect 6634 10906 6690 10908
rect 6714 10906 6770 10908
rect 6794 10906 6850 10908
rect 6554 10854 6600 10906
rect 6600 10854 6610 10906
rect 6634 10854 6664 10906
rect 6664 10854 6676 10906
rect 6676 10854 6690 10906
rect 6714 10854 6728 10906
rect 6728 10854 6740 10906
rect 6740 10854 6770 10906
rect 6794 10854 6804 10906
rect 6804 10854 6850 10906
rect 6554 10852 6610 10854
rect 6634 10852 6690 10854
rect 6714 10852 6770 10854
rect 6794 10852 6850 10854
rect 9353 12538 9409 12540
rect 9433 12538 9489 12540
rect 9513 12538 9569 12540
rect 9593 12538 9649 12540
rect 9353 12486 9399 12538
rect 9399 12486 9409 12538
rect 9433 12486 9463 12538
rect 9463 12486 9475 12538
rect 9475 12486 9489 12538
rect 9513 12486 9527 12538
rect 9527 12486 9539 12538
rect 9539 12486 9569 12538
rect 9593 12486 9603 12538
rect 9603 12486 9649 12538
rect 9353 12484 9409 12486
rect 9433 12484 9489 12486
rect 9513 12484 9569 12486
rect 9593 12484 9649 12486
rect 9353 11450 9409 11452
rect 9433 11450 9489 11452
rect 9513 11450 9569 11452
rect 9593 11450 9649 11452
rect 9353 11398 9399 11450
rect 9399 11398 9409 11450
rect 9433 11398 9463 11450
rect 9463 11398 9475 11450
rect 9475 11398 9489 11450
rect 9513 11398 9527 11450
rect 9527 11398 9539 11450
rect 9539 11398 9569 11450
rect 9593 11398 9603 11450
rect 9603 11398 9649 11450
rect 9353 11396 9409 11398
rect 9433 11396 9489 11398
rect 9513 11396 9569 11398
rect 9593 11396 9649 11398
rect 6554 9818 6610 9820
rect 6634 9818 6690 9820
rect 6714 9818 6770 9820
rect 6794 9818 6850 9820
rect 6554 9766 6600 9818
rect 6600 9766 6610 9818
rect 6634 9766 6664 9818
rect 6664 9766 6676 9818
rect 6676 9766 6690 9818
rect 6714 9766 6728 9818
rect 6728 9766 6740 9818
rect 6740 9766 6770 9818
rect 6794 9766 6804 9818
rect 6804 9766 6850 9818
rect 6554 9764 6610 9766
rect 6634 9764 6690 9766
rect 6714 9764 6770 9766
rect 6794 9764 6850 9766
rect 3755 8186 3811 8188
rect 3835 8186 3891 8188
rect 3915 8186 3971 8188
rect 3995 8186 4051 8188
rect 3755 8134 3801 8186
rect 3801 8134 3811 8186
rect 3835 8134 3865 8186
rect 3865 8134 3877 8186
rect 3877 8134 3891 8186
rect 3915 8134 3929 8186
rect 3929 8134 3941 8186
rect 3941 8134 3971 8186
rect 3995 8134 4005 8186
rect 4005 8134 4051 8186
rect 3755 8132 3811 8134
rect 3835 8132 3891 8134
rect 3915 8132 3971 8134
rect 3995 8132 4051 8134
rect 4894 8492 4950 8528
rect 4894 8472 4896 8492
rect 4896 8472 4948 8492
rect 4948 8472 4950 8492
rect 3755 7098 3811 7100
rect 3835 7098 3891 7100
rect 3915 7098 3971 7100
rect 3995 7098 4051 7100
rect 3755 7046 3801 7098
rect 3801 7046 3811 7098
rect 3835 7046 3865 7098
rect 3865 7046 3877 7098
rect 3877 7046 3891 7098
rect 3915 7046 3929 7098
rect 3929 7046 3941 7098
rect 3941 7046 3971 7098
rect 3995 7046 4005 7098
rect 4005 7046 4051 7098
rect 3755 7044 3811 7046
rect 3835 7044 3891 7046
rect 3915 7044 3971 7046
rect 3995 7044 4051 7046
rect 6554 8730 6610 8732
rect 6634 8730 6690 8732
rect 6714 8730 6770 8732
rect 6794 8730 6850 8732
rect 6554 8678 6600 8730
rect 6600 8678 6610 8730
rect 6634 8678 6664 8730
rect 6664 8678 6676 8730
rect 6676 8678 6690 8730
rect 6714 8678 6728 8730
rect 6728 8678 6740 8730
rect 6740 8678 6770 8730
rect 6794 8678 6804 8730
rect 6804 8678 6850 8730
rect 6554 8676 6610 8678
rect 6634 8676 6690 8678
rect 6714 8676 6770 8678
rect 6794 8676 6850 8678
rect 9353 10362 9409 10364
rect 9433 10362 9489 10364
rect 9513 10362 9569 10364
rect 9593 10362 9649 10364
rect 9353 10310 9399 10362
rect 9399 10310 9409 10362
rect 9433 10310 9463 10362
rect 9463 10310 9475 10362
rect 9475 10310 9489 10362
rect 9513 10310 9527 10362
rect 9527 10310 9539 10362
rect 9539 10310 9569 10362
rect 9593 10310 9603 10362
rect 9603 10310 9649 10362
rect 9353 10308 9409 10310
rect 9433 10308 9489 10310
rect 9513 10308 9569 10310
rect 9593 10308 9649 10310
rect 6554 7642 6610 7644
rect 6634 7642 6690 7644
rect 6714 7642 6770 7644
rect 6794 7642 6850 7644
rect 6554 7590 6600 7642
rect 6600 7590 6610 7642
rect 6634 7590 6664 7642
rect 6664 7590 6676 7642
rect 6676 7590 6690 7642
rect 6714 7590 6728 7642
rect 6728 7590 6740 7642
rect 6740 7590 6770 7642
rect 6794 7590 6804 7642
rect 6804 7590 6850 7642
rect 6554 7588 6610 7590
rect 6634 7588 6690 7590
rect 6714 7588 6770 7590
rect 6794 7588 6850 7590
rect 6554 6554 6610 6556
rect 6634 6554 6690 6556
rect 6714 6554 6770 6556
rect 6794 6554 6850 6556
rect 6554 6502 6600 6554
rect 6600 6502 6610 6554
rect 6634 6502 6664 6554
rect 6664 6502 6676 6554
rect 6676 6502 6690 6554
rect 6714 6502 6728 6554
rect 6728 6502 6740 6554
rect 6740 6502 6770 6554
rect 6794 6502 6804 6554
rect 6804 6502 6850 6554
rect 6554 6500 6610 6502
rect 6634 6500 6690 6502
rect 6714 6500 6770 6502
rect 6794 6500 6850 6502
rect 3755 6010 3811 6012
rect 3835 6010 3891 6012
rect 3915 6010 3971 6012
rect 3995 6010 4051 6012
rect 3755 5958 3801 6010
rect 3801 5958 3811 6010
rect 3835 5958 3865 6010
rect 3865 5958 3877 6010
rect 3877 5958 3891 6010
rect 3915 5958 3929 6010
rect 3929 5958 3941 6010
rect 3941 5958 3971 6010
rect 3995 5958 4005 6010
rect 4005 5958 4051 6010
rect 3755 5956 3811 5958
rect 3835 5956 3891 5958
rect 3915 5956 3971 5958
rect 3995 5956 4051 5958
rect 6554 5466 6610 5468
rect 6634 5466 6690 5468
rect 6714 5466 6770 5468
rect 6794 5466 6850 5468
rect 6554 5414 6600 5466
rect 6600 5414 6610 5466
rect 6634 5414 6664 5466
rect 6664 5414 6676 5466
rect 6676 5414 6690 5466
rect 6714 5414 6728 5466
rect 6728 5414 6740 5466
rect 6740 5414 6770 5466
rect 6794 5414 6804 5466
rect 6804 5414 6850 5466
rect 6554 5412 6610 5414
rect 6634 5412 6690 5414
rect 6714 5412 6770 5414
rect 6794 5412 6850 5414
rect 3755 4922 3811 4924
rect 3835 4922 3891 4924
rect 3915 4922 3971 4924
rect 3995 4922 4051 4924
rect 3755 4870 3801 4922
rect 3801 4870 3811 4922
rect 3835 4870 3865 4922
rect 3865 4870 3877 4922
rect 3877 4870 3891 4922
rect 3915 4870 3929 4922
rect 3929 4870 3941 4922
rect 3941 4870 3971 4922
rect 3995 4870 4005 4922
rect 4005 4870 4051 4922
rect 3755 4868 3811 4870
rect 3835 4868 3891 4870
rect 3915 4868 3971 4870
rect 3995 4868 4051 4870
rect 9353 9274 9409 9276
rect 9433 9274 9489 9276
rect 9513 9274 9569 9276
rect 9593 9274 9649 9276
rect 9353 9222 9399 9274
rect 9399 9222 9409 9274
rect 9433 9222 9463 9274
rect 9463 9222 9475 9274
rect 9475 9222 9489 9274
rect 9513 9222 9527 9274
rect 9527 9222 9539 9274
rect 9539 9222 9569 9274
rect 9593 9222 9603 9274
rect 9603 9222 9649 9274
rect 9353 9220 9409 9222
rect 9433 9220 9489 9222
rect 9513 9220 9569 9222
rect 9593 9220 9649 9222
rect 9353 8186 9409 8188
rect 9433 8186 9489 8188
rect 9513 8186 9569 8188
rect 9593 8186 9649 8188
rect 9353 8134 9399 8186
rect 9399 8134 9409 8186
rect 9433 8134 9463 8186
rect 9463 8134 9475 8186
rect 9475 8134 9489 8186
rect 9513 8134 9527 8186
rect 9527 8134 9539 8186
rect 9539 8134 9569 8186
rect 9593 8134 9603 8186
rect 9603 8134 9649 8186
rect 9353 8132 9409 8134
rect 9433 8132 9489 8134
rect 9513 8132 9569 8134
rect 9593 8132 9649 8134
rect 9353 7098 9409 7100
rect 9433 7098 9489 7100
rect 9513 7098 9569 7100
rect 9593 7098 9649 7100
rect 9353 7046 9399 7098
rect 9399 7046 9409 7098
rect 9433 7046 9463 7098
rect 9463 7046 9475 7098
rect 9475 7046 9489 7098
rect 9513 7046 9527 7098
rect 9527 7046 9539 7098
rect 9539 7046 9569 7098
rect 9593 7046 9603 7098
rect 9603 7046 9649 7098
rect 9353 7044 9409 7046
rect 9433 7044 9489 7046
rect 9513 7044 9569 7046
rect 9593 7044 9649 7046
rect 9353 6010 9409 6012
rect 9433 6010 9489 6012
rect 9513 6010 9569 6012
rect 9593 6010 9649 6012
rect 9353 5958 9399 6010
rect 9399 5958 9409 6010
rect 9433 5958 9463 6010
rect 9463 5958 9475 6010
rect 9475 5958 9489 6010
rect 9513 5958 9527 6010
rect 9527 5958 9539 6010
rect 9539 5958 9569 6010
rect 9593 5958 9603 6010
rect 9603 5958 9649 6010
rect 9353 5956 9409 5958
rect 9433 5956 9489 5958
rect 9513 5956 9569 5958
rect 9593 5956 9649 5958
rect 9353 4922 9409 4924
rect 9433 4922 9489 4924
rect 9513 4922 9569 4924
rect 9593 4922 9649 4924
rect 9353 4870 9399 4922
rect 9399 4870 9409 4922
rect 9433 4870 9463 4922
rect 9463 4870 9475 4922
rect 9475 4870 9489 4922
rect 9513 4870 9527 4922
rect 9527 4870 9539 4922
rect 9539 4870 9569 4922
rect 9593 4870 9603 4922
rect 9603 4870 9649 4922
rect 9353 4868 9409 4870
rect 9433 4868 9489 4870
rect 9513 4868 9569 4870
rect 9593 4868 9649 4870
rect 12152 20698 12208 20700
rect 12232 20698 12288 20700
rect 12312 20698 12368 20700
rect 12392 20698 12448 20700
rect 12152 20646 12198 20698
rect 12198 20646 12208 20698
rect 12232 20646 12262 20698
rect 12262 20646 12274 20698
rect 12274 20646 12288 20698
rect 12312 20646 12326 20698
rect 12326 20646 12338 20698
rect 12338 20646 12368 20698
rect 12392 20646 12402 20698
rect 12402 20646 12448 20698
rect 12152 20644 12208 20646
rect 12232 20644 12288 20646
rect 12312 20644 12368 20646
rect 12392 20644 12448 20646
rect 12162 20440 12218 20496
rect 12152 19610 12208 19612
rect 12232 19610 12288 19612
rect 12312 19610 12368 19612
rect 12392 19610 12448 19612
rect 12152 19558 12198 19610
rect 12198 19558 12208 19610
rect 12232 19558 12262 19610
rect 12262 19558 12274 19610
rect 12274 19558 12288 19610
rect 12312 19558 12326 19610
rect 12326 19558 12338 19610
rect 12338 19558 12368 19610
rect 12392 19558 12402 19610
rect 12402 19558 12448 19610
rect 12152 19556 12208 19558
rect 12232 19556 12288 19558
rect 12312 19556 12368 19558
rect 12392 19556 12448 19558
rect 12152 18522 12208 18524
rect 12232 18522 12288 18524
rect 12312 18522 12368 18524
rect 12392 18522 12448 18524
rect 12152 18470 12198 18522
rect 12198 18470 12208 18522
rect 12232 18470 12262 18522
rect 12262 18470 12274 18522
rect 12274 18470 12288 18522
rect 12312 18470 12326 18522
rect 12326 18470 12338 18522
rect 12338 18470 12368 18522
rect 12392 18470 12402 18522
rect 12402 18470 12448 18522
rect 12152 18468 12208 18470
rect 12232 18468 12288 18470
rect 12312 18468 12368 18470
rect 12392 18468 12448 18470
rect 12622 20304 12678 20360
rect 12152 17434 12208 17436
rect 12232 17434 12288 17436
rect 12312 17434 12368 17436
rect 12392 17434 12448 17436
rect 12152 17382 12198 17434
rect 12198 17382 12208 17434
rect 12232 17382 12262 17434
rect 12262 17382 12274 17434
rect 12274 17382 12288 17434
rect 12312 17382 12326 17434
rect 12326 17382 12338 17434
rect 12338 17382 12368 17434
rect 12392 17382 12402 17434
rect 12402 17382 12448 17434
rect 12152 17380 12208 17382
rect 12232 17380 12288 17382
rect 12312 17380 12368 17382
rect 12392 17380 12448 17382
rect 12152 16346 12208 16348
rect 12232 16346 12288 16348
rect 12312 16346 12368 16348
rect 12392 16346 12448 16348
rect 12152 16294 12198 16346
rect 12198 16294 12208 16346
rect 12232 16294 12262 16346
rect 12262 16294 12274 16346
rect 12274 16294 12288 16346
rect 12312 16294 12326 16346
rect 12326 16294 12338 16346
rect 12338 16294 12368 16346
rect 12392 16294 12402 16346
rect 12402 16294 12448 16346
rect 12152 16292 12208 16294
rect 12232 16292 12288 16294
rect 12312 16292 12368 16294
rect 12392 16292 12448 16294
rect 12152 15258 12208 15260
rect 12232 15258 12288 15260
rect 12312 15258 12368 15260
rect 12392 15258 12448 15260
rect 12152 15206 12198 15258
rect 12198 15206 12208 15258
rect 12232 15206 12262 15258
rect 12262 15206 12274 15258
rect 12274 15206 12288 15258
rect 12312 15206 12326 15258
rect 12326 15206 12338 15258
rect 12338 15206 12368 15258
rect 12392 15206 12402 15258
rect 12402 15206 12448 15258
rect 12152 15204 12208 15206
rect 12232 15204 12288 15206
rect 12312 15204 12368 15206
rect 12392 15204 12448 15206
rect 12152 14170 12208 14172
rect 12232 14170 12288 14172
rect 12312 14170 12368 14172
rect 12392 14170 12448 14172
rect 12152 14118 12198 14170
rect 12198 14118 12208 14170
rect 12232 14118 12262 14170
rect 12262 14118 12274 14170
rect 12274 14118 12288 14170
rect 12312 14118 12326 14170
rect 12326 14118 12338 14170
rect 12338 14118 12368 14170
rect 12392 14118 12402 14170
rect 12402 14118 12448 14170
rect 12152 14116 12208 14118
rect 12232 14116 12288 14118
rect 12312 14116 12368 14118
rect 12392 14116 12448 14118
rect 12152 13082 12208 13084
rect 12232 13082 12288 13084
rect 12312 13082 12368 13084
rect 12392 13082 12448 13084
rect 12152 13030 12198 13082
rect 12198 13030 12208 13082
rect 12232 13030 12262 13082
rect 12262 13030 12274 13082
rect 12274 13030 12288 13082
rect 12312 13030 12326 13082
rect 12326 13030 12338 13082
rect 12338 13030 12368 13082
rect 12392 13030 12402 13082
rect 12402 13030 12448 13082
rect 12152 13028 12208 13030
rect 12232 13028 12288 13030
rect 12312 13028 12368 13030
rect 12392 13028 12448 13030
rect 12152 11994 12208 11996
rect 12232 11994 12288 11996
rect 12312 11994 12368 11996
rect 12392 11994 12448 11996
rect 12152 11942 12198 11994
rect 12198 11942 12208 11994
rect 12232 11942 12262 11994
rect 12262 11942 12274 11994
rect 12274 11942 12288 11994
rect 12312 11942 12326 11994
rect 12326 11942 12338 11994
rect 12338 11942 12368 11994
rect 12392 11942 12402 11994
rect 12402 11942 12448 11994
rect 12152 11940 12208 11942
rect 12232 11940 12288 11942
rect 12312 11940 12368 11942
rect 12392 11940 12448 11942
rect 13726 21800 13782 21856
rect 12990 18808 13046 18864
rect 13726 19932 13728 19952
rect 13728 19932 13780 19952
rect 13780 19932 13782 19952
rect 13726 19896 13782 19932
rect 13450 18808 13506 18864
rect 13358 18672 13414 18728
rect 13910 17876 13966 17912
rect 13910 17856 13912 17876
rect 13912 17856 13964 17876
rect 13964 17856 13966 17876
rect 14951 22330 15007 22332
rect 15031 22330 15087 22332
rect 15111 22330 15167 22332
rect 15191 22330 15247 22332
rect 14951 22278 14997 22330
rect 14997 22278 15007 22330
rect 15031 22278 15061 22330
rect 15061 22278 15073 22330
rect 15073 22278 15087 22330
rect 15111 22278 15125 22330
rect 15125 22278 15137 22330
rect 15137 22278 15167 22330
rect 15191 22278 15201 22330
rect 15201 22278 15247 22330
rect 14951 22276 15007 22278
rect 15031 22276 15087 22278
rect 15111 22276 15167 22278
rect 15191 22276 15247 22278
rect 14646 21392 14702 21448
rect 15014 21664 15070 21720
rect 14951 21242 15007 21244
rect 15031 21242 15087 21244
rect 15111 21242 15167 21244
rect 15191 21242 15247 21244
rect 14951 21190 14997 21242
rect 14997 21190 15007 21242
rect 15031 21190 15061 21242
rect 15061 21190 15073 21242
rect 15073 21190 15087 21242
rect 15111 21190 15125 21242
rect 15125 21190 15137 21242
rect 15137 21190 15167 21242
rect 15191 21190 15201 21242
rect 15201 21190 15247 21242
rect 14951 21188 15007 21190
rect 15031 21188 15087 21190
rect 15111 21188 15167 21190
rect 15191 21188 15247 21190
rect 14738 20984 14794 21040
rect 14646 20712 14702 20768
rect 15658 21684 15714 21720
rect 15658 21664 15660 21684
rect 15660 21664 15712 21684
rect 15712 21664 15714 21684
rect 15474 21256 15530 21312
rect 15658 21120 15714 21176
rect 15934 21800 15990 21856
rect 15658 20712 15714 20768
rect 12152 10906 12208 10908
rect 12232 10906 12288 10908
rect 12312 10906 12368 10908
rect 12392 10906 12448 10908
rect 12152 10854 12198 10906
rect 12198 10854 12208 10906
rect 12232 10854 12262 10906
rect 12262 10854 12274 10906
rect 12274 10854 12288 10906
rect 12312 10854 12326 10906
rect 12326 10854 12338 10906
rect 12338 10854 12368 10906
rect 12392 10854 12402 10906
rect 12402 10854 12448 10906
rect 12152 10852 12208 10854
rect 12232 10852 12288 10854
rect 12312 10852 12368 10854
rect 12392 10852 12448 10854
rect 12152 9818 12208 9820
rect 12232 9818 12288 9820
rect 12312 9818 12368 9820
rect 12392 9818 12448 9820
rect 12152 9766 12198 9818
rect 12198 9766 12208 9818
rect 12232 9766 12262 9818
rect 12262 9766 12274 9818
rect 12274 9766 12288 9818
rect 12312 9766 12326 9818
rect 12326 9766 12338 9818
rect 12338 9766 12368 9818
rect 12392 9766 12402 9818
rect 12402 9766 12448 9818
rect 12152 9764 12208 9766
rect 12232 9764 12288 9766
rect 12312 9764 12368 9766
rect 12392 9764 12448 9766
rect 14094 13404 14096 13424
rect 14096 13404 14148 13424
rect 14148 13404 14150 13424
rect 14094 13368 14150 13404
rect 12152 8730 12208 8732
rect 12232 8730 12288 8732
rect 12312 8730 12368 8732
rect 12392 8730 12448 8732
rect 12152 8678 12198 8730
rect 12198 8678 12208 8730
rect 12232 8678 12262 8730
rect 12262 8678 12274 8730
rect 12274 8678 12288 8730
rect 12312 8678 12326 8730
rect 12326 8678 12338 8730
rect 12338 8678 12368 8730
rect 12392 8678 12402 8730
rect 12402 8678 12448 8730
rect 12152 8676 12208 8678
rect 12232 8676 12288 8678
rect 12312 8676 12368 8678
rect 12392 8676 12448 8678
rect 12152 7642 12208 7644
rect 12232 7642 12288 7644
rect 12312 7642 12368 7644
rect 12392 7642 12448 7644
rect 12152 7590 12198 7642
rect 12198 7590 12208 7642
rect 12232 7590 12262 7642
rect 12262 7590 12274 7642
rect 12274 7590 12288 7642
rect 12312 7590 12326 7642
rect 12326 7590 12338 7642
rect 12338 7590 12368 7642
rect 12392 7590 12402 7642
rect 12402 7590 12448 7642
rect 12152 7588 12208 7590
rect 12232 7588 12288 7590
rect 12312 7588 12368 7590
rect 12392 7588 12448 7590
rect 6554 4378 6610 4380
rect 6634 4378 6690 4380
rect 6714 4378 6770 4380
rect 6794 4378 6850 4380
rect 6554 4326 6600 4378
rect 6600 4326 6610 4378
rect 6634 4326 6664 4378
rect 6664 4326 6676 4378
rect 6676 4326 6690 4378
rect 6714 4326 6728 4378
rect 6728 4326 6740 4378
rect 6740 4326 6770 4378
rect 6794 4326 6804 4378
rect 6804 4326 6850 4378
rect 6554 4324 6610 4326
rect 6634 4324 6690 4326
rect 6714 4324 6770 4326
rect 6794 4324 6850 4326
rect 3755 3834 3811 3836
rect 3835 3834 3891 3836
rect 3915 3834 3971 3836
rect 3995 3834 4051 3836
rect 3755 3782 3801 3834
rect 3801 3782 3811 3834
rect 3835 3782 3865 3834
rect 3865 3782 3877 3834
rect 3877 3782 3891 3834
rect 3915 3782 3929 3834
rect 3929 3782 3941 3834
rect 3941 3782 3971 3834
rect 3995 3782 4005 3834
rect 4005 3782 4051 3834
rect 3755 3780 3811 3782
rect 3835 3780 3891 3782
rect 3915 3780 3971 3782
rect 3995 3780 4051 3782
rect 9353 3834 9409 3836
rect 9433 3834 9489 3836
rect 9513 3834 9569 3836
rect 9593 3834 9649 3836
rect 9353 3782 9399 3834
rect 9399 3782 9409 3834
rect 9433 3782 9463 3834
rect 9463 3782 9475 3834
rect 9475 3782 9489 3834
rect 9513 3782 9527 3834
rect 9527 3782 9539 3834
rect 9539 3782 9569 3834
rect 9593 3782 9603 3834
rect 9603 3782 9649 3834
rect 9353 3780 9409 3782
rect 9433 3780 9489 3782
rect 9513 3780 9569 3782
rect 9593 3780 9649 3782
rect 6554 3290 6610 3292
rect 6634 3290 6690 3292
rect 6714 3290 6770 3292
rect 6794 3290 6850 3292
rect 6554 3238 6600 3290
rect 6600 3238 6610 3290
rect 6634 3238 6664 3290
rect 6664 3238 6676 3290
rect 6676 3238 6690 3290
rect 6714 3238 6728 3290
rect 6728 3238 6740 3290
rect 6740 3238 6770 3290
rect 6794 3238 6804 3290
rect 6804 3238 6850 3290
rect 6554 3236 6610 3238
rect 6634 3236 6690 3238
rect 6714 3236 6770 3238
rect 6794 3236 6850 3238
rect 1398 3032 1454 3088
rect 12152 6554 12208 6556
rect 12232 6554 12288 6556
rect 12312 6554 12368 6556
rect 12392 6554 12448 6556
rect 12152 6502 12198 6554
rect 12198 6502 12208 6554
rect 12232 6502 12262 6554
rect 12262 6502 12274 6554
rect 12274 6502 12288 6554
rect 12312 6502 12326 6554
rect 12326 6502 12338 6554
rect 12338 6502 12368 6554
rect 12392 6502 12402 6554
rect 12402 6502 12448 6554
rect 12152 6500 12208 6502
rect 12232 6500 12288 6502
rect 12312 6500 12368 6502
rect 12392 6500 12448 6502
rect 12152 5466 12208 5468
rect 12232 5466 12288 5468
rect 12312 5466 12368 5468
rect 12392 5466 12448 5468
rect 12152 5414 12198 5466
rect 12198 5414 12208 5466
rect 12232 5414 12262 5466
rect 12262 5414 12274 5466
rect 12274 5414 12288 5466
rect 12312 5414 12326 5466
rect 12326 5414 12338 5466
rect 12338 5414 12368 5466
rect 12392 5414 12402 5466
rect 12402 5414 12448 5466
rect 12152 5412 12208 5414
rect 12232 5412 12288 5414
rect 12312 5412 12368 5414
rect 12392 5412 12448 5414
rect 14951 20154 15007 20156
rect 15031 20154 15087 20156
rect 15111 20154 15167 20156
rect 15191 20154 15247 20156
rect 14951 20102 14997 20154
rect 14997 20102 15007 20154
rect 15031 20102 15061 20154
rect 15061 20102 15073 20154
rect 15073 20102 15087 20154
rect 15111 20102 15125 20154
rect 15125 20102 15137 20154
rect 15137 20102 15167 20154
rect 15191 20102 15201 20154
rect 15201 20102 15247 20154
rect 14951 20100 15007 20102
rect 15031 20100 15087 20102
rect 15111 20100 15167 20102
rect 15191 20100 15247 20102
rect 14951 19066 15007 19068
rect 15031 19066 15087 19068
rect 15111 19066 15167 19068
rect 15191 19066 15247 19068
rect 14951 19014 14997 19066
rect 14997 19014 15007 19066
rect 15031 19014 15061 19066
rect 15061 19014 15073 19066
rect 15073 19014 15087 19066
rect 15111 19014 15125 19066
rect 15125 19014 15137 19066
rect 15137 19014 15167 19066
rect 15191 19014 15201 19066
rect 15201 19014 15247 19066
rect 14951 19012 15007 19014
rect 15031 19012 15087 19014
rect 15111 19012 15167 19014
rect 15191 19012 15247 19014
rect 14951 17978 15007 17980
rect 15031 17978 15087 17980
rect 15111 17978 15167 17980
rect 15191 17978 15247 17980
rect 14951 17926 14997 17978
rect 14997 17926 15007 17978
rect 15031 17926 15061 17978
rect 15061 17926 15073 17978
rect 15073 17926 15087 17978
rect 15111 17926 15125 17978
rect 15125 17926 15137 17978
rect 15137 17926 15167 17978
rect 15191 17926 15201 17978
rect 15201 17926 15247 17978
rect 14951 17924 15007 17926
rect 15031 17924 15087 17926
rect 15111 17924 15167 17926
rect 15191 17924 15247 17926
rect 14951 16890 15007 16892
rect 15031 16890 15087 16892
rect 15111 16890 15167 16892
rect 15191 16890 15247 16892
rect 14951 16838 14997 16890
rect 14997 16838 15007 16890
rect 15031 16838 15061 16890
rect 15061 16838 15073 16890
rect 15073 16838 15087 16890
rect 15111 16838 15125 16890
rect 15125 16838 15137 16890
rect 15137 16838 15167 16890
rect 15191 16838 15201 16890
rect 15201 16838 15247 16890
rect 14951 16836 15007 16838
rect 15031 16836 15087 16838
rect 15111 16836 15167 16838
rect 15191 16836 15247 16838
rect 15658 19352 15714 19408
rect 16302 21664 16358 21720
rect 14951 15802 15007 15804
rect 15031 15802 15087 15804
rect 15111 15802 15167 15804
rect 15191 15802 15247 15804
rect 14951 15750 14997 15802
rect 14997 15750 15007 15802
rect 15031 15750 15061 15802
rect 15061 15750 15073 15802
rect 15073 15750 15087 15802
rect 15111 15750 15125 15802
rect 15125 15750 15137 15802
rect 15137 15750 15167 15802
rect 15191 15750 15201 15802
rect 15201 15750 15247 15802
rect 14951 15748 15007 15750
rect 15031 15748 15087 15750
rect 15111 15748 15167 15750
rect 15191 15748 15247 15750
rect 16486 21664 16542 21720
rect 16762 21256 16818 21312
rect 16486 21120 16542 21176
rect 16394 20304 16450 20360
rect 17222 21800 17278 21856
rect 17222 21256 17278 21312
rect 17130 21120 17186 21176
rect 17038 20440 17094 20496
rect 17406 22072 17462 22128
rect 17750 21786 17806 21788
rect 17830 21786 17886 21788
rect 17910 21786 17966 21788
rect 17990 21786 18046 21788
rect 17750 21734 17796 21786
rect 17796 21734 17806 21786
rect 17830 21734 17860 21786
rect 17860 21734 17872 21786
rect 17872 21734 17886 21786
rect 17910 21734 17924 21786
rect 17924 21734 17936 21786
rect 17936 21734 17966 21786
rect 17990 21734 18000 21786
rect 18000 21734 18046 21786
rect 17750 21732 17806 21734
rect 17830 21732 17886 21734
rect 17910 21732 17966 21734
rect 17990 21732 18046 21734
rect 17866 21292 17868 21312
rect 17868 21292 17920 21312
rect 17920 21292 17922 21312
rect 17866 21256 17922 21292
rect 18418 21120 18474 21176
rect 18142 20984 18198 21040
rect 17750 20698 17806 20700
rect 17830 20698 17886 20700
rect 17910 20698 17966 20700
rect 17990 20698 18046 20700
rect 17750 20646 17796 20698
rect 17796 20646 17806 20698
rect 17830 20646 17860 20698
rect 17860 20646 17872 20698
rect 17872 20646 17886 20698
rect 17910 20646 17924 20698
rect 17924 20646 17936 20698
rect 17936 20646 17966 20698
rect 17990 20646 18000 20698
rect 18000 20646 18046 20698
rect 17750 20644 17806 20646
rect 17830 20644 17886 20646
rect 17910 20644 17966 20646
rect 17990 20644 18046 20646
rect 18050 19896 18106 19952
rect 17314 17584 17370 17640
rect 16578 14900 16580 14920
rect 16580 14900 16632 14920
rect 16632 14900 16634 14920
rect 16578 14864 16634 14900
rect 14951 14714 15007 14716
rect 15031 14714 15087 14716
rect 15111 14714 15167 14716
rect 15191 14714 15247 14716
rect 14951 14662 14997 14714
rect 14997 14662 15007 14714
rect 15031 14662 15061 14714
rect 15061 14662 15073 14714
rect 15073 14662 15087 14714
rect 15111 14662 15125 14714
rect 15125 14662 15137 14714
rect 15137 14662 15167 14714
rect 15191 14662 15201 14714
rect 15201 14662 15247 14714
rect 14951 14660 15007 14662
rect 15031 14660 15087 14662
rect 15111 14660 15167 14662
rect 15191 14660 15247 14662
rect 14738 14340 14794 14376
rect 14738 14320 14740 14340
rect 14740 14320 14792 14340
rect 14792 14320 14794 14340
rect 14951 13626 15007 13628
rect 15031 13626 15087 13628
rect 15111 13626 15167 13628
rect 15191 13626 15247 13628
rect 14951 13574 14997 13626
rect 14997 13574 15007 13626
rect 15031 13574 15061 13626
rect 15061 13574 15073 13626
rect 15073 13574 15087 13626
rect 15111 13574 15125 13626
rect 15125 13574 15137 13626
rect 15137 13574 15167 13626
rect 15191 13574 15201 13626
rect 15201 13574 15247 13626
rect 14951 13572 15007 13574
rect 15031 13572 15087 13574
rect 15111 13572 15167 13574
rect 15191 13572 15247 13574
rect 14951 12538 15007 12540
rect 15031 12538 15087 12540
rect 15111 12538 15167 12540
rect 15191 12538 15247 12540
rect 14951 12486 14997 12538
rect 14997 12486 15007 12538
rect 15031 12486 15061 12538
rect 15061 12486 15073 12538
rect 15073 12486 15087 12538
rect 15111 12486 15125 12538
rect 15125 12486 15137 12538
rect 15137 12486 15167 12538
rect 15191 12486 15201 12538
rect 15201 12486 15247 12538
rect 14951 12484 15007 12486
rect 15031 12484 15087 12486
rect 15111 12484 15167 12486
rect 15191 12484 15247 12486
rect 16578 13232 16634 13288
rect 14462 7384 14518 7440
rect 14370 6180 14426 6216
rect 14370 6160 14372 6180
rect 14372 6160 14424 6180
rect 14424 6160 14426 6180
rect 18602 22072 18658 22128
rect 18510 20440 18566 20496
rect 17750 19610 17806 19612
rect 17830 19610 17886 19612
rect 17910 19610 17966 19612
rect 17990 19610 18046 19612
rect 17750 19558 17796 19610
rect 17796 19558 17806 19610
rect 17830 19558 17860 19610
rect 17860 19558 17872 19610
rect 17872 19558 17886 19610
rect 17910 19558 17924 19610
rect 17924 19558 17936 19610
rect 17936 19558 17966 19610
rect 17990 19558 18000 19610
rect 18000 19558 18046 19610
rect 17750 19556 17806 19558
rect 17830 19556 17886 19558
rect 17910 19556 17966 19558
rect 17990 19556 18046 19558
rect 18602 19760 18658 19816
rect 20549 22330 20605 22332
rect 20629 22330 20685 22332
rect 20709 22330 20765 22332
rect 20789 22330 20845 22332
rect 20549 22278 20595 22330
rect 20595 22278 20605 22330
rect 20629 22278 20659 22330
rect 20659 22278 20671 22330
rect 20671 22278 20685 22330
rect 20709 22278 20723 22330
rect 20723 22278 20735 22330
rect 20735 22278 20765 22330
rect 20789 22278 20799 22330
rect 20799 22278 20845 22330
rect 20549 22276 20605 22278
rect 20629 22276 20685 22278
rect 20709 22276 20765 22278
rect 20789 22276 20845 22278
rect 20534 22072 20590 22128
rect 17750 18522 17806 18524
rect 17830 18522 17886 18524
rect 17910 18522 17966 18524
rect 17990 18522 18046 18524
rect 17750 18470 17796 18522
rect 17796 18470 17806 18522
rect 17830 18470 17860 18522
rect 17860 18470 17872 18522
rect 17872 18470 17886 18522
rect 17910 18470 17924 18522
rect 17924 18470 17936 18522
rect 17936 18470 17966 18522
rect 17990 18470 18000 18522
rect 18000 18470 18046 18522
rect 17750 18468 17806 18470
rect 17830 18468 17886 18470
rect 17910 18468 17966 18470
rect 17990 18468 18046 18470
rect 18878 19216 18934 19272
rect 18602 18536 18658 18592
rect 17750 17434 17806 17436
rect 17830 17434 17886 17436
rect 17910 17434 17966 17436
rect 17990 17434 18046 17436
rect 17750 17382 17796 17434
rect 17796 17382 17806 17434
rect 17830 17382 17860 17434
rect 17860 17382 17872 17434
rect 17872 17382 17886 17434
rect 17910 17382 17924 17434
rect 17924 17382 17936 17434
rect 17936 17382 17966 17434
rect 17990 17382 18000 17434
rect 18000 17382 18046 17434
rect 17750 17380 17806 17382
rect 17830 17380 17886 17382
rect 17910 17380 17966 17382
rect 17990 17380 18046 17382
rect 18510 17448 18566 17504
rect 17750 16346 17806 16348
rect 17830 16346 17886 16348
rect 17910 16346 17966 16348
rect 17990 16346 18046 16348
rect 17750 16294 17796 16346
rect 17796 16294 17806 16346
rect 17830 16294 17860 16346
rect 17860 16294 17872 16346
rect 17872 16294 17886 16346
rect 17910 16294 17924 16346
rect 17924 16294 17936 16346
rect 17936 16294 17966 16346
rect 17990 16294 18000 16346
rect 18000 16294 18046 16346
rect 17750 16292 17806 16294
rect 17830 16292 17886 16294
rect 17910 16292 17966 16294
rect 17990 16292 18046 16294
rect 18510 16632 18566 16688
rect 18878 18128 18934 18184
rect 17750 15258 17806 15260
rect 17830 15258 17886 15260
rect 17910 15258 17966 15260
rect 17990 15258 18046 15260
rect 17750 15206 17796 15258
rect 17796 15206 17806 15258
rect 17830 15206 17860 15258
rect 17860 15206 17872 15258
rect 17872 15206 17886 15258
rect 17910 15206 17924 15258
rect 17924 15206 17936 15258
rect 17936 15206 17966 15258
rect 17990 15206 18000 15258
rect 18000 15206 18046 15258
rect 17750 15204 17806 15206
rect 17830 15204 17886 15206
rect 17910 15204 17966 15206
rect 17990 15204 18046 15206
rect 17750 14170 17806 14172
rect 17830 14170 17886 14172
rect 17910 14170 17966 14172
rect 17990 14170 18046 14172
rect 17750 14118 17796 14170
rect 17796 14118 17806 14170
rect 17830 14118 17860 14170
rect 17860 14118 17872 14170
rect 17872 14118 17886 14170
rect 17910 14118 17924 14170
rect 17924 14118 17936 14170
rect 17936 14118 17966 14170
rect 17990 14118 18000 14170
rect 18000 14118 18046 14170
rect 17750 14116 17806 14118
rect 17830 14116 17886 14118
rect 17910 14116 17966 14118
rect 17990 14116 18046 14118
rect 17750 13082 17806 13084
rect 17830 13082 17886 13084
rect 17910 13082 17966 13084
rect 17990 13082 18046 13084
rect 17750 13030 17796 13082
rect 17796 13030 17806 13082
rect 17830 13030 17860 13082
rect 17860 13030 17872 13082
rect 17872 13030 17886 13082
rect 17910 13030 17924 13082
rect 17924 13030 17936 13082
rect 17936 13030 17966 13082
rect 17990 13030 18000 13082
rect 18000 13030 18046 13082
rect 17750 13028 17806 13030
rect 17830 13028 17886 13030
rect 17910 13028 17966 13030
rect 17990 13028 18046 13030
rect 14951 11450 15007 11452
rect 15031 11450 15087 11452
rect 15111 11450 15167 11452
rect 15191 11450 15247 11452
rect 14951 11398 14997 11450
rect 14997 11398 15007 11450
rect 15031 11398 15061 11450
rect 15061 11398 15073 11450
rect 15073 11398 15087 11450
rect 15111 11398 15125 11450
rect 15125 11398 15137 11450
rect 15137 11398 15167 11450
rect 15191 11398 15201 11450
rect 15201 11398 15247 11450
rect 14951 11396 15007 11398
rect 15031 11396 15087 11398
rect 15111 11396 15167 11398
rect 15191 11396 15247 11398
rect 14951 10362 15007 10364
rect 15031 10362 15087 10364
rect 15111 10362 15167 10364
rect 15191 10362 15247 10364
rect 14951 10310 14997 10362
rect 14997 10310 15007 10362
rect 15031 10310 15061 10362
rect 15061 10310 15073 10362
rect 15073 10310 15087 10362
rect 15111 10310 15125 10362
rect 15125 10310 15137 10362
rect 15137 10310 15167 10362
rect 15191 10310 15201 10362
rect 15201 10310 15247 10362
rect 14951 10308 15007 10310
rect 15031 10308 15087 10310
rect 15111 10308 15167 10310
rect 15191 10308 15247 10310
rect 14951 9274 15007 9276
rect 15031 9274 15087 9276
rect 15111 9274 15167 9276
rect 15191 9274 15247 9276
rect 14951 9222 14997 9274
rect 14997 9222 15007 9274
rect 15031 9222 15061 9274
rect 15061 9222 15073 9274
rect 15073 9222 15087 9274
rect 15111 9222 15125 9274
rect 15125 9222 15137 9274
rect 15137 9222 15167 9274
rect 15191 9222 15201 9274
rect 15201 9222 15247 9274
rect 14951 9220 15007 9222
rect 15031 9220 15087 9222
rect 15111 9220 15167 9222
rect 15191 9220 15247 9222
rect 14951 8186 15007 8188
rect 15031 8186 15087 8188
rect 15111 8186 15167 8188
rect 15191 8186 15247 8188
rect 14951 8134 14997 8186
rect 14997 8134 15007 8186
rect 15031 8134 15061 8186
rect 15061 8134 15073 8186
rect 15073 8134 15087 8186
rect 15111 8134 15125 8186
rect 15125 8134 15137 8186
rect 15137 8134 15167 8186
rect 15191 8134 15201 8186
rect 15201 8134 15247 8186
rect 14951 8132 15007 8134
rect 15031 8132 15087 8134
rect 15111 8132 15167 8134
rect 15191 8132 15247 8134
rect 14951 7098 15007 7100
rect 15031 7098 15087 7100
rect 15111 7098 15167 7100
rect 15191 7098 15247 7100
rect 14951 7046 14997 7098
rect 14997 7046 15007 7098
rect 15031 7046 15061 7098
rect 15061 7046 15073 7098
rect 15073 7046 15087 7098
rect 15111 7046 15125 7098
rect 15125 7046 15137 7098
rect 15137 7046 15167 7098
rect 15191 7046 15201 7098
rect 15201 7046 15247 7098
rect 14951 7044 15007 7046
rect 15031 7044 15087 7046
rect 15111 7044 15167 7046
rect 15191 7044 15247 7046
rect 16578 10104 16634 10160
rect 14951 6010 15007 6012
rect 15031 6010 15087 6012
rect 15111 6010 15167 6012
rect 15191 6010 15247 6012
rect 14951 5958 14997 6010
rect 14997 5958 15007 6010
rect 15031 5958 15061 6010
rect 15061 5958 15073 6010
rect 15073 5958 15087 6010
rect 15111 5958 15125 6010
rect 15125 5958 15137 6010
rect 15137 5958 15167 6010
rect 15191 5958 15201 6010
rect 15201 5958 15247 6010
rect 14951 5956 15007 5958
rect 15031 5956 15087 5958
rect 15111 5956 15167 5958
rect 15191 5956 15247 5958
rect 12152 4378 12208 4380
rect 12232 4378 12288 4380
rect 12312 4378 12368 4380
rect 12392 4378 12448 4380
rect 12152 4326 12198 4378
rect 12198 4326 12208 4378
rect 12232 4326 12262 4378
rect 12262 4326 12274 4378
rect 12274 4326 12288 4378
rect 12312 4326 12326 4378
rect 12326 4326 12338 4378
rect 12338 4326 12368 4378
rect 12392 4326 12402 4378
rect 12402 4326 12448 4378
rect 12152 4324 12208 4326
rect 12232 4324 12288 4326
rect 12312 4324 12368 4326
rect 12392 4324 12448 4326
rect 13726 4120 13782 4176
rect 14951 4922 15007 4924
rect 15031 4922 15087 4924
rect 15111 4922 15167 4924
rect 15191 4922 15247 4924
rect 14951 4870 14997 4922
rect 14997 4870 15007 4922
rect 15031 4870 15061 4922
rect 15061 4870 15073 4922
rect 15073 4870 15087 4922
rect 15111 4870 15125 4922
rect 15125 4870 15137 4922
rect 15137 4870 15167 4922
rect 15191 4870 15201 4922
rect 15201 4870 15247 4922
rect 14951 4868 15007 4870
rect 15031 4868 15087 4870
rect 15111 4868 15167 4870
rect 15191 4868 15247 4870
rect 14951 3834 15007 3836
rect 15031 3834 15087 3836
rect 15111 3834 15167 3836
rect 15191 3834 15247 3836
rect 14951 3782 14997 3834
rect 14997 3782 15007 3834
rect 15031 3782 15061 3834
rect 15061 3782 15073 3834
rect 15073 3782 15087 3834
rect 15111 3782 15125 3834
rect 15125 3782 15137 3834
rect 15137 3782 15167 3834
rect 15191 3782 15201 3834
rect 15201 3782 15247 3834
rect 14951 3780 15007 3782
rect 15031 3780 15087 3782
rect 15111 3780 15167 3782
rect 15191 3780 15247 3782
rect 15566 3576 15622 3632
rect 16486 8336 16542 8392
rect 16394 6296 16450 6352
rect 16946 7248 17002 7304
rect 17222 6704 17278 6760
rect 17130 6296 17186 6352
rect 17038 6160 17094 6216
rect 12152 3290 12208 3292
rect 12232 3290 12288 3292
rect 12312 3290 12368 3292
rect 12392 3290 12448 3292
rect 12152 3238 12198 3290
rect 12198 3238 12208 3290
rect 12232 3238 12262 3290
rect 12262 3238 12274 3290
rect 12274 3238 12288 3290
rect 12312 3238 12326 3290
rect 12326 3238 12338 3290
rect 12338 3238 12368 3290
rect 12392 3238 12402 3290
rect 12402 3238 12448 3290
rect 12152 3236 12208 3238
rect 12232 3236 12288 3238
rect 12312 3236 12368 3238
rect 12392 3236 12448 3238
rect 3755 2746 3811 2748
rect 3835 2746 3891 2748
rect 3915 2746 3971 2748
rect 3995 2746 4051 2748
rect 3755 2694 3801 2746
rect 3801 2694 3811 2746
rect 3835 2694 3865 2746
rect 3865 2694 3877 2746
rect 3877 2694 3891 2746
rect 3915 2694 3929 2746
rect 3929 2694 3941 2746
rect 3941 2694 3971 2746
rect 3995 2694 4005 2746
rect 4005 2694 4051 2746
rect 3755 2692 3811 2694
rect 3835 2692 3891 2694
rect 3915 2692 3971 2694
rect 3995 2692 4051 2694
rect 9353 2746 9409 2748
rect 9433 2746 9489 2748
rect 9513 2746 9569 2748
rect 9593 2746 9649 2748
rect 9353 2694 9399 2746
rect 9399 2694 9409 2746
rect 9433 2694 9463 2746
rect 9463 2694 9475 2746
rect 9475 2694 9489 2746
rect 9513 2694 9527 2746
rect 9527 2694 9539 2746
rect 9539 2694 9569 2746
rect 9593 2694 9603 2746
rect 9603 2694 9649 2746
rect 9353 2692 9409 2694
rect 9433 2692 9489 2694
rect 9513 2692 9569 2694
rect 9593 2692 9649 2694
rect 14951 2746 15007 2748
rect 15031 2746 15087 2748
rect 15111 2746 15167 2748
rect 15191 2746 15247 2748
rect 14951 2694 14997 2746
rect 14997 2694 15007 2746
rect 15031 2694 15061 2746
rect 15061 2694 15073 2746
rect 15073 2694 15087 2746
rect 15111 2694 15125 2746
rect 15125 2694 15137 2746
rect 15137 2694 15167 2746
rect 15191 2694 15201 2746
rect 15201 2694 15247 2746
rect 14951 2692 15007 2694
rect 15031 2692 15087 2694
rect 15111 2692 15167 2694
rect 15191 2692 15247 2694
rect 16302 3440 16358 3496
rect 18878 15544 18934 15600
rect 18234 12144 18290 12200
rect 18510 12688 18566 12744
rect 17750 11994 17806 11996
rect 17830 11994 17886 11996
rect 17910 11994 17966 11996
rect 17990 11994 18046 11996
rect 17750 11942 17796 11994
rect 17796 11942 17806 11994
rect 17830 11942 17860 11994
rect 17860 11942 17872 11994
rect 17872 11942 17886 11994
rect 17910 11942 17924 11994
rect 17924 11942 17936 11994
rect 17936 11942 17966 11994
rect 17990 11942 18000 11994
rect 18000 11942 18046 11994
rect 17750 11940 17806 11942
rect 17830 11940 17886 11942
rect 17910 11940 17966 11942
rect 17990 11940 18046 11942
rect 18878 12280 18934 12336
rect 18786 11600 18842 11656
rect 17750 10906 17806 10908
rect 17830 10906 17886 10908
rect 17910 10906 17966 10908
rect 17990 10906 18046 10908
rect 17750 10854 17796 10906
rect 17796 10854 17806 10906
rect 17830 10854 17860 10906
rect 17860 10854 17872 10906
rect 17872 10854 17886 10906
rect 17910 10854 17924 10906
rect 17924 10854 17936 10906
rect 17936 10854 17966 10906
rect 17990 10854 18000 10906
rect 18000 10854 18046 10906
rect 17750 10852 17806 10854
rect 17830 10852 17886 10854
rect 17910 10852 17966 10854
rect 17990 10852 18046 10854
rect 18050 9968 18106 10024
rect 17750 9818 17806 9820
rect 17830 9818 17886 9820
rect 17910 9818 17966 9820
rect 17990 9818 18046 9820
rect 17750 9766 17796 9818
rect 17796 9766 17806 9818
rect 17830 9766 17860 9818
rect 17860 9766 17872 9818
rect 17872 9766 17886 9818
rect 17910 9766 17924 9818
rect 17924 9766 17936 9818
rect 17936 9766 17966 9818
rect 17990 9766 18000 9818
rect 18000 9766 18046 9818
rect 17750 9764 17806 9766
rect 17830 9764 17886 9766
rect 17910 9764 17966 9766
rect 17990 9764 18046 9766
rect 18050 8880 18106 8936
rect 17750 8730 17806 8732
rect 17830 8730 17886 8732
rect 17910 8730 17966 8732
rect 17990 8730 18046 8732
rect 17750 8678 17796 8730
rect 17796 8678 17806 8730
rect 17830 8678 17860 8730
rect 17860 8678 17872 8730
rect 17872 8678 17886 8730
rect 17910 8678 17924 8730
rect 17924 8678 17936 8730
rect 17936 8678 17966 8730
rect 17990 8678 18000 8730
rect 18000 8678 18046 8730
rect 17750 8676 17806 8678
rect 17830 8676 17886 8678
rect 17910 8676 17966 8678
rect 17990 8676 18046 8678
rect 18418 9968 18474 10024
rect 18418 9832 18474 9888
rect 17750 7642 17806 7644
rect 17830 7642 17886 7644
rect 17910 7642 17966 7644
rect 17990 7642 18046 7644
rect 17750 7590 17796 7642
rect 17796 7590 17806 7642
rect 17830 7590 17860 7642
rect 17860 7590 17872 7642
rect 17872 7590 17886 7642
rect 17910 7590 17924 7642
rect 17924 7590 17936 7642
rect 17936 7590 17966 7642
rect 17990 7590 18000 7642
rect 18000 7590 18046 7642
rect 17750 7588 17806 7590
rect 17830 7588 17886 7590
rect 17910 7588 17966 7590
rect 17990 7588 18046 7590
rect 17750 6554 17806 6556
rect 17830 6554 17886 6556
rect 17910 6554 17966 6556
rect 17990 6554 18046 6556
rect 17750 6502 17796 6554
rect 17796 6502 17806 6554
rect 17830 6502 17860 6554
rect 17860 6502 17872 6554
rect 17872 6502 17886 6554
rect 17910 6502 17924 6554
rect 17924 6502 17936 6554
rect 17936 6502 17966 6554
rect 17990 6502 18000 6554
rect 18000 6502 18046 6554
rect 17750 6500 17806 6502
rect 17830 6500 17886 6502
rect 17910 6500 17966 6502
rect 17990 6500 18046 6502
rect 17750 5466 17806 5468
rect 17830 5466 17886 5468
rect 17910 5466 17966 5468
rect 17990 5466 18046 5468
rect 17750 5414 17796 5466
rect 17796 5414 17806 5466
rect 17830 5414 17860 5466
rect 17860 5414 17872 5466
rect 17872 5414 17886 5466
rect 17910 5414 17924 5466
rect 17924 5414 17936 5466
rect 17936 5414 17966 5466
rect 17990 5414 18000 5466
rect 18000 5414 18046 5466
rect 17750 5412 17806 5414
rect 17830 5412 17886 5414
rect 17910 5412 17966 5414
rect 17990 5412 18046 5414
rect 16670 3032 16726 3088
rect 19062 17756 19064 17776
rect 19064 17756 19116 17776
rect 19116 17756 19118 17776
rect 19062 17720 19118 17756
rect 19982 19352 20038 19408
rect 19154 15952 19210 16008
rect 19154 15544 19210 15600
rect 19430 16088 19486 16144
rect 19706 18128 19762 18184
rect 19062 12824 19118 12880
rect 18970 9968 19026 10024
rect 18878 9832 18934 9888
rect 18786 9696 18842 9752
rect 19338 13096 19394 13152
rect 20074 18808 20130 18864
rect 20994 21392 21050 21448
rect 20549 21242 20605 21244
rect 20629 21242 20685 21244
rect 20709 21242 20765 21244
rect 20789 21242 20845 21244
rect 20549 21190 20595 21242
rect 20595 21190 20605 21242
rect 20629 21190 20659 21242
rect 20659 21190 20671 21242
rect 20671 21190 20685 21242
rect 20709 21190 20723 21242
rect 20723 21190 20735 21242
rect 20735 21190 20765 21242
rect 20789 21190 20799 21242
rect 20799 21190 20845 21242
rect 20549 21188 20605 21190
rect 20629 21188 20685 21190
rect 20709 21188 20765 21190
rect 20789 21188 20845 21190
rect 20810 20984 20866 21040
rect 20549 20154 20605 20156
rect 20629 20154 20685 20156
rect 20709 20154 20765 20156
rect 20789 20154 20845 20156
rect 20549 20102 20595 20154
rect 20595 20102 20605 20154
rect 20629 20102 20659 20154
rect 20659 20102 20671 20154
rect 20671 20102 20685 20154
rect 20709 20102 20723 20154
rect 20723 20102 20735 20154
rect 20735 20102 20765 20154
rect 20789 20102 20799 20154
rect 20799 20102 20845 20154
rect 20549 20100 20605 20102
rect 20629 20100 20685 20102
rect 20709 20100 20765 20102
rect 20789 20100 20845 20102
rect 20902 19796 20904 19816
rect 20904 19796 20956 19816
rect 20956 19796 20958 19816
rect 20902 19760 20958 19796
rect 21822 21972 21824 21992
rect 21824 21972 21876 21992
rect 21876 21972 21878 21992
rect 21822 21936 21878 21972
rect 21362 20848 21418 20904
rect 22466 21528 22522 21584
rect 22650 21528 22706 21584
rect 23018 20984 23074 21040
rect 22190 20712 22246 20768
rect 23018 20440 23074 20496
rect 20549 19066 20605 19068
rect 20629 19066 20685 19068
rect 20709 19066 20765 19068
rect 20789 19066 20845 19068
rect 20549 19014 20595 19066
rect 20595 19014 20605 19066
rect 20629 19014 20659 19066
rect 20659 19014 20671 19066
rect 20671 19014 20685 19066
rect 20709 19014 20723 19066
rect 20723 19014 20735 19066
rect 20735 19014 20765 19066
rect 20789 19014 20799 19066
rect 20799 19014 20845 19066
rect 20549 19012 20605 19014
rect 20629 19012 20685 19014
rect 20709 19012 20765 19014
rect 20789 19012 20845 19014
rect 20810 18844 20812 18864
rect 20812 18844 20864 18864
rect 20864 18844 20866 18864
rect 20810 18808 20866 18844
rect 20549 17978 20605 17980
rect 20629 17978 20685 17980
rect 20709 17978 20765 17980
rect 20789 17978 20845 17980
rect 20549 17926 20595 17978
rect 20595 17926 20605 17978
rect 20629 17926 20659 17978
rect 20659 17926 20671 17978
rect 20671 17926 20685 17978
rect 20709 17926 20723 17978
rect 20723 17926 20735 17978
rect 20735 17926 20765 17978
rect 20789 17926 20799 17978
rect 20799 17926 20845 17978
rect 20549 17924 20605 17926
rect 20629 17924 20685 17926
rect 20709 17924 20765 17926
rect 20789 17924 20845 17926
rect 20902 17448 20958 17504
rect 20549 16890 20605 16892
rect 20629 16890 20685 16892
rect 20709 16890 20765 16892
rect 20789 16890 20845 16892
rect 20549 16838 20595 16890
rect 20595 16838 20605 16890
rect 20629 16838 20659 16890
rect 20659 16838 20671 16890
rect 20671 16838 20685 16890
rect 20709 16838 20723 16890
rect 20723 16838 20735 16890
rect 20735 16838 20765 16890
rect 20789 16838 20799 16890
rect 20799 16838 20845 16890
rect 20549 16836 20605 16838
rect 20629 16836 20685 16838
rect 20709 16836 20765 16838
rect 20789 16836 20845 16838
rect 20549 15802 20605 15804
rect 20629 15802 20685 15804
rect 20709 15802 20765 15804
rect 20789 15802 20845 15804
rect 20549 15750 20595 15802
rect 20595 15750 20605 15802
rect 20629 15750 20659 15802
rect 20659 15750 20671 15802
rect 20671 15750 20685 15802
rect 20709 15750 20723 15802
rect 20723 15750 20735 15802
rect 20735 15750 20765 15802
rect 20789 15750 20799 15802
rect 20799 15750 20845 15802
rect 20549 15748 20605 15750
rect 20629 15748 20685 15750
rect 20709 15748 20765 15750
rect 20789 15748 20845 15750
rect 20549 14714 20605 14716
rect 20629 14714 20685 14716
rect 20709 14714 20765 14716
rect 20789 14714 20845 14716
rect 20549 14662 20595 14714
rect 20595 14662 20605 14714
rect 20629 14662 20659 14714
rect 20659 14662 20671 14714
rect 20671 14662 20685 14714
rect 20709 14662 20723 14714
rect 20723 14662 20735 14714
rect 20735 14662 20765 14714
rect 20789 14662 20799 14714
rect 20799 14662 20845 14714
rect 20549 14660 20605 14662
rect 20629 14660 20685 14662
rect 20709 14660 20765 14662
rect 20789 14660 20845 14662
rect 21086 14864 21142 14920
rect 20994 14320 21050 14376
rect 20549 13626 20605 13628
rect 20629 13626 20685 13628
rect 20709 13626 20765 13628
rect 20789 13626 20845 13628
rect 20549 13574 20595 13626
rect 20595 13574 20605 13626
rect 20629 13574 20659 13626
rect 20659 13574 20671 13626
rect 20671 13574 20685 13626
rect 20709 13574 20723 13626
rect 20723 13574 20735 13626
rect 20735 13574 20765 13626
rect 20789 13574 20799 13626
rect 20799 13574 20845 13626
rect 20549 13572 20605 13574
rect 20629 13572 20685 13574
rect 20709 13572 20765 13574
rect 20789 13572 20845 13574
rect 20718 13232 20774 13288
rect 19338 11736 19394 11792
rect 19338 10648 19394 10704
rect 19338 9968 19394 10024
rect 19246 9832 19302 9888
rect 19154 9560 19210 9616
rect 19062 9424 19118 9480
rect 19614 11192 19670 11248
rect 19614 9016 19670 9072
rect 17750 4378 17806 4380
rect 17830 4378 17886 4380
rect 17910 4378 17966 4380
rect 17990 4378 18046 4380
rect 17750 4326 17796 4378
rect 17796 4326 17806 4378
rect 17830 4326 17860 4378
rect 17860 4326 17872 4378
rect 17872 4326 17886 4378
rect 17910 4326 17924 4378
rect 17924 4326 17936 4378
rect 17936 4326 17966 4378
rect 17990 4326 18000 4378
rect 18000 4326 18046 4378
rect 17750 4324 17806 4326
rect 17830 4324 17886 4326
rect 17910 4324 17966 4326
rect 17990 4324 18046 4326
rect 17750 3290 17806 3292
rect 17830 3290 17886 3292
rect 17910 3290 17966 3292
rect 17990 3290 18046 3292
rect 17750 3238 17796 3290
rect 17796 3238 17806 3290
rect 17830 3238 17860 3290
rect 17860 3238 17872 3290
rect 17872 3238 17886 3290
rect 17910 3238 17924 3290
rect 17924 3238 17936 3290
rect 17936 3238 17966 3290
rect 17990 3238 18000 3290
rect 18000 3238 18046 3290
rect 17750 3236 17806 3238
rect 17830 3236 17886 3238
rect 17910 3236 17966 3238
rect 17990 3236 18046 3238
rect 19338 8472 19394 8528
rect 20549 12538 20605 12540
rect 20629 12538 20685 12540
rect 20709 12538 20765 12540
rect 20789 12538 20845 12540
rect 20549 12486 20595 12538
rect 20595 12486 20605 12538
rect 20629 12486 20659 12538
rect 20659 12486 20671 12538
rect 20671 12486 20685 12538
rect 20709 12486 20723 12538
rect 20723 12486 20735 12538
rect 20735 12486 20765 12538
rect 20789 12486 20799 12538
rect 20799 12486 20845 12538
rect 20549 12484 20605 12486
rect 20629 12484 20685 12486
rect 20709 12484 20765 12486
rect 20789 12484 20845 12486
rect 22374 18808 22430 18864
rect 21546 15952 21602 16008
rect 20549 11450 20605 11452
rect 20629 11450 20685 11452
rect 20709 11450 20765 11452
rect 20789 11450 20845 11452
rect 20549 11398 20595 11450
rect 20595 11398 20605 11450
rect 20629 11398 20659 11450
rect 20659 11398 20671 11450
rect 20671 11398 20685 11450
rect 20709 11398 20723 11450
rect 20723 11398 20735 11450
rect 20735 11398 20765 11450
rect 20789 11398 20799 11450
rect 20799 11398 20845 11450
rect 20549 11396 20605 11398
rect 20629 11396 20685 11398
rect 20709 11396 20765 11398
rect 20789 11396 20845 11398
rect 19522 7112 19578 7168
rect 19430 6976 19486 7032
rect 19798 6976 19854 7032
rect 19430 6452 19486 6488
rect 19430 6432 19432 6452
rect 19432 6432 19484 6452
rect 19484 6432 19486 6452
rect 19982 6976 20038 7032
rect 19890 6432 19946 6488
rect 19430 6024 19486 6080
rect 19798 6024 19854 6080
rect 19614 4800 19670 4856
rect 20166 8744 20222 8800
rect 20549 10362 20605 10364
rect 20629 10362 20685 10364
rect 20709 10362 20765 10364
rect 20789 10362 20845 10364
rect 20549 10310 20595 10362
rect 20595 10310 20605 10362
rect 20629 10310 20659 10362
rect 20659 10310 20671 10362
rect 20671 10310 20685 10362
rect 20709 10310 20723 10362
rect 20723 10310 20735 10362
rect 20735 10310 20765 10362
rect 20789 10310 20799 10362
rect 20799 10310 20845 10362
rect 20549 10308 20605 10310
rect 20629 10308 20685 10310
rect 20709 10308 20765 10310
rect 20789 10308 20845 10310
rect 20549 9274 20605 9276
rect 20629 9274 20685 9276
rect 20709 9274 20765 9276
rect 20789 9274 20845 9276
rect 20549 9222 20595 9274
rect 20595 9222 20605 9274
rect 20629 9222 20659 9274
rect 20659 9222 20671 9274
rect 20671 9222 20685 9274
rect 20709 9222 20723 9274
rect 20723 9222 20735 9274
rect 20735 9222 20765 9274
rect 20789 9222 20799 9274
rect 20799 9222 20845 9274
rect 20549 9220 20605 9222
rect 20629 9220 20685 9222
rect 20709 9220 20765 9222
rect 20789 9220 20845 9222
rect 21362 12144 21418 12200
rect 21362 11056 21418 11112
rect 20718 8880 20774 8936
rect 21270 10124 21326 10160
rect 21270 10104 21272 10124
rect 21272 10104 21324 10124
rect 21324 10104 21326 10124
rect 22650 19216 22706 19272
rect 23018 19896 23074 19952
rect 22098 13368 22154 13424
rect 22006 13132 22008 13152
rect 22008 13132 22060 13152
rect 22060 13132 22062 13152
rect 22006 13096 22062 13132
rect 20074 5616 20130 5672
rect 20549 8186 20605 8188
rect 20629 8186 20685 8188
rect 20709 8186 20765 8188
rect 20789 8186 20845 8188
rect 20549 8134 20595 8186
rect 20595 8134 20605 8186
rect 20629 8134 20659 8186
rect 20659 8134 20671 8186
rect 20671 8134 20685 8186
rect 20709 8134 20723 8186
rect 20723 8134 20735 8186
rect 20735 8134 20765 8186
rect 20789 8134 20799 8186
rect 20799 8134 20845 8186
rect 20549 8132 20605 8134
rect 20629 8132 20685 8134
rect 20709 8132 20765 8134
rect 20789 8132 20845 8134
rect 20549 7098 20605 7100
rect 20629 7098 20685 7100
rect 20709 7098 20765 7100
rect 20789 7098 20845 7100
rect 20549 7046 20595 7098
rect 20595 7046 20605 7098
rect 20629 7046 20659 7098
rect 20659 7046 20671 7098
rect 20671 7046 20685 7098
rect 20709 7046 20723 7098
rect 20723 7046 20735 7098
rect 20735 7046 20765 7098
rect 20789 7046 20799 7098
rect 20799 7046 20845 7098
rect 20549 7044 20605 7046
rect 20629 7044 20685 7046
rect 20709 7044 20765 7046
rect 20789 7044 20845 7046
rect 21178 8336 21234 8392
rect 20549 6010 20605 6012
rect 20629 6010 20685 6012
rect 20709 6010 20765 6012
rect 20789 6010 20845 6012
rect 20549 5958 20595 6010
rect 20595 5958 20605 6010
rect 20629 5958 20659 6010
rect 20659 5958 20671 6010
rect 20671 5958 20685 6010
rect 20709 5958 20723 6010
rect 20723 5958 20735 6010
rect 20735 5958 20765 6010
rect 20789 5958 20799 6010
rect 20799 5958 20845 6010
rect 20549 5956 20605 5958
rect 20629 5956 20685 5958
rect 20709 5956 20765 5958
rect 20789 5956 20845 5958
rect 20442 5616 20498 5672
rect 20549 4922 20605 4924
rect 20629 4922 20685 4924
rect 20709 4922 20765 4924
rect 20789 4922 20845 4924
rect 20549 4870 20595 4922
rect 20595 4870 20605 4922
rect 20629 4870 20659 4922
rect 20659 4870 20671 4922
rect 20671 4870 20685 4922
rect 20709 4870 20723 4922
rect 20723 4870 20735 4922
rect 20735 4870 20765 4922
rect 20789 4870 20799 4922
rect 20799 4870 20845 4922
rect 20549 4868 20605 4870
rect 20629 4868 20685 4870
rect 20709 4868 20765 4870
rect 20789 4868 20845 4870
rect 20534 4664 20590 4720
rect 20549 3834 20605 3836
rect 20629 3834 20685 3836
rect 20709 3834 20765 3836
rect 20789 3834 20845 3836
rect 20549 3782 20595 3834
rect 20595 3782 20605 3834
rect 20629 3782 20659 3834
rect 20659 3782 20671 3834
rect 20671 3782 20685 3834
rect 20709 3782 20723 3834
rect 20723 3782 20735 3834
rect 20735 3782 20765 3834
rect 20789 3782 20799 3834
rect 20799 3782 20845 3834
rect 20549 3780 20605 3782
rect 20629 3780 20685 3782
rect 20709 3780 20765 3782
rect 20789 3780 20845 3782
rect 21270 6604 21272 6624
rect 21272 6604 21324 6624
rect 21324 6604 21326 6624
rect 21270 6568 21326 6604
rect 21270 6024 21326 6080
rect 19706 3052 19762 3088
rect 19706 3032 19708 3052
rect 19708 3032 19760 3052
rect 19760 3032 19762 3052
rect 20994 3032 21050 3088
rect 21546 7404 21602 7440
rect 21546 7384 21548 7404
rect 21548 7384 21600 7404
rect 21600 7384 21602 7404
rect 21454 6296 21510 6352
rect 21546 6024 21602 6080
rect 21362 4392 21418 4448
rect 21454 4120 21510 4176
rect 22466 9832 22522 9888
rect 22374 8744 22430 8800
rect 21914 6568 21970 6624
rect 22098 6432 22154 6488
rect 23018 19352 23074 19408
rect 23018 18808 23074 18864
rect 23018 18264 23074 18320
rect 22926 17856 22982 17912
rect 23202 17720 23258 17776
rect 23110 17584 23166 17640
rect 22742 9696 22798 9752
rect 23202 15000 23258 15056
rect 23110 14456 23166 14512
rect 23202 13368 23258 13424
rect 23478 13912 23534 13968
rect 23110 9424 23166 9480
rect 22650 8492 22706 8528
rect 22650 8472 22652 8492
rect 22652 8472 22704 8492
rect 22704 8472 22706 8492
rect 22466 6740 22468 6760
rect 22468 6740 22520 6760
rect 22520 6740 22522 6760
rect 22466 6704 22522 6740
rect 22558 3612 22560 3632
rect 22560 3612 22612 3632
rect 22612 3612 22614 3632
rect 22558 3576 22614 3612
rect 22374 3440 22430 3496
rect 23018 7928 23074 7984
rect 23018 7384 23074 7440
rect 22834 6296 22890 6352
rect 23018 6840 23074 6896
rect 23018 5752 23074 5808
rect 23018 5208 23074 5264
rect 23018 4664 23074 4720
rect 23386 6160 23442 6216
rect 23018 4120 23074 4176
rect 23018 3576 23074 3632
rect 23018 3032 23074 3088
rect 20549 2746 20605 2748
rect 20629 2746 20685 2748
rect 20709 2746 20765 2748
rect 20789 2746 20845 2748
rect 20549 2694 20595 2746
rect 20595 2694 20605 2746
rect 20629 2694 20659 2746
rect 20659 2694 20671 2746
rect 20671 2694 20685 2746
rect 20709 2694 20723 2746
rect 20723 2694 20735 2746
rect 20735 2694 20765 2746
rect 20789 2694 20799 2746
rect 20799 2694 20845 2746
rect 20549 2692 20605 2694
rect 20629 2692 20685 2694
rect 20709 2692 20765 2694
rect 20789 2692 20845 2694
rect 23662 11600 23718 11656
rect 23018 2488 23074 2544
rect 6554 2202 6610 2204
rect 6634 2202 6690 2204
rect 6714 2202 6770 2204
rect 6794 2202 6850 2204
rect 6554 2150 6600 2202
rect 6600 2150 6610 2202
rect 6634 2150 6664 2202
rect 6664 2150 6676 2202
rect 6676 2150 6690 2202
rect 6714 2150 6728 2202
rect 6728 2150 6740 2202
rect 6740 2150 6770 2202
rect 6794 2150 6804 2202
rect 6804 2150 6850 2202
rect 6554 2148 6610 2150
rect 6634 2148 6690 2150
rect 6714 2148 6770 2150
rect 6794 2148 6850 2150
rect 12152 2202 12208 2204
rect 12232 2202 12288 2204
rect 12312 2202 12368 2204
rect 12392 2202 12448 2204
rect 12152 2150 12198 2202
rect 12198 2150 12208 2202
rect 12232 2150 12262 2202
rect 12262 2150 12274 2202
rect 12274 2150 12288 2202
rect 12312 2150 12326 2202
rect 12326 2150 12338 2202
rect 12338 2150 12368 2202
rect 12392 2150 12402 2202
rect 12402 2150 12448 2202
rect 12152 2148 12208 2150
rect 12232 2148 12288 2150
rect 12312 2148 12368 2150
rect 12392 2148 12448 2150
rect 17750 2202 17806 2204
rect 17830 2202 17886 2204
rect 17910 2202 17966 2204
rect 17990 2202 18046 2204
rect 17750 2150 17796 2202
rect 17796 2150 17806 2202
rect 17830 2150 17860 2202
rect 17860 2150 17872 2202
rect 17872 2150 17886 2202
rect 17910 2150 17924 2202
rect 17924 2150 17936 2202
rect 17936 2150 17966 2202
rect 17990 2150 18000 2202
rect 18000 2150 18046 2202
rect 17750 2148 17806 2150
rect 17830 2148 17886 2150
rect 17910 2148 17966 2150
rect 17990 2148 18046 2150
<< metal3 >>
rect 3745 22336 4061 22337
rect 3745 22272 3751 22336
rect 3815 22272 3831 22336
rect 3895 22272 3911 22336
rect 3975 22272 3991 22336
rect 4055 22272 4061 22336
rect 3745 22271 4061 22272
rect 9343 22336 9659 22337
rect 9343 22272 9349 22336
rect 9413 22272 9429 22336
rect 9493 22272 9509 22336
rect 9573 22272 9589 22336
rect 9653 22272 9659 22336
rect 9343 22271 9659 22272
rect 14941 22336 15257 22337
rect 14941 22272 14947 22336
rect 15011 22272 15027 22336
rect 15091 22272 15107 22336
rect 15171 22272 15187 22336
rect 15251 22272 15257 22336
rect 14941 22271 15257 22272
rect 20539 22336 20855 22337
rect 20539 22272 20545 22336
rect 20609 22272 20625 22336
rect 20689 22272 20705 22336
rect 20769 22272 20785 22336
rect 20849 22272 20855 22336
rect 20539 22271 20855 22272
rect 16430 22068 16436 22132
rect 16500 22130 16506 22132
rect 17401 22130 17467 22133
rect 18597 22130 18663 22133
rect 16500 22070 16866 22130
rect 16500 22068 16506 22070
rect 11237 21994 11303 21997
rect 16806 21994 16866 22070
rect 17401 22128 18663 22130
rect 17401 22072 17406 22128
rect 17462 22072 18602 22128
rect 18658 22072 18663 22128
rect 17401 22070 18663 22072
rect 17401 22067 17467 22070
rect 18597 22067 18663 22070
rect 20529 22130 20595 22133
rect 23800 22130 24600 22160
rect 20529 22128 24600 22130
rect 20529 22072 20534 22128
rect 20590 22072 24600 22128
rect 20529 22070 24600 22072
rect 20529 22067 20595 22070
rect 23800 22040 24600 22070
rect 21817 21994 21883 21997
rect 11237 21992 16682 21994
rect 11237 21936 11242 21992
rect 11298 21936 16682 21992
rect 11237 21934 16682 21936
rect 16806 21992 21883 21994
rect 16806 21936 21822 21992
rect 21878 21936 21883 21992
rect 16806 21934 21883 21936
rect 11237 21931 11303 21934
rect 7097 21858 7163 21861
rect 10041 21858 10107 21861
rect 7097 21856 10107 21858
rect 7097 21800 7102 21856
rect 7158 21800 10046 21856
rect 10102 21800 10107 21856
rect 7097 21798 10107 21800
rect 7097 21795 7163 21798
rect 10041 21795 10107 21798
rect 13721 21858 13787 21861
rect 15929 21858 15995 21861
rect 13721 21856 15995 21858
rect 13721 21800 13726 21856
rect 13782 21800 15934 21856
rect 15990 21800 15995 21856
rect 13721 21798 15995 21800
rect 16622 21858 16682 21934
rect 21817 21931 21883 21934
rect 17217 21858 17283 21861
rect 16622 21856 17283 21858
rect 16622 21800 17222 21856
rect 17278 21800 17283 21856
rect 16622 21798 17283 21800
rect 13721 21795 13787 21798
rect 15929 21795 15995 21798
rect 17217 21795 17283 21798
rect 6544 21792 6860 21793
rect 6544 21728 6550 21792
rect 6614 21728 6630 21792
rect 6694 21728 6710 21792
rect 6774 21728 6790 21792
rect 6854 21728 6860 21792
rect 6544 21727 6860 21728
rect 12142 21792 12458 21793
rect 12142 21728 12148 21792
rect 12212 21728 12228 21792
rect 12292 21728 12308 21792
rect 12372 21728 12388 21792
rect 12452 21728 12458 21792
rect 12142 21727 12458 21728
rect 17740 21792 18056 21793
rect 17740 21728 17746 21792
rect 17810 21728 17826 21792
rect 17890 21728 17906 21792
rect 17970 21728 17986 21792
rect 18050 21728 18056 21792
rect 17740 21727 18056 21728
rect 8385 21722 8451 21725
rect 9213 21722 9279 21725
rect 10777 21722 10843 21725
rect 15009 21722 15075 21725
rect 15653 21722 15719 21725
rect 16297 21722 16363 21725
rect 8385 21720 11162 21722
rect 8385 21664 8390 21720
rect 8446 21664 9218 21720
rect 9274 21664 10782 21720
rect 10838 21664 11162 21720
rect 8385 21662 11162 21664
rect 8385 21659 8451 21662
rect 9213 21659 9279 21662
rect 10777 21659 10843 21662
rect 3969 21586 4035 21589
rect 10869 21586 10935 21589
rect 3969 21584 10935 21586
rect 3969 21528 3974 21584
rect 4030 21528 10874 21584
rect 10930 21528 10935 21584
rect 3969 21526 10935 21528
rect 11102 21586 11162 21662
rect 15009 21720 16363 21722
rect 15009 21664 15014 21720
rect 15070 21664 15658 21720
rect 15714 21664 16302 21720
rect 16358 21664 16363 21720
rect 15009 21662 16363 21664
rect 15009 21659 15075 21662
rect 15653 21659 15719 21662
rect 16297 21659 16363 21662
rect 16481 21722 16547 21725
rect 16481 21720 16682 21722
rect 16481 21664 16486 21720
rect 16542 21664 16682 21720
rect 16481 21662 16682 21664
rect 16481 21659 16547 21662
rect 16430 21586 16436 21588
rect 11102 21526 16436 21586
rect 3969 21523 4035 21526
rect 10869 21523 10935 21526
rect 16430 21524 16436 21526
rect 16500 21524 16506 21588
rect 16622 21586 16682 21662
rect 22461 21586 22527 21589
rect 16622 21584 22527 21586
rect 16622 21528 22466 21584
rect 22522 21528 22527 21584
rect 16622 21526 22527 21528
rect 22461 21523 22527 21526
rect 22645 21586 22711 21589
rect 23800 21586 24600 21616
rect 22645 21584 24600 21586
rect 22645 21528 22650 21584
rect 22706 21528 24600 21584
rect 22645 21526 24600 21528
rect 22645 21523 22711 21526
rect 23800 21496 24600 21526
rect 0 21360 800 21480
rect 4337 21450 4403 21453
rect 14641 21450 14707 21453
rect 20989 21450 21055 21453
rect 4337 21448 14707 21450
rect 4337 21392 4342 21448
rect 4398 21392 14646 21448
rect 14702 21392 14707 21448
rect 4337 21390 14707 21392
rect 4337 21387 4403 21390
rect 14641 21387 14707 21390
rect 14782 21448 21055 21450
rect 14782 21392 20994 21448
rect 21050 21392 21055 21448
rect 14782 21390 21055 21392
rect 4245 21314 4311 21317
rect 7373 21314 7439 21317
rect 13854 21314 13860 21316
rect 4245 21312 7439 21314
rect 4245 21256 4250 21312
rect 4306 21256 7378 21312
rect 7434 21256 7439 21312
rect 4245 21254 7439 21256
rect 4245 21251 4311 21254
rect 7373 21251 7439 21254
rect 12390 21254 13860 21314
rect 3745 21248 4061 21249
rect 3745 21184 3751 21248
rect 3815 21184 3831 21248
rect 3895 21184 3911 21248
rect 3975 21184 3991 21248
rect 4055 21184 4061 21248
rect 3745 21183 4061 21184
rect 9343 21248 9659 21249
rect 9343 21184 9349 21248
rect 9413 21184 9429 21248
rect 9493 21184 9509 21248
rect 9573 21184 9589 21248
rect 9653 21184 9659 21248
rect 9343 21183 9659 21184
rect 2773 21042 2839 21045
rect 8385 21042 8451 21045
rect 12390 21042 12450 21254
rect 13854 21252 13860 21254
rect 13924 21314 13930 21316
rect 14782 21314 14842 21390
rect 20989 21387 21055 21390
rect 13924 21254 14842 21314
rect 15469 21314 15535 21317
rect 16757 21314 16823 21317
rect 15469 21312 16823 21314
rect 15469 21256 15474 21312
rect 15530 21256 16762 21312
rect 16818 21256 16823 21312
rect 15469 21254 16823 21256
rect 13924 21252 13930 21254
rect 15469 21251 15535 21254
rect 16757 21251 16823 21254
rect 17217 21314 17283 21317
rect 17861 21314 17927 21317
rect 17217 21312 17927 21314
rect 17217 21256 17222 21312
rect 17278 21256 17866 21312
rect 17922 21256 17927 21312
rect 17217 21254 17927 21256
rect 17217 21251 17283 21254
rect 17861 21251 17927 21254
rect 14941 21248 15257 21249
rect 14941 21184 14947 21248
rect 15011 21184 15027 21248
rect 15091 21184 15107 21248
rect 15171 21184 15187 21248
rect 15251 21184 15257 21248
rect 14941 21183 15257 21184
rect 20539 21248 20855 21249
rect 20539 21184 20545 21248
rect 20609 21184 20625 21248
rect 20689 21184 20705 21248
rect 20769 21184 20785 21248
rect 20849 21184 20855 21248
rect 20539 21183 20855 21184
rect 15653 21178 15719 21181
rect 16481 21178 16547 21181
rect 15653 21176 16547 21178
rect 15653 21120 15658 21176
rect 15714 21120 16486 21176
rect 16542 21120 16547 21176
rect 15653 21118 16547 21120
rect 15653 21115 15719 21118
rect 16481 21115 16547 21118
rect 17125 21178 17191 21181
rect 18413 21178 18479 21181
rect 17125 21176 18479 21178
rect 17125 21120 17130 21176
rect 17186 21120 18418 21176
rect 18474 21120 18479 21176
rect 17125 21118 18479 21120
rect 17125 21115 17191 21118
rect 18413 21115 18479 21118
rect 2773 21040 12450 21042
rect 2773 20984 2778 21040
rect 2834 20984 8390 21040
rect 8446 20984 12450 21040
rect 2773 20982 12450 20984
rect 14733 21042 14799 21045
rect 18137 21042 18203 21045
rect 20805 21042 20871 21045
rect 14733 21040 20871 21042
rect 14733 20984 14738 21040
rect 14794 20984 18142 21040
rect 18198 20984 20810 21040
rect 20866 20984 20871 21040
rect 14733 20982 20871 20984
rect 2773 20979 2839 20982
rect 8385 20979 8451 20982
rect 14733 20979 14799 20982
rect 18137 20979 18203 20982
rect 20805 20979 20871 20982
rect 23013 21042 23079 21045
rect 23800 21042 24600 21072
rect 23013 21040 24600 21042
rect 23013 20984 23018 21040
rect 23074 20984 24600 21040
rect 23013 20982 24600 20984
rect 23013 20979 23079 20982
rect 23800 20952 24600 20982
rect 3693 20906 3759 20909
rect 11145 20906 11211 20909
rect 21357 20906 21423 20909
rect 3693 20904 7482 20906
rect 3693 20848 3698 20904
rect 3754 20848 7482 20904
rect 3693 20846 7482 20848
rect 3693 20843 3759 20846
rect 7422 20770 7482 20846
rect 11145 20904 21423 20906
rect 11145 20848 11150 20904
rect 11206 20848 21362 20904
rect 21418 20848 21423 20904
rect 11145 20846 21423 20848
rect 11145 20843 11211 20846
rect 21357 20843 21423 20846
rect 11237 20770 11303 20773
rect 7422 20768 11303 20770
rect 7422 20712 11242 20768
rect 11298 20712 11303 20768
rect 7422 20710 11303 20712
rect 11237 20707 11303 20710
rect 14641 20770 14707 20773
rect 15653 20770 15719 20773
rect 14641 20768 15719 20770
rect 14641 20712 14646 20768
rect 14702 20712 15658 20768
rect 15714 20712 15719 20768
rect 14641 20710 15719 20712
rect 14641 20707 14707 20710
rect 15653 20707 15719 20710
rect 21030 20708 21036 20772
rect 21100 20770 21106 20772
rect 22185 20770 22251 20773
rect 21100 20768 22251 20770
rect 21100 20712 22190 20768
rect 22246 20712 22251 20768
rect 21100 20710 22251 20712
rect 21100 20708 21106 20710
rect 22185 20707 22251 20710
rect 6544 20704 6860 20705
rect 6544 20640 6550 20704
rect 6614 20640 6630 20704
rect 6694 20640 6710 20704
rect 6774 20640 6790 20704
rect 6854 20640 6860 20704
rect 6544 20639 6860 20640
rect 12142 20704 12458 20705
rect 12142 20640 12148 20704
rect 12212 20640 12228 20704
rect 12292 20640 12308 20704
rect 12372 20640 12388 20704
rect 12452 20640 12458 20704
rect 12142 20639 12458 20640
rect 17740 20704 18056 20705
rect 17740 20640 17746 20704
rect 17810 20640 17826 20704
rect 17890 20640 17906 20704
rect 17970 20640 17986 20704
rect 18050 20640 18056 20704
rect 17740 20639 18056 20640
rect 3877 20498 3943 20501
rect 11145 20498 11211 20501
rect 3877 20496 11211 20498
rect 3877 20440 3882 20496
rect 3938 20440 11150 20496
rect 11206 20440 11211 20496
rect 3877 20438 11211 20440
rect 3877 20435 3943 20438
rect 11145 20435 11211 20438
rect 12157 20498 12223 20501
rect 17033 20498 17099 20501
rect 18505 20498 18571 20501
rect 12157 20496 18571 20498
rect 12157 20440 12162 20496
rect 12218 20440 17038 20496
rect 17094 20440 18510 20496
rect 18566 20440 18571 20496
rect 12157 20438 18571 20440
rect 12157 20435 12223 20438
rect 17033 20435 17099 20438
rect 18505 20435 18571 20438
rect 23013 20498 23079 20501
rect 23800 20498 24600 20528
rect 23013 20496 24600 20498
rect 23013 20440 23018 20496
rect 23074 20440 24600 20496
rect 23013 20438 24600 20440
rect 23013 20435 23079 20438
rect 23800 20408 24600 20438
rect 12617 20362 12683 20365
rect 16389 20362 16455 20365
rect 12617 20360 16455 20362
rect 12617 20304 12622 20360
rect 12678 20304 16394 20360
rect 16450 20304 16455 20360
rect 12617 20302 16455 20304
rect 12617 20299 12683 20302
rect 16389 20299 16455 20302
rect 3745 20160 4061 20161
rect 3745 20096 3751 20160
rect 3815 20096 3831 20160
rect 3895 20096 3911 20160
rect 3975 20096 3991 20160
rect 4055 20096 4061 20160
rect 3745 20095 4061 20096
rect 9343 20160 9659 20161
rect 9343 20096 9349 20160
rect 9413 20096 9429 20160
rect 9493 20096 9509 20160
rect 9573 20096 9589 20160
rect 9653 20096 9659 20160
rect 9343 20095 9659 20096
rect 14941 20160 15257 20161
rect 14941 20096 14947 20160
rect 15011 20096 15027 20160
rect 15091 20096 15107 20160
rect 15171 20096 15187 20160
rect 15251 20096 15257 20160
rect 14941 20095 15257 20096
rect 20539 20160 20855 20161
rect 20539 20096 20545 20160
rect 20609 20096 20625 20160
rect 20689 20096 20705 20160
rect 20769 20096 20785 20160
rect 20849 20096 20855 20160
rect 20539 20095 20855 20096
rect 11973 19954 12039 19957
rect 13721 19954 13787 19957
rect 18045 19954 18111 19957
rect 11973 19952 13554 19954
rect 11973 19896 11978 19952
rect 12034 19896 13554 19952
rect 11973 19894 13554 19896
rect 11973 19891 12039 19894
rect 4429 19818 4495 19821
rect 9489 19818 9555 19821
rect 4429 19816 9555 19818
rect 4429 19760 4434 19816
rect 4490 19760 9494 19816
rect 9550 19760 9555 19816
rect 4429 19758 9555 19760
rect 4429 19755 4495 19758
rect 9489 19755 9555 19758
rect 11421 19818 11487 19821
rect 13494 19818 13554 19894
rect 13721 19952 18111 19954
rect 13721 19896 13726 19952
rect 13782 19896 18050 19952
rect 18106 19896 18111 19952
rect 13721 19894 18111 19896
rect 13721 19891 13787 19894
rect 18045 19891 18111 19894
rect 23013 19954 23079 19957
rect 23800 19954 24600 19984
rect 23013 19952 24600 19954
rect 23013 19896 23018 19952
rect 23074 19896 24600 19952
rect 23013 19894 24600 19896
rect 23013 19891 23079 19894
rect 23800 19864 24600 19894
rect 18597 19818 18663 19821
rect 11421 19816 13370 19818
rect 11421 19760 11426 19816
rect 11482 19760 13370 19816
rect 11421 19758 13370 19760
rect 13494 19816 18663 19818
rect 13494 19760 18602 19816
rect 18658 19760 18663 19816
rect 13494 19758 18663 19760
rect 11421 19755 11487 19758
rect 6544 19616 6860 19617
rect 6544 19552 6550 19616
rect 6614 19552 6630 19616
rect 6694 19552 6710 19616
rect 6774 19552 6790 19616
rect 6854 19552 6860 19616
rect 6544 19551 6860 19552
rect 12142 19616 12458 19617
rect 12142 19552 12148 19616
rect 12212 19552 12228 19616
rect 12292 19552 12308 19616
rect 12372 19552 12388 19616
rect 12452 19552 12458 19616
rect 12142 19551 12458 19552
rect 11789 19546 11855 19549
rect 9262 19544 11855 19546
rect 9262 19488 11794 19544
rect 11850 19488 11855 19544
rect 9262 19486 11855 19488
rect 13310 19546 13370 19758
rect 18597 19755 18663 19758
rect 20897 19818 20963 19821
rect 21582 19818 21588 19820
rect 20897 19816 21588 19818
rect 20897 19760 20902 19816
rect 20958 19760 21588 19816
rect 20897 19758 21588 19760
rect 20897 19755 20963 19758
rect 21582 19756 21588 19758
rect 21652 19756 21658 19820
rect 17740 19616 18056 19617
rect 17740 19552 17746 19616
rect 17810 19552 17826 19616
rect 17890 19552 17906 19616
rect 17970 19552 17986 19616
rect 18050 19552 18056 19616
rect 17740 19551 18056 19552
rect 13310 19486 17602 19546
rect 2681 19410 2747 19413
rect 9262 19410 9322 19486
rect 11789 19483 11855 19486
rect 2681 19408 9322 19410
rect 2681 19352 2686 19408
rect 2742 19352 9322 19408
rect 2681 19350 9322 19352
rect 9489 19410 9555 19413
rect 15653 19410 15719 19413
rect 9489 19408 15719 19410
rect 9489 19352 9494 19408
rect 9550 19352 15658 19408
rect 15714 19352 15719 19408
rect 9489 19350 15719 19352
rect 17542 19410 17602 19486
rect 19977 19410 20043 19413
rect 17542 19408 20043 19410
rect 17542 19352 19982 19408
rect 20038 19352 20043 19408
rect 17542 19350 20043 19352
rect 2681 19347 2747 19350
rect 9489 19347 9555 19350
rect 15653 19347 15719 19350
rect 19977 19347 20043 19350
rect 23013 19410 23079 19413
rect 23800 19410 24600 19440
rect 23013 19408 24600 19410
rect 23013 19352 23018 19408
rect 23074 19352 24600 19408
rect 23013 19350 24600 19352
rect 23013 19347 23079 19350
rect 23800 19320 24600 19350
rect 18873 19274 18939 19277
rect 22645 19274 22711 19277
rect 18873 19272 22711 19274
rect 18873 19216 18878 19272
rect 18934 19216 22650 19272
rect 22706 19216 22711 19272
rect 18873 19214 22711 19216
rect 18873 19211 18939 19214
rect 22645 19211 22711 19214
rect 3745 19072 4061 19073
rect 3745 19008 3751 19072
rect 3815 19008 3831 19072
rect 3895 19008 3911 19072
rect 3975 19008 3991 19072
rect 4055 19008 4061 19072
rect 3745 19007 4061 19008
rect 9343 19072 9659 19073
rect 9343 19008 9349 19072
rect 9413 19008 9429 19072
rect 9493 19008 9509 19072
rect 9573 19008 9589 19072
rect 9653 19008 9659 19072
rect 9343 19007 9659 19008
rect 14941 19072 15257 19073
rect 14941 19008 14947 19072
rect 15011 19008 15027 19072
rect 15091 19008 15107 19072
rect 15171 19008 15187 19072
rect 15251 19008 15257 19072
rect 14941 19007 15257 19008
rect 20539 19072 20855 19073
rect 20539 19008 20545 19072
rect 20609 19008 20625 19072
rect 20689 19008 20705 19072
rect 20769 19008 20785 19072
rect 20849 19008 20855 19072
rect 20539 19007 20855 19008
rect 12985 18866 13051 18869
rect 13445 18866 13511 18869
rect 12985 18864 13511 18866
rect 12985 18808 12990 18864
rect 13046 18808 13450 18864
rect 13506 18808 13511 18864
rect 12985 18806 13511 18808
rect 12985 18803 13051 18806
rect 13445 18803 13511 18806
rect 20069 18866 20135 18869
rect 20805 18866 20871 18869
rect 22369 18866 22435 18869
rect 20069 18864 22435 18866
rect 20069 18808 20074 18864
rect 20130 18808 20810 18864
rect 20866 18808 22374 18864
rect 22430 18808 22435 18864
rect 20069 18806 22435 18808
rect 20069 18803 20135 18806
rect 20805 18803 20871 18806
rect 22369 18803 22435 18806
rect 23013 18866 23079 18869
rect 23800 18866 24600 18896
rect 23013 18864 24600 18866
rect 23013 18808 23018 18864
rect 23074 18808 24600 18864
rect 23013 18806 24600 18808
rect 23013 18803 23079 18806
rect 23800 18776 24600 18806
rect 2681 18730 2747 18733
rect 13353 18730 13419 18733
rect 2681 18728 13419 18730
rect 2681 18672 2686 18728
rect 2742 18672 13358 18728
rect 13414 18672 13419 18728
rect 2681 18670 13419 18672
rect 2681 18667 2747 18670
rect 13353 18667 13419 18670
rect 18597 18594 18663 18597
rect 21030 18594 21036 18596
rect 18597 18592 21036 18594
rect 18597 18536 18602 18592
rect 18658 18536 21036 18592
rect 18597 18534 21036 18536
rect 18597 18531 18663 18534
rect 21030 18532 21036 18534
rect 21100 18532 21106 18596
rect 6544 18528 6860 18529
rect 6544 18464 6550 18528
rect 6614 18464 6630 18528
rect 6694 18464 6710 18528
rect 6774 18464 6790 18528
rect 6854 18464 6860 18528
rect 6544 18463 6860 18464
rect 12142 18528 12458 18529
rect 12142 18464 12148 18528
rect 12212 18464 12228 18528
rect 12292 18464 12308 18528
rect 12372 18464 12388 18528
rect 12452 18464 12458 18528
rect 12142 18463 12458 18464
rect 17740 18528 18056 18529
rect 17740 18464 17746 18528
rect 17810 18464 17826 18528
rect 17890 18464 17906 18528
rect 17970 18464 17986 18528
rect 18050 18464 18056 18528
rect 17740 18463 18056 18464
rect 23013 18322 23079 18325
rect 23800 18322 24600 18352
rect 23013 18320 24600 18322
rect 23013 18264 23018 18320
rect 23074 18264 24600 18320
rect 23013 18262 24600 18264
rect 23013 18259 23079 18262
rect 23800 18232 24600 18262
rect 18873 18186 18939 18189
rect 19701 18186 19767 18189
rect 18873 18184 19767 18186
rect 18873 18128 18878 18184
rect 18934 18128 19706 18184
rect 19762 18128 19767 18184
rect 18873 18126 19767 18128
rect 18873 18123 18939 18126
rect 19701 18123 19767 18126
rect 3745 17984 4061 17985
rect 3745 17920 3751 17984
rect 3815 17920 3831 17984
rect 3895 17920 3911 17984
rect 3975 17920 3991 17984
rect 4055 17920 4061 17984
rect 3745 17919 4061 17920
rect 9343 17984 9659 17985
rect 9343 17920 9349 17984
rect 9413 17920 9429 17984
rect 9493 17920 9509 17984
rect 9573 17920 9589 17984
rect 9653 17920 9659 17984
rect 9343 17919 9659 17920
rect 14941 17984 15257 17985
rect 14941 17920 14947 17984
rect 15011 17920 15027 17984
rect 15091 17920 15107 17984
rect 15171 17920 15187 17984
rect 15251 17920 15257 17984
rect 14941 17919 15257 17920
rect 20539 17984 20855 17985
rect 20539 17920 20545 17984
rect 20609 17920 20625 17984
rect 20689 17920 20705 17984
rect 20769 17920 20785 17984
rect 20849 17920 20855 17984
rect 20539 17919 20855 17920
rect 13905 17916 13971 17917
rect 13854 17852 13860 17916
rect 13924 17914 13971 17916
rect 22921 17914 22987 17917
rect 13924 17912 14016 17914
rect 13966 17856 14016 17912
rect 13924 17854 14016 17856
rect 22050 17912 22987 17914
rect 22050 17856 22926 17912
rect 22982 17856 22987 17912
rect 22050 17854 22987 17856
rect 13924 17852 13971 17854
rect 13905 17851 13971 17852
rect 19057 17778 19123 17781
rect 22050 17778 22110 17854
rect 22921 17851 22987 17854
rect 19057 17776 22110 17778
rect 19057 17720 19062 17776
rect 19118 17720 22110 17776
rect 19057 17718 22110 17720
rect 23197 17778 23263 17781
rect 23800 17778 24600 17808
rect 23197 17776 24600 17778
rect 23197 17720 23202 17776
rect 23258 17720 24600 17776
rect 23197 17718 24600 17720
rect 19057 17715 19123 17718
rect 23197 17715 23263 17718
rect 23800 17688 24600 17718
rect 17309 17642 17375 17645
rect 23105 17642 23171 17645
rect 17309 17640 23171 17642
rect 17309 17584 17314 17640
rect 17370 17584 23110 17640
rect 23166 17584 23171 17640
rect 17309 17582 23171 17584
rect 17309 17579 17375 17582
rect 23105 17579 23171 17582
rect 18505 17506 18571 17509
rect 20897 17506 20963 17509
rect 18505 17504 22110 17506
rect 18505 17448 18510 17504
rect 18566 17448 20902 17504
rect 20958 17448 22110 17504
rect 18505 17446 22110 17448
rect 18505 17443 18571 17446
rect 20897 17443 20963 17446
rect 6544 17440 6860 17441
rect 6544 17376 6550 17440
rect 6614 17376 6630 17440
rect 6694 17376 6710 17440
rect 6774 17376 6790 17440
rect 6854 17376 6860 17440
rect 6544 17375 6860 17376
rect 12142 17440 12458 17441
rect 12142 17376 12148 17440
rect 12212 17376 12228 17440
rect 12292 17376 12308 17440
rect 12372 17376 12388 17440
rect 12452 17376 12458 17440
rect 12142 17375 12458 17376
rect 17740 17440 18056 17441
rect 17740 17376 17746 17440
rect 17810 17376 17826 17440
rect 17890 17376 17906 17440
rect 17970 17376 17986 17440
rect 18050 17376 18056 17440
rect 17740 17375 18056 17376
rect 22050 17234 22110 17446
rect 23800 17234 24600 17264
rect 22050 17174 24600 17234
rect 23800 17144 24600 17174
rect 3745 16896 4061 16897
rect 3745 16832 3751 16896
rect 3815 16832 3831 16896
rect 3895 16832 3911 16896
rect 3975 16832 3991 16896
rect 4055 16832 4061 16896
rect 3745 16831 4061 16832
rect 9343 16896 9659 16897
rect 9343 16832 9349 16896
rect 9413 16832 9429 16896
rect 9493 16832 9509 16896
rect 9573 16832 9589 16896
rect 9653 16832 9659 16896
rect 9343 16831 9659 16832
rect 14941 16896 15257 16897
rect 14941 16832 14947 16896
rect 15011 16832 15027 16896
rect 15091 16832 15107 16896
rect 15171 16832 15187 16896
rect 15251 16832 15257 16896
rect 14941 16831 15257 16832
rect 20539 16896 20855 16897
rect 20539 16832 20545 16896
rect 20609 16832 20625 16896
rect 20689 16832 20705 16896
rect 20769 16832 20785 16896
rect 20849 16832 20855 16896
rect 20539 16831 20855 16832
rect 18505 16690 18571 16693
rect 23800 16690 24600 16720
rect 18505 16688 24600 16690
rect 18505 16632 18510 16688
rect 18566 16632 24600 16688
rect 18505 16630 24600 16632
rect 18505 16627 18571 16630
rect 23800 16600 24600 16630
rect 2405 16418 2471 16421
rect 6085 16418 6151 16421
rect 6269 16418 6335 16421
rect 2405 16416 6335 16418
rect 2405 16360 2410 16416
rect 2466 16360 6090 16416
rect 6146 16360 6274 16416
rect 6330 16360 6335 16416
rect 2405 16358 6335 16360
rect 2405 16355 2471 16358
rect 6085 16355 6151 16358
rect 6269 16355 6335 16358
rect 6544 16352 6860 16353
rect 6544 16288 6550 16352
rect 6614 16288 6630 16352
rect 6694 16288 6710 16352
rect 6774 16288 6790 16352
rect 6854 16288 6860 16352
rect 6544 16287 6860 16288
rect 12142 16352 12458 16353
rect 12142 16288 12148 16352
rect 12212 16288 12228 16352
rect 12292 16288 12308 16352
rect 12372 16288 12388 16352
rect 12452 16288 12458 16352
rect 12142 16287 12458 16288
rect 17740 16352 18056 16353
rect 17740 16288 17746 16352
rect 17810 16288 17826 16352
rect 17890 16288 17906 16352
rect 17970 16288 17986 16352
rect 18050 16288 18056 16352
rect 17740 16287 18056 16288
rect 19425 16146 19491 16149
rect 23800 16146 24600 16176
rect 19425 16144 24600 16146
rect 19425 16088 19430 16144
rect 19486 16088 24600 16144
rect 19425 16086 24600 16088
rect 19425 16083 19491 16086
rect 23800 16056 24600 16086
rect 19149 16010 19215 16013
rect 21541 16010 21607 16013
rect 19149 16008 21607 16010
rect 19149 15952 19154 16008
rect 19210 15952 21546 16008
rect 21602 15952 21607 16008
rect 19149 15950 21607 15952
rect 19149 15947 19215 15950
rect 21541 15947 21607 15950
rect 3745 15808 4061 15809
rect 3745 15744 3751 15808
rect 3815 15744 3831 15808
rect 3895 15744 3911 15808
rect 3975 15744 3991 15808
rect 4055 15744 4061 15808
rect 3745 15743 4061 15744
rect 9343 15808 9659 15809
rect 9343 15744 9349 15808
rect 9413 15744 9429 15808
rect 9493 15744 9509 15808
rect 9573 15744 9589 15808
rect 9653 15744 9659 15808
rect 9343 15743 9659 15744
rect 14941 15808 15257 15809
rect 14941 15744 14947 15808
rect 15011 15744 15027 15808
rect 15091 15744 15107 15808
rect 15171 15744 15187 15808
rect 15251 15744 15257 15808
rect 14941 15743 15257 15744
rect 20539 15808 20855 15809
rect 20539 15744 20545 15808
rect 20609 15744 20625 15808
rect 20689 15744 20705 15808
rect 20769 15744 20785 15808
rect 20849 15744 20855 15808
rect 20539 15743 20855 15744
rect 18873 15604 18939 15605
rect 18822 15602 18828 15604
rect 18782 15542 18828 15602
rect 18892 15600 18939 15604
rect 18934 15544 18939 15600
rect 18822 15540 18828 15542
rect 18892 15540 18939 15544
rect 18873 15539 18939 15540
rect 19149 15602 19215 15605
rect 23800 15602 24600 15632
rect 19149 15600 24600 15602
rect 19149 15544 19154 15600
rect 19210 15544 24600 15600
rect 19149 15542 24600 15544
rect 19149 15539 19215 15542
rect 23800 15512 24600 15542
rect 3233 15466 3299 15469
rect 8661 15466 8727 15469
rect 3233 15464 8727 15466
rect 3233 15408 3238 15464
rect 3294 15408 8666 15464
rect 8722 15408 8727 15464
rect 3233 15406 8727 15408
rect 3233 15403 3299 15406
rect 8661 15403 8727 15406
rect 0 15330 800 15360
rect 1485 15330 1551 15333
rect 0 15328 1551 15330
rect 0 15272 1490 15328
rect 1546 15272 1551 15328
rect 0 15270 1551 15272
rect 0 15240 800 15270
rect 1485 15267 1551 15270
rect 6544 15264 6860 15265
rect 6544 15200 6550 15264
rect 6614 15200 6630 15264
rect 6694 15200 6710 15264
rect 6774 15200 6790 15264
rect 6854 15200 6860 15264
rect 6544 15199 6860 15200
rect 12142 15264 12458 15265
rect 12142 15200 12148 15264
rect 12212 15200 12228 15264
rect 12292 15200 12308 15264
rect 12372 15200 12388 15264
rect 12452 15200 12458 15264
rect 12142 15199 12458 15200
rect 17740 15264 18056 15265
rect 17740 15200 17746 15264
rect 17810 15200 17826 15264
rect 17890 15200 17906 15264
rect 17970 15200 17986 15264
rect 18050 15200 18056 15264
rect 17740 15199 18056 15200
rect 23197 15058 23263 15061
rect 23800 15058 24600 15088
rect 23197 15056 24600 15058
rect 23197 15000 23202 15056
rect 23258 15000 24600 15056
rect 23197 14998 24600 15000
rect 23197 14995 23263 14998
rect 23800 14968 24600 14998
rect 16573 14922 16639 14925
rect 21081 14922 21147 14925
rect 16573 14920 21147 14922
rect 16573 14864 16578 14920
rect 16634 14864 21086 14920
rect 21142 14864 21147 14920
rect 16573 14862 21147 14864
rect 16573 14859 16639 14862
rect 21081 14859 21147 14862
rect 3745 14720 4061 14721
rect 3745 14656 3751 14720
rect 3815 14656 3831 14720
rect 3895 14656 3911 14720
rect 3975 14656 3991 14720
rect 4055 14656 4061 14720
rect 3745 14655 4061 14656
rect 9343 14720 9659 14721
rect 9343 14656 9349 14720
rect 9413 14656 9429 14720
rect 9493 14656 9509 14720
rect 9573 14656 9589 14720
rect 9653 14656 9659 14720
rect 9343 14655 9659 14656
rect 14941 14720 15257 14721
rect 14941 14656 14947 14720
rect 15011 14656 15027 14720
rect 15091 14656 15107 14720
rect 15171 14656 15187 14720
rect 15251 14656 15257 14720
rect 14941 14655 15257 14656
rect 20539 14720 20855 14721
rect 20539 14656 20545 14720
rect 20609 14656 20625 14720
rect 20689 14656 20705 14720
rect 20769 14656 20785 14720
rect 20849 14656 20855 14720
rect 20539 14655 20855 14656
rect 23105 14514 23171 14517
rect 23800 14514 24600 14544
rect 23105 14512 24600 14514
rect 23105 14456 23110 14512
rect 23166 14456 24600 14512
rect 23105 14454 24600 14456
rect 23105 14451 23171 14454
rect 23800 14424 24600 14454
rect 14733 14378 14799 14381
rect 20989 14378 21055 14381
rect 14733 14376 21055 14378
rect 14733 14320 14738 14376
rect 14794 14320 20994 14376
rect 21050 14320 21055 14376
rect 14733 14318 21055 14320
rect 14733 14315 14799 14318
rect 20989 14315 21055 14318
rect 6544 14176 6860 14177
rect 6544 14112 6550 14176
rect 6614 14112 6630 14176
rect 6694 14112 6710 14176
rect 6774 14112 6790 14176
rect 6854 14112 6860 14176
rect 6544 14111 6860 14112
rect 12142 14176 12458 14177
rect 12142 14112 12148 14176
rect 12212 14112 12228 14176
rect 12292 14112 12308 14176
rect 12372 14112 12388 14176
rect 12452 14112 12458 14176
rect 12142 14111 12458 14112
rect 17740 14176 18056 14177
rect 17740 14112 17746 14176
rect 17810 14112 17826 14176
rect 17890 14112 17906 14176
rect 17970 14112 17986 14176
rect 18050 14112 18056 14176
rect 17740 14111 18056 14112
rect 5625 13970 5691 13973
rect 6545 13970 6611 13973
rect 5625 13968 6611 13970
rect 5625 13912 5630 13968
rect 5686 13912 6550 13968
rect 6606 13912 6611 13968
rect 5625 13910 6611 13912
rect 5625 13907 5691 13910
rect 6545 13907 6611 13910
rect 23473 13970 23539 13973
rect 23800 13970 24600 14000
rect 23473 13968 24600 13970
rect 23473 13912 23478 13968
rect 23534 13912 24600 13968
rect 23473 13910 24600 13912
rect 23473 13907 23539 13910
rect 23800 13880 24600 13910
rect 4429 13834 4495 13837
rect 8385 13834 8451 13837
rect 4429 13832 8451 13834
rect 4429 13776 4434 13832
rect 4490 13776 8390 13832
rect 8446 13776 8451 13832
rect 4429 13774 8451 13776
rect 4429 13771 4495 13774
rect 8385 13771 8451 13774
rect 3745 13632 4061 13633
rect 3745 13568 3751 13632
rect 3815 13568 3831 13632
rect 3895 13568 3911 13632
rect 3975 13568 3991 13632
rect 4055 13568 4061 13632
rect 3745 13567 4061 13568
rect 9343 13632 9659 13633
rect 9343 13568 9349 13632
rect 9413 13568 9429 13632
rect 9493 13568 9509 13632
rect 9573 13568 9589 13632
rect 9653 13568 9659 13632
rect 9343 13567 9659 13568
rect 14941 13632 15257 13633
rect 14941 13568 14947 13632
rect 15011 13568 15027 13632
rect 15091 13568 15107 13632
rect 15171 13568 15187 13632
rect 15251 13568 15257 13632
rect 14941 13567 15257 13568
rect 20539 13632 20855 13633
rect 20539 13568 20545 13632
rect 20609 13568 20625 13632
rect 20689 13568 20705 13632
rect 20769 13568 20785 13632
rect 20849 13568 20855 13632
rect 20539 13567 20855 13568
rect 14089 13426 14155 13429
rect 22093 13426 22159 13429
rect 14089 13424 22159 13426
rect 14089 13368 14094 13424
rect 14150 13368 22098 13424
rect 22154 13368 22159 13424
rect 14089 13366 22159 13368
rect 14089 13363 14155 13366
rect 22093 13363 22159 13366
rect 23197 13426 23263 13429
rect 23800 13426 24600 13456
rect 23197 13424 24600 13426
rect 23197 13368 23202 13424
rect 23258 13368 24600 13424
rect 23197 13366 24600 13368
rect 23197 13363 23263 13366
rect 23800 13336 24600 13366
rect 16573 13290 16639 13293
rect 20713 13290 20779 13293
rect 16573 13288 20779 13290
rect 16573 13232 16578 13288
rect 16634 13232 20718 13288
rect 20774 13232 20779 13288
rect 16573 13230 20779 13232
rect 16573 13227 16639 13230
rect 20713 13227 20779 13230
rect 19333 13154 19399 13157
rect 22001 13154 22067 13157
rect 19333 13152 22067 13154
rect 19333 13096 19338 13152
rect 19394 13096 22006 13152
rect 22062 13096 22067 13152
rect 19333 13094 22067 13096
rect 19333 13091 19399 13094
rect 22001 13091 22067 13094
rect 6544 13088 6860 13089
rect 6544 13024 6550 13088
rect 6614 13024 6630 13088
rect 6694 13024 6710 13088
rect 6774 13024 6790 13088
rect 6854 13024 6860 13088
rect 6544 13023 6860 13024
rect 12142 13088 12458 13089
rect 12142 13024 12148 13088
rect 12212 13024 12228 13088
rect 12292 13024 12308 13088
rect 12372 13024 12388 13088
rect 12452 13024 12458 13088
rect 12142 13023 12458 13024
rect 17740 13088 18056 13089
rect 17740 13024 17746 13088
rect 17810 13024 17826 13088
rect 17890 13024 17906 13088
rect 17970 13024 17986 13088
rect 18050 13024 18056 13088
rect 17740 13023 18056 13024
rect 19057 12882 19123 12885
rect 19190 12882 19196 12884
rect 19057 12880 19196 12882
rect 19057 12824 19062 12880
rect 19118 12824 19196 12880
rect 19057 12822 19196 12824
rect 19057 12819 19123 12822
rect 19190 12820 19196 12822
rect 19260 12820 19266 12884
rect 23800 12882 24600 12912
rect 22050 12822 24600 12882
rect 18505 12746 18571 12749
rect 22050 12746 22110 12822
rect 23800 12792 24600 12822
rect 18505 12744 22110 12746
rect 18505 12688 18510 12744
rect 18566 12688 22110 12744
rect 18505 12686 22110 12688
rect 18505 12683 18571 12686
rect 3745 12544 4061 12545
rect 3745 12480 3751 12544
rect 3815 12480 3831 12544
rect 3895 12480 3911 12544
rect 3975 12480 3991 12544
rect 4055 12480 4061 12544
rect 3745 12479 4061 12480
rect 9343 12544 9659 12545
rect 9343 12480 9349 12544
rect 9413 12480 9429 12544
rect 9493 12480 9509 12544
rect 9573 12480 9589 12544
rect 9653 12480 9659 12544
rect 9343 12479 9659 12480
rect 14941 12544 15257 12545
rect 14941 12480 14947 12544
rect 15011 12480 15027 12544
rect 15091 12480 15107 12544
rect 15171 12480 15187 12544
rect 15251 12480 15257 12544
rect 14941 12479 15257 12480
rect 20539 12544 20855 12545
rect 20539 12480 20545 12544
rect 20609 12480 20625 12544
rect 20689 12480 20705 12544
rect 20769 12480 20785 12544
rect 20849 12480 20855 12544
rect 20539 12479 20855 12480
rect 18873 12338 18939 12341
rect 23800 12338 24600 12368
rect 18873 12336 24600 12338
rect 18873 12280 18878 12336
rect 18934 12280 24600 12336
rect 18873 12278 24600 12280
rect 18873 12275 18939 12278
rect 23800 12248 24600 12278
rect 18229 12202 18295 12205
rect 21357 12202 21423 12205
rect 18229 12200 21423 12202
rect 18229 12144 18234 12200
rect 18290 12144 21362 12200
rect 21418 12144 21423 12200
rect 18229 12142 21423 12144
rect 18229 12139 18295 12142
rect 21357 12139 21423 12142
rect 6544 12000 6860 12001
rect 6544 11936 6550 12000
rect 6614 11936 6630 12000
rect 6694 11936 6710 12000
rect 6774 11936 6790 12000
rect 6854 11936 6860 12000
rect 6544 11935 6860 11936
rect 12142 12000 12458 12001
rect 12142 11936 12148 12000
rect 12212 11936 12228 12000
rect 12292 11936 12308 12000
rect 12372 11936 12388 12000
rect 12452 11936 12458 12000
rect 12142 11935 12458 11936
rect 17740 12000 18056 12001
rect 17740 11936 17746 12000
rect 17810 11936 17826 12000
rect 17890 11936 17906 12000
rect 17970 11936 17986 12000
rect 18050 11936 18056 12000
rect 17740 11935 18056 11936
rect 19333 11794 19399 11797
rect 23800 11794 24600 11824
rect 19333 11792 24600 11794
rect 19333 11736 19338 11792
rect 19394 11736 24600 11792
rect 19333 11734 24600 11736
rect 19333 11731 19399 11734
rect 23800 11704 24600 11734
rect 18781 11658 18847 11661
rect 23657 11658 23723 11661
rect 18781 11656 23723 11658
rect 18781 11600 18786 11656
rect 18842 11600 23662 11656
rect 23718 11600 23723 11656
rect 18781 11598 23723 11600
rect 18781 11595 18847 11598
rect 23657 11595 23723 11598
rect 3745 11456 4061 11457
rect 3745 11392 3751 11456
rect 3815 11392 3831 11456
rect 3895 11392 3911 11456
rect 3975 11392 3991 11456
rect 4055 11392 4061 11456
rect 3745 11391 4061 11392
rect 9343 11456 9659 11457
rect 9343 11392 9349 11456
rect 9413 11392 9429 11456
rect 9493 11392 9509 11456
rect 9573 11392 9589 11456
rect 9653 11392 9659 11456
rect 9343 11391 9659 11392
rect 14941 11456 15257 11457
rect 14941 11392 14947 11456
rect 15011 11392 15027 11456
rect 15091 11392 15107 11456
rect 15171 11392 15187 11456
rect 15251 11392 15257 11456
rect 14941 11391 15257 11392
rect 20539 11456 20855 11457
rect 20539 11392 20545 11456
rect 20609 11392 20625 11456
rect 20689 11392 20705 11456
rect 20769 11392 20785 11456
rect 20849 11392 20855 11456
rect 20539 11391 20855 11392
rect 19609 11250 19675 11253
rect 23800 11250 24600 11280
rect 19609 11248 24600 11250
rect 19609 11192 19614 11248
rect 19670 11192 24600 11248
rect 19609 11190 24600 11192
rect 19609 11187 19675 11190
rect 23800 11160 24600 11190
rect 21030 11052 21036 11116
rect 21100 11114 21106 11116
rect 21357 11114 21423 11117
rect 21100 11112 21423 11114
rect 21100 11056 21362 11112
rect 21418 11056 21423 11112
rect 21100 11054 21423 11056
rect 21100 11052 21106 11054
rect 21357 11051 21423 11054
rect 6544 10912 6860 10913
rect 6544 10848 6550 10912
rect 6614 10848 6630 10912
rect 6694 10848 6710 10912
rect 6774 10848 6790 10912
rect 6854 10848 6860 10912
rect 6544 10847 6860 10848
rect 12142 10912 12458 10913
rect 12142 10848 12148 10912
rect 12212 10848 12228 10912
rect 12292 10848 12308 10912
rect 12372 10848 12388 10912
rect 12452 10848 12458 10912
rect 12142 10847 12458 10848
rect 17740 10912 18056 10913
rect 17740 10848 17746 10912
rect 17810 10848 17826 10912
rect 17890 10848 17906 10912
rect 17970 10848 17986 10912
rect 18050 10848 18056 10912
rect 17740 10847 18056 10848
rect 19333 10706 19399 10709
rect 23800 10706 24600 10736
rect 19333 10704 24600 10706
rect 19333 10648 19338 10704
rect 19394 10648 24600 10704
rect 19333 10646 24600 10648
rect 19333 10643 19399 10646
rect 23800 10616 24600 10646
rect 3745 10368 4061 10369
rect 3745 10304 3751 10368
rect 3815 10304 3831 10368
rect 3895 10304 3911 10368
rect 3975 10304 3991 10368
rect 4055 10304 4061 10368
rect 3745 10303 4061 10304
rect 9343 10368 9659 10369
rect 9343 10304 9349 10368
rect 9413 10304 9429 10368
rect 9493 10304 9509 10368
rect 9573 10304 9589 10368
rect 9653 10304 9659 10368
rect 9343 10303 9659 10304
rect 14941 10368 15257 10369
rect 14941 10304 14947 10368
rect 15011 10304 15027 10368
rect 15091 10304 15107 10368
rect 15171 10304 15187 10368
rect 15251 10304 15257 10368
rect 14941 10303 15257 10304
rect 20539 10368 20855 10369
rect 20539 10304 20545 10368
rect 20609 10304 20625 10368
rect 20689 10304 20705 10368
rect 20769 10304 20785 10368
rect 20849 10304 20855 10368
rect 20539 10303 20855 10304
rect 16573 10162 16639 10165
rect 21265 10162 21331 10165
rect 23800 10162 24600 10192
rect 16573 10160 21331 10162
rect 16573 10104 16578 10160
rect 16634 10104 21270 10160
rect 21326 10104 21331 10160
rect 16573 10102 21331 10104
rect 16573 10099 16639 10102
rect 21265 10099 21331 10102
rect 22050 10102 24600 10162
rect 18045 10026 18111 10029
rect 18413 10026 18479 10029
rect 18965 10026 19031 10029
rect 18045 10024 18338 10026
rect 18045 9968 18050 10024
rect 18106 9968 18338 10024
rect 18045 9966 18338 9968
rect 18045 9963 18111 9966
rect 18278 9890 18338 9966
rect 18413 10024 19031 10026
rect 18413 9968 18418 10024
rect 18474 9968 18970 10024
rect 19026 9968 19031 10024
rect 18413 9966 19031 9968
rect 18413 9963 18479 9966
rect 18965 9963 19031 9966
rect 19333 10026 19399 10029
rect 22050 10026 22110 10102
rect 23800 10072 24600 10102
rect 19333 10024 22110 10026
rect 19333 9968 19338 10024
rect 19394 9968 22110 10024
rect 19333 9966 22110 9968
rect 19333 9963 19399 9966
rect 18413 9890 18479 9893
rect 18873 9892 18939 9893
rect 18278 9888 18479 9890
rect 18278 9832 18418 9888
rect 18474 9832 18479 9888
rect 18278 9830 18479 9832
rect 18413 9827 18479 9830
rect 18822 9828 18828 9892
rect 18892 9890 18939 9892
rect 19241 9890 19307 9893
rect 22461 9890 22527 9893
rect 18892 9888 18984 9890
rect 18934 9832 18984 9888
rect 18892 9830 18984 9832
rect 19241 9888 22527 9890
rect 19241 9832 19246 9888
rect 19302 9832 22466 9888
rect 22522 9832 22527 9888
rect 19241 9830 22527 9832
rect 18892 9828 18939 9830
rect 18873 9827 18939 9828
rect 19241 9827 19307 9830
rect 22461 9827 22527 9830
rect 6544 9824 6860 9825
rect 6544 9760 6550 9824
rect 6614 9760 6630 9824
rect 6694 9760 6710 9824
rect 6774 9760 6790 9824
rect 6854 9760 6860 9824
rect 6544 9759 6860 9760
rect 12142 9824 12458 9825
rect 12142 9760 12148 9824
rect 12212 9760 12228 9824
rect 12292 9760 12308 9824
rect 12372 9760 12388 9824
rect 12452 9760 12458 9824
rect 12142 9759 12458 9760
rect 17740 9824 18056 9825
rect 17740 9760 17746 9824
rect 17810 9760 17826 9824
rect 17890 9760 17906 9824
rect 17970 9760 17986 9824
rect 18050 9760 18056 9824
rect 17740 9759 18056 9760
rect 18781 9754 18847 9757
rect 22737 9754 22803 9757
rect 18781 9752 22803 9754
rect 18781 9696 18786 9752
rect 18842 9696 22742 9752
rect 22798 9696 22803 9752
rect 18781 9694 22803 9696
rect 18781 9691 18847 9694
rect 22737 9691 22803 9694
rect 19149 9618 19215 9621
rect 23800 9618 24600 9648
rect 19149 9616 24600 9618
rect 19149 9560 19154 9616
rect 19210 9560 24600 9616
rect 19149 9558 24600 9560
rect 19149 9555 19215 9558
rect 23800 9528 24600 9558
rect 19057 9482 19123 9485
rect 23105 9482 23171 9485
rect 19057 9480 23171 9482
rect 19057 9424 19062 9480
rect 19118 9424 23110 9480
rect 23166 9424 23171 9480
rect 19057 9422 23171 9424
rect 19057 9419 19123 9422
rect 23105 9419 23171 9422
rect 3745 9280 4061 9281
rect 0 9210 800 9240
rect 3745 9216 3751 9280
rect 3815 9216 3831 9280
rect 3895 9216 3911 9280
rect 3975 9216 3991 9280
rect 4055 9216 4061 9280
rect 3745 9215 4061 9216
rect 9343 9280 9659 9281
rect 9343 9216 9349 9280
rect 9413 9216 9429 9280
rect 9493 9216 9509 9280
rect 9573 9216 9589 9280
rect 9653 9216 9659 9280
rect 9343 9215 9659 9216
rect 14941 9280 15257 9281
rect 14941 9216 14947 9280
rect 15011 9216 15027 9280
rect 15091 9216 15107 9280
rect 15171 9216 15187 9280
rect 15251 9216 15257 9280
rect 14941 9215 15257 9216
rect 20539 9280 20855 9281
rect 20539 9216 20545 9280
rect 20609 9216 20625 9280
rect 20689 9216 20705 9280
rect 20769 9216 20785 9280
rect 20849 9216 20855 9280
rect 20539 9215 20855 9216
rect 1393 9210 1459 9213
rect 0 9208 1459 9210
rect 0 9152 1398 9208
rect 1454 9152 1459 9208
rect 0 9150 1459 9152
rect 0 9120 800 9150
rect 1393 9147 1459 9150
rect 19609 9074 19675 9077
rect 23800 9074 24600 9104
rect 19609 9072 24600 9074
rect 19609 9016 19614 9072
rect 19670 9016 24600 9072
rect 19609 9014 24600 9016
rect 19609 9011 19675 9014
rect 23800 8984 24600 9014
rect 18045 8938 18111 8941
rect 20713 8938 20779 8941
rect 18045 8936 20779 8938
rect 18045 8880 18050 8936
rect 18106 8880 20718 8936
rect 20774 8880 20779 8936
rect 18045 8878 20779 8880
rect 18045 8875 18111 8878
rect 20713 8875 20779 8878
rect 20161 8802 20227 8805
rect 22369 8802 22435 8805
rect 20161 8800 22435 8802
rect 20161 8744 20166 8800
rect 20222 8744 22374 8800
rect 22430 8744 22435 8800
rect 20161 8742 22435 8744
rect 20161 8739 20227 8742
rect 22369 8739 22435 8742
rect 6544 8736 6860 8737
rect 6544 8672 6550 8736
rect 6614 8672 6630 8736
rect 6694 8672 6710 8736
rect 6774 8672 6790 8736
rect 6854 8672 6860 8736
rect 6544 8671 6860 8672
rect 12142 8736 12458 8737
rect 12142 8672 12148 8736
rect 12212 8672 12228 8736
rect 12292 8672 12308 8736
rect 12372 8672 12388 8736
rect 12452 8672 12458 8736
rect 12142 8671 12458 8672
rect 17740 8736 18056 8737
rect 17740 8672 17746 8736
rect 17810 8672 17826 8736
rect 17890 8672 17906 8736
rect 17970 8672 17986 8736
rect 18050 8672 18056 8736
rect 17740 8671 18056 8672
rect 2957 8530 3023 8533
rect 4889 8530 4955 8533
rect 2957 8528 4955 8530
rect 2957 8472 2962 8528
rect 3018 8472 4894 8528
rect 4950 8472 4955 8528
rect 2957 8470 4955 8472
rect 2957 8467 3023 8470
rect 4889 8467 4955 8470
rect 19333 8530 19399 8533
rect 22645 8530 22711 8533
rect 23800 8530 24600 8560
rect 19333 8528 24600 8530
rect 19333 8472 19338 8528
rect 19394 8472 22650 8528
rect 22706 8472 24600 8528
rect 19333 8470 24600 8472
rect 19333 8467 19399 8470
rect 22645 8467 22711 8470
rect 23800 8440 24600 8470
rect 16481 8394 16547 8397
rect 21173 8394 21239 8397
rect 16481 8392 21239 8394
rect 16481 8336 16486 8392
rect 16542 8336 21178 8392
rect 21234 8336 21239 8392
rect 16481 8334 21239 8336
rect 16481 8331 16547 8334
rect 21173 8331 21239 8334
rect 3745 8192 4061 8193
rect 3745 8128 3751 8192
rect 3815 8128 3831 8192
rect 3895 8128 3911 8192
rect 3975 8128 3991 8192
rect 4055 8128 4061 8192
rect 3745 8127 4061 8128
rect 9343 8192 9659 8193
rect 9343 8128 9349 8192
rect 9413 8128 9429 8192
rect 9493 8128 9509 8192
rect 9573 8128 9589 8192
rect 9653 8128 9659 8192
rect 9343 8127 9659 8128
rect 14941 8192 15257 8193
rect 14941 8128 14947 8192
rect 15011 8128 15027 8192
rect 15091 8128 15107 8192
rect 15171 8128 15187 8192
rect 15251 8128 15257 8192
rect 14941 8127 15257 8128
rect 20539 8192 20855 8193
rect 20539 8128 20545 8192
rect 20609 8128 20625 8192
rect 20689 8128 20705 8192
rect 20769 8128 20785 8192
rect 20849 8128 20855 8192
rect 20539 8127 20855 8128
rect 23013 7986 23079 7989
rect 23800 7986 24600 8016
rect 23013 7984 24600 7986
rect 23013 7928 23018 7984
rect 23074 7928 24600 7984
rect 23013 7926 24600 7928
rect 23013 7923 23079 7926
rect 23800 7896 24600 7926
rect 6544 7648 6860 7649
rect 6544 7584 6550 7648
rect 6614 7584 6630 7648
rect 6694 7584 6710 7648
rect 6774 7584 6790 7648
rect 6854 7584 6860 7648
rect 6544 7583 6860 7584
rect 12142 7648 12458 7649
rect 12142 7584 12148 7648
rect 12212 7584 12228 7648
rect 12292 7584 12308 7648
rect 12372 7584 12388 7648
rect 12452 7584 12458 7648
rect 12142 7583 12458 7584
rect 17740 7648 18056 7649
rect 17740 7584 17746 7648
rect 17810 7584 17826 7648
rect 17890 7584 17906 7648
rect 17970 7584 17986 7648
rect 18050 7584 18056 7648
rect 17740 7583 18056 7584
rect 14457 7442 14523 7445
rect 21541 7444 21607 7445
rect 21214 7442 21220 7444
rect 14457 7440 21220 7442
rect 14457 7384 14462 7440
rect 14518 7384 21220 7440
rect 14457 7382 21220 7384
rect 14457 7379 14523 7382
rect 21214 7380 21220 7382
rect 21284 7380 21290 7444
rect 21541 7442 21588 7444
rect 21496 7440 21588 7442
rect 21496 7384 21546 7440
rect 21496 7382 21588 7384
rect 21541 7380 21588 7382
rect 21652 7380 21658 7444
rect 23013 7442 23079 7445
rect 23800 7442 24600 7472
rect 23013 7440 24600 7442
rect 23013 7384 23018 7440
rect 23074 7384 24600 7440
rect 23013 7382 24600 7384
rect 21541 7379 21607 7380
rect 23013 7379 23079 7382
rect 23800 7352 24600 7382
rect 16941 7306 17007 7309
rect 21030 7306 21036 7308
rect 16941 7304 21036 7306
rect 16941 7248 16946 7304
rect 17002 7248 21036 7304
rect 16941 7246 21036 7248
rect 16941 7243 17007 7246
rect 21030 7244 21036 7246
rect 21100 7244 21106 7308
rect 19517 7172 19583 7173
rect 19517 7170 19564 7172
rect 19472 7168 19564 7170
rect 19472 7112 19522 7168
rect 19472 7110 19564 7112
rect 19517 7108 19564 7110
rect 19628 7108 19634 7172
rect 19517 7107 19583 7108
rect 3745 7104 4061 7105
rect 3745 7040 3751 7104
rect 3815 7040 3831 7104
rect 3895 7040 3911 7104
rect 3975 7040 3991 7104
rect 4055 7040 4061 7104
rect 3745 7039 4061 7040
rect 9343 7104 9659 7105
rect 9343 7040 9349 7104
rect 9413 7040 9429 7104
rect 9493 7040 9509 7104
rect 9573 7040 9589 7104
rect 9653 7040 9659 7104
rect 9343 7039 9659 7040
rect 14941 7104 15257 7105
rect 14941 7040 14947 7104
rect 15011 7040 15027 7104
rect 15091 7040 15107 7104
rect 15171 7040 15187 7104
rect 15251 7040 15257 7104
rect 14941 7039 15257 7040
rect 20539 7104 20855 7105
rect 20539 7040 20545 7104
rect 20609 7040 20625 7104
rect 20689 7040 20705 7104
rect 20769 7040 20785 7104
rect 20849 7040 20855 7104
rect 20539 7039 20855 7040
rect 19425 7036 19491 7037
rect 19374 6972 19380 7036
rect 19444 7034 19491 7036
rect 19793 7034 19859 7037
rect 19977 7034 20043 7037
rect 19444 7032 19536 7034
rect 19486 6976 19536 7032
rect 19444 6974 19536 6976
rect 19793 7032 20043 7034
rect 19793 6976 19798 7032
rect 19854 6976 19982 7032
rect 20038 6976 20043 7032
rect 19793 6974 20043 6976
rect 19444 6972 19491 6974
rect 19425 6971 19491 6972
rect 19793 6971 19859 6974
rect 19977 6971 20043 6974
rect 23013 6898 23079 6901
rect 23800 6898 24600 6928
rect 23013 6896 24600 6898
rect 23013 6840 23018 6896
rect 23074 6840 24600 6896
rect 23013 6838 24600 6840
rect 23013 6835 23079 6838
rect 23800 6808 24600 6838
rect 17217 6762 17283 6765
rect 22461 6762 22527 6765
rect 17217 6760 22527 6762
rect 17217 6704 17222 6760
rect 17278 6704 22466 6760
rect 22522 6704 22527 6760
rect 17217 6702 22527 6704
rect 17217 6699 17283 6702
rect 22461 6699 22527 6702
rect 21265 6628 21331 6629
rect 21214 6564 21220 6628
rect 21284 6626 21331 6628
rect 21909 6626 21975 6629
rect 21284 6624 21975 6626
rect 21326 6568 21914 6624
rect 21970 6568 21975 6624
rect 21284 6566 21975 6568
rect 21284 6564 21331 6566
rect 21265 6563 21331 6564
rect 21909 6563 21975 6566
rect 6544 6560 6860 6561
rect 6544 6496 6550 6560
rect 6614 6496 6630 6560
rect 6694 6496 6710 6560
rect 6774 6496 6790 6560
rect 6854 6496 6860 6560
rect 6544 6495 6860 6496
rect 12142 6560 12458 6561
rect 12142 6496 12148 6560
rect 12212 6496 12228 6560
rect 12292 6496 12308 6560
rect 12372 6496 12388 6560
rect 12452 6496 12458 6560
rect 12142 6495 12458 6496
rect 17740 6560 18056 6561
rect 17740 6496 17746 6560
rect 17810 6496 17826 6560
rect 17890 6496 17906 6560
rect 17970 6496 17986 6560
rect 18050 6496 18056 6560
rect 17740 6495 18056 6496
rect 19425 6490 19491 6493
rect 19742 6490 19748 6492
rect 19425 6488 19748 6490
rect 19425 6432 19430 6488
rect 19486 6432 19748 6488
rect 19425 6430 19748 6432
rect 19425 6427 19491 6430
rect 19742 6428 19748 6430
rect 19812 6428 19818 6492
rect 19885 6490 19951 6493
rect 22093 6490 22159 6493
rect 19885 6488 22159 6490
rect 19885 6432 19890 6488
rect 19946 6432 22098 6488
rect 22154 6432 22159 6488
rect 19885 6430 22159 6432
rect 19885 6427 19951 6430
rect 22093 6427 22159 6430
rect 16389 6354 16455 6357
rect 17125 6354 17191 6357
rect 21449 6354 21515 6357
rect 16389 6352 21515 6354
rect 16389 6296 16394 6352
rect 16450 6296 17130 6352
rect 17186 6296 21454 6352
rect 21510 6296 21515 6352
rect 16389 6294 21515 6296
rect 16389 6291 16455 6294
rect 17125 6291 17191 6294
rect 21449 6291 21515 6294
rect 22829 6354 22895 6357
rect 23800 6354 24600 6384
rect 22829 6352 24600 6354
rect 22829 6296 22834 6352
rect 22890 6296 24600 6352
rect 22829 6294 24600 6296
rect 22829 6291 22895 6294
rect 23800 6264 24600 6294
rect 14365 6218 14431 6221
rect 17033 6218 17099 6221
rect 23381 6218 23447 6221
rect 14365 6216 23447 6218
rect 14365 6160 14370 6216
rect 14426 6160 17038 6216
rect 17094 6160 23386 6216
rect 23442 6160 23447 6216
rect 14365 6158 23447 6160
rect 14365 6155 14431 6158
rect 17033 6155 17099 6158
rect 23381 6155 23447 6158
rect 19425 6084 19491 6085
rect 19374 6082 19380 6084
rect 19334 6022 19380 6082
rect 19444 6080 19491 6084
rect 19486 6024 19491 6080
rect 19374 6020 19380 6022
rect 19444 6020 19491 6024
rect 19558 6020 19564 6084
rect 19628 6082 19634 6084
rect 19793 6082 19859 6085
rect 19628 6080 19859 6082
rect 19628 6024 19798 6080
rect 19854 6024 19859 6080
rect 19628 6022 19859 6024
rect 19628 6020 19634 6022
rect 19425 6019 19491 6020
rect 19793 6019 19859 6022
rect 21265 6082 21331 6085
rect 21541 6082 21607 6085
rect 21265 6080 21607 6082
rect 21265 6024 21270 6080
rect 21326 6024 21546 6080
rect 21602 6024 21607 6080
rect 21265 6022 21607 6024
rect 21265 6019 21331 6022
rect 21541 6019 21607 6022
rect 3745 6016 4061 6017
rect 3745 5952 3751 6016
rect 3815 5952 3831 6016
rect 3895 5952 3911 6016
rect 3975 5952 3991 6016
rect 4055 5952 4061 6016
rect 3745 5951 4061 5952
rect 9343 6016 9659 6017
rect 9343 5952 9349 6016
rect 9413 5952 9429 6016
rect 9493 5952 9509 6016
rect 9573 5952 9589 6016
rect 9653 5952 9659 6016
rect 9343 5951 9659 5952
rect 14941 6016 15257 6017
rect 14941 5952 14947 6016
rect 15011 5952 15027 6016
rect 15091 5952 15107 6016
rect 15171 5952 15187 6016
rect 15251 5952 15257 6016
rect 14941 5951 15257 5952
rect 20539 6016 20855 6017
rect 20539 5952 20545 6016
rect 20609 5952 20625 6016
rect 20689 5952 20705 6016
rect 20769 5952 20785 6016
rect 20849 5952 20855 6016
rect 20539 5951 20855 5952
rect 23013 5810 23079 5813
rect 23800 5810 24600 5840
rect 23013 5808 24600 5810
rect 23013 5752 23018 5808
rect 23074 5752 24600 5808
rect 23013 5750 24600 5752
rect 23013 5747 23079 5750
rect 23800 5720 24600 5750
rect 20069 5674 20135 5677
rect 20437 5674 20503 5677
rect 20069 5672 20503 5674
rect 20069 5616 20074 5672
rect 20130 5616 20442 5672
rect 20498 5616 20503 5672
rect 20069 5614 20503 5616
rect 20069 5611 20135 5614
rect 20437 5611 20503 5614
rect 6544 5472 6860 5473
rect 6544 5408 6550 5472
rect 6614 5408 6630 5472
rect 6694 5408 6710 5472
rect 6774 5408 6790 5472
rect 6854 5408 6860 5472
rect 6544 5407 6860 5408
rect 12142 5472 12458 5473
rect 12142 5408 12148 5472
rect 12212 5408 12228 5472
rect 12292 5408 12308 5472
rect 12372 5408 12388 5472
rect 12452 5408 12458 5472
rect 12142 5407 12458 5408
rect 17740 5472 18056 5473
rect 17740 5408 17746 5472
rect 17810 5408 17826 5472
rect 17890 5408 17906 5472
rect 17970 5408 17986 5472
rect 18050 5408 18056 5472
rect 17740 5407 18056 5408
rect 23013 5266 23079 5269
rect 23800 5266 24600 5296
rect 23013 5264 24600 5266
rect 23013 5208 23018 5264
rect 23074 5208 24600 5264
rect 23013 5206 24600 5208
rect 23013 5203 23079 5206
rect 23800 5176 24600 5206
rect 3745 4928 4061 4929
rect 3745 4864 3751 4928
rect 3815 4864 3831 4928
rect 3895 4864 3911 4928
rect 3975 4864 3991 4928
rect 4055 4864 4061 4928
rect 3745 4863 4061 4864
rect 9343 4928 9659 4929
rect 9343 4864 9349 4928
rect 9413 4864 9429 4928
rect 9493 4864 9509 4928
rect 9573 4864 9589 4928
rect 9653 4864 9659 4928
rect 9343 4863 9659 4864
rect 14941 4928 15257 4929
rect 14941 4864 14947 4928
rect 15011 4864 15027 4928
rect 15091 4864 15107 4928
rect 15171 4864 15187 4928
rect 15251 4864 15257 4928
rect 14941 4863 15257 4864
rect 20539 4928 20855 4929
rect 20539 4864 20545 4928
rect 20609 4864 20625 4928
rect 20689 4864 20705 4928
rect 20769 4864 20785 4928
rect 20849 4864 20855 4928
rect 20539 4863 20855 4864
rect 19609 4858 19675 4861
rect 19742 4858 19748 4860
rect 19609 4856 19748 4858
rect 19609 4800 19614 4856
rect 19670 4800 19748 4856
rect 19609 4798 19748 4800
rect 19609 4795 19675 4798
rect 19742 4796 19748 4798
rect 19812 4796 19818 4860
rect 19190 4660 19196 4724
rect 19260 4722 19266 4724
rect 20529 4722 20595 4725
rect 19260 4720 20595 4722
rect 19260 4664 20534 4720
rect 20590 4664 20595 4720
rect 19260 4662 20595 4664
rect 19260 4660 19266 4662
rect 20529 4659 20595 4662
rect 23013 4722 23079 4725
rect 23800 4722 24600 4752
rect 23013 4720 24600 4722
rect 23013 4664 23018 4720
rect 23074 4664 24600 4720
rect 23013 4662 24600 4664
rect 23013 4659 23079 4662
rect 23800 4632 24600 4662
rect 21214 4388 21220 4452
rect 21284 4450 21290 4452
rect 21357 4450 21423 4453
rect 21284 4448 21423 4450
rect 21284 4392 21362 4448
rect 21418 4392 21423 4448
rect 21284 4390 21423 4392
rect 21284 4388 21290 4390
rect 21357 4387 21423 4390
rect 6544 4384 6860 4385
rect 6544 4320 6550 4384
rect 6614 4320 6630 4384
rect 6694 4320 6710 4384
rect 6774 4320 6790 4384
rect 6854 4320 6860 4384
rect 6544 4319 6860 4320
rect 12142 4384 12458 4385
rect 12142 4320 12148 4384
rect 12212 4320 12228 4384
rect 12292 4320 12308 4384
rect 12372 4320 12388 4384
rect 12452 4320 12458 4384
rect 12142 4319 12458 4320
rect 17740 4384 18056 4385
rect 17740 4320 17746 4384
rect 17810 4320 17826 4384
rect 17890 4320 17906 4384
rect 17970 4320 17986 4384
rect 18050 4320 18056 4384
rect 17740 4319 18056 4320
rect 13721 4178 13787 4181
rect 21449 4178 21515 4181
rect 13721 4176 21515 4178
rect 13721 4120 13726 4176
rect 13782 4120 21454 4176
rect 21510 4120 21515 4176
rect 13721 4118 21515 4120
rect 13721 4115 13787 4118
rect 21449 4115 21515 4118
rect 23013 4178 23079 4181
rect 23800 4178 24600 4208
rect 23013 4176 24600 4178
rect 23013 4120 23018 4176
rect 23074 4120 24600 4176
rect 23013 4118 24600 4120
rect 23013 4115 23079 4118
rect 23800 4088 24600 4118
rect 3745 3840 4061 3841
rect 3745 3776 3751 3840
rect 3815 3776 3831 3840
rect 3895 3776 3911 3840
rect 3975 3776 3991 3840
rect 4055 3776 4061 3840
rect 3745 3775 4061 3776
rect 9343 3840 9659 3841
rect 9343 3776 9349 3840
rect 9413 3776 9429 3840
rect 9493 3776 9509 3840
rect 9573 3776 9589 3840
rect 9653 3776 9659 3840
rect 9343 3775 9659 3776
rect 14941 3840 15257 3841
rect 14941 3776 14947 3840
rect 15011 3776 15027 3840
rect 15091 3776 15107 3840
rect 15171 3776 15187 3840
rect 15251 3776 15257 3840
rect 14941 3775 15257 3776
rect 20539 3840 20855 3841
rect 20539 3776 20545 3840
rect 20609 3776 20625 3840
rect 20689 3776 20705 3840
rect 20769 3776 20785 3840
rect 20849 3776 20855 3840
rect 20539 3775 20855 3776
rect 15561 3634 15627 3637
rect 22553 3634 22619 3637
rect 15561 3632 22619 3634
rect 15561 3576 15566 3632
rect 15622 3576 22558 3632
rect 22614 3576 22619 3632
rect 15561 3574 22619 3576
rect 15561 3571 15627 3574
rect 22553 3571 22619 3574
rect 23013 3634 23079 3637
rect 23800 3634 24600 3664
rect 23013 3632 24600 3634
rect 23013 3576 23018 3632
rect 23074 3576 24600 3632
rect 23013 3574 24600 3576
rect 23013 3571 23079 3574
rect 23800 3544 24600 3574
rect 16297 3498 16363 3501
rect 22369 3498 22435 3501
rect 16297 3496 22435 3498
rect 16297 3440 16302 3496
rect 16358 3440 22374 3496
rect 22430 3440 22435 3496
rect 16297 3438 22435 3440
rect 16297 3435 16363 3438
rect 22369 3435 22435 3438
rect 6544 3296 6860 3297
rect 6544 3232 6550 3296
rect 6614 3232 6630 3296
rect 6694 3232 6710 3296
rect 6774 3232 6790 3296
rect 6854 3232 6860 3296
rect 6544 3231 6860 3232
rect 12142 3296 12458 3297
rect 12142 3232 12148 3296
rect 12212 3232 12228 3296
rect 12292 3232 12308 3296
rect 12372 3232 12388 3296
rect 12452 3232 12458 3296
rect 12142 3231 12458 3232
rect 17740 3296 18056 3297
rect 17740 3232 17746 3296
rect 17810 3232 17826 3296
rect 17890 3232 17906 3296
rect 17970 3232 17986 3296
rect 18050 3232 18056 3296
rect 17740 3231 18056 3232
rect 0 3090 800 3120
rect 1393 3090 1459 3093
rect 0 3088 1459 3090
rect 0 3032 1398 3088
rect 1454 3032 1459 3088
rect 0 3030 1459 3032
rect 0 3000 800 3030
rect 1393 3027 1459 3030
rect 16665 3090 16731 3093
rect 19701 3090 19767 3093
rect 20989 3090 21055 3093
rect 16665 3088 21055 3090
rect 16665 3032 16670 3088
rect 16726 3032 19706 3088
rect 19762 3032 20994 3088
rect 21050 3032 21055 3088
rect 16665 3030 21055 3032
rect 16665 3027 16731 3030
rect 19701 3027 19767 3030
rect 20989 3027 21055 3030
rect 23013 3090 23079 3093
rect 23800 3090 24600 3120
rect 23013 3088 24600 3090
rect 23013 3032 23018 3088
rect 23074 3032 24600 3088
rect 23013 3030 24600 3032
rect 23013 3027 23079 3030
rect 23800 3000 24600 3030
rect 3745 2752 4061 2753
rect 3745 2688 3751 2752
rect 3815 2688 3831 2752
rect 3895 2688 3911 2752
rect 3975 2688 3991 2752
rect 4055 2688 4061 2752
rect 3745 2687 4061 2688
rect 9343 2752 9659 2753
rect 9343 2688 9349 2752
rect 9413 2688 9429 2752
rect 9493 2688 9509 2752
rect 9573 2688 9589 2752
rect 9653 2688 9659 2752
rect 9343 2687 9659 2688
rect 14941 2752 15257 2753
rect 14941 2688 14947 2752
rect 15011 2688 15027 2752
rect 15091 2688 15107 2752
rect 15171 2688 15187 2752
rect 15251 2688 15257 2752
rect 14941 2687 15257 2688
rect 20539 2752 20855 2753
rect 20539 2688 20545 2752
rect 20609 2688 20625 2752
rect 20689 2688 20705 2752
rect 20769 2688 20785 2752
rect 20849 2688 20855 2752
rect 20539 2687 20855 2688
rect 23013 2546 23079 2549
rect 23800 2546 24600 2576
rect 23013 2544 24600 2546
rect 23013 2488 23018 2544
rect 23074 2488 24600 2544
rect 23013 2486 24600 2488
rect 23013 2483 23079 2486
rect 23800 2456 24600 2486
rect 6544 2208 6860 2209
rect 6544 2144 6550 2208
rect 6614 2144 6630 2208
rect 6694 2144 6710 2208
rect 6774 2144 6790 2208
rect 6854 2144 6860 2208
rect 6544 2143 6860 2144
rect 12142 2208 12458 2209
rect 12142 2144 12148 2208
rect 12212 2144 12228 2208
rect 12292 2144 12308 2208
rect 12372 2144 12388 2208
rect 12452 2144 12458 2208
rect 12142 2143 12458 2144
rect 17740 2208 18056 2209
rect 17740 2144 17746 2208
rect 17810 2144 17826 2208
rect 17890 2144 17906 2208
rect 17970 2144 17986 2208
rect 18050 2144 18056 2208
rect 17740 2143 18056 2144
<< via3 >>
rect 3751 22332 3815 22336
rect 3751 22276 3755 22332
rect 3755 22276 3811 22332
rect 3811 22276 3815 22332
rect 3751 22272 3815 22276
rect 3831 22332 3895 22336
rect 3831 22276 3835 22332
rect 3835 22276 3891 22332
rect 3891 22276 3895 22332
rect 3831 22272 3895 22276
rect 3911 22332 3975 22336
rect 3911 22276 3915 22332
rect 3915 22276 3971 22332
rect 3971 22276 3975 22332
rect 3911 22272 3975 22276
rect 3991 22332 4055 22336
rect 3991 22276 3995 22332
rect 3995 22276 4051 22332
rect 4051 22276 4055 22332
rect 3991 22272 4055 22276
rect 9349 22332 9413 22336
rect 9349 22276 9353 22332
rect 9353 22276 9409 22332
rect 9409 22276 9413 22332
rect 9349 22272 9413 22276
rect 9429 22332 9493 22336
rect 9429 22276 9433 22332
rect 9433 22276 9489 22332
rect 9489 22276 9493 22332
rect 9429 22272 9493 22276
rect 9509 22332 9573 22336
rect 9509 22276 9513 22332
rect 9513 22276 9569 22332
rect 9569 22276 9573 22332
rect 9509 22272 9573 22276
rect 9589 22332 9653 22336
rect 9589 22276 9593 22332
rect 9593 22276 9649 22332
rect 9649 22276 9653 22332
rect 9589 22272 9653 22276
rect 14947 22332 15011 22336
rect 14947 22276 14951 22332
rect 14951 22276 15007 22332
rect 15007 22276 15011 22332
rect 14947 22272 15011 22276
rect 15027 22332 15091 22336
rect 15027 22276 15031 22332
rect 15031 22276 15087 22332
rect 15087 22276 15091 22332
rect 15027 22272 15091 22276
rect 15107 22332 15171 22336
rect 15107 22276 15111 22332
rect 15111 22276 15167 22332
rect 15167 22276 15171 22332
rect 15107 22272 15171 22276
rect 15187 22332 15251 22336
rect 15187 22276 15191 22332
rect 15191 22276 15247 22332
rect 15247 22276 15251 22332
rect 15187 22272 15251 22276
rect 20545 22332 20609 22336
rect 20545 22276 20549 22332
rect 20549 22276 20605 22332
rect 20605 22276 20609 22332
rect 20545 22272 20609 22276
rect 20625 22332 20689 22336
rect 20625 22276 20629 22332
rect 20629 22276 20685 22332
rect 20685 22276 20689 22332
rect 20625 22272 20689 22276
rect 20705 22332 20769 22336
rect 20705 22276 20709 22332
rect 20709 22276 20765 22332
rect 20765 22276 20769 22332
rect 20705 22272 20769 22276
rect 20785 22332 20849 22336
rect 20785 22276 20789 22332
rect 20789 22276 20845 22332
rect 20845 22276 20849 22332
rect 20785 22272 20849 22276
rect 16436 22068 16500 22132
rect 6550 21788 6614 21792
rect 6550 21732 6554 21788
rect 6554 21732 6610 21788
rect 6610 21732 6614 21788
rect 6550 21728 6614 21732
rect 6630 21788 6694 21792
rect 6630 21732 6634 21788
rect 6634 21732 6690 21788
rect 6690 21732 6694 21788
rect 6630 21728 6694 21732
rect 6710 21788 6774 21792
rect 6710 21732 6714 21788
rect 6714 21732 6770 21788
rect 6770 21732 6774 21788
rect 6710 21728 6774 21732
rect 6790 21788 6854 21792
rect 6790 21732 6794 21788
rect 6794 21732 6850 21788
rect 6850 21732 6854 21788
rect 6790 21728 6854 21732
rect 12148 21788 12212 21792
rect 12148 21732 12152 21788
rect 12152 21732 12208 21788
rect 12208 21732 12212 21788
rect 12148 21728 12212 21732
rect 12228 21788 12292 21792
rect 12228 21732 12232 21788
rect 12232 21732 12288 21788
rect 12288 21732 12292 21788
rect 12228 21728 12292 21732
rect 12308 21788 12372 21792
rect 12308 21732 12312 21788
rect 12312 21732 12368 21788
rect 12368 21732 12372 21788
rect 12308 21728 12372 21732
rect 12388 21788 12452 21792
rect 12388 21732 12392 21788
rect 12392 21732 12448 21788
rect 12448 21732 12452 21788
rect 12388 21728 12452 21732
rect 17746 21788 17810 21792
rect 17746 21732 17750 21788
rect 17750 21732 17806 21788
rect 17806 21732 17810 21788
rect 17746 21728 17810 21732
rect 17826 21788 17890 21792
rect 17826 21732 17830 21788
rect 17830 21732 17886 21788
rect 17886 21732 17890 21788
rect 17826 21728 17890 21732
rect 17906 21788 17970 21792
rect 17906 21732 17910 21788
rect 17910 21732 17966 21788
rect 17966 21732 17970 21788
rect 17906 21728 17970 21732
rect 17986 21788 18050 21792
rect 17986 21732 17990 21788
rect 17990 21732 18046 21788
rect 18046 21732 18050 21788
rect 17986 21728 18050 21732
rect 16436 21524 16500 21588
rect 3751 21244 3815 21248
rect 3751 21188 3755 21244
rect 3755 21188 3811 21244
rect 3811 21188 3815 21244
rect 3751 21184 3815 21188
rect 3831 21244 3895 21248
rect 3831 21188 3835 21244
rect 3835 21188 3891 21244
rect 3891 21188 3895 21244
rect 3831 21184 3895 21188
rect 3911 21244 3975 21248
rect 3911 21188 3915 21244
rect 3915 21188 3971 21244
rect 3971 21188 3975 21244
rect 3911 21184 3975 21188
rect 3991 21244 4055 21248
rect 3991 21188 3995 21244
rect 3995 21188 4051 21244
rect 4051 21188 4055 21244
rect 3991 21184 4055 21188
rect 9349 21244 9413 21248
rect 9349 21188 9353 21244
rect 9353 21188 9409 21244
rect 9409 21188 9413 21244
rect 9349 21184 9413 21188
rect 9429 21244 9493 21248
rect 9429 21188 9433 21244
rect 9433 21188 9489 21244
rect 9489 21188 9493 21244
rect 9429 21184 9493 21188
rect 9509 21244 9573 21248
rect 9509 21188 9513 21244
rect 9513 21188 9569 21244
rect 9569 21188 9573 21244
rect 9509 21184 9573 21188
rect 9589 21244 9653 21248
rect 9589 21188 9593 21244
rect 9593 21188 9649 21244
rect 9649 21188 9653 21244
rect 9589 21184 9653 21188
rect 13860 21252 13924 21316
rect 14947 21244 15011 21248
rect 14947 21188 14951 21244
rect 14951 21188 15007 21244
rect 15007 21188 15011 21244
rect 14947 21184 15011 21188
rect 15027 21244 15091 21248
rect 15027 21188 15031 21244
rect 15031 21188 15087 21244
rect 15087 21188 15091 21244
rect 15027 21184 15091 21188
rect 15107 21244 15171 21248
rect 15107 21188 15111 21244
rect 15111 21188 15167 21244
rect 15167 21188 15171 21244
rect 15107 21184 15171 21188
rect 15187 21244 15251 21248
rect 15187 21188 15191 21244
rect 15191 21188 15247 21244
rect 15247 21188 15251 21244
rect 15187 21184 15251 21188
rect 20545 21244 20609 21248
rect 20545 21188 20549 21244
rect 20549 21188 20605 21244
rect 20605 21188 20609 21244
rect 20545 21184 20609 21188
rect 20625 21244 20689 21248
rect 20625 21188 20629 21244
rect 20629 21188 20685 21244
rect 20685 21188 20689 21244
rect 20625 21184 20689 21188
rect 20705 21244 20769 21248
rect 20705 21188 20709 21244
rect 20709 21188 20765 21244
rect 20765 21188 20769 21244
rect 20705 21184 20769 21188
rect 20785 21244 20849 21248
rect 20785 21188 20789 21244
rect 20789 21188 20845 21244
rect 20845 21188 20849 21244
rect 20785 21184 20849 21188
rect 21036 20708 21100 20772
rect 6550 20700 6614 20704
rect 6550 20644 6554 20700
rect 6554 20644 6610 20700
rect 6610 20644 6614 20700
rect 6550 20640 6614 20644
rect 6630 20700 6694 20704
rect 6630 20644 6634 20700
rect 6634 20644 6690 20700
rect 6690 20644 6694 20700
rect 6630 20640 6694 20644
rect 6710 20700 6774 20704
rect 6710 20644 6714 20700
rect 6714 20644 6770 20700
rect 6770 20644 6774 20700
rect 6710 20640 6774 20644
rect 6790 20700 6854 20704
rect 6790 20644 6794 20700
rect 6794 20644 6850 20700
rect 6850 20644 6854 20700
rect 6790 20640 6854 20644
rect 12148 20700 12212 20704
rect 12148 20644 12152 20700
rect 12152 20644 12208 20700
rect 12208 20644 12212 20700
rect 12148 20640 12212 20644
rect 12228 20700 12292 20704
rect 12228 20644 12232 20700
rect 12232 20644 12288 20700
rect 12288 20644 12292 20700
rect 12228 20640 12292 20644
rect 12308 20700 12372 20704
rect 12308 20644 12312 20700
rect 12312 20644 12368 20700
rect 12368 20644 12372 20700
rect 12308 20640 12372 20644
rect 12388 20700 12452 20704
rect 12388 20644 12392 20700
rect 12392 20644 12448 20700
rect 12448 20644 12452 20700
rect 12388 20640 12452 20644
rect 17746 20700 17810 20704
rect 17746 20644 17750 20700
rect 17750 20644 17806 20700
rect 17806 20644 17810 20700
rect 17746 20640 17810 20644
rect 17826 20700 17890 20704
rect 17826 20644 17830 20700
rect 17830 20644 17886 20700
rect 17886 20644 17890 20700
rect 17826 20640 17890 20644
rect 17906 20700 17970 20704
rect 17906 20644 17910 20700
rect 17910 20644 17966 20700
rect 17966 20644 17970 20700
rect 17906 20640 17970 20644
rect 17986 20700 18050 20704
rect 17986 20644 17990 20700
rect 17990 20644 18046 20700
rect 18046 20644 18050 20700
rect 17986 20640 18050 20644
rect 3751 20156 3815 20160
rect 3751 20100 3755 20156
rect 3755 20100 3811 20156
rect 3811 20100 3815 20156
rect 3751 20096 3815 20100
rect 3831 20156 3895 20160
rect 3831 20100 3835 20156
rect 3835 20100 3891 20156
rect 3891 20100 3895 20156
rect 3831 20096 3895 20100
rect 3911 20156 3975 20160
rect 3911 20100 3915 20156
rect 3915 20100 3971 20156
rect 3971 20100 3975 20156
rect 3911 20096 3975 20100
rect 3991 20156 4055 20160
rect 3991 20100 3995 20156
rect 3995 20100 4051 20156
rect 4051 20100 4055 20156
rect 3991 20096 4055 20100
rect 9349 20156 9413 20160
rect 9349 20100 9353 20156
rect 9353 20100 9409 20156
rect 9409 20100 9413 20156
rect 9349 20096 9413 20100
rect 9429 20156 9493 20160
rect 9429 20100 9433 20156
rect 9433 20100 9489 20156
rect 9489 20100 9493 20156
rect 9429 20096 9493 20100
rect 9509 20156 9573 20160
rect 9509 20100 9513 20156
rect 9513 20100 9569 20156
rect 9569 20100 9573 20156
rect 9509 20096 9573 20100
rect 9589 20156 9653 20160
rect 9589 20100 9593 20156
rect 9593 20100 9649 20156
rect 9649 20100 9653 20156
rect 9589 20096 9653 20100
rect 14947 20156 15011 20160
rect 14947 20100 14951 20156
rect 14951 20100 15007 20156
rect 15007 20100 15011 20156
rect 14947 20096 15011 20100
rect 15027 20156 15091 20160
rect 15027 20100 15031 20156
rect 15031 20100 15087 20156
rect 15087 20100 15091 20156
rect 15027 20096 15091 20100
rect 15107 20156 15171 20160
rect 15107 20100 15111 20156
rect 15111 20100 15167 20156
rect 15167 20100 15171 20156
rect 15107 20096 15171 20100
rect 15187 20156 15251 20160
rect 15187 20100 15191 20156
rect 15191 20100 15247 20156
rect 15247 20100 15251 20156
rect 15187 20096 15251 20100
rect 20545 20156 20609 20160
rect 20545 20100 20549 20156
rect 20549 20100 20605 20156
rect 20605 20100 20609 20156
rect 20545 20096 20609 20100
rect 20625 20156 20689 20160
rect 20625 20100 20629 20156
rect 20629 20100 20685 20156
rect 20685 20100 20689 20156
rect 20625 20096 20689 20100
rect 20705 20156 20769 20160
rect 20705 20100 20709 20156
rect 20709 20100 20765 20156
rect 20765 20100 20769 20156
rect 20705 20096 20769 20100
rect 20785 20156 20849 20160
rect 20785 20100 20789 20156
rect 20789 20100 20845 20156
rect 20845 20100 20849 20156
rect 20785 20096 20849 20100
rect 6550 19612 6614 19616
rect 6550 19556 6554 19612
rect 6554 19556 6610 19612
rect 6610 19556 6614 19612
rect 6550 19552 6614 19556
rect 6630 19612 6694 19616
rect 6630 19556 6634 19612
rect 6634 19556 6690 19612
rect 6690 19556 6694 19612
rect 6630 19552 6694 19556
rect 6710 19612 6774 19616
rect 6710 19556 6714 19612
rect 6714 19556 6770 19612
rect 6770 19556 6774 19612
rect 6710 19552 6774 19556
rect 6790 19612 6854 19616
rect 6790 19556 6794 19612
rect 6794 19556 6850 19612
rect 6850 19556 6854 19612
rect 6790 19552 6854 19556
rect 12148 19612 12212 19616
rect 12148 19556 12152 19612
rect 12152 19556 12208 19612
rect 12208 19556 12212 19612
rect 12148 19552 12212 19556
rect 12228 19612 12292 19616
rect 12228 19556 12232 19612
rect 12232 19556 12288 19612
rect 12288 19556 12292 19612
rect 12228 19552 12292 19556
rect 12308 19612 12372 19616
rect 12308 19556 12312 19612
rect 12312 19556 12368 19612
rect 12368 19556 12372 19612
rect 12308 19552 12372 19556
rect 12388 19612 12452 19616
rect 12388 19556 12392 19612
rect 12392 19556 12448 19612
rect 12448 19556 12452 19612
rect 12388 19552 12452 19556
rect 21588 19756 21652 19820
rect 17746 19612 17810 19616
rect 17746 19556 17750 19612
rect 17750 19556 17806 19612
rect 17806 19556 17810 19612
rect 17746 19552 17810 19556
rect 17826 19612 17890 19616
rect 17826 19556 17830 19612
rect 17830 19556 17886 19612
rect 17886 19556 17890 19612
rect 17826 19552 17890 19556
rect 17906 19612 17970 19616
rect 17906 19556 17910 19612
rect 17910 19556 17966 19612
rect 17966 19556 17970 19612
rect 17906 19552 17970 19556
rect 17986 19612 18050 19616
rect 17986 19556 17990 19612
rect 17990 19556 18046 19612
rect 18046 19556 18050 19612
rect 17986 19552 18050 19556
rect 3751 19068 3815 19072
rect 3751 19012 3755 19068
rect 3755 19012 3811 19068
rect 3811 19012 3815 19068
rect 3751 19008 3815 19012
rect 3831 19068 3895 19072
rect 3831 19012 3835 19068
rect 3835 19012 3891 19068
rect 3891 19012 3895 19068
rect 3831 19008 3895 19012
rect 3911 19068 3975 19072
rect 3911 19012 3915 19068
rect 3915 19012 3971 19068
rect 3971 19012 3975 19068
rect 3911 19008 3975 19012
rect 3991 19068 4055 19072
rect 3991 19012 3995 19068
rect 3995 19012 4051 19068
rect 4051 19012 4055 19068
rect 3991 19008 4055 19012
rect 9349 19068 9413 19072
rect 9349 19012 9353 19068
rect 9353 19012 9409 19068
rect 9409 19012 9413 19068
rect 9349 19008 9413 19012
rect 9429 19068 9493 19072
rect 9429 19012 9433 19068
rect 9433 19012 9489 19068
rect 9489 19012 9493 19068
rect 9429 19008 9493 19012
rect 9509 19068 9573 19072
rect 9509 19012 9513 19068
rect 9513 19012 9569 19068
rect 9569 19012 9573 19068
rect 9509 19008 9573 19012
rect 9589 19068 9653 19072
rect 9589 19012 9593 19068
rect 9593 19012 9649 19068
rect 9649 19012 9653 19068
rect 9589 19008 9653 19012
rect 14947 19068 15011 19072
rect 14947 19012 14951 19068
rect 14951 19012 15007 19068
rect 15007 19012 15011 19068
rect 14947 19008 15011 19012
rect 15027 19068 15091 19072
rect 15027 19012 15031 19068
rect 15031 19012 15087 19068
rect 15087 19012 15091 19068
rect 15027 19008 15091 19012
rect 15107 19068 15171 19072
rect 15107 19012 15111 19068
rect 15111 19012 15167 19068
rect 15167 19012 15171 19068
rect 15107 19008 15171 19012
rect 15187 19068 15251 19072
rect 15187 19012 15191 19068
rect 15191 19012 15247 19068
rect 15247 19012 15251 19068
rect 15187 19008 15251 19012
rect 20545 19068 20609 19072
rect 20545 19012 20549 19068
rect 20549 19012 20605 19068
rect 20605 19012 20609 19068
rect 20545 19008 20609 19012
rect 20625 19068 20689 19072
rect 20625 19012 20629 19068
rect 20629 19012 20685 19068
rect 20685 19012 20689 19068
rect 20625 19008 20689 19012
rect 20705 19068 20769 19072
rect 20705 19012 20709 19068
rect 20709 19012 20765 19068
rect 20765 19012 20769 19068
rect 20705 19008 20769 19012
rect 20785 19068 20849 19072
rect 20785 19012 20789 19068
rect 20789 19012 20845 19068
rect 20845 19012 20849 19068
rect 20785 19008 20849 19012
rect 21036 18532 21100 18596
rect 6550 18524 6614 18528
rect 6550 18468 6554 18524
rect 6554 18468 6610 18524
rect 6610 18468 6614 18524
rect 6550 18464 6614 18468
rect 6630 18524 6694 18528
rect 6630 18468 6634 18524
rect 6634 18468 6690 18524
rect 6690 18468 6694 18524
rect 6630 18464 6694 18468
rect 6710 18524 6774 18528
rect 6710 18468 6714 18524
rect 6714 18468 6770 18524
rect 6770 18468 6774 18524
rect 6710 18464 6774 18468
rect 6790 18524 6854 18528
rect 6790 18468 6794 18524
rect 6794 18468 6850 18524
rect 6850 18468 6854 18524
rect 6790 18464 6854 18468
rect 12148 18524 12212 18528
rect 12148 18468 12152 18524
rect 12152 18468 12208 18524
rect 12208 18468 12212 18524
rect 12148 18464 12212 18468
rect 12228 18524 12292 18528
rect 12228 18468 12232 18524
rect 12232 18468 12288 18524
rect 12288 18468 12292 18524
rect 12228 18464 12292 18468
rect 12308 18524 12372 18528
rect 12308 18468 12312 18524
rect 12312 18468 12368 18524
rect 12368 18468 12372 18524
rect 12308 18464 12372 18468
rect 12388 18524 12452 18528
rect 12388 18468 12392 18524
rect 12392 18468 12448 18524
rect 12448 18468 12452 18524
rect 12388 18464 12452 18468
rect 17746 18524 17810 18528
rect 17746 18468 17750 18524
rect 17750 18468 17806 18524
rect 17806 18468 17810 18524
rect 17746 18464 17810 18468
rect 17826 18524 17890 18528
rect 17826 18468 17830 18524
rect 17830 18468 17886 18524
rect 17886 18468 17890 18524
rect 17826 18464 17890 18468
rect 17906 18524 17970 18528
rect 17906 18468 17910 18524
rect 17910 18468 17966 18524
rect 17966 18468 17970 18524
rect 17906 18464 17970 18468
rect 17986 18524 18050 18528
rect 17986 18468 17990 18524
rect 17990 18468 18046 18524
rect 18046 18468 18050 18524
rect 17986 18464 18050 18468
rect 3751 17980 3815 17984
rect 3751 17924 3755 17980
rect 3755 17924 3811 17980
rect 3811 17924 3815 17980
rect 3751 17920 3815 17924
rect 3831 17980 3895 17984
rect 3831 17924 3835 17980
rect 3835 17924 3891 17980
rect 3891 17924 3895 17980
rect 3831 17920 3895 17924
rect 3911 17980 3975 17984
rect 3911 17924 3915 17980
rect 3915 17924 3971 17980
rect 3971 17924 3975 17980
rect 3911 17920 3975 17924
rect 3991 17980 4055 17984
rect 3991 17924 3995 17980
rect 3995 17924 4051 17980
rect 4051 17924 4055 17980
rect 3991 17920 4055 17924
rect 9349 17980 9413 17984
rect 9349 17924 9353 17980
rect 9353 17924 9409 17980
rect 9409 17924 9413 17980
rect 9349 17920 9413 17924
rect 9429 17980 9493 17984
rect 9429 17924 9433 17980
rect 9433 17924 9489 17980
rect 9489 17924 9493 17980
rect 9429 17920 9493 17924
rect 9509 17980 9573 17984
rect 9509 17924 9513 17980
rect 9513 17924 9569 17980
rect 9569 17924 9573 17980
rect 9509 17920 9573 17924
rect 9589 17980 9653 17984
rect 9589 17924 9593 17980
rect 9593 17924 9649 17980
rect 9649 17924 9653 17980
rect 9589 17920 9653 17924
rect 14947 17980 15011 17984
rect 14947 17924 14951 17980
rect 14951 17924 15007 17980
rect 15007 17924 15011 17980
rect 14947 17920 15011 17924
rect 15027 17980 15091 17984
rect 15027 17924 15031 17980
rect 15031 17924 15087 17980
rect 15087 17924 15091 17980
rect 15027 17920 15091 17924
rect 15107 17980 15171 17984
rect 15107 17924 15111 17980
rect 15111 17924 15167 17980
rect 15167 17924 15171 17980
rect 15107 17920 15171 17924
rect 15187 17980 15251 17984
rect 15187 17924 15191 17980
rect 15191 17924 15247 17980
rect 15247 17924 15251 17980
rect 15187 17920 15251 17924
rect 20545 17980 20609 17984
rect 20545 17924 20549 17980
rect 20549 17924 20605 17980
rect 20605 17924 20609 17980
rect 20545 17920 20609 17924
rect 20625 17980 20689 17984
rect 20625 17924 20629 17980
rect 20629 17924 20685 17980
rect 20685 17924 20689 17980
rect 20625 17920 20689 17924
rect 20705 17980 20769 17984
rect 20705 17924 20709 17980
rect 20709 17924 20765 17980
rect 20765 17924 20769 17980
rect 20705 17920 20769 17924
rect 20785 17980 20849 17984
rect 20785 17924 20789 17980
rect 20789 17924 20845 17980
rect 20845 17924 20849 17980
rect 20785 17920 20849 17924
rect 13860 17912 13924 17916
rect 13860 17856 13910 17912
rect 13910 17856 13924 17912
rect 13860 17852 13924 17856
rect 6550 17436 6614 17440
rect 6550 17380 6554 17436
rect 6554 17380 6610 17436
rect 6610 17380 6614 17436
rect 6550 17376 6614 17380
rect 6630 17436 6694 17440
rect 6630 17380 6634 17436
rect 6634 17380 6690 17436
rect 6690 17380 6694 17436
rect 6630 17376 6694 17380
rect 6710 17436 6774 17440
rect 6710 17380 6714 17436
rect 6714 17380 6770 17436
rect 6770 17380 6774 17436
rect 6710 17376 6774 17380
rect 6790 17436 6854 17440
rect 6790 17380 6794 17436
rect 6794 17380 6850 17436
rect 6850 17380 6854 17436
rect 6790 17376 6854 17380
rect 12148 17436 12212 17440
rect 12148 17380 12152 17436
rect 12152 17380 12208 17436
rect 12208 17380 12212 17436
rect 12148 17376 12212 17380
rect 12228 17436 12292 17440
rect 12228 17380 12232 17436
rect 12232 17380 12288 17436
rect 12288 17380 12292 17436
rect 12228 17376 12292 17380
rect 12308 17436 12372 17440
rect 12308 17380 12312 17436
rect 12312 17380 12368 17436
rect 12368 17380 12372 17436
rect 12308 17376 12372 17380
rect 12388 17436 12452 17440
rect 12388 17380 12392 17436
rect 12392 17380 12448 17436
rect 12448 17380 12452 17436
rect 12388 17376 12452 17380
rect 17746 17436 17810 17440
rect 17746 17380 17750 17436
rect 17750 17380 17806 17436
rect 17806 17380 17810 17436
rect 17746 17376 17810 17380
rect 17826 17436 17890 17440
rect 17826 17380 17830 17436
rect 17830 17380 17886 17436
rect 17886 17380 17890 17436
rect 17826 17376 17890 17380
rect 17906 17436 17970 17440
rect 17906 17380 17910 17436
rect 17910 17380 17966 17436
rect 17966 17380 17970 17436
rect 17906 17376 17970 17380
rect 17986 17436 18050 17440
rect 17986 17380 17990 17436
rect 17990 17380 18046 17436
rect 18046 17380 18050 17436
rect 17986 17376 18050 17380
rect 3751 16892 3815 16896
rect 3751 16836 3755 16892
rect 3755 16836 3811 16892
rect 3811 16836 3815 16892
rect 3751 16832 3815 16836
rect 3831 16892 3895 16896
rect 3831 16836 3835 16892
rect 3835 16836 3891 16892
rect 3891 16836 3895 16892
rect 3831 16832 3895 16836
rect 3911 16892 3975 16896
rect 3911 16836 3915 16892
rect 3915 16836 3971 16892
rect 3971 16836 3975 16892
rect 3911 16832 3975 16836
rect 3991 16892 4055 16896
rect 3991 16836 3995 16892
rect 3995 16836 4051 16892
rect 4051 16836 4055 16892
rect 3991 16832 4055 16836
rect 9349 16892 9413 16896
rect 9349 16836 9353 16892
rect 9353 16836 9409 16892
rect 9409 16836 9413 16892
rect 9349 16832 9413 16836
rect 9429 16892 9493 16896
rect 9429 16836 9433 16892
rect 9433 16836 9489 16892
rect 9489 16836 9493 16892
rect 9429 16832 9493 16836
rect 9509 16892 9573 16896
rect 9509 16836 9513 16892
rect 9513 16836 9569 16892
rect 9569 16836 9573 16892
rect 9509 16832 9573 16836
rect 9589 16892 9653 16896
rect 9589 16836 9593 16892
rect 9593 16836 9649 16892
rect 9649 16836 9653 16892
rect 9589 16832 9653 16836
rect 14947 16892 15011 16896
rect 14947 16836 14951 16892
rect 14951 16836 15007 16892
rect 15007 16836 15011 16892
rect 14947 16832 15011 16836
rect 15027 16892 15091 16896
rect 15027 16836 15031 16892
rect 15031 16836 15087 16892
rect 15087 16836 15091 16892
rect 15027 16832 15091 16836
rect 15107 16892 15171 16896
rect 15107 16836 15111 16892
rect 15111 16836 15167 16892
rect 15167 16836 15171 16892
rect 15107 16832 15171 16836
rect 15187 16892 15251 16896
rect 15187 16836 15191 16892
rect 15191 16836 15247 16892
rect 15247 16836 15251 16892
rect 15187 16832 15251 16836
rect 20545 16892 20609 16896
rect 20545 16836 20549 16892
rect 20549 16836 20605 16892
rect 20605 16836 20609 16892
rect 20545 16832 20609 16836
rect 20625 16892 20689 16896
rect 20625 16836 20629 16892
rect 20629 16836 20685 16892
rect 20685 16836 20689 16892
rect 20625 16832 20689 16836
rect 20705 16892 20769 16896
rect 20705 16836 20709 16892
rect 20709 16836 20765 16892
rect 20765 16836 20769 16892
rect 20705 16832 20769 16836
rect 20785 16892 20849 16896
rect 20785 16836 20789 16892
rect 20789 16836 20845 16892
rect 20845 16836 20849 16892
rect 20785 16832 20849 16836
rect 6550 16348 6614 16352
rect 6550 16292 6554 16348
rect 6554 16292 6610 16348
rect 6610 16292 6614 16348
rect 6550 16288 6614 16292
rect 6630 16348 6694 16352
rect 6630 16292 6634 16348
rect 6634 16292 6690 16348
rect 6690 16292 6694 16348
rect 6630 16288 6694 16292
rect 6710 16348 6774 16352
rect 6710 16292 6714 16348
rect 6714 16292 6770 16348
rect 6770 16292 6774 16348
rect 6710 16288 6774 16292
rect 6790 16348 6854 16352
rect 6790 16292 6794 16348
rect 6794 16292 6850 16348
rect 6850 16292 6854 16348
rect 6790 16288 6854 16292
rect 12148 16348 12212 16352
rect 12148 16292 12152 16348
rect 12152 16292 12208 16348
rect 12208 16292 12212 16348
rect 12148 16288 12212 16292
rect 12228 16348 12292 16352
rect 12228 16292 12232 16348
rect 12232 16292 12288 16348
rect 12288 16292 12292 16348
rect 12228 16288 12292 16292
rect 12308 16348 12372 16352
rect 12308 16292 12312 16348
rect 12312 16292 12368 16348
rect 12368 16292 12372 16348
rect 12308 16288 12372 16292
rect 12388 16348 12452 16352
rect 12388 16292 12392 16348
rect 12392 16292 12448 16348
rect 12448 16292 12452 16348
rect 12388 16288 12452 16292
rect 17746 16348 17810 16352
rect 17746 16292 17750 16348
rect 17750 16292 17806 16348
rect 17806 16292 17810 16348
rect 17746 16288 17810 16292
rect 17826 16348 17890 16352
rect 17826 16292 17830 16348
rect 17830 16292 17886 16348
rect 17886 16292 17890 16348
rect 17826 16288 17890 16292
rect 17906 16348 17970 16352
rect 17906 16292 17910 16348
rect 17910 16292 17966 16348
rect 17966 16292 17970 16348
rect 17906 16288 17970 16292
rect 17986 16348 18050 16352
rect 17986 16292 17990 16348
rect 17990 16292 18046 16348
rect 18046 16292 18050 16348
rect 17986 16288 18050 16292
rect 3751 15804 3815 15808
rect 3751 15748 3755 15804
rect 3755 15748 3811 15804
rect 3811 15748 3815 15804
rect 3751 15744 3815 15748
rect 3831 15804 3895 15808
rect 3831 15748 3835 15804
rect 3835 15748 3891 15804
rect 3891 15748 3895 15804
rect 3831 15744 3895 15748
rect 3911 15804 3975 15808
rect 3911 15748 3915 15804
rect 3915 15748 3971 15804
rect 3971 15748 3975 15804
rect 3911 15744 3975 15748
rect 3991 15804 4055 15808
rect 3991 15748 3995 15804
rect 3995 15748 4051 15804
rect 4051 15748 4055 15804
rect 3991 15744 4055 15748
rect 9349 15804 9413 15808
rect 9349 15748 9353 15804
rect 9353 15748 9409 15804
rect 9409 15748 9413 15804
rect 9349 15744 9413 15748
rect 9429 15804 9493 15808
rect 9429 15748 9433 15804
rect 9433 15748 9489 15804
rect 9489 15748 9493 15804
rect 9429 15744 9493 15748
rect 9509 15804 9573 15808
rect 9509 15748 9513 15804
rect 9513 15748 9569 15804
rect 9569 15748 9573 15804
rect 9509 15744 9573 15748
rect 9589 15804 9653 15808
rect 9589 15748 9593 15804
rect 9593 15748 9649 15804
rect 9649 15748 9653 15804
rect 9589 15744 9653 15748
rect 14947 15804 15011 15808
rect 14947 15748 14951 15804
rect 14951 15748 15007 15804
rect 15007 15748 15011 15804
rect 14947 15744 15011 15748
rect 15027 15804 15091 15808
rect 15027 15748 15031 15804
rect 15031 15748 15087 15804
rect 15087 15748 15091 15804
rect 15027 15744 15091 15748
rect 15107 15804 15171 15808
rect 15107 15748 15111 15804
rect 15111 15748 15167 15804
rect 15167 15748 15171 15804
rect 15107 15744 15171 15748
rect 15187 15804 15251 15808
rect 15187 15748 15191 15804
rect 15191 15748 15247 15804
rect 15247 15748 15251 15804
rect 15187 15744 15251 15748
rect 20545 15804 20609 15808
rect 20545 15748 20549 15804
rect 20549 15748 20605 15804
rect 20605 15748 20609 15804
rect 20545 15744 20609 15748
rect 20625 15804 20689 15808
rect 20625 15748 20629 15804
rect 20629 15748 20685 15804
rect 20685 15748 20689 15804
rect 20625 15744 20689 15748
rect 20705 15804 20769 15808
rect 20705 15748 20709 15804
rect 20709 15748 20765 15804
rect 20765 15748 20769 15804
rect 20705 15744 20769 15748
rect 20785 15804 20849 15808
rect 20785 15748 20789 15804
rect 20789 15748 20845 15804
rect 20845 15748 20849 15804
rect 20785 15744 20849 15748
rect 18828 15600 18892 15604
rect 18828 15544 18878 15600
rect 18878 15544 18892 15600
rect 18828 15540 18892 15544
rect 6550 15260 6614 15264
rect 6550 15204 6554 15260
rect 6554 15204 6610 15260
rect 6610 15204 6614 15260
rect 6550 15200 6614 15204
rect 6630 15260 6694 15264
rect 6630 15204 6634 15260
rect 6634 15204 6690 15260
rect 6690 15204 6694 15260
rect 6630 15200 6694 15204
rect 6710 15260 6774 15264
rect 6710 15204 6714 15260
rect 6714 15204 6770 15260
rect 6770 15204 6774 15260
rect 6710 15200 6774 15204
rect 6790 15260 6854 15264
rect 6790 15204 6794 15260
rect 6794 15204 6850 15260
rect 6850 15204 6854 15260
rect 6790 15200 6854 15204
rect 12148 15260 12212 15264
rect 12148 15204 12152 15260
rect 12152 15204 12208 15260
rect 12208 15204 12212 15260
rect 12148 15200 12212 15204
rect 12228 15260 12292 15264
rect 12228 15204 12232 15260
rect 12232 15204 12288 15260
rect 12288 15204 12292 15260
rect 12228 15200 12292 15204
rect 12308 15260 12372 15264
rect 12308 15204 12312 15260
rect 12312 15204 12368 15260
rect 12368 15204 12372 15260
rect 12308 15200 12372 15204
rect 12388 15260 12452 15264
rect 12388 15204 12392 15260
rect 12392 15204 12448 15260
rect 12448 15204 12452 15260
rect 12388 15200 12452 15204
rect 17746 15260 17810 15264
rect 17746 15204 17750 15260
rect 17750 15204 17806 15260
rect 17806 15204 17810 15260
rect 17746 15200 17810 15204
rect 17826 15260 17890 15264
rect 17826 15204 17830 15260
rect 17830 15204 17886 15260
rect 17886 15204 17890 15260
rect 17826 15200 17890 15204
rect 17906 15260 17970 15264
rect 17906 15204 17910 15260
rect 17910 15204 17966 15260
rect 17966 15204 17970 15260
rect 17906 15200 17970 15204
rect 17986 15260 18050 15264
rect 17986 15204 17990 15260
rect 17990 15204 18046 15260
rect 18046 15204 18050 15260
rect 17986 15200 18050 15204
rect 3751 14716 3815 14720
rect 3751 14660 3755 14716
rect 3755 14660 3811 14716
rect 3811 14660 3815 14716
rect 3751 14656 3815 14660
rect 3831 14716 3895 14720
rect 3831 14660 3835 14716
rect 3835 14660 3891 14716
rect 3891 14660 3895 14716
rect 3831 14656 3895 14660
rect 3911 14716 3975 14720
rect 3911 14660 3915 14716
rect 3915 14660 3971 14716
rect 3971 14660 3975 14716
rect 3911 14656 3975 14660
rect 3991 14716 4055 14720
rect 3991 14660 3995 14716
rect 3995 14660 4051 14716
rect 4051 14660 4055 14716
rect 3991 14656 4055 14660
rect 9349 14716 9413 14720
rect 9349 14660 9353 14716
rect 9353 14660 9409 14716
rect 9409 14660 9413 14716
rect 9349 14656 9413 14660
rect 9429 14716 9493 14720
rect 9429 14660 9433 14716
rect 9433 14660 9489 14716
rect 9489 14660 9493 14716
rect 9429 14656 9493 14660
rect 9509 14716 9573 14720
rect 9509 14660 9513 14716
rect 9513 14660 9569 14716
rect 9569 14660 9573 14716
rect 9509 14656 9573 14660
rect 9589 14716 9653 14720
rect 9589 14660 9593 14716
rect 9593 14660 9649 14716
rect 9649 14660 9653 14716
rect 9589 14656 9653 14660
rect 14947 14716 15011 14720
rect 14947 14660 14951 14716
rect 14951 14660 15007 14716
rect 15007 14660 15011 14716
rect 14947 14656 15011 14660
rect 15027 14716 15091 14720
rect 15027 14660 15031 14716
rect 15031 14660 15087 14716
rect 15087 14660 15091 14716
rect 15027 14656 15091 14660
rect 15107 14716 15171 14720
rect 15107 14660 15111 14716
rect 15111 14660 15167 14716
rect 15167 14660 15171 14716
rect 15107 14656 15171 14660
rect 15187 14716 15251 14720
rect 15187 14660 15191 14716
rect 15191 14660 15247 14716
rect 15247 14660 15251 14716
rect 15187 14656 15251 14660
rect 20545 14716 20609 14720
rect 20545 14660 20549 14716
rect 20549 14660 20605 14716
rect 20605 14660 20609 14716
rect 20545 14656 20609 14660
rect 20625 14716 20689 14720
rect 20625 14660 20629 14716
rect 20629 14660 20685 14716
rect 20685 14660 20689 14716
rect 20625 14656 20689 14660
rect 20705 14716 20769 14720
rect 20705 14660 20709 14716
rect 20709 14660 20765 14716
rect 20765 14660 20769 14716
rect 20705 14656 20769 14660
rect 20785 14716 20849 14720
rect 20785 14660 20789 14716
rect 20789 14660 20845 14716
rect 20845 14660 20849 14716
rect 20785 14656 20849 14660
rect 6550 14172 6614 14176
rect 6550 14116 6554 14172
rect 6554 14116 6610 14172
rect 6610 14116 6614 14172
rect 6550 14112 6614 14116
rect 6630 14172 6694 14176
rect 6630 14116 6634 14172
rect 6634 14116 6690 14172
rect 6690 14116 6694 14172
rect 6630 14112 6694 14116
rect 6710 14172 6774 14176
rect 6710 14116 6714 14172
rect 6714 14116 6770 14172
rect 6770 14116 6774 14172
rect 6710 14112 6774 14116
rect 6790 14172 6854 14176
rect 6790 14116 6794 14172
rect 6794 14116 6850 14172
rect 6850 14116 6854 14172
rect 6790 14112 6854 14116
rect 12148 14172 12212 14176
rect 12148 14116 12152 14172
rect 12152 14116 12208 14172
rect 12208 14116 12212 14172
rect 12148 14112 12212 14116
rect 12228 14172 12292 14176
rect 12228 14116 12232 14172
rect 12232 14116 12288 14172
rect 12288 14116 12292 14172
rect 12228 14112 12292 14116
rect 12308 14172 12372 14176
rect 12308 14116 12312 14172
rect 12312 14116 12368 14172
rect 12368 14116 12372 14172
rect 12308 14112 12372 14116
rect 12388 14172 12452 14176
rect 12388 14116 12392 14172
rect 12392 14116 12448 14172
rect 12448 14116 12452 14172
rect 12388 14112 12452 14116
rect 17746 14172 17810 14176
rect 17746 14116 17750 14172
rect 17750 14116 17806 14172
rect 17806 14116 17810 14172
rect 17746 14112 17810 14116
rect 17826 14172 17890 14176
rect 17826 14116 17830 14172
rect 17830 14116 17886 14172
rect 17886 14116 17890 14172
rect 17826 14112 17890 14116
rect 17906 14172 17970 14176
rect 17906 14116 17910 14172
rect 17910 14116 17966 14172
rect 17966 14116 17970 14172
rect 17906 14112 17970 14116
rect 17986 14172 18050 14176
rect 17986 14116 17990 14172
rect 17990 14116 18046 14172
rect 18046 14116 18050 14172
rect 17986 14112 18050 14116
rect 3751 13628 3815 13632
rect 3751 13572 3755 13628
rect 3755 13572 3811 13628
rect 3811 13572 3815 13628
rect 3751 13568 3815 13572
rect 3831 13628 3895 13632
rect 3831 13572 3835 13628
rect 3835 13572 3891 13628
rect 3891 13572 3895 13628
rect 3831 13568 3895 13572
rect 3911 13628 3975 13632
rect 3911 13572 3915 13628
rect 3915 13572 3971 13628
rect 3971 13572 3975 13628
rect 3911 13568 3975 13572
rect 3991 13628 4055 13632
rect 3991 13572 3995 13628
rect 3995 13572 4051 13628
rect 4051 13572 4055 13628
rect 3991 13568 4055 13572
rect 9349 13628 9413 13632
rect 9349 13572 9353 13628
rect 9353 13572 9409 13628
rect 9409 13572 9413 13628
rect 9349 13568 9413 13572
rect 9429 13628 9493 13632
rect 9429 13572 9433 13628
rect 9433 13572 9489 13628
rect 9489 13572 9493 13628
rect 9429 13568 9493 13572
rect 9509 13628 9573 13632
rect 9509 13572 9513 13628
rect 9513 13572 9569 13628
rect 9569 13572 9573 13628
rect 9509 13568 9573 13572
rect 9589 13628 9653 13632
rect 9589 13572 9593 13628
rect 9593 13572 9649 13628
rect 9649 13572 9653 13628
rect 9589 13568 9653 13572
rect 14947 13628 15011 13632
rect 14947 13572 14951 13628
rect 14951 13572 15007 13628
rect 15007 13572 15011 13628
rect 14947 13568 15011 13572
rect 15027 13628 15091 13632
rect 15027 13572 15031 13628
rect 15031 13572 15087 13628
rect 15087 13572 15091 13628
rect 15027 13568 15091 13572
rect 15107 13628 15171 13632
rect 15107 13572 15111 13628
rect 15111 13572 15167 13628
rect 15167 13572 15171 13628
rect 15107 13568 15171 13572
rect 15187 13628 15251 13632
rect 15187 13572 15191 13628
rect 15191 13572 15247 13628
rect 15247 13572 15251 13628
rect 15187 13568 15251 13572
rect 20545 13628 20609 13632
rect 20545 13572 20549 13628
rect 20549 13572 20605 13628
rect 20605 13572 20609 13628
rect 20545 13568 20609 13572
rect 20625 13628 20689 13632
rect 20625 13572 20629 13628
rect 20629 13572 20685 13628
rect 20685 13572 20689 13628
rect 20625 13568 20689 13572
rect 20705 13628 20769 13632
rect 20705 13572 20709 13628
rect 20709 13572 20765 13628
rect 20765 13572 20769 13628
rect 20705 13568 20769 13572
rect 20785 13628 20849 13632
rect 20785 13572 20789 13628
rect 20789 13572 20845 13628
rect 20845 13572 20849 13628
rect 20785 13568 20849 13572
rect 6550 13084 6614 13088
rect 6550 13028 6554 13084
rect 6554 13028 6610 13084
rect 6610 13028 6614 13084
rect 6550 13024 6614 13028
rect 6630 13084 6694 13088
rect 6630 13028 6634 13084
rect 6634 13028 6690 13084
rect 6690 13028 6694 13084
rect 6630 13024 6694 13028
rect 6710 13084 6774 13088
rect 6710 13028 6714 13084
rect 6714 13028 6770 13084
rect 6770 13028 6774 13084
rect 6710 13024 6774 13028
rect 6790 13084 6854 13088
rect 6790 13028 6794 13084
rect 6794 13028 6850 13084
rect 6850 13028 6854 13084
rect 6790 13024 6854 13028
rect 12148 13084 12212 13088
rect 12148 13028 12152 13084
rect 12152 13028 12208 13084
rect 12208 13028 12212 13084
rect 12148 13024 12212 13028
rect 12228 13084 12292 13088
rect 12228 13028 12232 13084
rect 12232 13028 12288 13084
rect 12288 13028 12292 13084
rect 12228 13024 12292 13028
rect 12308 13084 12372 13088
rect 12308 13028 12312 13084
rect 12312 13028 12368 13084
rect 12368 13028 12372 13084
rect 12308 13024 12372 13028
rect 12388 13084 12452 13088
rect 12388 13028 12392 13084
rect 12392 13028 12448 13084
rect 12448 13028 12452 13084
rect 12388 13024 12452 13028
rect 17746 13084 17810 13088
rect 17746 13028 17750 13084
rect 17750 13028 17806 13084
rect 17806 13028 17810 13084
rect 17746 13024 17810 13028
rect 17826 13084 17890 13088
rect 17826 13028 17830 13084
rect 17830 13028 17886 13084
rect 17886 13028 17890 13084
rect 17826 13024 17890 13028
rect 17906 13084 17970 13088
rect 17906 13028 17910 13084
rect 17910 13028 17966 13084
rect 17966 13028 17970 13084
rect 17906 13024 17970 13028
rect 17986 13084 18050 13088
rect 17986 13028 17990 13084
rect 17990 13028 18046 13084
rect 18046 13028 18050 13084
rect 17986 13024 18050 13028
rect 19196 12820 19260 12884
rect 3751 12540 3815 12544
rect 3751 12484 3755 12540
rect 3755 12484 3811 12540
rect 3811 12484 3815 12540
rect 3751 12480 3815 12484
rect 3831 12540 3895 12544
rect 3831 12484 3835 12540
rect 3835 12484 3891 12540
rect 3891 12484 3895 12540
rect 3831 12480 3895 12484
rect 3911 12540 3975 12544
rect 3911 12484 3915 12540
rect 3915 12484 3971 12540
rect 3971 12484 3975 12540
rect 3911 12480 3975 12484
rect 3991 12540 4055 12544
rect 3991 12484 3995 12540
rect 3995 12484 4051 12540
rect 4051 12484 4055 12540
rect 3991 12480 4055 12484
rect 9349 12540 9413 12544
rect 9349 12484 9353 12540
rect 9353 12484 9409 12540
rect 9409 12484 9413 12540
rect 9349 12480 9413 12484
rect 9429 12540 9493 12544
rect 9429 12484 9433 12540
rect 9433 12484 9489 12540
rect 9489 12484 9493 12540
rect 9429 12480 9493 12484
rect 9509 12540 9573 12544
rect 9509 12484 9513 12540
rect 9513 12484 9569 12540
rect 9569 12484 9573 12540
rect 9509 12480 9573 12484
rect 9589 12540 9653 12544
rect 9589 12484 9593 12540
rect 9593 12484 9649 12540
rect 9649 12484 9653 12540
rect 9589 12480 9653 12484
rect 14947 12540 15011 12544
rect 14947 12484 14951 12540
rect 14951 12484 15007 12540
rect 15007 12484 15011 12540
rect 14947 12480 15011 12484
rect 15027 12540 15091 12544
rect 15027 12484 15031 12540
rect 15031 12484 15087 12540
rect 15087 12484 15091 12540
rect 15027 12480 15091 12484
rect 15107 12540 15171 12544
rect 15107 12484 15111 12540
rect 15111 12484 15167 12540
rect 15167 12484 15171 12540
rect 15107 12480 15171 12484
rect 15187 12540 15251 12544
rect 15187 12484 15191 12540
rect 15191 12484 15247 12540
rect 15247 12484 15251 12540
rect 15187 12480 15251 12484
rect 20545 12540 20609 12544
rect 20545 12484 20549 12540
rect 20549 12484 20605 12540
rect 20605 12484 20609 12540
rect 20545 12480 20609 12484
rect 20625 12540 20689 12544
rect 20625 12484 20629 12540
rect 20629 12484 20685 12540
rect 20685 12484 20689 12540
rect 20625 12480 20689 12484
rect 20705 12540 20769 12544
rect 20705 12484 20709 12540
rect 20709 12484 20765 12540
rect 20765 12484 20769 12540
rect 20705 12480 20769 12484
rect 20785 12540 20849 12544
rect 20785 12484 20789 12540
rect 20789 12484 20845 12540
rect 20845 12484 20849 12540
rect 20785 12480 20849 12484
rect 6550 11996 6614 12000
rect 6550 11940 6554 11996
rect 6554 11940 6610 11996
rect 6610 11940 6614 11996
rect 6550 11936 6614 11940
rect 6630 11996 6694 12000
rect 6630 11940 6634 11996
rect 6634 11940 6690 11996
rect 6690 11940 6694 11996
rect 6630 11936 6694 11940
rect 6710 11996 6774 12000
rect 6710 11940 6714 11996
rect 6714 11940 6770 11996
rect 6770 11940 6774 11996
rect 6710 11936 6774 11940
rect 6790 11996 6854 12000
rect 6790 11940 6794 11996
rect 6794 11940 6850 11996
rect 6850 11940 6854 11996
rect 6790 11936 6854 11940
rect 12148 11996 12212 12000
rect 12148 11940 12152 11996
rect 12152 11940 12208 11996
rect 12208 11940 12212 11996
rect 12148 11936 12212 11940
rect 12228 11996 12292 12000
rect 12228 11940 12232 11996
rect 12232 11940 12288 11996
rect 12288 11940 12292 11996
rect 12228 11936 12292 11940
rect 12308 11996 12372 12000
rect 12308 11940 12312 11996
rect 12312 11940 12368 11996
rect 12368 11940 12372 11996
rect 12308 11936 12372 11940
rect 12388 11996 12452 12000
rect 12388 11940 12392 11996
rect 12392 11940 12448 11996
rect 12448 11940 12452 11996
rect 12388 11936 12452 11940
rect 17746 11996 17810 12000
rect 17746 11940 17750 11996
rect 17750 11940 17806 11996
rect 17806 11940 17810 11996
rect 17746 11936 17810 11940
rect 17826 11996 17890 12000
rect 17826 11940 17830 11996
rect 17830 11940 17886 11996
rect 17886 11940 17890 11996
rect 17826 11936 17890 11940
rect 17906 11996 17970 12000
rect 17906 11940 17910 11996
rect 17910 11940 17966 11996
rect 17966 11940 17970 11996
rect 17906 11936 17970 11940
rect 17986 11996 18050 12000
rect 17986 11940 17990 11996
rect 17990 11940 18046 11996
rect 18046 11940 18050 11996
rect 17986 11936 18050 11940
rect 3751 11452 3815 11456
rect 3751 11396 3755 11452
rect 3755 11396 3811 11452
rect 3811 11396 3815 11452
rect 3751 11392 3815 11396
rect 3831 11452 3895 11456
rect 3831 11396 3835 11452
rect 3835 11396 3891 11452
rect 3891 11396 3895 11452
rect 3831 11392 3895 11396
rect 3911 11452 3975 11456
rect 3911 11396 3915 11452
rect 3915 11396 3971 11452
rect 3971 11396 3975 11452
rect 3911 11392 3975 11396
rect 3991 11452 4055 11456
rect 3991 11396 3995 11452
rect 3995 11396 4051 11452
rect 4051 11396 4055 11452
rect 3991 11392 4055 11396
rect 9349 11452 9413 11456
rect 9349 11396 9353 11452
rect 9353 11396 9409 11452
rect 9409 11396 9413 11452
rect 9349 11392 9413 11396
rect 9429 11452 9493 11456
rect 9429 11396 9433 11452
rect 9433 11396 9489 11452
rect 9489 11396 9493 11452
rect 9429 11392 9493 11396
rect 9509 11452 9573 11456
rect 9509 11396 9513 11452
rect 9513 11396 9569 11452
rect 9569 11396 9573 11452
rect 9509 11392 9573 11396
rect 9589 11452 9653 11456
rect 9589 11396 9593 11452
rect 9593 11396 9649 11452
rect 9649 11396 9653 11452
rect 9589 11392 9653 11396
rect 14947 11452 15011 11456
rect 14947 11396 14951 11452
rect 14951 11396 15007 11452
rect 15007 11396 15011 11452
rect 14947 11392 15011 11396
rect 15027 11452 15091 11456
rect 15027 11396 15031 11452
rect 15031 11396 15087 11452
rect 15087 11396 15091 11452
rect 15027 11392 15091 11396
rect 15107 11452 15171 11456
rect 15107 11396 15111 11452
rect 15111 11396 15167 11452
rect 15167 11396 15171 11452
rect 15107 11392 15171 11396
rect 15187 11452 15251 11456
rect 15187 11396 15191 11452
rect 15191 11396 15247 11452
rect 15247 11396 15251 11452
rect 15187 11392 15251 11396
rect 20545 11452 20609 11456
rect 20545 11396 20549 11452
rect 20549 11396 20605 11452
rect 20605 11396 20609 11452
rect 20545 11392 20609 11396
rect 20625 11452 20689 11456
rect 20625 11396 20629 11452
rect 20629 11396 20685 11452
rect 20685 11396 20689 11452
rect 20625 11392 20689 11396
rect 20705 11452 20769 11456
rect 20705 11396 20709 11452
rect 20709 11396 20765 11452
rect 20765 11396 20769 11452
rect 20705 11392 20769 11396
rect 20785 11452 20849 11456
rect 20785 11396 20789 11452
rect 20789 11396 20845 11452
rect 20845 11396 20849 11452
rect 20785 11392 20849 11396
rect 21036 11052 21100 11116
rect 6550 10908 6614 10912
rect 6550 10852 6554 10908
rect 6554 10852 6610 10908
rect 6610 10852 6614 10908
rect 6550 10848 6614 10852
rect 6630 10908 6694 10912
rect 6630 10852 6634 10908
rect 6634 10852 6690 10908
rect 6690 10852 6694 10908
rect 6630 10848 6694 10852
rect 6710 10908 6774 10912
rect 6710 10852 6714 10908
rect 6714 10852 6770 10908
rect 6770 10852 6774 10908
rect 6710 10848 6774 10852
rect 6790 10908 6854 10912
rect 6790 10852 6794 10908
rect 6794 10852 6850 10908
rect 6850 10852 6854 10908
rect 6790 10848 6854 10852
rect 12148 10908 12212 10912
rect 12148 10852 12152 10908
rect 12152 10852 12208 10908
rect 12208 10852 12212 10908
rect 12148 10848 12212 10852
rect 12228 10908 12292 10912
rect 12228 10852 12232 10908
rect 12232 10852 12288 10908
rect 12288 10852 12292 10908
rect 12228 10848 12292 10852
rect 12308 10908 12372 10912
rect 12308 10852 12312 10908
rect 12312 10852 12368 10908
rect 12368 10852 12372 10908
rect 12308 10848 12372 10852
rect 12388 10908 12452 10912
rect 12388 10852 12392 10908
rect 12392 10852 12448 10908
rect 12448 10852 12452 10908
rect 12388 10848 12452 10852
rect 17746 10908 17810 10912
rect 17746 10852 17750 10908
rect 17750 10852 17806 10908
rect 17806 10852 17810 10908
rect 17746 10848 17810 10852
rect 17826 10908 17890 10912
rect 17826 10852 17830 10908
rect 17830 10852 17886 10908
rect 17886 10852 17890 10908
rect 17826 10848 17890 10852
rect 17906 10908 17970 10912
rect 17906 10852 17910 10908
rect 17910 10852 17966 10908
rect 17966 10852 17970 10908
rect 17906 10848 17970 10852
rect 17986 10908 18050 10912
rect 17986 10852 17990 10908
rect 17990 10852 18046 10908
rect 18046 10852 18050 10908
rect 17986 10848 18050 10852
rect 3751 10364 3815 10368
rect 3751 10308 3755 10364
rect 3755 10308 3811 10364
rect 3811 10308 3815 10364
rect 3751 10304 3815 10308
rect 3831 10364 3895 10368
rect 3831 10308 3835 10364
rect 3835 10308 3891 10364
rect 3891 10308 3895 10364
rect 3831 10304 3895 10308
rect 3911 10364 3975 10368
rect 3911 10308 3915 10364
rect 3915 10308 3971 10364
rect 3971 10308 3975 10364
rect 3911 10304 3975 10308
rect 3991 10364 4055 10368
rect 3991 10308 3995 10364
rect 3995 10308 4051 10364
rect 4051 10308 4055 10364
rect 3991 10304 4055 10308
rect 9349 10364 9413 10368
rect 9349 10308 9353 10364
rect 9353 10308 9409 10364
rect 9409 10308 9413 10364
rect 9349 10304 9413 10308
rect 9429 10364 9493 10368
rect 9429 10308 9433 10364
rect 9433 10308 9489 10364
rect 9489 10308 9493 10364
rect 9429 10304 9493 10308
rect 9509 10364 9573 10368
rect 9509 10308 9513 10364
rect 9513 10308 9569 10364
rect 9569 10308 9573 10364
rect 9509 10304 9573 10308
rect 9589 10364 9653 10368
rect 9589 10308 9593 10364
rect 9593 10308 9649 10364
rect 9649 10308 9653 10364
rect 9589 10304 9653 10308
rect 14947 10364 15011 10368
rect 14947 10308 14951 10364
rect 14951 10308 15007 10364
rect 15007 10308 15011 10364
rect 14947 10304 15011 10308
rect 15027 10364 15091 10368
rect 15027 10308 15031 10364
rect 15031 10308 15087 10364
rect 15087 10308 15091 10364
rect 15027 10304 15091 10308
rect 15107 10364 15171 10368
rect 15107 10308 15111 10364
rect 15111 10308 15167 10364
rect 15167 10308 15171 10364
rect 15107 10304 15171 10308
rect 15187 10364 15251 10368
rect 15187 10308 15191 10364
rect 15191 10308 15247 10364
rect 15247 10308 15251 10364
rect 15187 10304 15251 10308
rect 20545 10364 20609 10368
rect 20545 10308 20549 10364
rect 20549 10308 20605 10364
rect 20605 10308 20609 10364
rect 20545 10304 20609 10308
rect 20625 10364 20689 10368
rect 20625 10308 20629 10364
rect 20629 10308 20685 10364
rect 20685 10308 20689 10364
rect 20625 10304 20689 10308
rect 20705 10364 20769 10368
rect 20705 10308 20709 10364
rect 20709 10308 20765 10364
rect 20765 10308 20769 10364
rect 20705 10304 20769 10308
rect 20785 10364 20849 10368
rect 20785 10308 20789 10364
rect 20789 10308 20845 10364
rect 20845 10308 20849 10364
rect 20785 10304 20849 10308
rect 18828 9888 18892 9892
rect 18828 9832 18878 9888
rect 18878 9832 18892 9888
rect 18828 9828 18892 9832
rect 6550 9820 6614 9824
rect 6550 9764 6554 9820
rect 6554 9764 6610 9820
rect 6610 9764 6614 9820
rect 6550 9760 6614 9764
rect 6630 9820 6694 9824
rect 6630 9764 6634 9820
rect 6634 9764 6690 9820
rect 6690 9764 6694 9820
rect 6630 9760 6694 9764
rect 6710 9820 6774 9824
rect 6710 9764 6714 9820
rect 6714 9764 6770 9820
rect 6770 9764 6774 9820
rect 6710 9760 6774 9764
rect 6790 9820 6854 9824
rect 6790 9764 6794 9820
rect 6794 9764 6850 9820
rect 6850 9764 6854 9820
rect 6790 9760 6854 9764
rect 12148 9820 12212 9824
rect 12148 9764 12152 9820
rect 12152 9764 12208 9820
rect 12208 9764 12212 9820
rect 12148 9760 12212 9764
rect 12228 9820 12292 9824
rect 12228 9764 12232 9820
rect 12232 9764 12288 9820
rect 12288 9764 12292 9820
rect 12228 9760 12292 9764
rect 12308 9820 12372 9824
rect 12308 9764 12312 9820
rect 12312 9764 12368 9820
rect 12368 9764 12372 9820
rect 12308 9760 12372 9764
rect 12388 9820 12452 9824
rect 12388 9764 12392 9820
rect 12392 9764 12448 9820
rect 12448 9764 12452 9820
rect 12388 9760 12452 9764
rect 17746 9820 17810 9824
rect 17746 9764 17750 9820
rect 17750 9764 17806 9820
rect 17806 9764 17810 9820
rect 17746 9760 17810 9764
rect 17826 9820 17890 9824
rect 17826 9764 17830 9820
rect 17830 9764 17886 9820
rect 17886 9764 17890 9820
rect 17826 9760 17890 9764
rect 17906 9820 17970 9824
rect 17906 9764 17910 9820
rect 17910 9764 17966 9820
rect 17966 9764 17970 9820
rect 17906 9760 17970 9764
rect 17986 9820 18050 9824
rect 17986 9764 17990 9820
rect 17990 9764 18046 9820
rect 18046 9764 18050 9820
rect 17986 9760 18050 9764
rect 3751 9276 3815 9280
rect 3751 9220 3755 9276
rect 3755 9220 3811 9276
rect 3811 9220 3815 9276
rect 3751 9216 3815 9220
rect 3831 9276 3895 9280
rect 3831 9220 3835 9276
rect 3835 9220 3891 9276
rect 3891 9220 3895 9276
rect 3831 9216 3895 9220
rect 3911 9276 3975 9280
rect 3911 9220 3915 9276
rect 3915 9220 3971 9276
rect 3971 9220 3975 9276
rect 3911 9216 3975 9220
rect 3991 9276 4055 9280
rect 3991 9220 3995 9276
rect 3995 9220 4051 9276
rect 4051 9220 4055 9276
rect 3991 9216 4055 9220
rect 9349 9276 9413 9280
rect 9349 9220 9353 9276
rect 9353 9220 9409 9276
rect 9409 9220 9413 9276
rect 9349 9216 9413 9220
rect 9429 9276 9493 9280
rect 9429 9220 9433 9276
rect 9433 9220 9489 9276
rect 9489 9220 9493 9276
rect 9429 9216 9493 9220
rect 9509 9276 9573 9280
rect 9509 9220 9513 9276
rect 9513 9220 9569 9276
rect 9569 9220 9573 9276
rect 9509 9216 9573 9220
rect 9589 9276 9653 9280
rect 9589 9220 9593 9276
rect 9593 9220 9649 9276
rect 9649 9220 9653 9276
rect 9589 9216 9653 9220
rect 14947 9276 15011 9280
rect 14947 9220 14951 9276
rect 14951 9220 15007 9276
rect 15007 9220 15011 9276
rect 14947 9216 15011 9220
rect 15027 9276 15091 9280
rect 15027 9220 15031 9276
rect 15031 9220 15087 9276
rect 15087 9220 15091 9276
rect 15027 9216 15091 9220
rect 15107 9276 15171 9280
rect 15107 9220 15111 9276
rect 15111 9220 15167 9276
rect 15167 9220 15171 9276
rect 15107 9216 15171 9220
rect 15187 9276 15251 9280
rect 15187 9220 15191 9276
rect 15191 9220 15247 9276
rect 15247 9220 15251 9276
rect 15187 9216 15251 9220
rect 20545 9276 20609 9280
rect 20545 9220 20549 9276
rect 20549 9220 20605 9276
rect 20605 9220 20609 9276
rect 20545 9216 20609 9220
rect 20625 9276 20689 9280
rect 20625 9220 20629 9276
rect 20629 9220 20685 9276
rect 20685 9220 20689 9276
rect 20625 9216 20689 9220
rect 20705 9276 20769 9280
rect 20705 9220 20709 9276
rect 20709 9220 20765 9276
rect 20765 9220 20769 9276
rect 20705 9216 20769 9220
rect 20785 9276 20849 9280
rect 20785 9220 20789 9276
rect 20789 9220 20845 9276
rect 20845 9220 20849 9276
rect 20785 9216 20849 9220
rect 6550 8732 6614 8736
rect 6550 8676 6554 8732
rect 6554 8676 6610 8732
rect 6610 8676 6614 8732
rect 6550 8672 6614 8676
rect 6630 8732 6694 8736
rect 6630 8676 6634 8732
rect 6634 8676 6690 8732
rect 6690 8676 6694 8732
rect 6630 8672 6694 8676
rect 6710 8732 6774 8736
rect 6710 8676 6714 8732
rect 6714 8676 6770 8732
rect 6770 8676 6774 8732
rect 6710 8672 6774 8676
rect 6790 8732 6854 8736
rect 6790 8676 6794 8732
rect 6794 8676 6850 8732
rect 6850 8676 6854 8732
rect 6790 8672 6854 8676
rect 12148 8732 12212 8736
rect 12148 8676 12152 8732
rect 12152 8676 12208 8732
rect 12208 8676 12212 8732
rect 12148 8672 12212 8676
rect 12228 8732 12292 8736
rect 12228 8676 12232 8732
rect 12232 8676 12288 8732
rect 12288 8676 12292 8732
rect 12228 8672 12292 8676
rect 12308 8732 12372 8736
rect 12308 8676 12312 8732
rect 12312 8676 12368 8732
rect 12368 8676 12372 8732
rect 12308 8672 12372 8676
rect 12388 8732 12452 8736
rect 12388 8676 12392 8732
rect 12392 8676 12448 8732
rect 12448 8676 12452 8732
rect 12388 8672 12452 8676
rect 17746 8732 17810 8736
rect 17746 8676 17750 8732
rect 17750 8676 17806 8732
rect 17806 8676 17810 8732
rect 17746 8672 17810 8676
rect 17826 8732 17890 8736
rect 17826 8676 17830 8732
rect 17830 8676 17886 8732
rect 17886 8676 17890 8732
rect 17826 8672 17890 8676
rect 17906 8732 17970 8736
rect 17906 8676 17910 8732
rect 17910 8676 17966 8732
rect 17966 8676 17970 8732
rect 17906 8672 17970 8676
rect 17986 8732 18050 8736
rect 17986 8676 17990 8732
rect 17990 8676 18046 8732
rect 18046 8676 18050 8732
rect 17986 8672 18050 8676
rect 3751 8188 3815 8192
rect 3751 8132 3755 8188
rect 3755 8132 3811 8188
rect 3811 8132 3815 8188
rect 3751 8128 3815 8132
rect 3831 8188 3895 8192
rect 3831 8132 3835 8188
rect 3835 8132 3891 8188
rect 3891 8132 3895 8188
rect 3831 8128 3895 8132
rect 3911 8188 3975 8192
rect 3911 8132 3915 8188
rect 3915 8132 3971 8188
rect 3971 8132 3975 8188
rect 3911 8128 3975 8132
rect 3991 8188 4055 8192
rect 3991 8132 3995 8188
rect 3995 8132 4051 8188
rect 4051 8132 4055 8188
rect 3991 8128 4055 8132
rect 9349 8188 9413 8192
rect 9349 8132 9353 8188
rect 9353 8132 9409 8188
rect 9409 8132 9413 8188
rect 9349 8128 9413 8132
rect 9429 8188 9493 8192
rect 9429 8132 9433 8188
rect 9433 8132 9489 8188
rect 9489 8132 9493 8188
rect 9429 8128 9493 8132
rect 9509 8188 9573 8192
rect 9509 8132 9513 8188
rect 9513 8132 9569 8188
rect 9569 8132 9573 8188
rect 9509 8128 9573 8132
rect 9589 8188 9653 8192
rect 9589 8132 9593 8188
rect 9593 8132 9649 8188
rect 9649 8132 9653 8188
rect 9589 8128 9653 8132
rect 14947 8188 15011 8192
rect 14947 8132 14951 8188
rect 14951 8132 15007 8188
rect 15007 8132 15011 8188
rect 14947 8128 15011 8132
rect 15027 8188 15091 8192
rect 15027 8132 15031 8188
rect 15031 8132 15087 8188
rect 15087 8132 15091 8188
rect 15027 8128 15091 8132
rect 15107 8188 15171 8192
rect 15107 8132 15111 8188
rect 15111 8132 15167 8188
rect 15167 8132 15171 8188
rect 15107 8128 15171 8132
rect 15187 8188 15251 8192
rect 15187 8132 15191 8188
rect 15191 8132 15247 8188
rect 15247 8132 15251 8188
rect 15187 8128 15251 8132
rect 20545 8188 20609 8192
rect 20545 8132 20549 8188
rect 20549 8132 20605 8188
rect 20605 8132 20609 8188
rect 20545 8128 20609 8132
rect 20625 8188 20689 8192
rect 20625 8132 20629 8188
rect 20629 8132 20685 8188
rect 20685 8132 20689 8188
rect 20625 8128 20689 8132
rect 20705 8188 20769 8192
rect 20705 8132 20709 8188
rect 20709 8132 20765 8188
rect 20765 8132 20769 8188
rect 20705 8128 20769 8132
rect 20785 8188 20849 8192
rect 20785 8132 20789 8188
rect 20789 8132 20845 8188
rect 20845 8132 20849 8188
rect 20785 8128 20849 8132
rect 6550 7644 6614 7648
rect 6550 7588 6554 7644
rect 6554 7588 6610 7644
rect 6610 7588 6614 7644
rect 6550 7584 6614 7588
rect 6630 7644 6694 7648
rect 6630 7588 6634 7644
rect 6634 7588 6690 7644
rect 6690 7588 6694 7644
rect 6630 7584 6694 7588
rect 6710 7644 6774 7648
rect 6710 7588 6714 7644
rect 6714 7588 6770 7644
rect 6770 7588 6774 7644
rect 6710 7584 6774 7588
rect 6790 7644 6854 7648
rect 6790 7588 6794 7644
rect 6794 7588 6850 7644
rect 6850 7588 6854 7644
rect 6790 7584 6854 7588
rect 12148 7644 12212 7648
rect 12148 7588 12152 7644
rect 12152 7588 12208 7644
rect 12208 7588 12212 7644
rect 12148 7584 12212 7588
rect 12228 7644 12292 7648
rect 12228 7588 12232 7644
rect 12232 7588 12288 7644
rect 12288 7588 12292 7644
rect 12228 7584 12292 7588
rect 12308 7644 12372 7648
rect 12308 7588 12312 7644
rect 12312 7588 12368 7644
rect 12368 7588 12372 7644
rect 12308 7584 12372 7588
rect 12388 7644 12452 7648
rect 12388 7588 12392 7644
rect 12392 7588 12448 7644
rect 12448 7588 12452 7644
rect 12388 7584 12452 7588
rect 17746 7644 17810 7648
rect 17746 7588 17750 7644
rect 17750 7588 17806 7644
rect 17806 7588 17810 7644
rect 17746 7584 17810 7588
rect 17826 7644 17890 7648
rect 17826 7588 17830 7644
rect 17830 7588 17886 7644
rect 17886 7588 17890 7644
rect 17826 7584 17890 7588
rect 17906 7644 17970 7648
rect 17906 7588 17910 7644
rect 17910 7588 17966 7644
rect 17966 7588 17970 7644
rect 17906 7584 17970 7588
rect 17986 7644 18050 7648
rect 17986 7588 17990 7644
rect 17990 7588 18046 7644
rect 18046 7588 18050 7644
rect 17986 7584 18050 7588
rect 21220 7380 21284 7444
rect 21588 7440 21652 7444
rect 21588 7384 21602 7440
rect 21602 7384 21652 7440
rect 21588 7380 21652 7384
rect 21036 7244 21100 7308
rect 19564 7168 19628 7172
rect 19564 7112 19578 7168
rect 19578 7112 19628 7168
rect 19564 7108 19628 7112
rect 3751 7100 3815 7104
rect 3751 7044 3755 7100
rect 3755 7044 3811 7100
rect 3811 7044 3815 7100
rect 3751 7040 3815 7044
rect 3831 7100 3895 7104
rect 3831 7044 3835 7100
rect 3835 7044 3891 7100
rect 3891 7044 3895 7100
rect 3831 7040 3895 7044
rect 3911 7100 3975 7104
rect 3911 7044 3915 7100
rect 3915 7044 3971 7100
rect 3971 7044 3975 7100
rect 3911 7040 3975 7044
rect 3991 7100 4055 7104
rect 3991 7044 3995 7100
rect 3995 7044 4051 7100
rect 4051 7044 4055 7100
rect 3991 7040 4055 7044
rect 9349 7100 9413 7104
rect 9349 7044 9353 7100
rect 9353 7044 9409 7100
rect 9409 7044 9413 7100
rect 9349 7040 9413 7044
rect 9429 7100 9493 7104
rect 9429 7044 9433 7100
rect 9433 7044 9489 7100
rect 9489 7044 9493 7100
rect 9429 7040 9493 7044
rect 9509 7100 9573 7104
rect 9509 7044 9513 7100
rect 9513 7044 9569 7100
rect 9569 7044 9573 7100
rect 9509 7040 9573 7044
rect 9589 7100 9653 7104
rect 9589 7044 9593 7100
rect 9593 7044 9649 7100
rect 9649 7044 9653 7100
rect 9589 7040 9653 7044
rect 14947 7100 15011 7104
rect 14947 7044 14951 7100
rect 14951 7044 15007 7100
rect 15007 7044 15011 7100
rect 14947 7040 15011 7044
rect 15027 7100 15091 7104
rect 15027 7044 15031 7100
rect 15031 7044 15087 7100
rect 15087 7044 15091 7100
rect 15027 7040 15091 7044
rect 15107 7100 15171 7104
rect 15107 7044 15111 7100
rect 15111 7044 15167 7100
rect 15167 7044 15171 7100
rect 15107 7040 15171 7044
rect 15187 7100 15251 7104
rect 15187 7044 15191 7100
rect 15191 7044 15247 7100
rect 15247 7044 15251 7100
rect 15187 7040 15251 7044
rect 20545 7100 20609 7104
rect 20545 7044 20549 7100
rect 20549 7044 20605 7100
rect 20605 7044 20609 7100
rect 20545 7040 20609 7044
rect 20625 7100 20689 7104
rect 20625 7044 20629 7100
rect 20629 7044 20685 7100
rect 20685 7044 20689 7100
rect 20625 7040 20689 7044
rect 20705 7100 20769 7104
rect 20705 7044 20709 7100
rect 20709 7044 20765 7100
rect 20765 7044 20769 7100
rect 20705 7040 20769 7044
rect 20785 7100 20849 7104
rect 20785 7044 20789 7100
rect 20789 7044 20845 7100
rect 20845 7044 20849 7100
rect 20785 7040 20849 7044
rect 19380 7032 19444 7036
rect 19380 6976 19430 7032
rect 19430 6976 19444 7032
rect 19380 6972 19444 6976
rect 21220 6624 21284 6628
rect 21220 6568 21270 6624
rect 21270 6568 21284 6624
rect 21220 6564 21284 6568
rect 6550 6556 6614 6560
rect 6550 6500 6554 6556
rect 6554 6500 6610 6556
rect 6610 6500 6614 6556
rect 6550 6496 6614 6500
rect 6630 6556 6694 6560
rect 6630 6500 6634 6556
rect 6634 6500 6690 6556
rect 6690 6500 6694 6556
rect 6630 6496 6694 6500
rect 6710 6556 6774 6560
rect 6710 6500 6714 6556
rect 6714 6500 6770 6556
rect 6770 6500 6774 6556
rect 6710 6496 6774 6500
rect 6790 6556 6854 6560
rect 6790 6500 6794 6556
rect 6794 6500 6850 6556
rect 6850 6500 6854 6556
rect 6790 6496 6854 6500
rect 12148 6556 12212 6560
rect 12148 6500 12152 6556
rect 12152 6500 12208 6556
rect 12208 6500 12212 6556
rect 12148 6496 12212 6500
rect 12228 6556 12292 6560
rect 12228 6500 12232 6556
rect 12232 6500 12288 6556
rect 12288 6500 12292 6556
rect 12228 6496 12292 6500
rect 12308 6556 12372 6560
rect 12308 6500 12312 6556
rect 12312 6500 12368 6556
rect 12368 6500 12372 6556
rect 12308 6496 12372 6500
rect 12388 6556 12452 6560
rect 12388 6500 12392 6556
rect 12392 6500 12448 6556
rect 12448 6500 12452 6556
rect 12388 6496 12452 6500
rect 17746 6556 17810 6560
rect 17746 6500 17750 6556
rect 17750 6500 17806 6556
rect 17806 6500 17810 6556
rect 17746 6496 17810 6500
rect 17826 6556 17890 6560
rect 17826 6500 17830 6556
rect 17830 6500 17886 6556
rect 17886 6500 17890 6556
rect 17826 6496 17890 6500
rect 17906 6556 17970 6560
rect 17906 6500 17910 6556
rect 17910 6500 17966 6556
rect 17966 6500 17970 6556
rect 17906 6496 17970 6500
rect 17986 6556 18050 6560
rect 17986 6500 17990 6556
rect 17990 6500 18046 6556
rect 18046 6500 18050 6556
rect 17986 6496 18050 6500
rect 19748 6428 19812 6492
rect 19380 6080 19444 6084
rect 19380 6024 19430 6080
rect 19430 6024 19444 6080
rect 19380 6020 19444 6024
rect 19564 6020 19628 6084
rect 3751 6012 3815 6016
rect 3751 5956 3755 6012
rect 3755 5956 3811 6012
rect 3811 5956 3815 6012
rect 3751 5952 3815 5956
rect 3831 6012 3895 6016
rect 3831 5956 3835 6012
rect 3835 5956 3891 6012
rect 3891 5956 3895 6012
rect 3831 5952 3895 5956
rect 3911 6012 3975 6016
rect 3911 5956 3915 6012
rect 3915 5956 3971 6012
rect 3971 5956 3975 6012
rect 3911 5952 3975 5956
rect 3991 6012 4055 6016
rect 3991 5956 3995 6012
rect 3995 5956 4051 6012
rect 4051 5956 4055 6012
rect 3991 5952 4055 5956
rect 9349 6012 9413 6016
rect 9349 5956 9353 6012
rect 9353 5956 9409 6012
rect 9409 5956 9413 6012
rect 9349 5952 9413 5956
rect 9429 6012 9493 6016
rect 9429 5956 9433 6012
rect 9433 5956 9489 6012
rect 9489 5956 9493 6012
rect 9429 5952 9493 5956
rect 9509 6012 9573 6016
rect 9509 5956 9513 6012
rect 9513 5956 9569 6012
rect 9569 5956 9573 6012
rect 9509 5952 9573 5956
rect 9589 6012 9653 6016
rect 9589 5956 9593 6012
rect 9593 5956 9649 6012
rect 9649 5956 9653 6012
rect 9589 5952 9653 5956
rect 14947 6012 15011 6016
rect 14947 5956 14951 6012
rect 14951 5956 15007 6012
rect 15007 5956 15011 6012
rect 14947 5952 15011 5956
rect 15027 6012 15091 6016
rect 15027 5956 15031 6012
rect 15031 5956 15087 6012
rect 15087 5956 15091 6012
rect 15027 5952 15091 5956
rect 15107 6012 15171 6016
rect 15107 5956 15111 6012
rect 15111 5956 15167 6012
rect 15167 5956 15171 6012
rect 15107 5952 15171 5956
rect 15187 6012 15251 6016
rect 15187 5956 15191 6012
rect 15191 5956 15247 6012
rect 15247 5956 15251 6012
rect 15187 5952 15251 5956
rect 20545 6012 20609 6016
rect 20545 5956 20549 6012
rect 20549 5956 20605 6012
rect 20605 5956 20609 6012
rect 20545 5952 20609 5956
rect 20625 6012 20689 6016
rect 20625 5956 20629 6012
rect 20629 5956 20685 6012
rect 20685 5956 20689 6012
rect 20625 5952 20689 5956
rect 20705 6012 20769 6016
rect 20705 5956 20709 6012
rect 20709 5956 20765 6012
rect 20765 5956 20769 6012
rect 20705 5952 20769 5956
rect 20785 6012 20849 6016
rect 20785 5956 20789 6012
rect 20789 5956 20845 6012
rect 20845 5956 20849 6012
rect 20785 5952 20849 5956
rect 6550 5468 6614 5472
rect 6550 5412 6554 5468
rect 6554 5412 6610 5468
rect 6610 5412 6614 5468
rect 6550 5408 6614 5412
rect 6630 5468 6694 5472
rect 6630 5412 6634 5468
rect 6634 5412 6690 5468
rect 6690 5412 6694 5468
rect 6630 5408 6694 5412
rect 6710 5468 6774 5472
rect 6710 5412 6714 5468
rect 6714 5412 6770 5468
rect 6770 5412 6774 5468
rect 6710 5408 6774 5412
rect 6790 5468 6854 5472
rect 6790 5412 6794 5468
rect 6794 5412 6850 5468
rect 6850 5412 6854 5468
rect 6790 5408 6854 5412
rect 12148 5468 12212 5472
rect 12148 5412 12152 5468
rect 12152 5412 12208 5468
rect 12208 5412 12212 5468
rect 12148 5408 12212 5412
rect 12228 5468 12292 5472
rect 12228 5412 12232 5468
rect 12232 5412 12288 5468
rect 12288 5412 12292 5468
rect 12228 5408 12292 5412
rect 12308 5468 12372 5472
rect 12308 5412 12312 5468
rect 12312 5412 12368 5468
rect 12368 5412 12372 5468
rect 12308 5408 12372 5412
rect 12388 5468 12452 5472
rect 12388 5412 12392 5468
rect 12392 5412 12448 5468
rect 12448 5412 12452 5468
rect 12388 5408 12452 5412
rect 17746 5468 17810 5472
rect 17746 5412 17750 5468
rect 17750 5412 17806 5468
rect 17806 5412 17810 5468
rect 17746 5408 17810 5412
rect 17826 5468 17890 5472
rect 17826 5412 17830 5468
rect 17830 5412 17886 5468
rect 17886 5412 17890 5468
rect 17826 5408 17890 5412
rect 17906 5468 17970 5472
rect 17906 5412 17910 5468
rect 17910 5412 17966 5468
rect 17966 5412 17970 5468
rect 17906 5408 17970 5412
rect 17986 5468 18050 5472
rect 17986 5412 17990 5468
rect 17990 5412 18046 5468
rect 18046 5412 18050 5468
rect 17986 5408 18050 5412
rect 3751 4924 3815 4928
rect 3751 4868 3755 4924
rect 3755 4868 3811 4924
rect 3811 4868 3815 4924
rect 3751 4864 3815 4868
rect 3831 4924 3895 4928
rect 3831 4868 3835 4924
rect 3835 4868 3891 4924
rect 3891 4868 3895 4924
rect 3831 4864 3895 4868
rect 3911 4924 3975 4928
rect 3911 4868 3915 4924
rect 3915 4868 3971 4924
rect 3971 4868 3975 4924
rect 3911 4864 3975 4868
rect 3991 4924 4055 4928
rect 3991 4868 3995 4924
rect 3995 4868 4051 4924
rect 4051 4868 4055 4924
rect 3991 4864 4055 4868
rect 9349 4924 9413 4928
rect 9349 4868 9353 4924
rect 9353 4868 9409 4924
rect 9409 4868 9413 4924
rect 9349 4864 9413 4868
rect 9429 4924 9493 4928
rect 9429 4868 9433 4924
rect 9433 4868 9489 4924
rect 9489 4868 9493 4924
rect 9429 4864 9493 4868
rect 9509 4924 9573 4928
rect 9509 4868 9513 4924
rect 9513 4868 9569 4924
rect 9569 4868 9573 4924
rect 9509 4864 9573 4868
rect 9589 4924 9653 4928
rect 9589 4868 9593 4924
rect 9593 4868 9649 4924
rect 9649 4868 9653 4924
rect 9589 4864 9653 4868
rect 14947 4924 15011 4928
rect 14947 4868 14951 4924
rect 14951 4868 15007 4924
rect 15007 4868 15011 4924
rect 14947 4864 15011 4868
rect 15027 4924 15091 4928
rect 15027 4868 15031 4924
rect 15031 4868 15087 4924
rect 15087 4868 15091 4924
rect 15027 4864 15091 4868
rect 15107 4924 15171 4928
rect 15107 4868 15111 4924
rect 15111 4868 15167 4924
rect 15167 4868 15171 4924
rect 15107 4864 15171 4868
rect 15187 4924 15251 4928
rect 15187 4868 15191 4924
rect 15191 4868 15247 4924
rect 15247 4868 15251 4924
rect 15187 4864 15251 4868
rect 20545 4924 20609 4928
rect 20545 4868 20549 4924
rect 20549 4868 20605 4924
rect 20605 4868 20609 4924
rect 20545 4864 20609 4868
rect 20625 4924 20689 4928
rect 20625 4868 20629 4924
rect 20629 4868 20685 4924
rect 20685 4868 20689 4924
rect 20625 4864 20689 4868
rect 20705 4924 20769 4928
rect 20705 4868 20709 4924
rect 20709 4868 20765 4924
rect 20765 4868 20769 4924
rect 20705 4864 20769 4868
rect 20785 4924 20849 4928
rect 20785 4868 20789 4924
rect 20789 4868 20845 4924
rect 20845 4868 20849 4924
rect 20785 4864 20849 4868
rect 19748 4796 19812 4860
rect 19196 4660 19260 4724
rect 21220 4388 21284 4452
rect 6550 4380 6614 4384
rect 6550 4324 6554 4380
rect 6554 4324 6610 4380
rect 6610 4324 6614 4380
rect 6550 4320 6614 4324
rect 6630 4380 6694 4384
rect 6630 4324 6634 4380
rect 6634 4324 6690 4380
rect 6690 4324 6694 4380
rect 6630 4320 6694 4324
rect 6710 4380 6774 4384
rect 6710 4324 6714 4380
rect 6714 4324 6770 4380
rect 6770 4324 6774 4380
rect 6710 4320 6774 4324
rect 6790 4380 6854 4384
rect 6790 4324 6794 4380
rect 6794 4324 6850 4380
rect 6850 4324 6854 4380
rect 6790 4320 6854 4324
rect 12148 4380 12212 4384
rect 12148 4324 12152 4380
rect 12152 4324 12208 4380
rect 12208 4324 12212 4380
rect 12148 4320 12212 4324
rect 12228 4380 12292 4384
rect 12228 4324 12232 4380
rect 12232 4324 12288 4380
rect 12288 4324 12292 4380
rect 12228 4320 12292 4324
rect 12308 4380 12372 4384
rect 12308 4324 12312 4380
rect 12312 4324 12368 4380
rect 12368 4324 12372 4380
rect 12308 4320 12372 4324
rect 12388 4380 12452 4384
rect 12388 4324 12392 4380
rect 12392 4324 12448 4380
rect 12448 4324 12452 4380
rect 12388 4320 12452 4324
rect 17746 4380 17810 4384
rect 17746 4324 17750 4380
rect 17750 4324 17806 4380
rect 17806 4324 17810 4380
rect 17746 4320 17810 4324
rect 17826 4380 17890 4384
rect 17826 4324 17830 4380
rect 17830 4324 17886 4380
rect 17886 4324 17890 4380
rect 17826 4320 17890 4324
rect 17906 4380 17970 4384
rect 17906 4324 17910 4380
rect 17910 4324 17966 4380
rect 17966 4324 17970 4380
rect 17906 4320 17970 4324
rect 17986 4380 18050 4384
rect 17986 4324 17990 4380
rect 17990 4324 18046 4380
rect 18046 4324 18050 4380
rect 17986 4320 18050 4324
rect 3751 3836 3815 3840
rect 3751 3780 3755 3836
rect 3755 3780 3811 3836
rect 3811 3780 3815 3836
rect 3751 3776 3815 3780
rect 3831 3836 3895 3840
rect 3831 3780 3835 3836
rect 3835 3780 3891 3836
rect 3891 3780 3895 3836
rect 3831 3776 3895 3780
rect 3911 3836 3975 3840
rect 3911 3780 3915 3836
rect 3915 3780 3971 3836
rect 3971 3780 3975 3836
rect 3911 3776 3975 3780
rect 3991 3836 4055 3840
rect 3991 3780 3995 3836
rect 3995 3780 4051 3836
rect 4051 3780 4055 3836
rect 3991 3776 4055 3780
rect 9349 3836 9413 3840
rect 9349 3780 9353 3836
rect 9353 3780 9409 3836
rect 9409 3780 9413 3836
rect 9349 3776 9413 3780
rect 9429 3836 9493 3840
rect 9429 3780 9433 3836
rect 9433 3780 9489 3836
rect 9489 3780 9493 3836
rect 9429 3776 9493 3780
rect 9509 3836 9573 3840
rect 9509 3780 9513 3836
rect 9513 3780 9569 3836
rect 9569 3780 9573 3836
rect 9509 3776 9573 3780
rect 9589 3836 9653 3840
rect 9589 3780 9593 3836
rect 9593 3780 9649 3836
rect 9649 3780 9653 3836
rect 9589 3776 9653 3780
rect 14947 3836 15011 3840
rect 14947 3780 14951 3836
rect 14951 3780 15007 3836
rect 15007 3780 15011 3836
rect 14947 3776 15011 3780
rect 15027 3836 15091 3840
rect 15027 3780 15031 3836
rect 15031 3780 15087 3836
rect 15087 3780 15091 3836
rect 15027 3776 15091 3780
rect 15107 3836 15171 3840
rect 15107 3780 15111 3836
rect 15111 3780 15167 3836
rect 15167 3780 15171 3836
rect 15107 3776 15171 3780
rect 15187 3836 15251 3840
rect 15187 3780 15191 3836
rect 15191 3780 15247 3836
rect 15247 3780 15251 3836
rect 15187 3776 15251 3780
rect 20545 3836 20609 3840
rect 20545 3780 20549 3836
rect 20549 3780 20605 3836
rect 20605 3780 20609 3836
rect 20545 3776 20609 3780
rect 20625 3836 20689 3840
rect 20625 3780 20629 3836
rect 20629 3780 20685 3836
rect 20685 3780 20689 3836
rect 20625 3776 20689 3780
rect 20705 3836 20769 3840
rect 20705 3780 20709 3836
rect 20709 3780 20765 3836
rect 20765 3780 20769 3836
rect 20705 3776 20769 3780
rect 20785 3836 20849 3840
rect 20785 3780 20789 3836
rect 20789 3780 20845 3836
rect 20845 3780 20849 3836
rect 20785 3776 20849 3780
rect 6550 3292 6614 3296
rect 6550 3236 6554 3292
rect 6554 3236 6610 3292
rect 6610 3236 6614 3292
rect 6550 3232 6614 3236
rect 6630 3292 6694 3296
rect 6630 3236 6634 3292
rect 6634 3236 6690 3292
rect 6690 3236 6694 3292
rect 6630 3232 6694 3236
rect 6710 3292 6774 3296
rect 6710 3236 6714 3292
rect 6714 3236 6770 3292
rect 6770 3236 6774 3292
rect 6710 3232 6774 3236
rect 6790 3292 6854 3296
rect 6790 3236 6794 3292
rect 6794 3236 6850 3292
rect 6850 3236 6854 3292
rect 6790 3232 6854 3236
rect 12148 3292 12212 3296
rect 12148 3236 12152 3292
rect 12152 3236 12208 3292
rect 12208 3236 12212 3292
rect 12148 3232 12212 3236
rect 12228 3292 12292 3296
rect 12228 3236 12232 3292
rect 12232 3236 12288 3292
rect 12288 3236 12292 3292
rect 12228 3232 12292 3236
rect 12308 3292 12372 3296
rect 12308 3236 12312 3292
rect 12312 3236 12368 3292
rect 12368 3236 12372 3292
rect 12308 3232 12372 3236
rect 12388 3292 12452 3296
rect 12388 3236 12392 3292
rect 12392 3236 12448 3292
rect 12448 3236 12452 3292
rect 12388 3232 12452 3236
rect 17746 3292 17810 3296
rect 17746 3236 17750 3292
rect 17750 3236 17806 3292
rect 17806 3236 17810 3292
rect 17746 3232 17810 3236
rect 17826 3292 17890 3296
rect 17826 3236 17830 3292
rect 17830 3236 17886 3292
rect 17886 3236 17890 3292
rect 17826 3232 17890 3236
rect 17906 3292 17970 3296
rect 17906 3236 17910 3292
rect 17910 3236 17966 3292
rect 17966 3236 17970 3292
rect 17906 3232 17970 3236
rect 17986 3292 18050 3296
rect 17986 3236 17990 3292
rect 17990 3236 18046 3292
rect 18046 3236 18050 3292
rect 17986 3232 18050 3236
rect 3751 2748 3815 2752
rect 3751 2692 3755 2748
rect 3755 2692 3811 2748
rect 3811 2692 3815 2748
rect 3751 2688 3815 2692
rect 3831 2748 3895 2752
rect 3831 2692 3835 2748
rect 3835 2692 3891 2748
rect 3891 2692 3895 2748
rect 3831 2688 3895 2692
rect 3911 2748 3975 2752
rect 3911 2692 3915 2748
rect 3915 2692 3971 2748
rect 3971 2692 3975 2748
rect 3911 2688 3975 2692
rect 3991 2748 4055 2752
rect 3991 2692 3995 2748
rect 3995 2692 4051 2748
rect 4051 2692 4055 2748
rect 3991 2688 4055 2692
rect 9349 2748 9413 2752
rect 9349 2692 9353 2748
rect 9353 2692 9409 2748
rect 9409 2692 9413 2748
rect 9349 2688 9413 2692
rect 9429 2748 9493 2752
rect 9429 2692 9433 2748
rect 9433 2692 9489 2748
rect 9489 2692 9493 2748
rect 9429 2688 9493 2692
rect 9509 2748 9573 2752
rect 9509 2692 9513 2748
rect 9513 2692 9569 2748
rect 9569 2692 9573 2748
rect 9509 2688 9573 2692
rect 9589 2748 9653 2752
rect 9589 2692 9593 2748
rect 9593 2692 9649 2748
rect 9649 2692 9653 2748
rect 9589 2688 9653 2692
rect 14947 2748 15011 2752
rect 14947 2692 14951 2748
rect 14951 2692 15007 2748
rect 15007 2692 15011 2748
rect 14947 2688 15011 2692
rect 15027 2748 15091 2752
rect 15027 2692 15031 2748
rect 15031 2692 15087 2748
rect 15087 2692 15091 2748
rect 15027 2688 15091 2692
rect 15107 2748 15171 2752
rect 15107 2692 15111 2748
rect 15111 2692 15167 2748
rect 15167 2692 15171 2748
rect 15107 2688 15171 2692
rect 15187 2748 15251 2752
rect 15187 2692 15191 2748
rect 15191 2692 15247 2748
rect 15247 2692 15251 2748
rect 15187 2688 15251 2692
rect 20545 2748 20609 2752
rect 20545 2692 20549 2748
rect 20549 2692 20605 2748
rect 20605 2692 20609 2748
rect 20545 2688 20609 2692
rect 20625 2748 20689 2752
rect 20625 2692 20629 2748
rect 20629 2692 20685 2748
rect 20685 2692 20689 2748
rect 20625 2688 20689 2692
rect 20705 2748 20769 2752
rect 20705 2692 20709 2748
rect 20709 2692 20765 2748
rect 20765 2692 20769 2748
rect 20705 2688 20769 2692
rect 20785 2748 20849 2752
rect 20785 2692 20789 2748
rect 20789 2692 20845 2748
rect 20845 2692 20849 2748
rect 20785 2688 20849 2692
rect 6550 2204 6614 2208
rect 6550 2148 6554 2204
rect 6554 2148 6610 2204
rect 6610 2148 6614 2204
rect 6550 2144 6614 2148
rect 6630 2204 6694 2208
rect 6630 2148 6634 2204
rect 6634 2148 6690 2204
rect 6690 2148 6694 2204
rect 6630 2144 6694 2148
rect 6710 2204 6774 2208
rect 6710 2148 6714 2204
rect 6714 2148 6770 2204
rect 6770 2148 6774 2204
rect 6710 2144 6774 2148
rect 6790 2204 6854 2208
rect 6790 2148 6794 2204
rect 6794 2148 6850 2204
rect 6850 2148 6854 2204
rect 6790 2144 6854 2148
rect 12148 2204 12212 2208
rect 12148 2148 12152 2204
rect 12152 2148 12208 2204
rect 12208 2148 12212 2204
rect 12148 2144 12212 2148
rect 12228 2204 12292 2208
rect 12228 2148 12232 2204
rect 12232 2148 12288 2204
rect 12288 2148 12292 2204
rect 12228 2144 12292 2148
rect 12308 2204 12372 2208
rect 12308 2148 12312 2204
rect 12312 2148 12368 2204
rect 12368 2148 12372 2204
rect 12308 2144 12372 2148
rect 12388 2204 12452 2208
rect 12388 2148 12392 2204
rect 12392 2148 12448 2204
rect 12448 2148 12452 2204
rect 12388 2144 12452 2148
rect 17746 2204 17810 2208
rect 17746 2148 17750 2204
rect 17750 2148 17806 2204
rect 17806 2148 17810 2204
rect 17746 2144 17810 2148
rect 17826 2204 17890 2208
rect 17826 2148 17830 2204
rect 17830 2148 17886 2204
rect 17886 2148 17890 2204
rect 17826 2144 17890 2148
rect 17906 2204 17970 2208
rect 17906 2148 17910 2204
rect 17910 2148 17966 2204
rect 17966 2148 17970 2204
rect 17906 2144 17970 2148
rect 17986 2204 18050 2208
rect 17986 2148 17990 2204
rect 17990 2148 18046 2204
rect 18046 2148 18050 2204
rect 17986 2144 18050 2148
<< metal4 >>
rect 3743 22336 4063 22352
rect 3743 22272 3751 22336
rect 3815 22272 3831 22336
rect 3895 22272 3911 22336
rect 3975 22272 3991 22336
rect 4055 22272 4063 22336
rect 3743 21248 4063 22272
rect 3743 21184 3751 21248
rect 3815 21184 3831 21248
rect 3895 21184 3911 21248
rect 3975 21184 3991 21248
rect 4055 21184 4063 21248
rect 3743 20160 4063 21184
rect 3743 20096 3751 20160
rect 3815 20096 3831 20160
rect 3895 20096 3911 20160
rect 3975 20096 3991 20160
rect 4055 20096 4063 20160
rect 3743 19072 4063 20096
rect 3743 19008 3751 19072
rect 3815 19008 3831 19072
rect 3895 19008 3911 19072
rect 3975 19008 3991 19072
rect 4055 19008 4063 19072
rect 3743 17984 4063 19008
rect 3743 17920 3751 17984
rect 3815 17920 3831 17984
rect 3895 17920 3911 17984
rect 3975 17920 3991 17984
rect 4055 17920 4063 17984
rect 3743 16896 4063 17920
rect 3743 16832 3751 16896
rect 3815 16832 3831 16896
rect 3895 16832 3911 16896
rect 3975 16832 3991 16896
rect 4055 16832 4063 16896
rect 3743 15808 4063 16832
rect 3743 15744 3751 15808
rect 3815 15744 3831 15808
rect 3895 15744 3911 15808
rect 3975 15744 3991 15808
rect 4055 15744 4063 15808
rect 3743 14720 4063 15744
rect 3743 14656 3751 14720
rect 3815 14656 3831 14720
rect 3895 14656 3911 14720
rect 3975 14656 3991 14720
rect 4055 14656 4063 14720
rect 3743 13632 4063 14656
rect 3743 13568 3751 13632
rect 3815 13568 3831 13632
rect 3895 13568 3911 13632
rect 3975 13568 3991 13632
rect 4055 13568 4063 13632
rect 3743 12544 4063 13568
rect 3743 12480 3751 12544
rect 3815 12480 3831 12544
rect 3895 12480 3911 12544
rect 3975 12480 3991 12544
rect 4055 12480 4063 12544
rect 3743 11456 4063 12480
rect 3743 11392 3751 11456
rect 3815 11392 3831 11456
rect 3895 11392 3911 11456
rect 3975 11392 3991 11456
rect 4055 11392 4063 11456
rect 3743 10368 4063 11392
rect 3743 10304 3751 10368
rect 3815 10304 3831 10368
rect 3895 10304 3911 10368
rect 3975 10304 3991 10368
rect 4055 10304 4063 10368
rect 3743 9280 4063 10304
rect 3743 9216 3751 9280
rect 3815 9216 3831 9280
rect 3895 9216 3911 9280
rect 3975 9216 3991 9280
rect 4055 9216 4063 9280
rect 3743 8192 4063 9216
rect 3743 8128 3751 8192
rect 3815 8128 3831 8192
rect 3895 8128 3911 8192
rect 3975 8128 3991 8192
rect 4055 8128 4063 8192
rect 3743 7104 4063 8128
rect 3743 7040 3751 7104
rect 3815 7040 3831 7104
rect 3895 7040 3911 7104
rect 3975 7040 3991 7104
rect 4055 7040 4063 7104
rect 3743 6016 4063 7040
rect 3743 5952 3751 6016
rect 3815 5952 3831 6016
rect 3895 5952 3911 6016
rect 3975 5952 3991 6016
rect 4055 5952 4063 6016
rect 3743 4928 4063 5952
rect 3743 4864 3751 4928
rect 3815 4864 3831 4928
rect 3895 4864 3911 4928
rect 3975 4864 3991 4928
rect 4055 4864 4063 4928
rect 3743 3840 4063 4864
rect 3743 3776 3751 3840
rect 3815 3776 3831 3840
rect 3895 3776 3911 3840
rect 3975 3776 3991 3840
rect 4055 3776 4063 3840
rect 3743 2752 4063 3776
rect 3743 2688 3751 2752
rect 3815 2688 3831 2752
rect 3895 2688 3911 2752
rect 3975 2688 3991 2752
rect 4055 2688 4063 2752
rect 3743 2128 4063 2688
rect 6542 21792 6862 22352
rect 6542 21728 6550 21792
rect 6614 21728 6630 21792
rect 6694 21728 6710 21792
rect 6774 21728 6790 21792
rect 6854 21728 6862 21792
rect 6542 20704 6862 21728
rect 6542 20640 6550 20704
rect 6614 20640 6630 20704
rect 6694 20640 6710 20704
rect 6774 20640 6790 20704
rect 6854 20640 6862 20704
rect 6542 19616 6862 20640
rect 6542 19552 6550 19616
rect 6614 19552 6630 19616
rect 6694 19552 6710 19616
rect 6774 19552 6790 19616
rect 6854 19552 6862 19616
rect 6542 18528 6862 19552
rect 6542 18464 6550 18528
rect 6614 18464 6630 18528
rect 6694 18464 6710 18528
rect 6774 18464 6790 18528
rect 6854 18464 6862 18528
rect 6542 17440 6862 18464
rect 6542 17376 6550 17440
rect 6614 17376 6630 17440
rect 6694 17376 6710 17440
rect 6774 17376 6790 17440
rect 6854 17376 6862 17440
rect 6542 16352 6862 17376
rect 6542 16288 6550 16352
rect 6614 16288 6630 16352
rect 6694 16288 6710 16352
rect 6774 16288 6790 16352
rect 6854 16288 6862 16352
rect 6542 15264 6862 16288
rect 6542 15200 6550 15264
rect 6614 15200 6630 15264
rect 6694 15200 6710 15264
rect 6774 15200 6790 15264
rect 6854 15200 6862 15264
rect 6542 14176 6862 15200
rect 6542 14112 6550 14176
rect 6614 14112 6630 14176
rect 6694 14112 6710 14176
rect 6774 14112 6790 14176
rect 6854 14112 6862 14176
rect 6542 13088 6862 14112
rect 6542 13024 6550 13088
rect 6614 13024 6630 13088
rect 6694 13024 6710 13088
rect 6774 13024 6790 13088
rect 6854 13024 6862 13088
rect 6542 12000 6862 13024
rect 6542 11936 6550 12000
rect 6614 11936 6630 12000
rect 6694 11936 6710 12000
rect 6774 11936 6790 12000
rect 6854 11936 6862 12000
rect 6542 10912 6862 11936
rect 6542 10848 6550 10912
rect 6614 10848 6630 10912
rect 6694 10848 6710 10912
rect 6774 10848 6790 10912
rect 6854 10848 6862 10912
rect 6542 9824 6862 10848
rect 6542 9760 6550 9824
rect 6614 9760 6630 9824
rect 6694 9760 6710 9824
rect 6774 9760 6790 9824
rect 6854 9760 6862 9824
rect 6542 8736 6862 9760
rect 6542 8672 6550 8736
rect 6614 8672 6630 8736
rect 6694 8672 6710 8736
rect 6774 8672 6790 8736
rect 6854 8672 6862 8736
rect 6542 7648 6862 8672
rect 6542 7584 6550 7648
rect 6614 7584 6630 7648
rect 6694 7584 6710 7648
rect 6774 7584 6790 7648
rect 6854 7584 6862 7648
rect 6542 6560 6862 7584
rect 6542 6496 6550 6560
rect 6614 6496 6630 6560
rect 6694 6496 6710 6560
rect 6774 6496 6790 6560
rect 6854 6496 6862 6560
rect 6542 5472 6862 6496
rect 6542 5408 6550 5472
rect 6614 5408 6630 5472
rect 6694 5408 6710 5472
rect 6774 5408 6790 5472
rect 6854 5408 6862 5472
rect 6542 4384 6862 5408
rect 6542 4320 6550 4384
rect 6614 4320 6630 4384
rect 6694 4320 6710 4384
rect 6774 4320 6790 4384
rect 6854 4320 6862 4384
rect 6542 3296 6862 4320
rect 6542 3232 6550 3296
rect 6614 3232 6630 3296
rect 6694 3232 6710 3296
rect 6774 3232 6790 3296
rect 6854 3232 6862 3296
rect 6542 2208 6862 3232
rect 6542 2144 6550 2208
rect 6614 2144 6630 2208
rect 6694 2144 6710 2208
rect 6774 2144 6790 2208
rect 6854 2144 6862 2208
rect 6542 2128 6862 2144
rect 9341 22336 9661 22352
rect 9341 22272 9349 22336
rect 9413 22272 9429 22336
rect 9493 22272 9509 22336
rect 9573 22272 9589 22336
rect 9653 22272 9661 22336
rect 9341 21248 9661 22272
rect 9341 21184 9349 21248
rect 9413 21184 9429 21248
rect 9493 21184 9509 21248
rect 9573 21184 9589 21248
rect 9653 21184 9661 21248
rect 9341 20160 9661 21184
rect 9341 20096 9349 20160
rect 9413 20096 9429 20160
rect 9493 20096 9509 20160
rect 9573 20096 9589 20160
rect 9653 20096 9661 20160
rect 9341 19072 9661 20096
rect 9341 19008 9349 19072
rect 9413 19008 9429 19072
rect 9493 19008 9509 19072
rect 9573 19008 9589 19072
rect 9653 19008 9661 19072
rect 9341 17984 9661 19008
rect 9341 17920 9349 17984
rect 9413 17920 9429 17984
rect 9493 17920 9509 17984
rect 9573 17920 9589 17984
rect 9653 17920 9661 17984
rect 9341 16896 9661 17920
rect 9341 16832 9349 16896
rect 9413 16832 9429 16896
rect 9493 16832 9509 16896
rect 9573 16832 9589 16896
rect 9653 16832 9661 16896
rect 9341 15808 9661 16832
rect 9341 15744 9349 15808
rect 9413 15744 9429 15808
rect 9493 15744 9509 15808
rect 9573 15744 9589 15808
rect 9653 15744 9661 15808
rect 9341 14720 9661 15744
rect 9341 14656 9349 14720
rect 9413 14656 9429 14720
rect 9493 14656 9509 14720
rect 9573 14656 9589 14720
rect 9653 14656 9661 14720
rect 9341 13632 9661 14656
rect 9341 13568 9349 13632
rect 9413 13568 9429 13632
rect 9493 13568 9509 13632
rect 9573 13568 9589 13632
rect 9653 13568 9661 13632
rect 9341 12544 9661 13568
rect 9341 12480 9349 12544
rect 9413 12480 9429 12544
rect 9493 12480 9509 12544
rect 9573 12480 9589 12544
rect 9653 12480 9661 12544
rect 9341 11456 9661 12480
rect 9341 11392 9349 11456
rect 9413 11392 9429 11456
rect 9493 11392 9509 11456
rect 9573 11392 9589 11456
rect 9653 11392 9661 11456
rect 9341 10368 9661 11392
rect 9341 10304 9349 10368
rect 9413 10304 9429 10368
rect 9493 10304 9509 10368
rect 9573 10304 9589 10368
rect 9653 10304 9661 10368
rect 9341 9280 9661 10304
rect 9341 9216 9349 9280
rect 9413 9216 9429 9280
rect 9493 9216 9509 9280
rect 9573 9216 9589 9280
rect 9653 9216 9661 9280
rect 9341 8192 9661 9216
rect 9341 8128 9349 8192
rect 9413 8128 9429 8192
rect 9493 8128 9509 8192
rect 9573 8128 9589 8192
rect 9653 8128 9661 8192
rect 9341 7104 9661 8128
rect 9341 7040 9349 7104
rect 9413 7040 9429 7104
rect 9493 7040 9509 7104
rect 9573 7040 9589 7104
rect 9653 7040 9661 7104
rect 9341 6016 9661 7040
rect 9341 5952 9349 6016
rect 9413 5952 9429 6016
rect 9493 5952 9509 6016
rect 9573 5952 9589 6016
rect 9653 5952 9661 6016
rect 9341 4928 9661 5952
rect 9341 4864 9349 4928
rect 9413 4864 9429 4928
rect 9493 4864 9509 4928
rect 9573 4864 9589 4928
rect 9653 4864 9661 4928
rect 9341 3840 9661 4864
rect 9341 3776 9349 3840
rect 9413 3776 9429 3840
rect 9493 3776 9509 3840
rect 9573 3776 9589 3840
rect 9653 3776 9661 3840
rect 9341 2752 9661 3776
rect 9341 2688 9349 2752
rect 9413 2688 9429 2752
rect 9493 2688 9509 2752
rect 9573 2688 9589 2752
rect 9653 2688 9661 2752
rect 9341 2128 9661 2688
rect 12140 21792 12460 22352
rect 12140 21728 12148 21792
rect 12212 21728 12228 21792
rect 12292 21728 12308 21792
rect 12372 21728 12388 21792
rect 12452 21728 12460 21792
rect 12140 20704 12460 21728
rect 14939 22336 15259 22352
rect 14939 22272 14947 22336
rect 15011 22272 15027 22336
rect 15091 22272 15107 22336
rect 15171 22272 15187 22336
rect 15251 22272 15259 22336
rect 13859 21316 13925 21317
rect 13859 21252 13860 21316
rect 13924 21252 13925 21316
rect 13859 21251 13925 21252
rect 12140 20640 12148 20704
rect 12212 20640 12228 20704
rect 12292 20640 12308 20704
rect 12372 20640 12388 20704
rect 12452 20640 12460 20704
rect 12140 19616 12460 20640
rect 12140 19552 12148 19616
rect 12212 19552 12228 19616
rect 12292 19552 12308 19616
rect 12372 19552 12388 19616
rect 12452 19552 12460 19616
rect 12140 18528 12460 19552
rect 12140 18464 12148 18528
rect 12212 18464 12228 18528
rect 12292 18464 12308 18528
rect 12372 18464 12388 18528
rect 12452 18464 12460 18528
rect 12140 17440 12460 18464
rect 13862 17917 13922 21251
rect 14939 21248 15259 22272
rect 16435 22132 16501 22133
rect 16435 22068 16436 22132
rect 16500 22068 16501 22132
rect 16435 22067 16501 22068
rect 16438 21589 16498 22067
rect 17738 21792 18058 22352
rect 17738 21728 17746 21792
rect 17810 21728 17826 21792
rect 17890 21728 17906 21792
rect 17970 21728 17986 21792
rect 18050 21728 18058 21792
rect 16435 21588 16501 21589
rect 16435 21524 16436 21588
rect 16500 21524 16501 21588
rect 16435 21523 16501 21524
rect 14939 21184 14947 21248
rect 15011 21184 15027 21248
rect 15091 21184 15107 21248
rect 15171 21184 15187 21248
rect 15251 21184 15259 21248
rect 14939 20160 15259 21184
rect 14939 20096 14947 20160
rect 15011 20096 15027 20160
rect 15091 20096 15107 20160
rect 15171 20096 15187 20160
rect 15251 20096 15259 20160
rect 14939 19072 15259 20096
rect 14939 19008 14947 19072
rect 15011 19008 15027 19072
rect 15091 19008 15107 19072
rect 15171 19008 15187 19072
rect 15251 19008 15259 19072
rect 14939 17984 15259 19008
rect 14939 17920 14947 17984
rect 15011 17920 15027 17984
rect 15091 17920 15107 17984
rect 15171 17920 15187 17984
rect 15251 17920 15259 17984
rect 13859 17916 13925 17917
rect 13859 17852 13860 17916
rect 13924 17852 13925 17916
rect 13859 17851 13925 17852
rect 12140 17376 12148 17440
rect 12212 17376 12228 17440
rect 12292 17376 12308 17440
rect 12372 17376 12388 17440
rect 12452 17376 12460 17440
rect 12140 16352 12460 17376
rect 12140 16288 12148 16352
rect 12212 16288 12228 16352
rect 12292 16288 12308 16352
rect 12372 16288 12388 16352
rect 12452 16288 12460 16352
rect 12140 15264 12460 16288
rect 12140 15200 12148 15264
rect 12212 15200 12228 15264
rect 12292 15200 12308 15264
rect 12372 15200 12388 15264
rect 12452 15200 12460 15264
rect 12140 14176 12460 15200
rect 12140 14112 12148 14176
rect 12212 14112 12228 14176
rect 12292 14112 12308 14176
rect 12372 14112 12388 14176
rect 12452 14112 12460 14176
rect 12140 13088 12460 14112
rect 12140 13024 12148 13088
rect 12212 13024 12228 13088
rect 12292 13024 12308 13088
rect 12372 13024 12388 13088
rect 12452 13024 12460 13088
rect 12140 12000 12460 13024
rect 12140 11936 12148 12000
rect 12212 11936 12228 12000
rect 12292 11936 12308 12000
rect 12372 11936 12388 12000
rect 12452 11936 12460 12000
rect 12140 10912 12460 11936
rect 12140 10848 12148 10912
rect 12212 10848 12228 10912
rect 12292 10848 12308 10912
rect 12372 10848 12388 10912
rect 12452 10848 12460 10912
rect 12140 9824 12460 10848
rect 12140 9760 12148 9824
rect 12212 9760 12228 9824
rect 12292 9760 12308 9824
rect 12372 9760 12388 9824
rect 12452 9760 12460 9824
rect 12140 8736 12460 9760
rect 12140 8672 12148 8736
rect 12212 8672 12228 8736
rect 12292 8672 12308 8736
rect 12372 8672 12388 8736
rect 12452 8672 12460 8736
rect 12140 7648 12460 8672
rect 12140 7584 12148 7648
rect 12212 7584 12228 7648
rect 12292 7584 12308 7648
rect 12372 7584 12388 7648
rect 12452 7584 12460 7648
rect 12140 6560 12460 7584
rect 12140 6496 12148 6560
rect 12212 6496 12228 6560
rect 12292 6496 12308 6560
rect 12372 6496 12388 6560
rect 12452 6496 12460 6560
rect 12140 5472 12460 6496
rect 12140 5408 12148 5472
rect 12212 5408 12228 5472
rect 12292 5408 12308 5472
rect 12372 5408 12388 5472
rect 12452 5408 12460 5472
rect 12140 4384 12460 5408
rect 12140 4320 12148 4384
rect 12212 4320 12228 4384
rect 12292 4320 12308 4384
rect 12372 4320 12388 4384
rect 12452 4320 12460 4384
rect 12140 3296 12460 4320
rect 12140 3232 12148 3296
rect 12212 3232 12228 3296
rect 12292 3232 12308 3296
rect 12372 3232 12388 3296
rect 12452 3232 12460 3296
rect 12140 2208 12460 3232
rect 12140 2144 12148 2208
rect 12212 2144 12228 2208
rect 12292 2144 12308 2208
rect 12372 2144 12388 2208
rect 12452 2144 12460 2208
rect 12140 2128 12460 2144
rect 14939 16896 15259 17920
rect 14939 16832 14947 16896
rect 15011 16832 15027 16896
rect 15091 16832 15107 16896
rect 15171 16832 15187 16896
rect 15251 16832 15259 16896
rect 14939 15808 15259 16832
rect 14939 15744 14947 15808
rect 15011 15744 15027 15808
rect 15091 15744 15107 15808
rect 15171 15744 15187 15808
rect 15251 15744 15259 15808
rect 14939 14720 15259 15744
rect 14939 14656 14947 14720
rect 15011 14656 15027 14720
rect 15091 14656 15107 14720
rect 15171 14656 15187 14720
rect 15251 14656 15259 14720
rect 14939 13632 15259 14656
rect 14939 13568 14947 13632
rect 15011 13568 15027 13632
rect 15091 13568 15107 13632
rect 15171 13568 15187 13632
rect 15251 13568 15259 13632
rect 14939 12544 15259 13568
rect 14939 12480 14947 12544
rect 15011 12480 15027 12544
rect 15091 12480 15107 12544
rect 15171 12480 15187 12544
rect 15251 12480 15259 12544
rect 14939 11456 15259 12480
rect 14939 11392 14947 11456
rect 15011 11392 15027 11456
rect 15091 11392 15107 11456
rect 15171 11392 15187 11456
rect 15251 11392 15259 11456
rect 14939 10368 15259 11392
rect 14939 10304 14947 10368
rect 15011 10304 15027 10368
rect 15091 10304 15107 10368
rect 15171 10304 15187 10368
rect 15251 10304 15259 10368
rect 14939 9280 15259 10304
rect 14939 9216 14947 9280
rect 15011 9216 15027 9280
rect 15091 9216 15107 9280
rect 15171 9216 15187 9280
rect 15251 9216 15259 9280
rect 14939 8192 15259 9216
rect 14939 8128 14947 8192
rect 15011 8128 15027 8192
rect 15091 8128 15107 8192
rect 15171 8128 15187 8192
rect 15251 8128 15259 8192
rect 14939 7104 15259 8128
rect 14939 7040 14947 7104
rect 15011 7040 15027 7104
rect 15091 7040 15107 7104
rect 15171 7040 15187 7104
rect 15251 7040 15259 7104
rect 14939 6016 15259 7040
rect 14939 5952 14947 6016
rect 15011 5952 15027 6016
rect 15091 5952 15107 6016
rect 15171 5952 15187 6016
rect 15251 5952 15259 6016
rect 14939 4928 15259 5952
rect 14939 4864 14947 4928
rect 15011 4864 15027 4928
rect 15091 4864 15107 4928
rect 15171 4864 15187 4928
rect 15251 4864 15259 4928
rect 14939 3840 15259 4864
rect 14939 3776 14947 3840
rect 15011 3776 15027 3840
rect 15091 3776 15107 3840
rect 15171 3776 15187 3840
rect 15251 3776 15259 3840
rect 14939 2752 15259 3776
rect 14939 2688 14947 2752
rect 15011 2688 15027 2752
rect 15091 2688 15107 2752
rect 15171 2688 15187 2752
rect 15251 2688 15259 2752
rect 14939 2128 15259 2688
rect 17738 20704 18058 21728
rect 17738 20640 17746 20704
rect 17810 20640 17826 20704
rect 17890 20640 17906 20704
rect 17970 20640 17986 20704
rect 18050 20640 18058 20704
rect 17738 19616 18058 20640
rect 17738 19552 17746 19616
rect 17810 19552 17826 19616
rect 17890 19552 17906 19616
rect 17970 19552 17986 19616
rect 18050 19552 18058 19616
rect 17738 18528 18058 19552
rect 17738 18464 17746 18528
rect 17810 18464 17826 18528
rect 17890 18464 17906 18528
rect 17970 18464 17986 18528
rect 18050 18464 18058 18528
rect 17738 17440 18058 18464
rect 17738 17376 17746 17440
rect 17810 17376 17826 17440
rect 17890 17376 17906 17440
rect 17970 17376 17986 17440
rect 18050 17376 18058 17440
rect 17738 16352 18058 17376
rect 17738 16288 17746 16352
rect 17810 16288 17826 16352
rect 17890 16288 17906 16352
rect 17970 16288 17986 16352
rect 18050 16288 18058 16352
rect 17738 15264 18058 16288
rect 20537 22336 20857 22352
rect 20537 22272 20545 22336
rect 20609 22272 20625 22336
rect 20689 22272 20705 22336
rect 20769 22272 20785 22336
rect 20849 22272 20857 22336
rect 20537 21248 20857 22272
rect 20537 21184 20545 21248
rect 20609 21184 20625 21248
rect 20689 21184 20705 21248
rect 20769 21184 20785 21248
rect 20849 21184 20857 21248
rect 20537 20160 20857 21184
rect 21035 20772 21101 20773
rect 21035 20708 21036 20772
rect 21100 20708 21101 20772
rect 21035 20707 21101 20708
rect 20537 20096 20545 20160
rect 20609 20096 20625 20160
rect 20689 20096 20705 20160
rect 20769 20096 20785 20160
rect 20849 20096 20857 20160
rect 20537 19072 20857 20096
rect 20537 19008 20545 19072
rect 20609 19008 20625 19072
rect 20689 19008 20705 19072
rect 20769 19008 20785 19072
rect 20849 19008 20857 19072
rect 20537 17984 20857 19008
rect 21038 18597 21098 20707
rect 21587 19820 21653 19821
rect 21587 19756 21588 19820
rect 21652 19756 21653 19820
rect 21587 19755 21653 19756
rect 21035 18596 21101 18597
rect 21035 18532 21036 18596
rect 21100 18532 21101 18596
rect 21035 18531 21101 18532
rect 20537 17920 20545 17984
rect 20609 17920 20625 17984
rect 20689 17920 20705 17984
rect 20769 17920 20785 17984
rect 20849 17920 20857 17984
rect 20537 16896 20857 17920
rect 20537 16832 20545 16896
rect 20609 16832 20625 16896
rect 20689 16832 20705 16896
rect 20769 16832 20785 16896
rect 20849 16832 20857 16896
rect 20537 15808 20857 16832
rect 20537 15744 20545 15808
rect 20609 15744 20625 15808
rect 20689 15744 20705 15808
rect 20769 15744 20785 15808
rect 20849 15744 20857 15808
rect 18827 15604 18893 15605
rect 18827 15540 18828 15604
rect 18892 15540 18893 15604
rect 18827 15539 18893 15540
rect 17738 15200 17746 15264
rect 17810 15200 17826 15264
rect 17890 15200 17906 15264
rect 17970 15200 17986 15264
rect 18050 15200 18058 15264
rect 17738 14176 18058 15200
rect 17738 14112 17746 14176
rect 17810 14112 17826 14176
rect 17890 14112 17906 14176
rect 17970 14112 17986 14176
rect 18050 14112 18058 14176
rect 17738 13088 18058 14112
rect 17738 13024 17746 13088
rect 17810 13024 17826 13088
rect 17890 13024 17906 13088
rect 17970 13024 17986 13088
rect 18050 13024 18058 13088
rect 17738 12000 18058 13024
rect 17738 11936 17746 12000
rect 17810 11936 17826 12000
rect 17890 11936 17906 12000
rect 17970 11936 17986 12000
rect 18050 11936 18058 12000
rect 17738 10912 18058 11936
rect 17738 10848 17746 10912
rect 17810 10848 17826 10912
rect 17890 10848 17906 10912
rect 17970 10848 17986 10912
rect 18050 10848 18058 10912
rect 17738 9824 18058 10848
rect 18830 9893 18890 15539
rect 20537 14720 20857 15744
rect 20537 14656 20545 14720
rect 20609 14656 20625 14720
rect 20689 14656 20705 14720
rect 20769 14656 20785 14720
rect 20849 14656 20857 14720
rect 20537 13632 20857 14656
rect 20537 13568 20545 13632
rect 20609 13568 20625 13632
rect 20689 13568 20705 13632
rect 20769 13568 20785 13632
rect 20849 13568 20857 13632
rect 19195 12884 19261 12885
rect 19195 12820 19196 12884
rect 19260 12820 19261 12884
rect 19195 12819 19261 12820
rect 18827 9892 18893 9893
rect 18827 9828 18828 9892
rect 18892 9828 18893 9892
rect 18827 9827 18893 9828
rect 17738 9760 17746 9824
rect 17810 9760 17826 9824
rect 17890 9760 17906 9824
rect 17970 9760 17986 9824
rect 18050 9760 18058 9824
rect 17738 8736 18058 9760
rect 17738 8672 17746 8736
rect 17810 8672 17826 8736
rect 17890 8672 17906 8736
rect 17970 8672 17986 8736
rect 18050 8672 18058 8736
rect 17738 7648 18058 8672
rect 17738 7584 17746 7648
rect 17810 7584 17826 7648
rect 17890 7584 17906 7648
rect 17970 7584 17986 7648
rect 18050 7584 18058 7648
rect 17738 6560 18058 7584
rect 17738 6496 17746 6560
rect 17810 6496 17826 6560
rect 17890 6496 17906 6560
rect 17970 6496 17986 6560
rect 18050 6496 18058 6560
rect 17738 5472 18058 6496
rect 17738 5408 17746 5472
rect 17810 5408 17826 5472
rect 17890 5408 17906 5472
rect 17970 5408 17986 5472
rect 18050 5408 18058 5472
rect 17738 4384 18058 5408
rect 19198 4725 19258 12819
rect 20537 12544 20857 13568
rect 20537 12480 20545 12544
rect 20609 12480 20625 12544
rect 20689 12480 20705 12544
rect 20769 12480 20785 12544
rect 20849 12480 20857 12544
rect 20537 11456 20857 12480
rect 20537 11392 20545 11456
rect 20609 11392 20625 11456
rect 20689 11392 20705 11456
rect 20769 11392 20785 11456
rect 20849 11392 20857 11456
rect 20537 10368 20857 11392
rect 21035 11116 21101 11117
rect 21035 11052 21036 11116
rect 21100 11052 21101 11116
rect 21035 11051 21101 11052
rect 20537 10304 20545 10368
rect 20609 10304 20625 10368
rect 20689 10304 20705 10368
rect 20769 10304 20785 10368
rect 20849 10304 20857 10368
rect 20537 9280 20857 10304
rect 20537 9216 20545 9280
rect 20609 9216 20625 9280
rect 20689 9216 20705 9280
rect 20769 9216 20785 9280
rect 20849 9216 20857 9280
rect 20537 8192 20857 9216
rect 20537 8128 20545 8192
rect 20609 8128 20625 8192
rect 20689 8128 20705 8192
rect 20769 8128 20785 8192
rect 20849 8128 20857 8192
rect 19563 7172 19629 7173
rect 19563 7108 19564 7172
rect 19628 7108 19629 7172
rect 19563 7107 19629 7108
rect 19379 7036 19445 7037
rect 19379 6972 19380 7036
rect 19444 6972 19445 7036
rect 19379 6971 19445 6972
rect 19382 6085 19442 6971
rect 19566 6085 19626 7107
rect 20537 7104 20857 8128
rect 21038 7309 21098 11051
rect 21590 7445 21650 19755
rect 21219 7444 21285 7445
rect 21219 7380 21220 7444
rect 21284 7380 21285 7444
rect 21219 7379 21285 7380
rect 21587 7444 21653 7445
rect 21587 7380 21588 7444
rect 21652 7380 21653 7444
rect 21587 7379 21653 7380
rect 21035 7308 21101 7309
rect 21035 7244 21036 7308
rect 21100 7244 21101 7308
rect 21035 7243 21101 7244
rect 20537 7040 20545 7104
rect 20609 7040 20625 7104
rect 20689 7040 20705 7104
rect 20769 7040 20785 7104
rect 20849 7040 20857 7104
rect 19747 6492 19813 6493
rect 19747 6428 19748 6492
rect 19812 6428 19813 6492
rect 19747 6427 19813 6428
rect 19379 6084 19445 6085
rect 19379 6020 19380 6084
rect 19444 6020 19445 6084
rect 19379 6019 19445 6020
rect 19563 6084 19629 6085
rect 19563 6020 19564 6084
rect 19628 6020 19629 6084
rect 19563 6019 19629 6020
rect 19750 4861 19810 6427
rect 20537 6016 20857 7040
rect 21222 6629 21282 7379
rect 21219 6628 21285 6629
rect 21219 6564 21220 6628
rect 21284 6564 21285 6628
rect 21219 6563 21285 6564
rect 20537 5952 20545 6016
rect 20609 5952 20625 6016
rect 20689 5952 20705 6016
rect 20769 5952 20785 6016
rect 20849 5952 20857 6016
rect 20537 4928 20857 5952
rect 20537 4864 20545 4928
rect 20609 4864 20625 4928
rect 20689 4864 20705 4928
rect 20769 4864 20785 4928
rect 20849 4864 20857 4928
rect 19747 4860 19813 4861
rect 19747 4796 19748 4860
rect 19812 4796 19813 4860
rect 19747 4795 19813 4796
rect 19195 4724 19261 4725
rect 19195 4660 19196 4724
rect 19260 4660 19261 4724
rect 19195 4659 19261 4660
rect 17738 4320 17746 4384
rect 17810 4320 17826 4384
rect 17890 4320 17906 4384
rect 17970 4320 17986 4384
rect 18050 4320 18058 4384
rect 17738 3296 18058 4320
rect 17738 3232 17746 3296
rect 17810 3232 17826 3296
rect 17890 3232 17906 3296
rect 17970 3232 17986 3296
rect 18050 3232 18058 3296
rect 17738 2208 18058 3232
rect 17738 2144 17746 2208
rect 17810 2144 17826 2208
rect 17890 2144 17906 2208
rect 17970 2144 17986 2208
rect 18050 2144 18058 2208
rect 17738 2128 18058 2144
rect 20537 3840 20857 4864
rect 21222 4453 21282 6563
rect 21219 4452 21285 4453
rect 21219 4388 21220 4452
rect 21284 4388 21285 4452
rect 21219 4387 21285 4388
rect 20537 3776 20545 3840
rect 20609 3776 20625 3840
rect 20689 3776 20705 3840
rect 20769 3776 20785 3840
rect 20849 3776 20857 3840
rect 20537 2752 20857 3776
rect 20537 2688 20545 2752
rect 20609 2688 20625 2752
rect 20689 2688 20705 2752
rect 20769 2688 20785 2752
rect 20849 2688 20857 2752
rect 20537 2128 20857 2688
use sky130_fd_sc_hd__diode_2  ANTENNA_Test_en_E_FTB01_A dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 21436 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Test_en_FTB00_A
timestamp 1649977179
transform 1 0 12420 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Test_en_W_FTB01_A
timestamp 1649977179
transform -1 0 2300 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__65__A
timestamp 1649977179
transform 1 0 11684 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__66__A
timestamp 1649977179
transform 1 0 8648 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__68__A
timestamp 1649977179
transform -1 0 11500 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__70__A
timestamp 1649977179
transform -1 0 22816 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__71__A
timestamp 1649977179
transform -1 0 14720 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__73__A
timestamp 1649977179
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__77__A
timestamp 1649977179
transform 1 0 2668 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__78__A
timestamp 1649977179
transform 1 0 3220 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__79__A
timestamp 1649977179
transform 1 0 3496 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__80__A
timestamp 1649977179
transform 1 0 4232 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__81__A
timestamp 1649977179
transform 1 0 3772 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1649977179
transform -1 0 12236 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1649977179
transform -1 0 21988 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1649977179
transform -1 0 1840 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1649977179
transform -1 0 12052 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1649977179
transform -1 0 17204 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1649977179
transform -1 0 19136 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1649977179
transform -1 0 16560 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1649977179
transform -1 0 16928 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1649977179
transform -1 0 18400 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1649977179
transform -1 0 17112 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1649977179
transform -1 0 18584 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1649977179
transform -1 0 18584 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1649977179
transform -1 0 18400 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1649977179
transform -1 0 23184 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1649977179
transform -1 0 16560 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1649977179
transform -1 0 18768 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1649977179
transform -1 0 17940 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1649977179
transform -1 0 18124 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1649977179
transform -1 0 14628 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1649977179
transform -1 0 22816 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1649977179
transform -1 0 5520 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1649977179
transform -1 0 10580 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1649977179
transform 1 0 12420 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1649977179
transform -1 0 14260 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1649977179
transform -1 0 17204 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1649977179
transform -1 0 17940 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1649977179
transform -1 0 14536 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1649977179
transform -1 0 6072 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1649977179
transform -1 0 6256 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1649977179
transform -1 0 11684 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1649977179
transform -1 0 6808 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1649977179
transform -1 0 7268 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1649977179
transform -1 0 8372 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1649977179
transform -1 0 8280 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1649977179
transform -1 0 10028 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1649977179
transform -1 0 9108 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1649977179
transform -1 0 11316 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1649977179
transform 1 0 13524 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 6532 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 4784 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4__CLK
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5__CLK
timestamp 1649977179
transform 1 0 6532 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6__CLK
timestamp 1649977179
transform 1 0 4968 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7__CLK
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8__CLK
timestamp 1649977179
transform 1 0 8280 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9__CLK
timestamp 1649977179
transform 1 0 8464 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10__CLK
timestamp 1649977179
transform 1 0 6992 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11__CLK
timestamp 1649977179
transform 1 0 6532 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12__CLK
timestamp 1649977179
transform 1 0 7176 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13__CLK
timestamp 1649977179
transform 1 0 7820 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14__CLK
timestamp 1649977179
transform 1 0 10672 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15__CLK
timestamp 1649977179
transform 1 0 11960 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16__CLK
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 4600 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 6532 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 9660 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 8464 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 11132 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11132 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 11408 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13064 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 9752 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 8280 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 10764 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 10948 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4__CLK
timestamp 1649977179
transform 1 0 12144 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5__CLK
timestamp 1649977179
transform 1 0 9844 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6__CLK
timestamp 1649977179
transform 1 0 9936 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7__CLK
timestamp 1649977179
transform 1 0 8188 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8__CLK
timestamp 1649977179
transform 1 0 6532 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9__CLK
timestamp 1649977179
transform 1 0 6624 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10__CLK
timestamp 1649977179
transform 1 0 6716 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11__CLK
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12__CLK
timestamp 1649977179
transform 1 0 8464 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13__CLK
timestamp 1649977179
transform 1 0 11408 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14__CLK
timestamp 1649977179
transform 1 0 10580 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15__CLK
timestamp 1649977179
transform 1 0 7820 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16__CLK
timestamp 1649977179
transform 1 0 7544 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 8464 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 6900 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 8188 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 9568 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11132 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 8924 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 7360 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 6992 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 6716 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 6348 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 6900 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4__CLK
timestamp 1649977179
transform 1 0 7820 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5__CLK
timestamp 1649977179
transform 1 0 8188 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6__CLK
timestamp 1649977179
transform 1 0 6532 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7__CLK
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8__CLK
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9__CLK
timestamp 1649977179
transform 1 0 7176 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10__CLK
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11__CLK
timestamp 1649977179
transform 1 0 6532 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12__CLK
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13__CLK
timestamp 1649977179
transform 1 0 6532 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14__CLK
timestamp 1649977179
transform 1 0 7084 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15__CLK
timestamp 1649977179
transform 1 0 6348 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16__CLK
timestamp 1649977179
transform 1 0 12420 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 12420 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13708 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 16100 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 14076 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 16100 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 16192 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 18584 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 18124 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 16284 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 13064 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 11960 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4__CLK
timestamp 1649977179
transform 1 0 12236 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5__CLK
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6__CLK
timestamp 1649977179
transform 1 0 12144 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7__CLK
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8__CLK
timestamp 1649977179
transform 1 0 12972 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9__CLK
timestamp 1649977179
transform 1 0 13156 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10__CLK
timestamp 1649977179
transform 1 0 13616 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11__CLK
timestamp 1649977179
transform 1 0 13708 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12__CLK
timestamp 1649977179
transform 1 0 13800 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13__CLK
timestamp 1649977179
transform 1 0 15548 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14__CLK
timestamp 1649977179
transform 1 0 15732 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15__CLK
timestamp 1649977179
transform 1 0 16376 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16__CLK
timestamp 1649977179
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 16100 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 16468 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 20424 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 20700 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 22632 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13524 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 16744 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
timestamp 1649977179
transform 1 0 9936 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
timestamp 1649977179
transform -1 0 9108 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
timestamp 1649977179
transform 1 0 9568 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
timestamp 1649977179
transform 1 0 9752 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 12972 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 10488 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 11684 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 9108 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4__CLK
timestamp 1649977179
transform 1 0 6716 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5__CLK
timestamp 1649977179
transform 1 0 7084 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6__CLK
timestamp 1649977179
transform 1 0 6808 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7__CLK
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8__CLK
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9__CLK
timestamp 1649977179
transform 1 0 9016 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10__CLK
timestamp 1649977179
transform 1 0 9292 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11__CLK
timestamp 1649977179
transform 1 0 10672 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12__CLK
timestamp 1649977179
transform 1 0 11500 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13__CLK
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14__CLK
timestamp 1649977179
transform 1 0 10488 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15__CLK
timestamp 1649977179
transform 1 0 9200 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16__CLK
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 17204 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 16836 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 16468 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 17296 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 16836 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 16652 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 14812 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1649977179
transform 1 0 13524 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13156 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13064 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 11500 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 11684 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4__CLK
timestamp 1649977179
transform 1 0 13064 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5__CLK
timestamp 1649977179
transform 1 0 14444 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6__CLK
timestamp 1649977179
transform 1 0 13340 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7__CLK
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8__CLK
timestamp 1649977179
transform 1 0 11776 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9__CLK
timestamp 1649977179
transform 1 0 13248 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10__CLK
timestamp 1649977179
transform 1 0 14076 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11__CLK
timestamp 1649977179
transform 1 0 15916 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12__CLK
timestamp 1649977179
transform 1 0 15916 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13__CLK
timestamp 1649977179
transform 1 0 14444 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14__CLK
timestamp 1649977179
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15__CLK
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16__CLK
timestamp 1649977179
transform 1 0 17572 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 17204 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 21528 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 22632 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 22632 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 16192 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 22632 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 15732 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 16100 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 17020 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 16192 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4__CLK
timestamp 1649977179
transform 1 0 14720 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5__CLK
timestamp 1649977179
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6__CLK
timestamp 1649977179
transform 1 0 17020 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7__CLK
timestamp 1649977179
transform 1 0 18492 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8__CLK
timestamp 1649977179
transform 1 0 18124 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9__CLK
timestamp 1649977179
transform 1 0 17756 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10__CLK
timestamp 1649977179
transform 1 0 18584 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11__CLK
timestamp 1649977179
transform 1 0 18124 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12__CLK
timestamp 1649977179
transform 1 0 18032 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13__CLK
timestamp 1649977179
transform 1 0 21528 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14__CLK
timestamp 1649977179
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15__CLK
timestamp 1649977179
transform 1 0 18768 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16__CLK
timestamp 1649977179
transform 1 0 18676 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 23000 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 20332 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 16836 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 19504 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 20332 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 22632 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 17112 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 14812 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 16284 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 16100 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 18124 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4__CLK
timestamp 1649977179
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5__CLK
timestamp 1649977179
transform 1 0 22632 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6__CLK
timestamp 1649977179
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7__CLK
timestamp 1649977179
transform 1 0 21160 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8__CLK
timestamp 1649977179
transform 1 0 23000 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9__CLK
timestamp 1649977179
transform 1 0 22724 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10__CLK
timestamp 1649977179
transform 1 0 18124 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11__CLK
timestamp 1649977179
transform 1 0 17572 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12__CLK
timestamp 1649977179
transform 1 0 17388 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13__CLK
timestamp 1649977179
transform 1 0 23000 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14__CLK
timestamp 1649977179
transform 1 0 14168 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15__CLK
timestamp 1649977179
transform 1 0 22632 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16__CLK
timestamp 1649977179
transform 1 0 16928 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 17112 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 18584 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 14260 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 17572 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 10948 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13892 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 17020 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 13156 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output38_A
timestamp 1649977179
transform 1 0 10672 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output50_A
timestamp 1649977179
transform -1 0 22908 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output54_A
timestamp 1649977179
transform -1 0 21804 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output56_A
timestamp 1649977179
transform -1 0 21988 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output60_A
timestamp 1649977179
transform -1 0 22816 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output68_A
timestamp 1649977179
transform -1 0 13984 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output70_A
timestamp 1649977179
transform -1 0 10948 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output72_A
timestamp 1649977179
transform -1 0 10764 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output74_A
timestamp 1649977179
transform -1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output76_A
timestamp 1649977179
transform -1 0 11132 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_E_FTB01_A
timestamp 1649977179
transform 1 0 22632 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1649977179
transform 1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_N_FTB01_A
timestamp 1649977179
transform 1 0 17388 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_S_FTB01_A
timestamp 1649977179
transform 1 0 21896 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_W_FTB01_A
timestamp 1649977179
transform -1 0 16836 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_repeater101_A
timestamp 1649977179
transform -1 0 16560 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_repeater103_A
timestamp 1649977179
transform 1 0 14260 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2116 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2576 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1649977179
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1649977179
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60
timestamp 1649977179
transform 1 0 6624 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72
timestamp 1649977179
transform 1 0 7728 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_97
timestamp 1649977179
transform 1 0 10028 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_106 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 10856 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1649977179
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1649977179
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1649977179
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1649977179
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_171
timestamp 1649977179
transform 1 0 16836 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_183
timestamp 1649977179
transform 1 0 17940 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 1649977179
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1649977179
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1649977179
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1649977179
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_225
timestamp 1649977179
transform 1 0 21804 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_231
timestamp 1649977179
transform 1 0 22356 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_237
timestamp 1649977179
transform 1 0 22908 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1649977179
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1649977179
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1649977179
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1649977179
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1649977179
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1649977179
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_69
timestamp 1649977179
transform 1 0 7452 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_77 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 8188 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_84
timestamp 1649977179
transform 1 0 8832 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_96
timestamp 1649977179
transform 1 0 9936 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_108
timestamp 1649977179
transform 1 0 11040 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1649977179
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1649977179
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1649977179
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_161
timestamp 1649977179
transform 1 0 15916 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_211
timestamp 1649977179
transform 1 0 20516 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1649977179
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_225
timestamp 1649977179
transform 1 0 21804 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6
timestamp 1649977179
transform 1 0 1656 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_18
timestamp 1649977179
transform 1 0 2760 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1649977179
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1649977179
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1649977179
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1649977179
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1649977179
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1649977179
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1649977179
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1649977179
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1649977179
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1649977179
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1649977179
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_153
timestamp 1649977179
transform 1 0 15180 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_157
timestamp 1649977179
transform 1 0 15548 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_187
timestamp 1649977179
transform 1 0 18308 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_217
timestamp 1649977179
transform 1 0 21068 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1649977179
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1649977179
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1649977179
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1649977179
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1649977179
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1649977179
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1649977179
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1649977179
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1649977179
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1649977179
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1649977179
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1649977179
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_149
timestamp 1649977179
transform 1 0 14812 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_164
timestamp 1649977179
transform 1 0 16192 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1649977179
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1649977179
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1649977179
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1649977179
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1649977179
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1649977179
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_65
timestamp 1649977179
transform 1 0 7084 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_73
timestamp 1649977179
transform 1 0 7820 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_87
timestamp 1649977179
transform 1 0 9108 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_99
timestamp 1649977179
transform 1 0 10212 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_111
timestamp 1649977179
transform 1 0 11316 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_125
timestamp 1649977179
transform 1 0 12604 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_137
timestamp 1649977179
transform 1 0 13708 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_153
timestamp 1649977179
transform 1 0 15180 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_188
timestamp 1649977179
transform 1 0 18400 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_192
timestamp 1649977179
transform 1 0 18768 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_235
timestamp 1649977179
transform 1 0 22724 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1649977179
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1649977179
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1649977179
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1649977179
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1649977179
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1649977179
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_69
timestamp 1649977179
transform 1 0 7452 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_73
timestamp 1649977179
transform 1 0 7820 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_94
timestamp 1649977179
transform 1 0 9752 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_106
timestamp 1649977179
transform 1 0 10856 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_113
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_117
timestamp 1649977179
transform 1 0 11868 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_127
timestamp 1649977179
transform 1 0 12788 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_139
timestamp 1649977179
transform 1 0 13892 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1649977179
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_187
timestamp 1649977179
transform 1 0 18308 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1649977179
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1649977179
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1649977179
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1649977179
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_65
timestamp 1649977179
transform 1 0 7084 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_98
timestamp 1649977179
transform 1 0 10120 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_6_128
timestamp 1649977179
transform 1 0 12880 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_134
timestamp 1649977179
transform 1 0 13432 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_192
timestamp 1649977179
transform 1 0 18768 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1649977179
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1649977179
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_39
timestamp 1649977179
transform 1 0 4692 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_59
timestamp 1649977179
transform 1 0 6532 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_133
timestamp 1649977179
transform 1 0 13340 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_148
timestamp 1649977179
transform 1 0 14720 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1649977179
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_187
timestamp 1649977179
transform 1 0 18308 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1649977179
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1649977179
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_29
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_37
timestamp 1649977179
transform 1 0 4508 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_42
timestamp 1649977179
transform 1 0 4968 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_61
timestamp 1649977179
transform 1 0 6716 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1649977179
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_87
timestamp 1649977179
transform 1 0 9108 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_120
timestamp 1649977179
transform 1 0 12144 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_141
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_222
timestamp 1649977179
transform 1 0 21528 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_15
timestamp 1649977179
transform 1 0 2484 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_23
timestamp 1649977179
transform 1 0 3220 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_106
timestamp 1649977179
transform 1 0 10856 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_109
timestamp 1649977179
transform 1 0 11132 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_113
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_138
timestamp 1649977179
transform 1 0 13800 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_143
timestamp 1649977179
transform 1 0 14260 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1649977179
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1649977179
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_3
timestamp 1649977179
transform 1 0 1380 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_9
timestamp 1649977179
transform 1 0 1932 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_29
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_35
timestamp 1649977179
transform 1 0 4324 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1649977179
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_189
timestamp 1649977179
transform 1 0 18492 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_3
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_61
timestamp 1649977179
transform 1 0 6716 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_115
timestamp 1649977179
transform 1 0 11684 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_134
timestamp 1649977179
transform 1 0 13432 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_142
timestamp 1649977179
transform 1 0 14168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_163
timestamp 1649977179
transform 1 0 16100 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_228
timestamp 1649977179
transform 1 0 22080 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_239
timestamp 1649977179
transform 1 0 23092 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_3
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_9
timestamp 1649977179
transform 1 0 1932 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_29
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_85
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_88
timestamp 1649977179
transform 1 0 9200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_135
timestamp 1649977179
transform 1 0 13524 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1649977179
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_141
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_149
timestamp 1649977179
transform 1 0 14812 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_8
timestamp 1649977179
transform 1 0 1840 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_14
timestamp 1649977179
transform 1 0 2392 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_59
timestamp 1649977179
transform 1 0 6532 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_147
timestamp 1649977179
transform 1 0 14628 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_151
timestamp 1649977179
transform 1 0 14996 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1649977179
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_3
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_11
timestamp 1649977179
transform 1 0 2116 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_44
timestamp 1649977179
transform 1 0 5152 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1649977179
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_93
timestamp 1649977179
transform 1 0 9660 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_132
timestamp 1649977179
transform 1 0 13248 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_138
timestamp 1649977179
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_141
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_178
timestamp 1649977179
transform 1 0 17480 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_227
timestamp 1649977179
transform 1 0 21988 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_15
timestamp 1649977179
transform 1 0 2484 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_15_24
timestamp 1649977179
transform 1 0 3312 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_39
timestamp 1649977179
transform 1 0 4692 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_57
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_63
timestamp 1649977179
transform 1 0 6900 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_117
timestamp 1649977179
transform 1 0 11868 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_209
timestamp 1649977179
transform 1 0 20332 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_15
timestamp 1649977179
transform 1 0 2484 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_29
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_33
timestamp 1649977179
transform 1 0 4140 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_43
timestamp 1649977179
transform 1 0 5060 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_79
timestamp 1649977179
transform 1 0 8372 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1649977179
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_85
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_104
timestamp 1649977179
transform 1 0 10672 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_143
timestamp 1649977179
transform 1 0 14260 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_189
timestamp 1649977179
transform 1 0 18492 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_192
timestamp 1649977179
transform 1 0 18768 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1649977179
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_15
timestamp 1649977179
transform 1 0 2484 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_61
timestamp 1649977179
transform 1 0 6716 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_69
timestamp 1649977179
transform 1 0 7452 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_17_106
timestamp 1649977179
transform 1 0 10856 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_133
timestamp 1649977179
transform 1 0 13340 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_145
timestamp 1649977179
transform 1 0 14444 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_165
timestamp 1649977179
transform 1 0 16284 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_169
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_3
timestamp 1649977179
transform 1 0 1380 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_9
timestamp 1649977179
transform 1 0 1932 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_75
timestamp 1649977179
transform 1 0 8004 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_79
timestamp 1649977179
transform 1 0 8372 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1649977179
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_85
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_90
timestamp 1649977179
transform 1 0 9384 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_94
timestamp 1649977179
transform 1 0 9752 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_117
timestamp 1649977179
transform 1 0 11868 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_123
timestamp 1649977179
transform 1 0 12420 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_143
timestamp 1649977179
transform 1 0 14260 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_147
timestamp 1649977179
transform 1 0 14628 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_150
timestamp 1649977179
transform 1 0 14904 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_162
timestamp 1649977179
transform 1 0 16008 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_183
timestamp 1649977179
transform 1 0 17940 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1649977179
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_46
timestamp 1649977179
transform 1 0 5336 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_54
timestamp 1649977179
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_59
timestamp 1649977179
transform 1 0 6532 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_63
timestamp 1649977179
transform 1 0 6900 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_113
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1649977179
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_3
timestamp 1649977179
transform 1 0 1380 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_7
timestamp 1649977179
transform 1 0 1748 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_13
timestamp 1649977179
transform 1 0 2300 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_25
timestamp 1649977179
transform 1 0 3404 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_29
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_75
timestamp 1649977179
transform 1 0 8004 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1649977179
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_101
timestamp 1649977179
transform 1 0 10396 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_122
timestamp 1649977179
transform 1 0 12328 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_134
timestamp 1649977179
transform 1 0 13432 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_239
timestamp 1649977179
transform 1 0 23092 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_3
timestamp 1649977179
transform 1 0 1380 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_11
timestamp 1649977179
transform 1 0 2116 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_79
timestamp 1649977179
transform 1 0 8372 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_131
timestamp 1649977179
transform 1 0 13156 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_151
timestamp 1649977179
transform 1 0 14996 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_171
timestamp 1649977179
transform 1 0 16836 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_175
timestamp 1649977179
transform 1 0 17204 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_3
timestamp 1649977179
transform 1 0 1380 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_38
timestamp 1649977179
transform 1 0 4600 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_56
timestamp 1649977179
transform 1 0 6256 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_75
timestamp 1649977179
transform 1 0 8004 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1649977179
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_85
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_109
timestamp 1649977179
transform 1 0 11132 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_22_114
timestamp 1649977179
transform 1 0 11592 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_120
timestamp 1649977179
transform 1 0 12144 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1649977179
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_175
timestamp 1649977179
transform 1 0 17204 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_183
timestamp 1649977179
transform 1 0 17940 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_222
timestamp 1649977179
transform 1 0 21528 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1649977179
transform 1 0 1380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_38
timestamp 1649977179
transform 1 0 4600 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_61
timestamp 1649977179
transform 1 0 6716 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_65
timestamp 1649977179
transform 1 0 7084 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_68
timestamp 1649977179
transform 1 0 7360 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_76
timestamp 1649977179
transform 1 0 8096 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_115
timestamp 1649977179
transform 1 0 11684 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_127
timestamp 1649977179
transform 1 0 12788 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1649977179
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_187
timestamp 1649977179
transform 1 0 18308 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_66
timestamp 1649977179
transform 1 0 7176 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1649977179
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_85
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_122
timestamp 1649977179
transform 1 0 12328 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_157
timestamp 1649977179
transform 1 0 15548 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_192
timestamp 1649977179
transform 1 0 18768 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_239
timestamp 1649977179
transform 1 0 23092 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_3
timestamp 1649977179
transform 1 0 1380 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_37
timestamp 1649977179
transform 1 0 4508 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_59
timestamp 1649977179
transform 1 0 6532 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_71
timestamp 1649977179
transform 1 0 7636 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1649977179
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_115
timestamp 1649977179
transform 1 0 11684 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_137
timestamp 1649977179
transform 1 0 13708 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_156
timestamp 1649977179
transform 1 0 15456 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_161
timestamp 1649977179
transform 1 0 15916 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_165
timestamp 1649977179
transform 1 0 16284 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_169
timestamp 1649977179
transform 1 0 16652 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_176
timestamp 1649977179
transform 1 0 17296 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1649977179
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_3
timestamp 1649977179
transform 1 0 1380 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_9
timestamp 1649977179
transform 1 0 1932 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_42
timestamp 1649977179
transform 1 0 4968 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_46
timestamp 1649977179
transform 1 0 5336 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_65
timestamp 1649977179
transform 1 0 7084 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_87
timestamp 1649977179
transform 1 0 9108 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_91
timestamp 1649977179
transform 1 0 9476 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_123
timestamp 1649977179
transform 1 0 12420 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_135
timestamp 1649977179
transform 1 0 13524 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1649977179
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_141
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_147
timestamp 1649977179
transform 1 0 14628 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_166
timestamp 1649977179
transform 1 0 16376 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1649977179
transform 1 0 1380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_7
timestamp 1649977179
transform 1 0 1748 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_23
timestamp 1649977179
transform 1 0 3220 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_33
timestamp 1649977179
transform 1 0 4140 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_37
timestamp 1649977179
transform 1 0 4508 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_59
timestamp 1649977179
transform 1 0 6532 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_63
timestamp 1649977179
transform 1 0 6900 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_113
timestamp 1649977179
transform 1 0 11500 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_143
timestamp 1649977179
transform 1 0 14260 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1649977179
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_3
timestamp 1649977179
transform 1 0 1380 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_72
timestamp 1649977179
transform 1 0 7728 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_76
timestamp 1649977179
transform 1 0 8096 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_79
timestamp 1649977179
transform 1 0 8372 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1649977179
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_85
timestamp 1649977179
transform 1 0 8924 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_125
timestamp 1649977179
transform 1 0 12604 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_135
timestamp 1649977179
transform 1 0 13524 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_189
timestamp 1649977179
transform 1 0 18492 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1649977179
transform 1 0 1380 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_7
timestamp 1649977179
transform 1 0 1748 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_95
timestamp 1649977179
transform 1 0 9844 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_113
timestamp 1649977179
transform 1 0 11500 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_217
timestamp 1649977179
transform 1 0 21068 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_3
timestamp 1649977179
transform 1 0 1380 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_18
timestamp 1649977179
transform 1 0 2760 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_29
timestamp 1649977179
transform 1 0 3772 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_87
timestamp 1649977179
transform 1 0 9108 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_111
timestamp 1649977179
transform 1 0 11316 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_143
timestamp 1649977179
transform 1 0 14260 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_192
timestamp 1649977179
transform 1 0 18768 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 1649977179
transform 1 0 1380 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_7
timestamp 1649977179
transform 1 0 1748 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_17
timestamp 1649977179
transform 1 0 2668 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_37
timestamp 1649977179
transform 1 0 4508 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1649977179
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_63
timestamp 1649977179
transform 1 0 6900 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_66
timestamp 1649977179
transform 1 0 7176 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_70
timestamp 1649977179
transform 1 0 7544 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1649977179
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1649977179
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_15
timestamp 1649977179
transform 1 0 2484 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1649977179
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_82
timestamp 1649977179
transform 1 0 8648 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_85
timestamp 1649977179
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_96
timestamp 1649977179
transform 1 0 9936 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_102
timestamp 1649977179
transform 1 0 10488 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_189
timestamp 1649977179
transform 1 0 18492 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1649977179
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1649977179
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_27
timestamp 1649977179
transform 1 0 3588 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_33
timestamp 1649977179
transform 1 0 4140 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_62
timestamp 1649977179
transform 1 0 6808 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_67
timestamp 1649977179
transform 1 0 7268 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_98
timestamp 1649977179
transform 1 0 10120 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_108
timestamp 1649977179
transform 1 0 11040 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1649977179
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_178
timestamp 1649977179
transform 1 0 17480 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1649977179
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_15
timestamp 1649977179
transform 1 0 2484 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_19
timestamp 1649977179
transform 1 0 2852 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_25
timestamp 1649977179
transform 1 0 3404 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_36
timestamp 1649977179
transform 1 0 4416 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_85
timestamp 1649977179
transform 1 0 8924 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_118
timestamp 1649977179
transform 1 0 11960 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_209
timestamp 1649977179
transform 1 0 20332 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_231
timestamp 1649977179
transform 1 0 22356 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_33
timestamp 1649977179
transform 1 0 4140 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_38
timestamp 1649977179
transform 1 0 4600 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_45
timestamp 1649977179
transform 1 0 5244 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_54
timestamp 1649977179
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_57
timestamp 1649977179
transform 1 0 6348 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_61
timestamp 1649977179
transform 1 0 6716 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_65
timestamp 1649977179
transform 1 0 7084 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_35_106
timestamp 1649977179
transform 1 0 10856 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_125
timestamp 1649977179
transform 1 0 12604 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1649977179
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_199
timestamp 1649977179
transform 1 0 19412 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_36_3
timestamp 1649977179
transform 1 0 1380 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_36_10
timestamp 1649977179
transform 1 0 2024 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_36_17
timestamp 1649977179
transform 1 0 2668 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_24
timestamp 1649977179
transform 1 0 3312 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_33
timestamp 1649977179
transform 1 0 4140 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_45
timestamp 1649977179
transform 1 0 5244 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_51
timestamp 1649977179
transform 1 0 5796 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_96
timestamp 1649977179
transform 1 0 9936 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_100
timestamp 1649977179
transform 1 0 10304 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_116
timestamp 1649977179
transform 1 0 11776 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_169
timestamp 1649977179
transform 1 0 16652 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1649977179
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_197
timestamp 1649977179
transform 1 0 19228 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_206
timestamp 1649977179
transform 1 0 20056 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_229
timestamp 1649977179
transform 1 0 22172 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 23460 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 23460 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 23460 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 23460 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 23460 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 23460 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 23460 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 23460 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 23460 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 23460 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 23460 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 23460 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 23460 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 23460 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 23460 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 23460 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 23460 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 23460 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 23460 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 23460 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 23460 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 23460 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 23460 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 23460 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 23460 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 23460 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 23460 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 23460 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1649977179
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1649977179
transform -1 0 23460 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1649977179
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1649977179
transform -1 0 23460 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1649977179
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1649977179
transform -1 0 23460 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1649977179
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1649977179
transform -1 0 23460 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1649977179
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1649977179
transform -1 0 23460 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1649977179
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1649977179
transform -1 0 23460 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1649977179
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1649977179
transform -1 0 23460 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1649977179
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1649977179
transform -1 0 23460 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1649977179
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1649977179
transform -1 0 23460 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1649977179
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1649977179
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1649977179
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1649977179
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1649977179
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1649977179
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1649977179
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1649977179
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1649977179
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1649977179
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1649977179
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1649977179
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1649977179
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1649977179
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1649977179
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1649977179
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1649977179
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1649977179
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1649977179
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1649977179
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1649977179
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1649977179
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1649977179
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1649977179
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1649977179
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1649977179
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1649977179
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1649977179
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1649977179
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1649977179
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1649977179
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1649977179
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1649977179
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1649977179
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1649977179
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1649977179
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1649977179
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1649977179
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1649977179
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1649977179
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1649977179
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1649977179
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1649977179
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1649977179
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1649977179
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1649977179
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1649977179
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1649977179
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1649977179
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1649977179
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1649977179
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1649977179
transform 1 0 6256 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1649977179
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1649977179
transform 1 0 11408 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1649977179
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1649977179
transform 1 0 16560 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1649977179
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1649977179
transform 1 0 21712 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  Test_en_E_FTB01 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 22540 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  Test_en_FTB00 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 11592 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Test_en_W_FTB01
timestamp 1649977179
transform 1 0 1840 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _65_
timestamp 1649977179
transform 1 0 18860 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _66_
timestamp 1649977179
transform 1 0 8372 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _67_
timestamp 1649977179
transform 1 0 22816 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _68_
timestamp 1649977179
transform -1 0 20332 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _69_
timestamp 1649977179
transform -1 0 19136 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _70_
timestamp 1649977179
transform -1 0 19136 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _71_
timestamp 1649977179
transform -1 0 14352 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _72_
timestamp 1649977179
transform -1 0 17664 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _73_
timestamp 1649977179
transform -1 0 17388 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _74_
timestamp 1649977179
transform -1 0 17112 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _75_
timestamp 1649977179
transform 1 0 2116 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _76_
timestamp 1649977179
transform 1 0 2668 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _77_
timestamp 1649977179
transform 1 0 2392 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _78_
timestamp 1649977179
transform 1 0 2944 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _79_
timestamp 1649977179
transform 1 0 3220 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _80_
timestamp 1649977179
transform 1 0 3956 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _81_
timestamp 1649977179
transform -1 0 3772 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _82_
timestamp 1649977179
transform 1 0 4968 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  clk_0_FTB00
timestamp 1649977179
transform -1 0 17480 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  grid_clb_104 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 6624 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 4784 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1649977179
transform 1 0 9292 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1649977179
transform 1 0 6808 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1649977179
transform -1 0 9660 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1649977179
transform -1 0 11408 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1649977179
transform 1 0 5520 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1649977179
transform 1 0 18308 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input2 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 23184 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1649977179
transform -1 0 1656 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1649977179
transform 1 0 18584 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1649977179
transform -1 0 18308 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1649977179
transform -1 0 18584 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1649977179
transform -1 0 19136 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1649977179
transform -1 0 19044 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1649977179
transform -1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1649977179
transform -1 0 19136 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1649977179
transform -1 0 19136 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1649977179
transform 1 0 22632 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1649977179
transform -1 0 23184 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1649977179
transform 1 0 22908 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1649977179
transform 1 0 22908 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1649977179
transform -1 0 19136 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1649977179
transform -1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1649977179
transform -1 0 17940 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1649977179
transform 1 0 20608 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1649977179
transform -1 0 19136 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1649977179
transform 1 0 5520 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1649977179
transform 1 0 11132 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1649977179
transform 1 0 11868 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1649977179
transform -1 0 13708 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1649977179
transform 1 0 15548 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1649977179
transform 1 0 15824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1649977179
transform 1 0 16100 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1649977179
transform 1 0 6348 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1649977179
transform 1 0 6808 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1649977179
transform 1 0 18768 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1649977179
transform 1 0 7268 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1649977179
transform 1 0 7544 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1649977179
transform 1 0 8280 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1649977179
transform 1 0 8556 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1649977179
transform 1 0 10028 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1649977179
transform 1 0 10580 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1649977179
transform 1 0 10856 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 16008 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1649977179
transform -1 0 9660 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2484 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1649977179
transform 1 0 2024 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1649977179
transform 1 0 2852 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1649977179
transform 1 0 2484 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1649977179
transform 1 0 2852 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1649977179
transform 1 0 3864 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1649977179
transform -1 0 3680 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1649977179
transform -1 0 2484 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1649977179
transform -1 0 2852 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1649977179
transform 1 0 2852 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1649977179
transform -1 0 3680 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1649977179
transform 1 0 2024 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1649977179
transform 1 0 2484 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1649977179
transform 1 0 1840 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1649977179
transform -1 0 2024 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1649977179
transform -1 0 2116 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1649977179
transform -1 0 2024 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1649977179
transform -1 0 2576 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1649977179
transform 1 0 3036 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1649977179
transform -1 0 2852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1649977179
transform 1 0 3956 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1649977179
transform -1 0 6072 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1649977179
transform -1 0 4600 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1649977179
transform 1 0 3312 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 4416 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 4416 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 4784 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 6532 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 3312 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1649977179
transform -1 0 6256 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1649977179
transform -1 0 4784 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1649977179
transform 1 0 3312 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1649977179
transform 1 0 4784 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1649977179
transform 1 0 6808 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1649977179
transform -1 0 8464 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1649977179
transform -1 0 6992 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1649977179
transform -1 0 6256 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1649977179
transform 1 0 4048 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1649977179
transform 1 0 6348 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1649977179
transform 1 0 9200 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1649977179
transform -1 0 11960 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1649977179
transform -1 0 6256 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 4784 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 4784 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1649977179
transform -1 0 3680 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__126
timestamp 1649977179
transform -1 0 4048 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1649977179
transform -1 0 4508 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 8188 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 6992 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 9660 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 11132 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 9936 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 13064 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1649977179
transform -1 0 9936 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0__127
timestamp 1649977179
transform 1 0 10028 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 9200 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1649977179
transform 1 0 8004 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0__128
timestamp 1649977179
transform 1 0 7820 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1649977179
transform 1 0 7360 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1649977179
transform 1 0 15180 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 14720 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0__129
timestamp 1649977179
transform 1 0 15824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1649977179
transform 1 0 8188 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1649977179
transform 1 0 10028 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1649977179
transform 1 0 2852 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1649977179
transform 1 0 4140 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1649977179
transform 1 0 4232 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1649977179
transform 1 0 3956 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1649977179
transform 1 0 4048 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1649977179
transform 1 0 3956 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1649977179
transform 1 0 3128 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1649977179
transform 1 0 2024 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1649977179
transform 1 0 3312 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1649977179
transform 1 0 3128 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1649977179
transform 1 0 2300 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1649977179
transform -1 0 2852 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1649977179
transform 1 0 2576 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1649977179
transform 1 0 2024 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1649977179
transform -1 0 3220 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1649977179
transform -1 0 3312 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1649977179
transform -1 0 2024 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1649977179
transform -1 0 1748 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1649977179
transform 1 0 2576 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1649977179
transform 1 0 2852 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1649977179
transform -1 0 2024 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1649977179
transform 1 0 6440 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1649977179
transform -1 0 5704 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1649977179
transform 1 0 4600 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1649977179
transform 1 0 4232 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1649977179
transform -1 0 6808 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 9844 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 7268 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 8464 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 9936 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1649977179
transform -1 0 9936 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1649977179
transform -1 0 9936 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1649977179
transform -1 0 8188 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1649977179
transform -1 0 6256 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1649977179
transform -1 0 6808 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1649977179
transform -1 0 6716 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1649977179
transform 1 0 4876 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1649977179
transform 1 0 6992 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1649977179
transform -1 0 11408 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1649977179
transform -1 0 10580 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1649977179
transform -1 0 7820 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1649977179
transform 1 0 6072 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 8464 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 6900 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1649977179
transform -1 0 3680 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1649977179
transform -1 0 5428 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__130
timestamp 1649977179
transform -1 0 4784 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 6716 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 7360 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 8464 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 10948 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 8832 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 7360 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1649977179
transform -1 0 9844 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 9108 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0__131
timestamp 1649977179
transform 1 0 10304 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1649977179
transform 1 0 10212 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0__132
timestamp 1649977179
transform 1 0 10580 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1649977179
transform 1 0 8372 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7360 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1649977179
transform -1 0 8004 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0__133
timestamp 1649977179
transform -1 0 7176 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1649977179
transform 1 0 14536 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1649977179
transform 1 0 17848 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1649977179
transform -1 0 4140 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1649977179
transform -1 0 2852 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1649977179
transform 1 0 2852 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1649977179
transform 1 0 2852 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1649977179
transform 1 0 2852 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1649977179
transform 1 0 3680 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1649977179
transform 1 0 2852 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1649977179
transform 1 0 3772 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1649977179
transform 1 0 3772 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1649977179
transform 1 0 2024 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1649977179
transform 1 0 2024 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1649977179
transform 1 0 2852 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1649977179
transform -1 0 2668 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1649977179
transform -1 0 2760 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1649977179
transform -1 0 12604 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1649977179
transform -1 0 12052 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1649977179
transform -1 0 13524 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1649977179
transform -1 0 12420 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1649977179
transform 1 0 2668 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1649977179
transform -1 0 2024 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1649977179
transform -1 0 1748 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1649977179
transform 1 0 2116 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1649977179
transform 1 0 4692 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1649977179
transform -1 0 4140 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1649977179
transform 1 0 6808 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1649977179
transform -1 0 11776 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1649977179
transform -1 0 11408 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 6992 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 5520 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 4600 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 5428 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1649977179
transform -1 0 7820 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1649977179
transform -1 0 8188 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1649977179
transform -1 0 6256 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1649977179
transform 1 0 4876 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1649977179
transform -1 0 6256 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1649977179
transform -1 0 7176 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1649977179
transform -1 0 6256 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1649977179
transform -1 0 5704 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1649977179
transform -1 0 6256 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1649977179
transform -1 0 6164 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1649977179
transform -1 0 6256 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1649977179
transform -1 0 5888 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1649977179
transform -1 0 12420 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 9936 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 12236 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1649977179
transform -1 0 12880 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__134
timestamp 1649977179
transform 1 0 16468 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1649977179
transform -1 0 16836 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 14628 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 12604 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14076 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14720 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 18584 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 18124 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1649977179
transform 1 0 16652 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0__135
timestamp 1649977179
transform 1 0 16744 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 15548 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1649977179
transform 1 0 17664 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1649977179
transform 1 0 17204 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0__136
timestamp 1649977179
transform 1 0 17572 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1649977179
transform 1 0 16836 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 16652 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0__105
timestamp 1649977179
transform -1 0 16560 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1649977179
transform 1 0 20884 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1649977179
transform 1 0 20424 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1649977179
transform 1 0 13248 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1649977179
transform 1 0 12972 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1649977179
transform -1 0 12236 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1649977179
transform -1 0 12420 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1649977179
transform 1 0 12236 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1649977179
transform 1 0 12696 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1649977179
transform 1 0 15548 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1649977179
transform 1 0 14352 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1649977179
transform -1 0 13708 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1649977179
transform 1 0 12880 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1649977179
transform 1 0 12052 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1649977179
transform 1 0 13708 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1649977179
transform -1 0 13432 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1649977179
transform -1 0 13524 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1649977179
transform -1 0 17572 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1649977179
transform 1 0 19136 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1649977179
transform -1 0 18860 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1649977179
transform 1 0 18032 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1649977179
transform 1 0 14076 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1649977179
transform -1 0 11776 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1649977179
transform -1 0 11776 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1649977179
transform 1 0 13708 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1649977179
transform -1 0 13984 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1649977179
transform -1 0 14076 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1649977179
transform 1 0 14260 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1649977179
transform 1 0 17480 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1649977179
transform 1 0 16008 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 16100 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 11592 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 12972 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 11960 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1649977179
transform -1 0 11408 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1649977179
transform -1 0 11316 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1649977179
transform 1 0 9016 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1649977179
transform 1 0 9936 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1649977179
transform 1 0 11040 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1649977179
transform 1 0 12144 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1649977179
transform -1 0 13708 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1649977179
transform 1 0 12512 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1649977179
transform -1 0 15456 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1649977179
transform -1 0 15824 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1649977179
transform 1 0 14076 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14352 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 15548 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1649977179
transform -1 0 18400 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__106
timestamp 1649977179
transform -1 0 19136 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1649977179
transform -1 0 20056 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 15824 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 16652 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 17296 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 19228 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 18952 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 18492 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1649977179
transform 1 0 21804 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 19504 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0__107
timestamp 1649977179
transform -1 0 20056 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1649977179
transform -1 0 21528 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1649977179
transform 1 0 21804 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0__108
timestamp 1649977179
transform -1 0 18584 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1649977179
transform -1 0 21160 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1649977179
transform -1 0 21344 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0__109
timestamp 1649977179
transform -1 0 13984 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1649977179
transform 1 0 20700 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1649977179
transform 1 0 20792 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1649977179
transform 1 0 9568 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1649977179
transform 1 0 8096 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1649977179
transform -1 0 8004 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1649977179
transform -1 0 8096 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1649977179
transform 1 0 8740 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1649977179
transform 1 0 10396 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1649977179
transform 1 0 9844 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1649977179
transform -1 0 8832 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1649977179
transform -1 0 8832 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1649977179
transform -1 0 8740 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1649977179
transform -1 0 9752 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1649977179
transform -1 0 16836 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1649977179
transform -1 0 16192 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1649977179
transform 1 0 21804 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1649977179
transform -1 0 21068 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1649977179
transform -1 0 19136 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1649977179
transform -1 0 21620 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1649977179
transform -1 0 13984 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1649977179
transform -1 0 15088 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1649977179
transform -1 0 15364 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1649977179
transform -1 0 15640 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1649977179
transform 1 0 18584 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1649977179
transform -1 0 23092 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1649977179
transform 1 0 22540 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1649977179
transform -1 0 20792 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1649977179
transform 1 0 21528 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 12972 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 9016 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 11592 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 8464 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1649977179
transform 1 0 6900 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1649977179
transform -1 0 8740 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1649977179
transform 1 0 5888 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1649977179
transform -1 0 8832 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1649977179
transform 1 0 7360 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1649977179
transform 1 0 7544 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1649977179
transform -1 0 9936 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1649977179
transform 1 0 8372 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1649977179
transform 1 0 10028 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1649977179
transform -1 0 11408 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1649977179
transform -1 0 10488 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1649977179
transform 1 0 7728 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1649977179
transform 1 0 12512 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 18860 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 20700 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1649977179
transform 1 0 21804 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__110
timestamp 1649977179
transform -1 0 18584 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1649977179
transform -1 0 21528 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14996 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 15640 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 17020 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 18860 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 16560 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 15088 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1649977179
transform -1 0 22356 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0__111
timestamp 1649977179
transform -1 0 18860 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 22356 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1649977179
transform -1 0 19228 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1649977179
transform -1 0 20884 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0__112
timestamp 1649977179
transform -1 0 20332 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1649977179
transform 1 0 20700 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1649977179
transform -1 0 21344 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0__113
timestamp 1649977179
transform 1 0 21804 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1649977179
transform 1 0 16652 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1649977179
transform -1 0 11224 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1649977179
transform -1 0 10580 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1649977179
transform 1 0 12328 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1649977179
transform 1 0 12052 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1649977179
transform 1 0 12328 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1649977179
transform 1 0 13156 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1649977179
transform -1 0 16468 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1649977179
transform 1 0 17664 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1649977179
transform -1 0 12052 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1649977179
transform -1 0 11408 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1649977179
transform -1 0 12788 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1649977179
transform -1 0 18400 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1649977179
transform 1 0 20240 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1649977179
transform -1 0 20240 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1649977179
transform 1 0 19964 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1649977179
transform -1 0 19964 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1649977179
transform 1 0 18584 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1649977179
transform -1 0 19412 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1649977179
transform -1 0 19136 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1649977179
transform -1 0 19504 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1649977179
transform -1 0 18860 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1649977179
transform -1 0 19136 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1649977179
transform 1 0 22264 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1649977179
transform -1 0 22632 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1649977179
transform 1 0 22540 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1649977179
transform -1 0 19136 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1649977179
transform -1 0 20884 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 12972 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 13064 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 11408 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 10028 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1649977179
transform 1 0 11592 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1649977179
transform -1 0 14444 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1649977179
transform -1 0 13156 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1649977179
transform 1 0 9936 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1649977179
transform 1 0 10948 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1649977179
transform -1 0 13248 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1649977179
transform 1 0 11960 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1649977179
transform 1 0 14444 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1649977179
transform 1 0 14628 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1649977179
transform -1 0 16376 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1649977179
transform 1 0 15088 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1649977179
transform 1 0 16652 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 18860 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 20700 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1649977179
transform 1 0 20056 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__114
timestamp 1649977179
transform -1 0 19136 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 19228 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 16652 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 18124 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 19228 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 19596 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 15732 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 16100 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1649977179
transform -1 0 18400 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1649977179
transform -1 0 20056 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0__115
timestamp 1649977179
transform -1 0 18768 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1649977179
transform -1 0 20056 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1649977179
transform -1 0 21712 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0__116
timestamp 1649977179
transform -1 0 21344 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1649977179
transform 1 0 15640 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 14812 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0__117
timestamp 1649977179
transform 1 0 15364 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1649977179
transform -1 0 18584 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1649977179
transform -1 0 20516 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1649977179
transform -1 0 22540 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1649977179
transform -1 0 22632 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1649977179
transform -1 0 21528 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1649977179
transform -1 0 21528 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1649977179
transform -1 0 22356 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1649977179
transform -1 0 21344 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1649977179
transform -1 0 21528 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1649977179
transform -1 0 21528 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1649977179
transform -1 0 22816 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1649977179
transform 1 0 21804 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1649977179
transform -1 0 23000 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1649977179
transform -1 0 22632 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1649977179
transform -1 0 22908 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1649977179
transform 1 0 22080 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1649977179
transform 1 0 21804 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1649977179
transform 1 0 22908 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1649977179
transform 1 0 21712 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1649977179
transform 1 0 21344 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1649977179
transform 1 0 22908 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1649977179
transform -1 0 22080 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1649977179
transform 1 0 22632 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1649977179
transform 1 0 22908 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1649977179
transform 1 0 22908 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1649977179
transform -1 0 23000 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1649977179
transform 1 0 22632 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1649977179
transform 1 0 22908 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1649977179
transform 1 0 21620 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 15088 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 17020 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 15548 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 12512 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1649977179
transform 1 0 13248 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1649977179
transform 1 0 14720 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1649977179
transform 1 0 15548 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1649977179
transform 1 0 17020 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1649977179
transform -1 0 18124 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1649977179
transform 1 0 16284 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1649977179
transform 1 0 19228 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1649977179
transform 1 0 19044 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1649977179
transform 1 0 19780 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1649977179
transform -1 0 20700 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1649977179
transform 1 0 19228 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1649977179
transform -1 0 20700 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1649977179
transform -1 0 19228 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 18308 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 22172 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1649977179
transform 1 0 20884 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 20700 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__118
timestamp 1649977179
transform 1 0 21068 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 19228 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 20700 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 19228 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 20700 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 19228 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 15640 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1649977179
transform -1 0 21528 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1649977179
transform -1 0 22632 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0__119
timestamp 1649977179
transform -1 0 22264 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1649977179
transform -1 0 21528 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1649977179
transform 1 0 21620 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0__120
timestamp 1649977179
transform 1 0 21988 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1649977179
transform 1 0 18400 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0__121
timestamp 1649977179
transform 1 0 18676 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 17480 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1649977179
transform -1 0 17572 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 17664 0 1 3264
box -38 -48 2062 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1649977179
transform -1 0 21528 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1649977179
transform -1 0 20700 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1649977179
transform -1 0 21528 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1649977179
transform -1 0 22356 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1649977179
transform -1 0 21712 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1649977179
transform -1 0 21528 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1649977179
transform 1 0 21804 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1649977179
transform 1 0 22356 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1649977179
transform -1 0 22632 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1649977179
transform 1 0 22356 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1649977179
transform 1 0 21620 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1649977179
transform -1 0 21712 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1649977179
transform -1 0 22632 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1649977179
transform 1 0 21804 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1649977179
transform -1 0 22632 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1649977179
transform -1 0 22816 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1649977179
transform -1 0 21712 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1649977179
transform -1 0 22908 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1649977179
transform 1 0 22632 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1649977179
transform 1 0 22448 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1649977179
transform -1 0 21712 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1649977179
transform -1 0 21436 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1649977179
transform -1 0 19136 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1649977179
transform -1 0 23000 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1649977179
transform -1 0 18860 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1649977179
transform 1 0 22816 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1649977179
transform 1 0 21528 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 13340 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 14628 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 16652 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1649977179
transform 1 0 18400 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1649977179
transform 1 0 19228 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1649977179
transform -1 0 20884 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1649977179
transform 1 0 19596 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1649977179
transform -1 0 20884 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1649977179
transform 1 0 17940 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1649977179
transform 1 0 19228 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1649977179
transform -1 0 20700 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1649977179
transform 1 0 19780 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1649977179
transform -1 0 22356 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1649977179
transform -1 0 20424 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1649977179
transform 1 0 18124 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1649977179
transform -1 0 19780 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 15640 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 18584 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1649977179
transform 1 0 22356 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__122
timestamp 1649977179
transform 1 0 21988 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 20884 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 16100 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 17848 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 9476 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 12420 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 15548 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 17020 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1649977179
transform -1 0 17480 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0__123
timestamp 1649977179
transform 1 0 18400 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1649977179
transform -1 0 17664 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1649977179
transform -1 0 12328 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0__124
timestamp 1649977179
transform 1 0 14444 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1649977179
transform -1 0 14444 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1649977179
transform -1 0 17480 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0__125
timestamp 1649977179
transform 1 0 18492 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 17480 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  output38 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 10672 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output39
timestamp 1649977179
transform -1 0 18768 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output40
timestamp 1649977179
transform 1 0 22816 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output41
timestamp 1649977179
transform -1 0 1748 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output42
timestamp 1649977179
transform -1 0 2576 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output43
timestamp 1649977179
transform 1 0 22816 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  output44
timestamp 1649977179
transform -1 0 18032 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output45
timestamp 1649977179
transform 1 0 20056 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output46
timestamp 1649977179
transform 1 0 22448 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output47
timestamp 1649977179
transform 1 0 1380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output48
timestamp 1649977179
transform 1 0 22816 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp 1649977179
transform 1 0 22816 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp 1649977179
transform 1 0 22816 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output51
timestamp 1649977179
transform 1 0 22816 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output52
timestamp 1649977179
transform 1 0 22816 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp 1649977179
transform 1 0 22816 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp 1649977179
transform 1 0 22816 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp 1649977179
transform 1 0 22816 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp 1649977179
transform 1 0 22816 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp 1649977179
transform 1 0 22816 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp 1649977179
transform 1 0 22816 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp 1649977179
transform 1 0 22816 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp 1649977179
transform 1 0 22816 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp 1649977179
transform 1 0 22448 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 1649977179
transform 1 0 22448 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp 1649977179
transform 1 0 20332 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1649977179
transform 1 0 19688 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1649977179
transform -1 0 1748 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1649977179
transform 1 0 20148 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 1649977179
transform -1 0 2116 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 1649977179
transform 1 0 21344 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 1649977179
transform -1 0 2024 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1649977179
transform 1 0 21804 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1649977179
transform -1 0 2668 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 1649977179
transform 1 0 22264 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1649977179
transform -1 0 3312 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1649977179
transform 1 0 22816 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1649977179
transform -1 0 4140 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1649977179
transform 1 0 21344 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1649977179
transform 1 0 4232 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1649977179
transform 1 0 19320 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1649977179
transform -1 0 5244 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_E_FTB01 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 22724 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 17848 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_N_FTB01
timestamp 1649977179
transform 1 0 18584 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_S_FTB01
timestamp 1649977179
transform 1 0 22080 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_W_FTB01
timestamp 1649977179
transform -1 0 16560 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  repeater80
timestamp 1649977179
transform 1 0 21252 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater81 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 20700 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  repeater82
timestamp 1649977179
transform -1 0 21620 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater83
timestamp 1649977179
transform 1 0 22080 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  repeater84
timestamp 1649977179
transform -1 0 13800 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater85
timestamp 1649977179
transform -1 0 16468 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater86
timestamp 1649977179
transform -1 0 9568 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater87
timestamp 1649977179
transform 1 0 11224 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  repeater88
timestamp 1649977179
transform -1 0 14168 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater89
timestamp 1649977179
transform -1 0 13984 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  repeater90
timestamp 1649977179
transform -1 0 4968 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater91
timestamp 1649977179
transform -1 0 3312 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  repeater92
timestamp 1649977179
transform -1 0 4876 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater93
timestamp 1649977179
transform -1 0 4600 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  repeater94
timestamp 1649977179
transform -1 0 4968 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater95
timestamp 1649977179
transform -1 0 5336 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  repeater96
timestamp 1649977179
transform 1 0 15272 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater97
timestamp 1649977179
transform 1 0 18032 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater98
timestamp 1649977179
transform 1 0 21344 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater99
timestamp 1649977179
transform 1 0 17940 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  repeater100
timestamp 1649977179
transform 1 0 14536 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater101
timestamp 1649977179
transform -1 0 15272 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater102
timestamp 1649977179
transform 1 0 17664 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater103
timestamp 1649977179
transform 1 0 14444 0 -1 5440
box -38 -48 406 592
<< labels >>
flabel metal2 s 17038 23800 17094 24600 0 FreeSans 224 90 0 0 SC_IN_TOP
port 0 nsew signal input
flabel metal2 s 10230 0 10286 800 0 FreeSans 224 90 0 0 SC_OUT_BOT
port 1 nsew signal tristate
flabel metal2 s 17682 23800 17738 24600 0 FreeSans 224 90 0 0 SC_OUT_TOP
port 2 nsew signal tristate
flabel metal3 s 23800 7896 24600 8016 0 FreeSans 480 0 0 0 Test_en_E_in
port 3 nsew signal input
flabel metal3 s 23800 7352 24600 7472 0 FreeSans 480 0 0 0 Test_en_E_out
port 4 nsew signal tristate
flabel metal3 s 0 21360 800 21480 0 FreeSans 480 0 0 0 Test_en_W_in
port 5 nsew signal input
flabel metal3 s 0 15240 800 15360 0 FreeSans 480 0 0 0 Test_en_W_out
port 6 nsew signal tristate
flabel metal4 s 6542 2128 6862 22352 0 FreeSans 1920 90 0 0 VGND
port 7 nsew ground bidirectional
flabel metal4 s 12140 2128 12460 22352 0 FreeSans 1920 90 0 0 VGND
port 7 nsew ground bidirectional
flabel metal4 s 17738 2128 18058 22352 0 FreeSans 1920 90 0 0 VGND
port 7 nsew ground bidirectional
flabel metal4 s 3743 2128 4063 22352 0 FreeSans 1920 90 0 0 VPWR
port 8 nsew power bidirectional
flabel metal4 s 9341 2128 9661 22352 0 FreeSans 1920 90 0 0 VPWR
port 8 nsew power bidirectional
flabel metal4 s 14939 2128 15259 22352 0 FreeSans 1920 90 0 0 VPWR
port 8 nsew power bidirectional
flabel metal4 s 20537 2128 20857 22352 0 FreeSans 1920 90 0 0 VPWR
port 8 nsew power bidirectional
flabel metal2 s 2134 0 2190 800 0 FreeSans 224 90 0 0 bottom_width_0_height_0__pin_50_
port 9 nsew signal tristate
flabel metal2 s 6182 0 6238 800 0 FreeSans 224 90 0 0 bottom_width_0_height_0__pin_51_
port 10 nsew signal tristate
flabel metal3 s 0 9120 800 9240 0 FreeSans 480 0 0 0 ccff_head
port 11 nsew signal input
flabel metal3 s 23800 6808 24600 6928 0 FreeSans 480 0 0 0 ccff_tail
port 12 nsew signal tristate
flabel metal2 s 18326 23800 18382 24600 0 FreeSans 224 90 0 0 clk_0_N_in
port 13 nsew signal input
flabel metal2 s 14278 0 14334 800 0 FreeSans 224 90 0 0 clk_0_S_in
port 14 nsew signal input
flabel metal3 s 23800 8984 24600 9104 0 FreeSans 480 0 0 0 prog_clk_0_E_out
port 15 nsew signal tristate
flabel metal3 s 23800 8440 24600 8560 0 FreeSans 480 0 0 0 prog_clk_0_N_in
port 16 nsew signal input
flabel metal2 s 18970 23800 19026 24600 0 FreeSans 224 90 0 0 prog_clk_0_N_out
port 17 nsew signal tristate
flabel metal2 s 18326 0 18382 800 0 FreeSans 224 90 0 0 prog_clk_0_S_in
port 18 nsew signal input
flabel metal2 s 22374 0 22430 800 0 FreeSans 224 90 0 0 prog_clk_0_S_out
port 19 nsew signal tristate
flabel metal3 s 0 3000 800 3120 0 FreeSans 480 0 0 0 prog_clk_0_W_out
port 20 nsew signal tristate
flabel metal3 s 23800 9528 24600 9648 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_16_
port 21 nsew signal input
flabel metal3 s 23800 10072 24600 10192 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_17_
port 22 nsew signal input
flabel metal3 s 23800 10616 24600 10736 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_18_
port 23 nsew signal input
flabel metal3 s 23800 11160 24600 11280 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_19_
port 24 nsew signal input
flabel metal3 s 23800 11704 24600 11824 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_20_
port 25 nsew signal input
flabel metal3 s 23800 12248 24600 12368 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_21_
port 26 nsew signal input
flabel metal3 s 23800 12792 24600 12912 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_22_
port 27 nsew signal input
flabel metal3 s 23800 13336 24600 13456 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_23_
port 28 nsew signal input
flabel metal3 s 23800 13880 24600 14000 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_24_
port 29 nsew signal input
flabel metal3 s 23800 14424 24600 14544 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_25_
port 30 nsew signal input
flabel metal3 s 23800 14968 24600 15088 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_26_
port 31 nsew signal input
flabel metal3 s 23800 15512 24600 15632 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_27_
port 32 nsew signal input
flabel metal3 s 23800 16056 24600 16176 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_28_
port 33 nsew signal input
flabel metal3 s 23800 16600 24600 16720 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_29_
port 34 nsew signal input
flabel metal3 s 23800 17144 24600 17264 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_30_
port 35 nsew signal input
flabel metal3 s 23800 17688 24600 17808 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_31_
port 36 nsew signal input
flabel metal3 s 23800 2456 24600 2576 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_42_lower
port 37 nsew signal tristate
flabel metal3 s 23800 18232 24600 18352 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_42_upper
port 38 nsew signal tristate
flabel metal3 s 23800 3000 24600 3120 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_43_lower
port 39 nsew signal tristate
flabel metal3 s 23800 18776 24600 18896 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_43_upper
port 40 nsew signal tristate
flabel metal3 s 23800 3544 24600 3664 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_44_lower
port 41 nsew signal tristate
flabel metal3 s 23800 19320 24600 19440 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_44_upper
port 42 nsew signal tristate
flabel metal3 s 23800 4088 24600 4208 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_45_lower
port 43 nsew signal tristate
flabel metal3 s 23800 19864 24600 19984 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_45_upper
port 44 nsew signal tristate
flabel metal3 s 23800 4632 24600 4752 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_46_lower
port 45 nsew signal tristate
flabel metal3 s 23800 20408 24600 20528 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_46_upper
port 46 nsew signal tristate
flabel metal3 s 23800 5176 24600 5296 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_47_lower
port 47 nsew signal tristate
flabel metal3 s 23800 20952 24600 21072 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_47_upper
port 48 nsew signal tristate
flabel metal3 s 23800 5720 24600 5840 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_48_lower
port 49 nsew signal tristate
flabel metal3 s 23800 21496 24600 21616 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_48_upper
port 50 nsew signal tristate
flabel metal3 s 23800 6264 24600 6384 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_49_lower
port 51 nsew signal tristate
flabel metal3 s 23800 22040 24600 22160 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_49_upper
port 52 nsew signal tristate
flabel metal2 s 5446 23800 5502 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_0_
port 53 nsew signal input
flabel metal2 s 11886 23800 11942 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_10_
port 54 nsew signal input
flabel metal2 s 12530 23800 12586 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_11_
port 55 nsew signal input
flabel metal2 s 13174 23800 13230 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_12_
port 56 nsew signal input
flabel metal2 s 13818 23800 13874 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_13_
port 57 nsew signal input
flabel metal2 s 14462 23800 14518 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_14_
port 58 nsew signal input
flabel metal2 s 15106 23800 15162 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_15_
port 59 nsew signal input
flabel metal2 s 6090 23800 6146 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_1_
port 60 nsew signal input
flabel metal2 s 6734 23800 6790 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_2_
port 61 nsew signal input
flabel metal2 s 15750 23800 15806 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_32_
port 62 nsew signal input
flabel metal2 s 16394 23800 16450 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_33_
port 63 nsew signal input
flabel metal2 s 19614 23800 19670 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_34_lower
port 64 nsew signal tristate
flabel metal2 s 294 23800 350 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_34_upper
port 65 nsew signal tristate
flabel metal2 s 20258 23800 20314 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_35_lower
port 66 nsew signal tristate
flabel metal2 s 938 23800 994 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_35_upper
port 67 nsew signal tristate
flabel metal2 s 20902 23800 20958 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_36_lower
port 68 nsew signal tristate
flabel metal2 s 1582 23800 1638 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_36_upper
port 69 nsew signal tristate
flabel metal2 s 21546 23800 21602 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_37_lower
port 70 nsew signal tristate
flabel metal2 s 2226 23800 2282 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_37_upper
port 71 nsew signal tristate
flabel metal2 s 22190 23800 22246 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_38_lower
port 72 nsew signal tristate
flabel metal2 s 2870 23800 2926 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_38_upper
port 73 nsew signal tristate
flabel metal2 s 22834 23800 22890 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_39_lower
port 74 nsew signal tristate
flabel metal2 s 3514 23800 3570 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_39_upper
port 75 nsew signal tristate
flabel metal2 s 7378 23800 7434 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_3_
port 76 nsew signal input
flabel metal2 s 23478 23800 23534 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_40_lower
port 77 nsew signal tristate
flabel metal2 s 4158 23800 4214 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_40_upper
port 78 nsew signal tristate
flabel metal2 s 24122 23800 24178 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_41_lower
port 79 nsew signal tristate
flabel metal2 s 4802 23800 4858 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_41_upper
port 80 nsew signal tristate
flabel metal2 s 8022 23800 8078 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_4_
port 81 nsew signal input
flabel metal2 s 8666 23800 8722 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_5_
port 82 nsew signal input
flabel metal2 s 9310 23800 9366 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_6_
port 83 nsew signal input
flabel metal2 s 9954 23800 10010 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_7_
port 84 nsew signal input
flabel metal2 s 10598 23800 10654 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_8_
port 85 nsew signal input
flabel metal2 s 11242 23800 11298 24600 0 FreeSans 224 90 0 0 top_width_0_height_0__pin_9_
port 86 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 24600 24600
<< end >>
