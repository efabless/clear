magic
tech sky130A
magscale 1 2
timestamp 1680090092
<< obsli1 >>
rect 368 2159 494592 540753
<< obsm1 >>
rect 368 2048 494592 540784
<< metal2 >>
rect 6734 542200 6790 543000
rect 11150 542200 11206 543000
rect 15566 542200 15622 543000
rect 19982 542200 20038 543000
rect 24398 542200 24454 543000
rect 28814 542200 28870 543000
rect 33230 542200 33286 543000
rect 37646 542200 37702 543000
rect 42062 542200 42118 543000
rect 46478 542200 46534 543000
rect 50894 542200 50950 543000
rect 55310 542200 55366 543000
rect 59726 542200 59782 543000
rect 64142 542200 64198 543000
rect 68558 542200 68614 543000
rect 72974 542200 73030 543000
rect 77390 542200 77446 543000
rect 81806 542200 81862 543000
rect 86222 542200 86278 543000
rect 90638 542200 90694 543000
rect 95054 542200 95110 543000
rect 99470 542200 99526 543000
rect 103886 542200 103942 543000
rect 108302 542200 108358 543000
rect 112718 542200 112774 543000
rect 117134 542200 117190 543000
rect 121550 542200 121606 543000
rect 125966 542200 126022 543000
rect 130382 542200 130438 543000
rect 134798 542200 134854 543000
rect 139214 542200 139270 543000
rect 143630 542200 143686 543000
rect 148046 542200 148102 543000
rect 152462 542200 152518 543000
rect 156878 542200 156934 543000
rect 161294 542200 161350 543000
rect 165710 542200 165766 543000
rect 170126 542200 170182 543000
rect 174542 542200 174598 543000
rect 178958 542200 179014 543000
rect 183374 542200 183430 543000
rect 187790 542200 187846 543000
rect 192206 542200 192262 543000
rect 196622 542200 196678 543000
rect 201038 542200 201094 543000
rect 205454 542200 205510 543000
rect 209870 542200 209926 543000
rect 214286 542200 214342 543000
rect 218702 542200 218758 543000
rect 223118 542200 223174 543000
rect 227534 542200 227590 543000
rect 231950 542200 232006 543000
rect 236366 542200 236422 543000
rect 240782 542200 240838 543000
rect 245198 542200 245254 543000
rect 249614 542200 249670 543000
rect 254030 542200 254086 543000
rect 258446 542200 258502 543000
rect 262862 542200 262918 543000
rect 267278 542200 267334 543000
rect 271694 542200 271750 543000
rect 276110 542200 276166 543000
rect 280526 542200 280582 543000
rect 284942 542200 284998 543000
rect 289358 542200 289414 543000
rect 293774 542200 293830 543000
rect 298190 542200 298246 543000
rect 302606 542200 302662 543000
rect 307022 542200 307078 543000
rect 311438 542200 311494 543000
rect 315854 542200 315910 543000
rect 320270 542200 320326 543000
rect 324686 542200 324742 543000
rect 329102 542200 329158 543000
rect 333518 542200 333574 543000
rect 337934 542200 337990 543000
rect 342350 542200 342406 543000
rect 346766 542200 346822 543000
rect 351182 542200 351238 543000
rect 355598 542200 355654 543000
rect 360014 542200 360070 543000
rect 364430 542200 364486 543000
rect 368846 542200 368902 543000
rect 373262 542200 373318 543000
rect 377678 542200 377734 543000
rect 382094 542200 382150 543000
rect 386510 542200 386566 543000
rect 390926 542200 390982 543000
rect 395342 542200 395398 543000
rect 399758 542200 399814 543000
rect 404174 542200 404230 543000
rect 408590 542200 408646 543000
rect 413006 542200 413062 543000
rect 417422 542200 417478 543000
rect 421838 542200 421894 543000
rect 426254 542200 426310 543000
rect 430670 542200 430726 543000
rect 435086 542200 435142 543000
rect 439502 542200 439558 543000
rect 443918 542200 443974 543000
rect 448334 542200 448390 543000
rect 452750 542200 452806 543000
rect 457166 542200 457222 543000
rect 461582 542200 461638 543000
rect 465998 542200 466054 543000
rect 470414 542200 470470 543000
rect 474830 542200 474886 543000
rect 479246 542200 479302 543000
rect 483662 542200 483718 543000
rect 488078 542200 488134 543000
rect 3974 0 4030 800
rect 9770 0 9826 800
rect 15566 0 15622 800
rect 21362 0 21418 800
rect 27158 0 27214 800
rect 32954 0 33010 800
rect 38750 0 38806 800
rect 44546 0 44602 800
rect 50342 0 50398 800
rect 56138 0 56194 800
rect 61934 0 61990 800
rect 67730 0 67786 800
rect 73526 0 73582 800
rect 79322 0 79378 800
rect 85118 0 85174 800
rect 90914 0 90970 800
rect 96710 0 96766 800
rect 102506 0 102562 800
rect 108302 0 108358 800
rect 114098 0 114154 800
rect 119894 0 119950 800
rect 125690 0 125746 800
rect 131486 0 131542 800
rect 137282 0 137338 800
rect 143078 0 143134 800
rect 148874 0 148930 800
rect 154670 0 154726 800
rect 160466 0 160522 800
rect 166262 0 166318 800
rect 172058 0 172114 800
rect 177854 0 177910 800
rect 183650 0 183706 800
rect 189446 0 189502 800
rect 195242 0 195298 800
rect 201038 0 201094 800
rect 206834 0 206890 800
rect 212630 0 212686 800
rect 218426 0 218482 800
rect 224222 0 224278 800
rect 230018 0 230074 800
rect 235814 0 235870 800
rect 241610 0 241666 800
rect 247406 0 247462 800
rect 253202 0 253258 800
rect 258998 0 259054 800
rect 264794 0 264850 800
rect 270590 0 270646 800
rect 276386 0 276442 800
rect 282182 0 282238 800
rect 287978 0 288034 800
rect 293774 0 293830 800
rect 299570 0 299626 800
rect 305366 0 305422 800
rect 311162 0 311218 800
rect 316958 0 317014 800
rect 322754 0 322810 800
rect 328550 0 328606 800
rect 334346 0 334402 800
rect 340142 0 340198 800
rect 345938 0 345994 800
rect 351734 0 351790 800
rect 357530 0 357586 800
rect 363326 0 363382 800
rect 369122 0 369178 800
rect 374918 0 374974 800
rect 380714 0 380770 800
rect 386510 0 386566 800
rect 392306 0 392362 800
rect 398102 0 398158 800
rect 403898 0 403954 800
rect 409694 0 409750 800
rect 415490 0 415546 800
rect 421286 0 421342 800
rect 427082 0 427138 800
rect 432878 0 432934 800
rect 438674 0 438730 800
rect 444470 0 444526 800
rect 450266 0 450322 800
rect 456062 0 456118 800
rect 461858 0 461914 800
rect 467654 0 467710 800
rect 473450 0 473506 800
rect 479246 0 479302 800
rect 485042 0 485098 800
rect 490838 0 490894 800
<< obsm2 >>
rect 756 542144 6678 542314
rect 6846 542144 11094 542314
rect 11262 542144 15510 542314
rect 15678 542144 19926 542314
rect 20094 542144 24342 542314
rect 24510 542144 28758 542314
rect 28926 542144 33174 542314
rect 33342 542144 37590 542314
rect 37758 542144 42006 542314
rect 42174 542144 46422 542314
rect 46590 542144 50838 542314
rect 51006 542144 55254 542314
rect 55422 542144 59670 542314
rect 59838 542144 64086 542314
rect 64254 542144 68502 542314
rect 68670 542144 72918 542314
rect 73086 542144 77334 542314
rect 77502 542144 81750 542314
rect 81918 542144 86166 542314
rect 86334 542144 90582 542314
rect 90750 542144 94998 542314
rect 95166 542144 99414 542314
rect 99582 542144 103830 542314
rect 103998 542144 108246 542314
rect 108414 542144 112662 542314
rect 112830 542144 117078 542314
rect 117246 542144 121494 542314
rect 121662 542144 125910 542314
rect 126078 542144 130326 542314
rect 130494 542144 134742 542314
rect 134910 542144 139158 542314
rect 139326 542144 143574 542314
rect 143742 542144 147990 542314
rect 148158 542144 152406 542314
rect 152574 542144 156822 542314
rect 156990 542144 161238 542314
rect 161406 542144 165654 542314
rect 165822 542144 170070 542314
rect 170238 542144 174486 542314
rect 174654 542144 178902 542314
rect 179070 542144 183318 542314
rect 183486 542144 187734 542314
rect 187902 542144 192150 542314
rect 192318 542144 196566 542314
rect 196734 542144 200982 542314
rect 201150 542144 205398 542314
rect 205566 542144 209814 542314
rect 209982 542144 214230 542314
rect 214398 542144 218646 542314
rect 218814 542144 223062 542314
rect 223230 542144 227478 542314
rect 227646 542144 231894 542314
rect 232062 542144 236310 542314
rect 236478 542144 240726 542314
rect 240894 542144 245142 542314
rect 245310 542144 249558 542314
rect 249726 542144 253974 542314
rect 254142 542144 258390 542314
rect 258558 542144 262806 542314
rect 262974 542144 267222 542314
rect 267390 542144 271638 542314
rect 271806 542144 276054 542314
rect 276222 542144 280470 542314
rect 280638 542144 284886 542314
rect 285054 542144 289302 542314
rect 289470 542144 293718 542314
rect 293886 542144 298134 542314
rect 298302 542144 302550 542314
rect 302718 542144 306966 542314
rect 307134 542144 311382 542314
rect 311550 542144 315798 542314
rect 315966 542144 320214 542314
rect 320382 542144 324630 542314
rect 324798 542144 329046 542314
rect 329214 542144 333462 542314
rect 333630 542144 337878 542314
rect 338046 542144 342294 542314
rect 342462 542144 346710 542314
rect 346878 542144 351126 542314
rect 351294 542144 355542 542314
rect 355710 542144 359958 542314
rect 360126 542144 364374 542314
rect 364542 542144 368790 542314
rect 368958 542144 373206 542314
rect 373374 542144 377622 542314
rect 377790 542144 382038 542314
rect 382206 542144 386454 542314
rect 386622 542144 390870 542314
rect 391038 542144 395286 542314
rect 395454 542144 399702 542314
rect 399870 542144 404118 542314
rect 404286 542144 408534 542314
rect 408702 542144 412950 542314
rect 413118 542144 417366 542314
rect 417534 542144 421782 542314
rect 421950 542144 426198 542314
rect 426366 542144 430614 542314
rect 430782 542144 435030 542314
rect 435198 542144 439446 542314
rect 439614 542144 443862 542314
rect 444030 542144 448278 542314
rect 448446 542144 452694 542314
rect 452862 542144 457110 542314
rect 457278 542144 461526 542314
rect 461694 542144 465942 542314
rect 466110 542144 470358 542314
rect 470526 542144 474774 542314
rect 474942 542144 479190 542314
rect 479358 542144 483606 542314
rect 483774 542144 488022 542314
rect 488190 542144 494204 542314
rect 756 856 494204 542144
rect 756 734 3918 856
rect 4086 734 9714 856
rect 9882 734 15510 856
rect 15678 734 21306 856
rect 21474 734 27102 856
rect 27270 734 32898 856
rect 33066 734 38694 856
rect 38862 734 44490 856
rect 44658 734 50286 856
rect 50454 734 56082 856
rect 56250 734 61878 856
rect 62046 734 67674 856
rect 67842 734 73470 856
rect 73638 734 79266 856
rect 79434 734 85062 856
rect 85230 734 90858 856
rect 91026 734 96654 856
rect 96822 734 102450 856
rect 102618 734 108246 856
rect 108414 734 114042 856
rect 114210 734 119838 856
rect 120006 734 125634 856
rect 125802 734 131430 856
rect 131598 734 137226 856
rect 137394 734 143022 856
rect 143190 734 148818 856
rect 148986 734 154614 856
rect 154782 734 160410 856
rect 160578 734 166206 856
rect 166374 734 172002 856
rect 172170 734 177798 856
rect 177966 734 183594 856
rect 183762 734 189390 856
rect 189558 734 195186 856
rect 195354 734 200982 856
rect 201150 734 206778 856
rect 206946 734 212574 856
rect 212742 734 218370 856
rect 218538 734 224166 856
rect 224334 734 229962 856
rect 230130 734 235758 856
rect 235926 734 241554 856
rect 241722 734 247350 856
rect 247518 734 253146 856
rect 253314 734 258942 856
rect 259110 734 264738 856
rect 264906 734 270534 856
rect 270702 734 276330 856
rect 276498 734 282126 856
rect 282294 734 287922 856
rect 288090 734 293718 856
rect 293886 734 299514 856
rect 299682 734 305310 856
rect 305478 734 311106 856
rect 311274 734 316902 856
rect 317070 734 322698 856
rect 322866 734 328494 856
rect 328662 734 334290 856
rect 334458 734 340086 856
rect 340254 734 345882 856
rect 346050 734 351678 856
rect 351846 734 357474 856
rect 357642 734 363270 856
rect 363438 734 369066 856
rect 369234 734 374862 856
rect 375030 734 380658 856
rect 380826 734 386454 856
rect 386622 734 392250 856
rect 392418 734 398046 856
rect 398214 734 403842 856
rect 404010 734 409638 856
rect 409806 734 415434 856
rect 415602 734 421230 856
rect 421398 734 427026 856
rect 427194 734 432822 856
rect 432990 734 438618 856
rect 438786 734 444414 856
rect 444582 734 450210 856
rect 450378 734 456006 856
rect 456174 734 461802 856
rect 461970 734 467598 856
rect 467766 734 473394 856
rect 473562 734 479190 856
rect 479358 734 484986 856
rect 485154 734 490782 856
rect 490950 734 494204 856
<< metal3 >>
rect 0 537888 800 538008
rect 494200 533944 495000 534064
rect 0 532448 800 532568
rect 494200 528640 495000 528760
rect 0 527008 800 527128
rect 494200 523336 495000 523456
rect 0 521568 800 521688
rect 494200 518032 495000 518152
rect 0 516128 800 516248
rect 494200 512728 495000 512848
rect 0 510688 800 510808
rect 494200 507424 495000 507544
rect 0 505248 800 505368
rect 494200 502120 495000 502240
rect 0 499808 800 499928
rect 494200 496816 495000 496936
rect 0 494368 800 494488
rect 494200 491512 495000 491632
rect 0 488928 800 489048
rect 494200 486208 495000 486328
rect 0 483488 800 483608
rect 494200 480904 495000 481024
rect 0 478048 800 478168
rect 494200 475600 495000 475720
rect 0 472608 800 472728
rect 494200 470296 495000 470416
rect 0 467168 800 467288
rect 494200 464992 495000 465112
rect 0 461728 800 461848
rect 494200 459688 495000 459808
rect 0 456288 800 456408
rect 494200 454384 495000 454504
rect 0 450848 800 450968
rect 494200 449080 495000 449200
rect 0 445408 800 445528
rect 494200 443776 495000 443896
rect 0 439968 800 440088
rect 494200 438472 495000 438592
rect 0 434528 800 434648
rect 494200 433168 495000 433288
rect 0 429088 800 429208
rect 494200 427864 495000 427984
rect 0 423648 800 423768
rect 494200 422560 495000 422680
rect 0 418208 800 418328
rect 494200 417256 495000 417376
rect 0 412768 800 412888
rect 494200 411952 495000 412072
rect 0 407328 800 407448
rect 494200 406648 495000 406768
rect 0 401888 800 402008
rect 494200 401344 495000 401464
rect 0 396448 800 396568
rect 494200 396040 495000 396160
rect 0 391008 800 391128
rect 494200 390736 495000 390856
rect 0 385568 800 385688
rect 494200 385432 495000 385552
rect 0 380128 800 380248
rect 494200 380128 495000 380248
rect 0 374688 800 374808
rect 494200 374824 495000 374944
rect 494200 369520 495000 369640
rect 0 369248 800 369368
rect 494200 364216 495000 364336
rect 0 363808 800 363928
rect 494200 358912 495000 359032
rect 0 358368 800 358488
rect 494200 353608 495000 353728
rect 0 352928 800 353048
rect 494200 348304 495000 348424
rect 0 347488 800 347608
rect 494200 343000 495000 343120
rect 0 342048 800 342168
rect 494200 337696 495000 337816
rect 0 336608 800 336728
rect 494200 332392 495000 332512
rect 0 331168 800 331288
rect 494200 327088 495000 327208
rect 0 325728 800 325848
rect 494200 321784 495000 321904
rect 0 320288 800 320408
rect 494200 316480 495000 316600
rect 0 314848 800 314968
rect 494200 311176 495000 311296
rect 0 309408 800 309528
rect 494200 305872 495000 305992
rect 0 303968 800 304088
rect 494200 300568 495000 300688
rect 0 298528 800 298648
rect 494200 295264 495000 295384
rect 0 293088 800 293208
rect 494200 289960 495000 290080
rect 0 287648 800 287768
rect 494200 284656 495000 284776
rect 0 282208 800 282328
rect 494200 279352 495000 279472
rect 0 276768 800 276888
rect 494200 274048 495000 274168
rect 0 271328 800 271448
rect 494200 268744 495000 268864
rect 0 265888 800 266008
rect 494200 263440 495000 263560
rect 0 260448 800 260568
rect 494200 258136 495000 258256
rect 0 255008 800 255128
rect 494200 252832 495000 252952
rect 0 249568 800 249688
rect 494200 247528 495000 247648
rect 0 244128 800 244248
rect 494200 242224 495000 242344
rect 0 238688 800 238808
rect 494200 236920 495000 237040
rect 0 233248 800 233368
rect 494200 231616 495000 231736
rect 0 227808 800 227928
rect 494200 226312 495000 226432
rect 0 222368 800 222488
rect 494200 221008 495000 221128
rect 0 216928 800 217048
rect 494200 215704 495000 215824
rect 0 211488 800 211608
rect 494200 210400 495000 210520
rect 0 206048 800 206168
rect 494200 205096 495000 205216
rect 0 200608 800 200728
rect 494200 199792 495000 199912
rect 0 195168 800 195288
rect 494200 194488 495000 194608
rect 0 189728 800 189848
rect 494200 189184 495000 189304
rect 0 184288 800 184408
rect 494200 183880 495000 184000
rect 0 178848 800 178968
rect 494200 178576 495000 178696
rect 0 173408 800 173528
rect 494200 173272 495000 173392
rect 0 167968 800 168088
rect 494200 167968 495000 168088
rect 0 162528 800 162648
rect 494200 162664 495000 162784
rect 494200 157360 495000 157480
rect 0 157088 800 157208
rect 494200 152056 495000 152176
rect 0 151648 800 151768
rect 494200 146752 495000 146872
rect 0 146208 800 146328
rect 494200 141448 495000 141568
rect 0 140768 800 140888
rect 494200 136144 495000 136264
rect 0 135328 800 135448
rect 494200 130840 495000 130960
rect 0 129888 800 130008
rect 494200 125536 495000 125656
rect 0 124448 800 124568
rect 494200 120232 495000 120352
rect 0 119008 800 119128
rect 494200 114928 495000 115048
rect 0 113568 800 113688
rect 494200 109624 495000 109744
rect 0 108128 800 108248
rect 494200 104320 495000 104440
rect 0 102688 800 102808
rect 494200 99016 495000 99136
rect 0 97248 800 97368
rect 494200 93712 495000 93832
rect 0 91808 800 91928
rect 494200 88408 495000 88528
rect 0 86368 800 86488
rect 494200 83104 495000 83224
rect 0 80928 800 81048
rect 494200 77800 495000 77920
rect 0 75488 800 75608
rect 494200 72496 495000 72616
rect 0 70048 800 70168
rect 494200 67192 495000 67312
rect 0 64608 800 64728
rect 494200 61888 495000 62008
rect 0 59168 800 59288
rect 494200 56584 495000 56704
rect 0 53728 800 53848
rect 494200 51280 495000 51400
rect 0 48288 800 48408
rect 494200 45976 495000 46096
rect 0 42848 800 42968
rect 494200 40672 495000 40792
rect 0 37408 800 37528
rect 494200 35368 495000 35488
rect 0 31968 800 32088
rect 494200 30064 495000 30184
rect 0 26528 800 26648
rect 494200 24760 495000 24880
rect 0 21088 800 21208
rect 494200 19456 495000 19576
rect 0 15648 800 15768
rect 494200 14152 495000 14272
rect 0 10208 800 10328
rect 494200 8848 495000 8968
rect 0 4768 800 4888
<< obsm3 >>
rect 798 538088 494200 540769
rect 880 537808 494200 538088
rect 798 534144 494200 537808
rect 798 533864 494120 534144
rect 798 532648 494200 533864
rect 880 532368 494200 532648
rect 798 528840 494200 532368
rect 798 528560 494120 528840
rect 798 527208 494200 528560
rect 880 526928 494200 527208
rect 798 523536 494200 526928
rect 798 523256 494120 523536
rect 798 521768 494200 523256
rect 880 521488 494200 521768
rect 798 518232 494200 521488
rect 798 517952 494120 518232
rect 798 516328 494200 517952
rect 880 516048 494200 516328
rect 798 512928 494200 516048
rect 798 512648 494120 512928
rect 798 510888 494200 512648
rect 880 510608 494200 510888
rect 798 507624 494200 510608
rect 798 507344 494120 507624
rect 798 505448 494200 507344
rect 880 505168 494200 505448
rect 798 502320 494200 505168
rect 798 502040 494120 502320
rect 798 500008 494200 502040
rect 880 499728 494200 500008
rect 798 497016 494200 499728
rect 798 496736 494120 497016
rect 798 494568 494200 496736
rect 880 494288 494200 494568
rect 798 491712 494200 494288
rect 798 491432 494120 491712
rect 798 489128 494200 491432
rect 880 488848 494200 489128
rect 798 486408 494200 488848
rect 798 486128 494120 486408
rect 798 483688 494200 486128
rect 880 483408 494200 483688
rect 798 481104 494200 483408
rect 798 480824 494120 481104
rect 798 478248 494200 480824
rect 880 477968 494200 478248
rect 798 475800 494200 477968
rect 798 475520 494120 475800
rect 798 472808 494200 475520
rect 880 472528 494200 472808
rect 798 470496 494200 472528
rect 798 470216 494120 470496
rect 798 467368 494200 470216
rect 880 467088 494200 467368
rect 798 465192 494200 467088
rect 798 464912 494120 465192
rect 798 461928 494200 464912
rect 880 461648 494200 461928
rect 798 459888 494200 461648
rect 798 459608 494120 459888
rect 798 456488 494200 459608
rect 880 456208 494200 456488
rect 798 454584 494200 456208
rect 798 454304 494120 454584
rect 798 451048 494200 454304
rect 880 450768 494200 451048
rect 798 449280 494200 450768
rect 798 449000 494120 449280
rect 798 445608 494200 449000
rect 880 445328 494200 445608
rect 798 443976 494200 445328
rect 798 443696 494120 443976
rect 798 440168 494200 443696
rect 880 439888 494200 440168
rect 798 438672 494200 439888
rect 798 438392 494120 438672
rect 798 434728 494200 438392
rect 880 434448 494200 434728
rect 798 433368 494200 434448
rect 798 433088 494120 433368
rect 798 429288 494200 433088
rect 880 429008 494200 429288
rect 798 428064 494200 429008
rect 798 427784 494120 428064
rect 798 423848 494200 427784
rect 880 423568 494200 423848
rect 798 422760 494200 423568
rect 798 422480 494120 422760
rect 798 418408 494200 422480
rect 880 418128 494200 418408
rect 798 417456 494200 418128
rect 798 417176 494120 417456
rect 798 412968 494200 417176
rect 880 412688 494200 412968
rect 798 412152 494200 412688
rect 798 411872 494120 412152
rect 798 407528 494200 411872
rect 880 407248 494200 407528
rect 798 406848 494200 407248
rect 798 406568 494120 406848
rect 798 402088 494200 406568
rect 880 401808 494200 402088
rect 798 401544 494200 401808
rect 798 401264 494120 401544
rect 798 396648 494200 401264
rect 880 396368 494200 396648
rect 798 396240 494200 396368
rect 798 395960 494120 396240
rect 798 391208 494200 395960
rect 880 390936 494200 391208
rect 880 390928 494120 390936
rect 798 390656 494120 390928
rect 798 385768 494200 390656
rect 880 385632 494200 385768
rect 880 385488 494120 385632
rect 798 385352 494120 385488
rect 798 380328 494200 385352
rect 880 380048 494120 380328
rect 798 375024 494200 380048
rect 798 374888 494120 375024
rect 880 374744 494120 374888
rect 880 374608 494200 374744
rect 798 369720 494200 374608
rect 798 369448 494120 369720
rect 880 369440 494120 369448
rect 880 369168 494200 369440
rect 798 364416 494200 369168
rect 798 364136 494120 364416
rect 798 364008 494200 364136
rect 880 363728 494200 364008
rect 798 359112 494200 363728
rect 798 358832 494120 359112
rect 798 358568 494200 358832
rect 880 358288 494200 358568
rect 798 353808 494200 358288
rect 798 353528 494120 353808
rect 798 353128 494200 353528
rect 880 352848 494200 353128
rect 798 348504 494200 352848
rect 798 348224 494120 348504
rect 798 347688 494200 348224
rect 880 347408 494200 347688
rect 798 343200 494200 347408
rect 798 342920 494120 343200
rect 798 342248 494200 342920
rect 880 341968 494200 342248
rect 798 337896 494200 341968
rect 798 337616 494120 337896
rect 798 336808 494200 337616
rect 880 336528 494200 336808
rect 798 332592 494200 336528
rect 798 332312 494120 332592
rect 798 331368 494200 332312
rect 880 331088 494200 331368
rect 798 327288 494200 331088
rect 798 327008 494120 327288
rect 798 325928 494200 327008
rect 880 325648 494200 325928
rect 798 321984 494200 325648
rect 798 321704 494120 321984
rect 798 320488 494200 321704
rect 880 320208 494200 320488
rect 798 316680 494200 320208
rect 798 316400 494120 316680
rect 798 315048 494200 316400
rect 880 314768 494200 315048
rect 798 311376 494200 314768
rect 798 311096 494120 311376
rect 798 309608 494200 311096
rect 880 309328 494200 309608
rect 798 306072 494200 309328
rect 798 305792 494120 306072
rect 798 304168 494200 305792
rect 880 303888 494200 304168
rect 798 300768 494200 303888
rect 798 300488 494120 300768
rect 798 298728 494200 300488
rect 880 298448 494200 298728
rect 798 295464 494200 298448
rect 798 295184 494120 295464
rect 798 293288 494200 295184
rect 880 293008 494200 293288
rect 798 290160 494200 293008
rect 798 289880 494120 290160
rect 798 287848 494200 289880
rect 880 287568 494200 287848
rect 798 284856 494200 287568
rect 798 284576 494120 284856
rect 798 282408 494200 284576
rect 880 282128 494200 282408
rect 798 279552 494200 282128
rect 798 279272 494120 279552
rect 798 276968 494200 279272
rect 880 276688 494200 276968
rect 798 274248 494200 276688
rect 798 273968 494120 274248
rect 798 271528 494200 273968
rect 880 271248 494200 271528
rect 798 268944 494200 271248
rect 798 268664 494120 268944
rect 798 266088 494200 268664
rect 880 265808 494200 266088
rect 798 263640 494200 265808
rect 798 263360 494120 263640
rect 798 260648 494200 263360
rect 880 260368 494200 260648
rect 798 258336 494200 260368
rect 798 258056 494120 258336
rect 798 255208 494200 258056
rect 880 254928 494200 255208
rect 798 253032 494200 254928
rect 798 252752 494120 253032
rect 798 249768 494200 252752
rect 880 249488 494200 249768
rect 798 247728 494200 249488
rect 798 247448 494120 247728
rect 798 244328 494200 247448
rect 880 244048 494200 244328
rect 798 242424 494200 244048
rect 798 242144 494120 242424
rect 798 238888 494200 242144
rect 880 238608 494200 238888
rect 798 237120 494200 238608
rect 798 236840 494120 237120
rect 798 233448 494200 236840
rect 880 233168 494200 233448
rect 798 231816 494200 233168
rect 798 231536 494120 231816
rect 798 228008 494200 231536
rect 880 227728 494200 228008
rect 798 226512 494200 227728
rect 798 226232 494120 226512
rect 798 222568 494200 226232
rect 880 222288 494200 222568
rect 798 221208 494200 222288
rect 798 220928 494120 221208
rect 798 217128 494200 220928
rect 880 216848 494200 217128
rect 798 215904 494200 216848
rect 798 215624 494120 215904
rect 798 211688 494200 215624
rect 880 211408 494200 211688
rect 798 210600 494200 211408
rect 798 210320 494120 210600
rect 798 206248 494200 210320
rect 880 205968 494200 206248
rect 798 205296 494200 205968
rect 798 205016 494120 205296
rect 798 200808 494200 205016
rect 880 200528 494200 200808
rect 798 199992 494200 200528
rect 798 199712 494120 199992
rect 798 195368 494200 199712
rect 880 195088 494200 195368
rect 798 194688 494200 195088
rect 798 194408 494120 194688
rect 798 189928 494200 194408
rect 880 189648 494200 189928
rect 798 189384 494200 189648
rect 798 189104 494120 189384
rect 798 184488 494200 189104
rect 880 184208 494200 184488
rect 798 184080 494200 184208
rect 798 183800 494120 184080
rect 798 179048 494200 183800
rect 880 178776 494200 179048
rect 880 178768 494120 178776
rect 798 178496 494120 178768
rect 798 173608 494200 178496
rect 880 173472 494200 173608
rect 880 173328 494120 173472
rect 798 173192 494120 173328
rect 798 168168 494200 173192
rect 880 167888 494120 168168
rect 798 162864 494200 167888
rect 798 162728 494120 162864
rect 880 162584 494120 162728
rect 880 162448 494200 162584
rect 798 157560 494200 162448
rect 798 157288 494120 157560
rect 880 157280 494120 157288
rect 880 157008 494200 157280
rect 798 152256 494200 157008
rect 798 151976 494120 152256
rect 798 151848 494200 151976
rect 880 151568 494200 151848
rect 798 146952 494200 151568
rect 798 146672 494120 146952
rect 798 146408 494200 146672
rect 880 146128 494200 146408
rect 798 141648 494200 146128
rect 798 141368 494120 141648
rect 798 140968 494200 141368
rect 880 140688 494200 140968
rect 798 136344 494200 140688
rect 798 136064 494120 136344
rect 798 135528 494200 136064
rect 880 135248 494200 135528
rect 798 131040 494200 135248
rect 798 130760 494120 131040
rect 798 130088 494200 130760
rect 880 129808 494200 130088
rect 798 125736 494200 129808
rect 798 125456 494120 125736
rect 798 124648 494200 125456
rect 880 124368 494200 124648
rect 798 120432 494200 124368
rect 798 120152 494120 120432
rect 798 119208 494200 120152
rect 880 118928 494200 119208
rect 798 115128 494200 118928
rect 798 114848 494120 115128
rect 798 113768 494200 114848
rect 880 113488 494200 113768
rect 798 109824 494200 113488
rect 798 109544 494120 109824
rect 798 108328 494200 109544
rect 880 108048 494200 108328
rect 798 104520 494200 108048
rect 798 104240 494120 104520
rect 798 102888 494200 104240
rect 880 102608 494200 102888
rect 798 99216 494200 102608
rect 798 98936 494120 99216
rect 798 97448 494200 98936
rect 880 97168 494200 97448
rect 798 93912 494200 97168
rect 798 93632 494120 93912
rect 798 92008 494200 93632
rect 880 91728 494200 92008
rect 798 88608 494200 91728
rect 798 88328 494120 88608
rect 798 86568 494200 88328
rect 880 86288 494200 86568
rect 798 83304 494200 86288
rect 798 83024 494120 83304
rect 798 81128 494200 83024
rect 880 80848 494200 81128
rect 798 78000 494200 80848
rect 798 77720 494120 78000
rect 798 75688 494200 77720
rect 880 75408 494200 75688
rect 798 72696 494200 75408
rect 798 72416 494120 72696
rect 798 70248 494200 72416
rect 880 69968 494200 70248
rect 798 67392 494200 69968
rect 798 67112 494120 67392
rect 798 64808 494200 67112
rect 880 64528 494200 64808
rect 798 62088 494200 64528
rect 798 61808 494120 62088
rect 798 59368 494200 61808
rect 880 59088 494200 59368
rect 798 56784 494200 59088
rect 798 56504 494120 56784
rect 798 53928 494200 56504
rect 880 53648 494200 53928
rect 798 51480 494200 53648
rect 798 51200 494120 51480
rect 798 48488 494200 51200
rect 880 48208 494200 48488
rect 798 46176 494200 48208
rect 798 45896 494120 46176
rect 798 43048 494200 45896
rect 880 42768 494200 43048
rect 798 40872 494200 42768
rect 798 40592 494120 40872
rect 798 37608 494200 40592
rect 880 37328 494200 37608
rect 798 35568 494200 37328
rect 798 35288 494120 35568
rect 798 32168 494200 35288
rect 880 31888 494200 32168
rect 798 30264 494200 31888
rect 798 29984 494120 30264
rect 798 26728 494200 29984
rect 880 26448 494200 26728
rect 798 24960 494200 26448
rect 798 24680 494120 24960
rect 798 21288 494200 24680
rect 880 21008 494200 21288
rect 798 19656 494200 21008
rect 798 19376 494120 19656
rect 798 15848 494200 19376
rect 880 15568 494200 15848
rect 798 14352 494200 15568
rect 798 14072 494120 14352
rect 798 10408 494200 14072
rect 880 10128 494200 10408
rect 798 9048 494200 10128
rect 798 8768 494120 9048
rect 798 4968 494200 8768
rect 880 4688 494200 4968
rect 798 2143 494200 4688
<< metal4 >>
rect -2552 -744 -1592 543656
rect -1192 616 -232 542296
rect 1024 -744 1664 543656
rect 1984 -744 2624 543656
rect 12424 34273 13064 543656
rect 13384 536508 14024 543656
rect 23824 536508 24464 543656
rect 24784 508001 25424 543656
rect 13384 473508 14024 480068
rect 23824 473508 24464 479743
rect 24784 473017 25424 479743
rect 13384 410508 14024 417068
rect 23824 410508 24464 417068
rect 24784 410017 25424 417559
rect 13384 347508 14024 354068
rect 23824 347508 24464 354068
rect 24784 347017 25424 354559
rect 13384 284508 14024 291068
rect 23824 284508 24464 291068
rect 24784 284017 25424 291559
rect 13384 221508 14024 228068
rect 23824 221508 24464 228068
rect 24784 221017 25424 228559
rect 13384 158508 14024 165068
rect 23824 158508 24464 165068
rect 24784 158017 25424 165559
rect 13384 95508 14024 102068
rect 23824 95508 24464 102068
rect 24784 95017 25424 102559
rect 13384 34273 14024 39068
rect 23824 34273 24464 39068
rect 24784 34273 25424 39559
rect 12424 -744 13064 9415
rect 13384 -744 14024 6068
rect 23824 -744 24464 6068
rect 24784 -744 25424 9415
rect 35224 -744 35864 543656
rect 36184 -744 36824 543656
rect 46624 536508 47264 543656
rect 47584 533977 48224 543656
rect 58024 533977 58664 543656
rect 58984 533977 59624 543656
rect 69424 533977 70064 543656
rect 70384 533977 71024 543656
rect 46624 473508 47264 480068
rect 47584 473017 48224 483687
rect 58024 473017 58664 483687
rect 58984 473017 59624 483687
rect 69424 473017 70064 483687
rect 70384 473017 71024 483687
rect 80824 473017 81464 543656
rect 81784 536508 82424 543656
rect 81784 473508 82424 480068
rect 46624 410508 47264 417068
rect 47584 410017 48224 418919
rect 58024 410017 58664 418919
rect 58984 410017 59624 418919
rect 69424 410017 70064 418919
rect 70384 410017 71024 418919
rect 80824 410017 81464 418919
rect 81784 410508 82424 417068
rect 46624 347508 47264 354068
rect 47584 347017 48224 355919
rect 58024 347017 58664 355919
rect 58984 347017 59624 355919
rect 69424 347017 70064 355919
rect 70384 347017 71024 355919
rect 80824 347017 81464 355919
rect 81784 347508 82424 354068
rect 46624 284508 47264 291068
rect 47584 284017 48224 292919
rect 58024 284017 58664 292919
rect 58984 284017 59624 292919
rect 69424 284017 70064 292919
rect 70384 284017 71024 292919
rect 80824 284017 81464 292919
rect 81784 284508 82424 291068
rect 46624 221508 47264 228068
rect 47584 221017 48224 229919
rect 58024 221017 58664 229919
rect 58984 221017 59624 229919
rect 69424 221017 70064 229919
rect 70384 221017 71024 229919
rect 80824 221017 81464 229919
rect 81784 221508 82424 228068
rect 46624 158508 47264 165068
rect 47584 158017 48224 166919
rect 58024 158017 58664 166919
rect 58984 158017 59624 166919
rect 69424 158017 70064 166919
rect 70384 158017 71024 166919
rect 80824 158017 81464 166919
rect 81784 158508 82424 165068
rect 46624 95508 47264 102068
rect 47584 95017 48224 103919
rect 58024 95017 58664 103919
rect 58984 95017 59624 103919
rect 69424 95017 70064 103919
rect 70384 95017 71024 103919
rect 80824 95017 81464 103919
rect 81784 95508 82424 102068
rect 46624 32588 47264 39068
rect 46624 -744 47264 6068
rect 47584 -744 48224 40919
rect 58024 32097 58664 40919
rect 58984 32097 59624 40919
rect 69424 32097 70064 40919
rect 70384 32097 71024 40919
rect 58024 -744 58664 12951
rect 58984 -744 59624 12951
rect 69424 -744 70064 12951
rect 70384 -744 71024 12951
rect 80824 -744 81464 40919
rect 81784 32588 82424 39068
rect 81784 -744 82424 6068
rect 92224 -744 92864 543656
rect 93184 -744 93824 543656
rect 103624 536508 104264 543656
rect 104584 533977 105224 543656
rect 115024 533977 115664 543656
rect 115984 533977 116624 543656
rect 126424 533977 127064 543656
rect 127384 533977 128024 543656
rect 103624 473508 104264 480068
rect 104584 473017 105224 483687
rect 115024 473017 115664 483687
rect 115984 473017 116624 483687
rect 126424 473017 127064 483687
rect 127384 473017 128024 483687
rect 137824 473017 138464 543656
rect 138784 536508 139424 543656
rect 138784 473508 139424 480068
rect 103624 410508 104264 417068
rect 104584 410017 105224 418919
rect 115024 410017 115664 418919
rect 115984 410017 116624 418919
rect 126424 410017 127064 418919
rect 127384 410017 128024 418919
rect 137824 410017 138464 418919
rect 138784 410508 139424 417068
rect 103624 347508 104264 354068
rect 104584 347017 105224 355919
rect 115024 347017 115664 355919
rect 115984 347017 116624 355919
rect 126424 347017 127064 355919
rect 127384 347017 128024 355919
rect 137824 347017 138464 355919
rect 138784 347508 139424 354068
rect 103624 284508 104264 291068
rect 104584 284017 105224 292919
rect 115024 284017 115664 292919
rect 115984 284017 116624 292919
rect 126424 284017 127064 292919
rect 127384 284017 128024 292919
rect 137824 284017 138464 292919
rect 138784 284508 139424 291068
rect 103624 221508 104264 228068
rect 104584 221017 105224 229919
rect 115024 221017 115664 229919
rect 115984 221017 116624 229919
rect 126424 221017 127064 229919
rect 127384 221017 128024 229919
rect 137824 221017 138464 229919
rect 138784 221508 139424 228068
rect 103624 158508 104264 165068
rect 104584 158017 105224 166919
rect 115024 158017 115664 166919
rect 115984 158017 116624 166919
rect 126424 158017 127064 166919
rect 127384 158017 128024 166919
rect 137824 158017 138464 166919
rect 138784 158508 139424 165068
rect 103624 95508 104264 102068
rect 104584 95017 105224 103919
rect 115024 95017 115664 103919
rect 115984 95017 116624 103919
rect 126424 95017 127064 103919
rect 127384 95017 128024 103919
rect 137824 95017 138464 103919
rect 138784 95508 139424 102068
rect 103624 32588 104264 39068
rect 103624 -744 104264 6068
rect 104584 -744 105224 40919
rect 115024 32097 115664 40919
rect 115984 32097 116624 40919
rect 126424 32097 127064 40919
rect 127384 32097 128024 40919
rect 115024 -744 115664 12951
rect 115984 -744 116624 12951
rect 126424 -744 127064 12951
rect 127384 -744 128024 12951
rect 137824 -744 138464 40919
rect 138784 32588 139424 39068
rect 138784 -744 139424 6068
rect 149224 -744 149864 543656
rect 150184 -744 150824 543656
rect 160624 536508 161264 543656
rect 161584 533977 162224 543656
rect 172024 533977 172664 543656
rect 172984 533977 173624 543656
rect 183424 533977 184064 543656
rect 184384 533977 185024 543656
rect 160624 473508 161264 480068
rect 161584 473017 162224 483687
rect 172024 473017 172664 483687
rect 172984 473017 173624 483687
rect 183424 473017 184064 483687
rect 184384 473017 185024 483687
rect 194824 473017 195464 543656
rect 195784 536508 196424 543656
rect 195784 473508 196424 480068
rect 160624 410508 161264 417068
rect 161584 410017 162224 418919
rect 172024 410017 172664 418919
rect 172984 410017 173624 418919
rect 183424 410017 184064 418919
rect 184384 410017 185024 418919
rect 194824 410017 195464 418919
rect 195784 410508 196424 417068
rect 160624 347508 161264 354068
rect 161584 347017 162224 355919
rect 172024 347017 172664 355919
rect 172984 347017 173624 355919
rect 183424 347017 184064 355919
rect 184384 347017 185024 355919
rect 194824 347017 195464 355919
rect 195784 347508 196424 354068
rect 160624 284508 161264 291068
rect 161584 284017 162224 292919
rect 172024 284017 172664 292919
rect 172984 284017 173624 292919
rect 183424 284017 184064 292919
rect 184384 284017 185024 292919
rect 194824 284017 195464 292919
rect 195784 284508 196424 291068
rect 160624 221508 161264 228068
rect 161584 221017 162224 229919
rect 172024 221017 172664 229919
rect 172984 221017 173624 229919
rect 183424 221017 184064 229919
rect 184384 221017 185024 229919
rect 194824 221017 195464 229919
rect 195784 221508 196424 228068
rect 160624 158508 161264 165068
rect 161584 158017 162224 166919
rect 172024 158017 172664 166919
rect 172984 158017 173624 166919
rect 183424 158017 184064 166919
rect 184384 158017 185024 166919
rect 194824 158017 195464 166919
rect 195784 158508 196424 165068
rect 160624 95508 161264 102068
rect 161584 95017 162224 103919
rect 172024 95017 172664 103919
rect 172984 95017 173624 103919
rect 183424 95017 184064 103919
rect 184384 95017 185024 103919
rect 194824 95017 195464 103919
rect 195784 95508 196424 102068
rect 160624 32588 161264 39068
rect 160624 -744 161264 6068
rect 161584 -744 162224 40919
rect 172024 32097 172664 40919
rect 172984 32097 173624 40919
rect 183424 32097 184064 40919
rect 184384 32097 185024 40919
rect 172024 -744 172664 12951
rect 172984 -744 173624 12951
rect 183424 -744 184064 12951
rect 184384 -744 185024 12951
rect 194824 -744 195464 40919
rect 195784 32588 196424 39068
rect 195784 -744 196424 6068
rect 206224 -744 206864 543656
rect 207184 -744 207824 543656
rect 217624 536508 218264 543656
rect 218584 533977 219224 543656
rect 229024 533977 229664 543656
rect 229984 533977 230624 543656
rect 240424 533977 241064 543656
rect 241384 533977 242024 543656
rect 217624 473508 218264 480068
rect 218584 473017 219224 483687
rect 229024 473017 229664 483687
rect 229984 473017 230624 483687
rect 240424 473017 241064 483687
rect 241384 473017 242024 483687
rect 251824 473017 252464 543656
rect 252784 536508 253424 543656
rect 252784 473508 253424 480068
rect 217624 410508 218264 417068
rect 218584 410017 219224 418919
rect 229024 410017 229664 418919
rect 229984 410017 230624 418919
rect 240424 410017 241064 418919
rect 241384 410017 242024 418919
rect 251824 410017 252464 418919
rect 252784 410508 253424 417068
rect 217624 347508 218264 354068
rect 218584 347017 219224 355919
rect 229024 347017 229664 355919
rect 229984 347017 230624 355919
rect 240424 347017 241064 355919
rect 241384 347017 242024 355919
rect 251824 347017 252464 355919
rect 252784 347508 253424 354068
rect 217624 284508 218264 291068
rect 218584 284017 219224 292919
rect 229024 284017 229664 292919
rect 229984 284017 230624 292919
rect 240424 284017 241064 292919
rect 241384 284017 242024 292919
rect 251824 284017 252464 292919
rect 252784 284508 253424 291068
rect 217624 221508 218264 228068
rect 218584 221017 219224 229919
rect 229024 221017 229664 229919
rect 229984 221017 230624 229919
rect 240424 221017 241064 229919
rect 241384 221017 242024 229919
rect 251824 221017 252464 229919
rect 252784 221508 253424 228068
rect 217624 158508 218264 165068
rect 218584 158017 219224 166919
rect 229024 158017 229664 166919
rect 229984 158017 230624 166919
rect 240424 158017 241064 166919
rect 241384 158017 242024 166919
rect 251824 158017 252464 166919
rect 252784 158508 253424 165068
rect 217624 95508 218264 102068
rect 218584 95017 219224 103919
rect 229024 95017 229664 103919
rect 229984 95017 230624 103919
rect 240424 95017 241064 103919
rect 241384 95017 242024 103919
rect 251824 95017 252464 103919
rect 252784 95508 253424 102068
rect 217624 32588 218264 39068
rect 217624 -744 218264 6068
rect 218584 -744 219224 40919
rect 229024 32097 229664 40919
rect 229984 32097 230624 40919
rect 240424 32097 241064 40919
rect 241384 32097 242024 40919
rect 229024 -744 229664 12951
rect 229984 -744 230624 12951
rect 240424 -744 241064 12951
rect 241384 -744 242024 12951
rect 251824 -744 252464 40919
rect 252784 32588 253424 39068
rect 252784 -744 253424 6068
rect 263224 -744 263864 543656
rect 264184 -744 264824 543656
rect 274624 536508 275264 543656
rect 275584 533977 276224 543656
rect 286024 533977 286664 543656
rect 286984 533977 287624 543656
rect 297424 533977 298064 543656
rect 298384 533977 299024 543656
rect 274624 473508 275264 480068
rect 275584 473017 276224 483687
rect 286024 473017 286664 483687
rect 286984 473017 287624 483687
rect 297424 473017 298064 483687
rect 298384 473017 299024 483687
rect 308824 473017 309464 543656
rect 309784 536508 310424 543656
rect 309784 473508 310424 480068
rect 274624 410508 275264 417068
rect 275584 410017 276224 418919
rect 286024 410017 286664 418919
rect 286984 410017 287624 418919
rect 297424 410017 298064 418919
rect 298384 410017 299024 418919
rect 308824 410017 309464 418919
rect 309784 410508 310424 417068
rect 274624 347508 275264 354068
rect 275584 347017 276224 355919
rect 286024 347017 286664 355919
rect 286984 347017 287624 355919
rect 297424 347017 298064 355919
rect 298384 347017 299024 355919
rect 308824 347017 309464 355919
rect 309784 347508 310424 354068
rect 274624 284508 275264 291068
rect 275584 284017 276224 292919
rect 286024 284017 286664 292919
rect 286984 284017 287624 292919
rect 297424 284017 298064 292919
rect 298384 284017 299024 292919
rect 308824 284017 309464 292919
rect 309784 284508 310424 291068
rect 274624 221508 275264 228068
rect 275584 221017 276224 229919
rect 286024 221017 286664 229919
rect 286984 221017 287624 229919
rect 297424 221017 298064 229919
rect 298384 221017 299024 229919
rect 308824 221017 309464 229919
rect 309784 221508 310424 228068
rect 274624 158508 275264 165068
rect 275584 158017 276224 166919
rect 286024 158017 286664 166919
rect 286984 158017 287624 166919
rect 297424 158017 298064 166919
rect 298384 158017 299024 166919
rect 308824 158017 309464 166919
rect 309784 158508 310424 165068
rect 274624 95508 275264 102068
rect 275584 95017 276224 103919
rect 286024 95017 286664 103919
rect 286984 95017 287624 103919
rect 297424 95017 298064 103919
rect 298384 95017 299024 103919
rect 308824 95017 309464 103919
rect 309784 95508 310424 102068
rect 274624 32588 275264 39068
rect 274624 -744 275264 6068
rect 275584 -744 276224 40919
rect 286024 32097 286664 40919
rect 286984 32097 287624 40919
rect 297424 32097 298064 40919
rect 298384 32097 299024 40919
rect 286024 -744 286664 12951
rect 286984 -744 287624 12951
rect 297424 -744 298064 12951
rect 298384 -744 299024 12951
rect 308824 -744 309464 40919
rect 309784 32588 310424 39068
rect 309784 -744 310424 6068
rect 320224 -744 320864 543656
rect 321184 -744 321824 543656
rect 331624 536508 332264 543656
rect 332584 533977 333224 543656
rect 343024 533977 343664 543656
rect 343984 533977 344624 543656
rect 354424 533977 355064 543656
rect 355384 533977 356024 543656
rect 331624 473508 332264 480068
rect 332584 473017 333224 483687
rect 343024 473017 343664 483687
rect 343984 473017 344624 483687
rect 354424 473017 355064 483687
rect 355384 473017 356024 483687
rect 365824 473017 366464 543656
rect 366784 536508 367424 543656
rect 366784 473508 367424 480068
rect 331624 410508 332264 417068
rect 332584 410017 333224 418919
rect 343024 410017 343664 418919
rect 343984 410017 344624 418919
rect 354424 410017 355064 418919
rect 355384 410017 356024 418919
rect 365824 410017 366464 418919
rect 366784 410508 367424 417068
rect 331624 347508 332264 354068
rect 332584 347017 333224 355919
rect 343024 347017 343664 355919
rect 343984 347017 344624 355919
rect 354424 347017 355064 355919
rect 355384 347017 356024 355919
rect 365824 347017 366464 355919
rect 366784 347508 367424 354068
rect 331624 284508 332264 291068
rect 332584 284017 333224 292919
rect 343024 284017 343664 292919
rect 343984 284017 344624 292919
rect 354424 284017 355064 292919
rect 355384 284017 356024 292919
rect 365824 284017 366464 292919
rect 366784 284508 367424 291068
rect 331624 221508 332264 228068
rect 332584 221017 333224 229919
rect 343024 221017 343664 229919
rect 343984 221017 344624 229919
rect 354424 221017 355064 229919
rect 355384 221017 356024 229919
rect 365824 221017 366464 229919
rect 366784 221508 367424 228068
rect 331624 158508 332264 165068
rect 332584 158017 333224 166919
rect 343024 158017 343664 166919
rect 343984 158017 344624 166919
rect 354424 158017 355064 166919
rect 355384 158017 356024 166919
rect 365824 158017 366464 166919
rect 366784 158508 367424 165068
rect 331624 95508 332264 102068
rect 332584 95017 333224 103919
rect 343024 95017 343664 103919
rect 343984 95017 344624 103919
rect 354424 95017 355064 103919
rect 355384 95017 356024 103919
rect 365824 95017 366464 103919
rect 366784 95508 367424 102068
rect 331624 32588 332264 39068
rect 331624 -744 332264 6068
rect 332584 -744 333224 40919
rect 343024 32097 343664 40919
rect 343984 32097 344624 40919
rect 354424 32097 355064 40919
rect 355384 32097 356024 40919
rect 343024 -744 343664 12951
rect 343984 -744 344624 12951
rect 354424 -744 355064 12951
rect 355384 -744 356024 12951
rect 365824 -744 366464 40919
rect 366784 32588 367424 39068
rect 366784 -744 367424 6068
rect 377224 -744 377864 543656
rect 378184 -744 378824 543656
rect 388624 536508 389264 543656
rect 389584 533977 390224 543656
rect 400024 533977 400664 543656
rect 400984 533977 401624 543656
rect 411424 533977 412064 543656
rect 412384 533977 413024 543656
rect 388624 473508 389264 480068
rect 389584 473017 390224 483687
rect 400024 473017 400664 483687
rect 400984 473017 401624 483687
rect 411424 473017 412064 483687
rect 412384 473017 413024 483687
rect 422824 473017 423464 543656
rect 423784 536508 424424 543656
rect 423784 473508 424424 480068
rect 388624 410508 389264 417068
rect 389584 410017 390224 418919
rect 400024 410017 400664 418919
rect 400984 410017 401624 418919
rect 411424 410017 412064 418919
rect 412384 410017 413024 418919
rect 422824 410017 423464 418919
rect 423784 410508 424424 417068
rect 388624 347508 389264 354068
rect 389584 347017 390224 355919
rect 400024 347017 400664 355919
rect 400984 347017 401624 355919
rect 411424 347017 412064 355919
rect 412384 347017 413024 355919
rect 422824 347017 423464 355919
rect 423784 347508 424424 354068
rect 388624 284508 389264 291068
rect 389584 284017 390224 292919
rect 400024 284017 400664 292919
rect 400984 284017 401624 292919
rect 411424 284017 412064 292919
rect 412384 284017 413024 292919
rect 422824 284017 423464 292919
rect 423784 284508 424424 291068
rect 388624 221508 389264 228068
rect 389584 221017 390224 229919
rect 400024 221017 400664 229919
rect 400984 221017 401624 229919
rect 411424 221017 412064 229919
rect 412384 221017 413024 229919
rect 422824 221017 423464 229919
rect 423784 221508 424424 228068
rect 388624 158508 389264 165068
rect 389584 158017 390224 166919
rect 400024 158017 400664 166919
rect 400984 158017 401624 166919
rect 411424 158017 412064 166919
rect 412384 158017 413024 166919
rect 422824 158017 423464 166919
rect 423784 158508 424424 165068
rect 388624 95508 389264 102068
rect 389584 95017 390224 103919
rect 400024 95017 400664 103919
rect 400984 95017 401624 103919
rect 411424 95017 412064 103919
rect 412384 95017 413024 103919
rect 422824 95017 423464 103919
rect 423784 95508 424424 102068
rect 388624 32588 389264 39068
rect 388624 -744 389264 6068
rect 389584 -744 390224 40919
rect 400024 32097 400664 40919
rect 400984 32097 401624 40919
rect 411424 32097 412064 40919
rect 412384 32097 413024 40919
rect 400024 -744 400664 12951
rect 400984 -744 401624 12951
rect 411424 -744 412064 12951
rect 412384 -744 413024 12951
rect 422824 -744 423464 40919
rect 423784 32588 424424 39068
rect 423784 -744 424424 6068
rect 434224 -744 434864 543656
rect 435184 -744 435824 543656
rect 445624 536508 446264 543656
rect 446584 536017 447224 543656
rect 457024 536017 457664 543656
rect 457984 536017 458624 543656
rect 468424 536017 469064 543656
rect 469384 536017 470024 543656
rect 479824 536017 480464 543656
rect 480784 536508 481424 543656
rect 445624 473508 446264 480068
rect 446584 473017 447224 480287
rect 457024 473017 457664 480287
rect 457984 473017 458624 480287
rect 468424 473017 469064 480287
rect 469384 473017 470024 480287
rect 479824 473017 480464 480287
rect 480784 473508 481424 480068
rect 445624 410508 446264 417068
rect 446584 410017 447224 417287
rect 457024 410017 457664 417287
rect 457984 410017 458624 417287
rect 468424 410017 469064 417287
rect 469384 410017 470024 417287
rect 479824 410017 480464 417287
rect 480784 410508 481424 417068
rect 445624 347508 446264 354068
rect 446584 347017 447224 354287
rect 457024 347017 457664 354287
rect 457984 347017 458624 354287
rect 468424 347017 469064 354287
rect 469384 347017 470024 354287
rect 479824 347017 480464 354287
rect 480784 347508 481424 354068
rect 445624 284508 446264 291068
rect 446584 284017 447224 291287
rect 457024 284017 457664 291287
rect 457984 284017 458624 291287
rect 468424 284017 469064 291287
rect 469384 284017 470024 291287
rect 479824 284017 480464 291287
rect 480784 284508 481424 291068
rect 445624 221508 446264 228068
rect 446584 221017 447224 228287
rect 457024 221017 457664 228287
rect 457984 221017 458624 228287
rect 468424 221017 469064 228287
rect 469384 221017 470024 228287
rect 479824 221017 480464 228287
rect 480784 221508 481424 228068
rect 445624 158508 446264 165068
rect 446584 158017 447224 165287
rect 457024 158017 457664 165287
rect 457984 158017 458624 165287
rect 468424 158017 469064 165287
rect 469384 158017 470024 165287
rect 479824 158017 480464 165287
rect 480784 158508 481424 165068
rect 445624 95508 446264 102068
rect 446584 95017 447224 102287
rect 457024 95017 457664 102287
rect 457984 95017 458624 102287
rect 468424 95017 469064 102287
rect 469384 95017 470024 102287
rect 479824 95017 480464 102287
rect 480784 95508 481424 102068
rect 445624 32588 446264 39068
rect 446584 31689 447224 39287
rect 457024 31689 457664 39287
rect 457984 31689 458624 39287
rect 445624 -744 446264 6068
rect 446584 -744 447224 13087
rect 457024 -744 457664 13087
rect 457984 -744 458624 13087
rect 468424 -744 469064 39287
rect 469384 -744 470024 39287
rect 479824 -744 480464 39287
rect 480784 32588 481424 39068
rect 480784 -744 481424 6068
rect 491224 -744 491864 543656
rect 492184 -744 492824 543656
rect 495192 616 496152 542296
rect 496552 -744 497512 543656
<< obsm4 >>
rect 8944 34193 12344 534448
rect 13144 507921 24704 534448
rect 25504 507921 35144 534448
rect 13144 480148 35144 507921
rect 13144 473428 13304 480148
rect 14104 479823 35144 480148
rect 14104 473428 23744 479823
rect 24544 473428 24704 479823
rect 13144 472937 24704 473428
rect 25504 472937 35144 479823
rect 13144 417639 35144 472937
rect 13144 417148 24704 417639
rect 13144 410428 13304 417148
rect 14104 410428 23744 417148
rect 24544 410428 24704 417148
rect 13144 409937 24704 410428
rect 25504 409937 35144 417639
rect 13144 354639 35144 409937
rect 13144 354148 24704 354639
rect 13144 347428 13304 354148
rect 14104 347428 23744 354148
rect 24544 347428 24704 354148
rect 13144 346937 24704 347428
rect 25504 346937 35144 354639
rect 13144 291639 35144 346937
rect 13144 291148 24704 291639
rect 13144 284428 13304 291148
rect 14104 284428 23744 291148
rect 24544 284428 24704 291148
rect 13144 283937 24704 284428
rect 25504 283937 35144 291639
rect 13144 228639 35144 283937
rect 13144 228148 24704 228639
rect 13144 221428 13304 228148
rect 14104 221428 23744 228148
rect 24544 221428 24704 228148
rect 13144 220937 24704 221428
rect 25504 220937 35144 228639
rect 13144 165639 35144 220937
rect 13144 165148 24704 165639
rect 13144 158428 13304 165148
rect 14104 158428 23744 165148
rect 24544 158428 24704 165148
rect 13144 157937 24704 158428
rect 25504 157937 35144 165639
rect 13144 102639 35144 157937
rect 13144 102148 24704 102639
rect 13144 95428 13304 102148
rect 14104 95428 23744 102148
rect 24544 95428 24704 102148
rect 13144 94937 24704 95428
rect 25504 94937 35144 102639
rect 13144 39639 35144 94937
rect 13144 39148 24704 39639
rect 13144 34193 13304 39148
rect 14104 34193 23744 39148
rect 24544 34193 24704 39148
rect 25504 34193 35144 39639
rect 8944 9495 35144 34193
rect 8944 8128 12344 9495
rect 13144 8128 24704 9495
rect 25504 8128 35144 9495
rect 35944 8128 36104 534448
rect 36904 533897 47504 534448
rect 48304 533897 57944 534448
rect 58744 533897 58904 534448
rect 59704 533897 69344 534448
rect 70144 533897 70304 534448
rect 71104 533897 80744 534448
rect 36904 483767 80744 533897
rect 36904 480148 47504 483767
rect 36904 473428 46544 480148
rect 47344 473428 47504 480148
rect 36904 472937 47504 473428
rect 48304 472937 57944 483767
rect 58744 472937 58904 483767
rect 59704 472937 69344 483767
rect 70144 472937 70304 483767
rect 71104 472937 80744 483767
rect 81544 480148 92144 534448
rect 81544 473428 81704 480148
rect 82504 473428 92144 480148
rect 81544 472937 92144 473428
rect 36904 418999 92144 472937
rect 36904 417148 47504 418999
rect 36904 410428 46544 417148
rect 47344 410428 47504 417148
rect 36904 409937 47504 410428
rect 48304 409937 57944 418999
rect 58744 409937 58904 418999
rect 59704 409937 69344 418999
rect 70144 409937 70304 418999
rect 71104 409937 80744 418999
rect 81544 417148 92144 418999
rect 81544 410428 81704 417148
rect 82504 410428 92144 417148
rect 81544 409937 92144 410428
rect 36904 355999 92144 409937
rect 36904 354148 47504 355999
rect 36904 347428 46544 354148
rect 47344 347428 47504 354148
rect 36904 346937 47504 347428
rect 48304 346937 57944 355999
rect 58744 346937 58904 355999
rect 59704 346937 69344 355999
rect 70144 346937 70304 355999
rect 71104 346937 80744 355999
rect 81544 354148 92144 355999
rect 81544 347428 81704 354148
rect 82504 347428 92144 354148
rect 81544 346937 92144 347428
rect 36904 292999 92144 346937
rect 36904 291148 47504 292999
rect 36904 284428 46544 291148
rect 47344 284428 47504 291148
rect 36904 283937 47504 284428
rect 48304 283937 57944 292999
rect 58744 283937 58904 292999
rect 59704 283937 69344 292999
rect 70144 283937 70304 292999
rect 71104 283937 80744 292999
rect 81544 291148 92144 292999
rect 81544 284428 81704 291148
rect 82504 284428 92144 291148
rect 81544 283937 92144 284428
rect 36904 229999 92144 283937
rect 36904 228148 47504 229999
rect 36904 221428 46544 228148
rect 47344 221428 47504 228148
rect 36904 220937 47504 221428
rect 48304 220937 57944 229999
rect 58744 220937 58904 229999
rect 59704 220937 69344 229999
rect 70144 220937 70304 229999
rect 71104 220937 80744 229999
rect 81544 228148 92144 229999
rect 81544 221428 81704 228148
rect 82504 221428 92144 228148
rect 81544 220937 92144 221428
rect 36904 166999 92144 220937
rect 36904 165148 47504 166999
rect 36904 158428 46544 165148
rect 47344 158428 47504 165148
rect 36904 157937 47504 158428
rect 48304 157937 57944 166999
rect 58744 157937 58904 166999
rect 59704 157937 69344 166999
rect 70144 157937 70304 166999
rect 71104 157937 80744 166999
rect 81544 165148 92144 166999
rect 81544 158428 81704 165148
rect 82504 158428 92144 165148
rect 81544 157937 92144 158428
rect 36904 103999 92144 157937
rect 36904 102148 47504 103999
rect 36904 95428 46544 102148
rect 47344 95428 47504 102148
rect 36904 94937 47504 95428
rect 48304 94937 57944 103999
rect 58744 94937 58904 103999
rect 59704 94937 69344 103999
rect 70144 94937 70304 103999
rect 71104 94937 80744 103999
rect 81544 102148 92144 103999
rect 81544 95428 81704 102148
rect 82504 95428 92144 102148
rect 81544 94937 92144 95428
rect 36904 40999 92144 94937
rect 36904 39148 47504 40999
rect 36904 32508 46544 39148
rect 47344 32508 47504 39148
rect 36904 8128 47504 32508
rect 48304 32017 57944 40999
rect 58744 32017 58904 40999
rect 59704 32017 69344 40999
rect 70144 32017 70304 40999
rect 71104 32017 80744 40999
rect 48304 13031 80744 32017
rect 48304 8128 57944 13031
rect 58744 8128 58904 13031
rect 59704 8128 69344 13031
rect 70144 8128 70304 13031
rect 71104 8128 80744 13031
rect 81544 39148 92144 40999
rect 81544 32508 81704 39148
rect 82504 32508 92144 39148
rect 81544 8128 92144 32508
rect 92944 8128 93104 534448
rect 93904 533897 104504 534448
rect 105304 533897 114944 534448
rect 115744 533897 115904 534448
rect 116704 533897 126344 534448
rect 127144 533897 127304 534448
rect 128104 533897 137744 534448
rect 93904 483767 137744 533897
rect 93904 480148 104504 483767
rect 93904 473428 103544 480148
rect 104344 473428 104504 480148
rect 93904 472937 104504 473428
rect 105304 472937 114944 483767
rect 115744 472937 115904 483767
rect 116704 472937 126344 483767
rect 127144 472937 127304 483767
rect 128104 472937 137744 483767
rect 138544 480148 149144 534448
rect 138544 473428 138704 480148
rect 139504 473428 149144 480148
rect 138544 472937 149144 473428
rect 93904 418999 149144 472937
rect 93904 417148 104504 418999
rect 93904 410428 103544 417148
rect 104344 410428 104504 417148
rect 93904 409937 104504 410428
rect 105304 409937 114944 418999
rect 115744 409937 115904 418999
rect 116704 409937 126344 418999
rect 127144 409937 127304 418999
rect 128104 409937 137744 418999
rect 138544 417148 149144 418999
rect 138544 410428 138704 417148
rect 139504 410428 149144 417148
rect 138544 409937 149144 410428
rect 93904 355999 149144 409937
rect 93904 354148 104504 355999
rect 93904 347428 103544 354148
rect 104344 347428 104504 354148
rect 93904 346937 104504 347428
rect 105304 346937 114944 355999
rect 115744 346937 115904 355999
rect 116704 346937 126344 355999
rect 127144 346937 127304 355999
rect 128104 346937 137744 355999
rect 138544 354148 149144 355999
rect 138544 347428 138704 354148
rect 139504 347428 149144 354148
rect 138544 346937 149144 347428
rect 93904 292999 149144 346937
rect 93904 291148 104504 292999
rect 93904 284428 103544 291148
rect 104344 284428 104504 291148
rect 93904 283937 104504 284428
rect 105304 283937 114944 292999
rect 115744 283937 115904 292999
rect 116704 283937 126344 292999
rect 127144 283937 127304 292999
rect 128104 283937 137744 292999
rect 138544 291148 149144 292999
rect 138544 284428 138704 291148
rect 139504 284428 149144 291148
rect 138544 283937 149144 284428
rect 93904 229999 149144 283937
rect 93904 228148 104504 229999
rect 93904 221428 103544 228148
rect 104344 221428 104504 228148
rect 93904 220937 104504 221428
rect 105304 220937 114944 229999
rect 115744 220937 115904 229999
rect 116704 220937 126344 229999
rect 127144 220937 127304 229999
rect 128104 220937 137744 229999
rect 138544 228148 149144 229999
rect 138544 221428 138704 228148
rect 139504 221428 149144 228148
rect 138544 220937 149144 221428
rect 93904 166999 149144 220937
rect 93904 165148 104504 166999
rect 93904 158428 103544 165148
rect 104344 158428 104504 165148
rect 93904 157937 104504 158428
rect 105304 157937 114944 166999
rect 115744 157937 115904 166999
rect 116704 157937 126344 166999
rect 127144 157937 127304 166999
rect 128104 157937 137744 166999
rect 138544 165148 149144 166999
rect 138544 158428 138704 165148
rect 139504 158428 149144 165148
rect 138544 157937 149144 158428
rect 93904 103999 149144 157937
rect 93904 102148 104504 103999
rect 93904 95428 103544 102148
rect 104344 95428 104504 102148
rect 93904 94937 104504 95428
rect 105304 94937 114944 103999
rect 115744 94937 115904 103999
rect 116704 94937 126344 103999
rect 127144 94937 127304 103999
rect 128104 94937 137744 103999
rect 138544 102148 149144 103999
rect 138544 95428 138704 102148
rect 139504 95428 149144 102148
rect 138544 94937 149144 95428
rect 93904 40999 149144 94937
rect 93904 39148 104504 40999
rect 93904 32508 103544 39148
rect 104344 32508 104504 39148
rect 93904 8128 104504 32508
rect 105304 32017 114944 40999
rect 115744 32017 115904 40999
rect 116704 32017 126344 40999
rect 127144 32017 127304 40999
rect 128104 32017 137744 40999
rect 105304 13031 137744 32017
rect 105304 8128 114944 13031
rect 115744 8128 115904 13031
rect 116704 8128 126344 13031
rect 127144 8128 127304 13031
rect 128104 8128 137744 13031
rect 138544 39148 149144 40999
rect 138544 32508 138704 39148
rect 139504 32508 149144 39148
rect 138544 8128 149144 32508
rect 149944 8128 150104 534448
rect 150904 533897 161504 534448
rect 162304 533897 171944 534448
rect 172744 533897 172904 534448
rect 173704 533897 183344 534448
rect 184144 533897 184304 534448
rect 185104 533897 194744 534448
rect 150904 483767 194744 533897
rect 150904 480148 161504 483767
rect 150904 473428 160544 480148
rect 161344 473428 161504 480148
rect 150904 472937 161504 473428
rect 162304 472937 171944 483767
rect 172744 472937 172904 483767
rect 173704 472937 183344 483767
rect 184144 472937 184304 483767
rect 185104 472937 194744 483767
rect 195544 480148 206144 534448
rect 195544 473428 195704 480148
rect 196504 473428 206144 480148
rect 195544 472937 206144 473428
rect 150904 418999 206144 472937
rect 150904 417148 161504 418999
rect 150904 410428 160544 417148
rect 161344 410428 161504 417148
rect 150904 409937 161504 410428
rect 162304 409937 171944 418999
rect 172744 409937 172904 418999
rect 173704 409937 183344 418999
rect 184144 409937 184304 418999
rect 185104 409937 194744 418999
rect 195544 417148 206144 418999
rect 195544 410428 195704 417148
rect 196504 410428 206144 417148
rect 195544 409937 206144 410428
rect 150904 355999 206144 409937
rect 150904 354148 161504 355999
rect 150904 347428 160544 354148
rect 161344 347428 161504 354148
rect 150904 346937 161504 347428
rect 162304 346937 171944 355999
rect 172744 346937 172904 355999
rect 173704 346937 183344 355999
rect 184144 346937 184304 355999
rect 185104 346937 194744 355999
rect 195544 354148 206144 355999
rect 195544 347428 195704 354148
rect 196504 347428 206144 354148
rect 195544 346937 206144 347428
rect 150904 292999 206144 346937
rect 150904 291148 161504 292999
rect 150904 284428 160544 291148
rect 161344 284428 161504 291148
rect 150904 283937 161504 284428
rect 162304 283937 171944 292999
rect 172744 283937 172904 292999
rect 173704 283937 183344 292999
rect 184144 283937 184304 292999
rect 185104 283937 194744 292999
rect 195544 291148 206144 292999
rect 195544 284428 195704 291148
rect 196504 284428 206144 291148
rect 195544 283937 206144 284428
rect 150904 229999 206144 283937
rect 150904 228148 161504 229999
rect 150904 221428 160544 228148
rect 161344 221428 161504 228148
rect 150904 220937 161504 221428
rect 162304 220937 171944 229999
rect 172744 220937 172904 229999
rect 173704 220937 183344 229999
rect 184144 220937 184304 229999
rect 185104 220937 194744 229999
rect 195544 228148 206144 229999
rect 195544 221428 195704 228148
rect 196504 221428 206144 228148
rect 195544 220937 206144 221428
rect 150904 166999 206144 220937
rect 150904 165148 161504 166999
rect 150904 158428 160544 165148
rect 161344 158428 161504 165148
rect 150904 157937 161504 158428
rect 162304 157937 171944 166999
rect 172744 157937 172904 166999
rect 173704 157937 183344 166999
rect 184144 157937 184304 166999
rect 185104 157937 194744 166999
rect 195544 165148 206144 166999
rect 195544 158428 195704 165148
rect 196504 158428 206144 165148
rect 195544 157937 206144 158428
rect 150904 103999 206144 157937
rect 150904 102148 161504 103999
rect 150904 95428 160544 102148
rect 161344 95428 161504 102148
rect 150904 94937 161504 95428
rect 162304 94937 171944 103999
rect 172744 94937 172904 103999
rect 173704 94937 183344 103999
rect 184144 94937 184304 103999
rect 185104 94937 194744 103999
rect 195544 102148 206144 103999
rect 195544 95428 195704 102148
rect 196504 95428 206144 102148
rect 195544 94937 206144 95428
rect 150904 40999 206144 94937
rect 150904 39148 161504 40999
rect 150904 32508 160544 39148
rect 161344 32508 161504 39148
rect 150904 8128 161504 32508
rect 162304 32017 171944 40999
rect 172744 32017 172904 40999
rect 173704 32017 183344 40999
rect 184144 32017 184304 40999
rect 185104 32017 194744 40999
rect 162304 13031 194744 32017
rect 162304 8128 171944 13031
rect 172744 8128 172904 13031
rect 173704 8128 183344 13031
rect 184144 8128 184304 13031
rect 185104 8128 194744 13031
rect 195544 39148 206144 40999
rect 195544 32508 195704 39148
rect 196504 32508 206144 39148
rect 195544 8128 206144 32508
rect 206944 8128 207104 534448
rect 207904 533897 218504 534448
rect 219304 533897 228944 534448
rect 229744 533897 229904 534448
rect 230704 533897 240344 534448
rect 241144 533897 241304 534448
rect 242104 533897 251744 534448
rect 207904 483767 251744 533897
rect 207904 480148 218504 483767
rect 207904 473428 217544 480148
rect 218344 473428 218504 480148
rect 207904 472937 218504 473428
rect 219304 472937 228944 483767
rect 229744 472937 229904 483767
rect 230704 472937 240344 483767
rect 241144 472937 241304 483767
rect 242104 472937 251744 483767
rect 252544 480148 263144 534448
rect 252544 473428 252704 480148
rect 253504 473428 263144 480148
rect 252544 472937 263144 473428
rect 207904 418999 263144 472937
rect 207904 417148 218504 418999
rect 207904 410428 217544 417148
rect 218344 410428 218504 417148
rect 207904 409937 218504 410428
rect 219304 409937 228944 418999
rect 229744 409937 229904 418999
rect 230704 409937 240344 418999
rect 241144 409937 241304 418999
rect 242104 409937 251744 418999
rect 252544 417148 263144 418999
rect 252544 410428 252704 417148
rect 253504 410428 263144 417148
rect 252544 409937 263144 410428
rect 207904 355999 263144 409937
rect 207904 354148 218504 355999
rect 207904 347428 217544 354148
rect 218344 347428 218504 354148
rect 207904 346937 218504 347428
rect 219304 346937 228944 355999
rect 229744 346937 229904 355999
rect 230704 346937 240344 355999
rect 241144 346937 241304 355999
rect 242104 346937 251744 355999
rect 252544 354148 263144 355999
rect 252544 347428 252704 354148
rect 253504 347428 263144 354148
rect 252544 346937 263144 347428
rect 207904 292999 263144 346937
rect 207904 291148 218504 292999
rect 207904 284428 217544 291148
rect 218344 284428 218504 291148
rect 207904 283937 218504 284428
rect 219304 283937 228944 292999
rect 229744 283937 229904 292999
rect 230704 283937 240344 292999
rect 241144 283937 241304 292999
rect 242104 283937 251744 292999
rect 252544 291148 263144 292999
rect 252544 284428 252704 291148
rect 253504 284428 263144 291148
rect 252544 283937 263144 284428
rect 207904 229999 263144 283937
rect 207904 228148 218504 229999
rect 207904 221428 217544 228148
rect 218344 221428 218504 228148
rect 207904 220937 218504 221428
rect 219304 220937 228944 229999
rect 229744 220937 229904 229999
rect 230704 220937 240344 229999
rect 241144 220937 241304 229999
rect 242104 220937 251744 229999
rect 252544 228148 263144 229999
rect 252544 221428 252704 228148
rect 253504 221428 263144 228148
rect 252544 220937 263144 221428
rect 207904 166999 263144 220937
rect 207904 165148 218504 166999
rect 207904 158428 217544 165148
rect 218344 158428 218504 165148
rect 207904 157937 218504 158428
rect 219304 157937 228944 166999
rect 229744 157937 229904 166999
rect 230704 157937 240344 166999
rect 241144 157937 241304 166999
rect 242104 157937 251744 166999
rect 252544 165148 263144 166999
rect 252544 158428 252704 165148
rect 253504 158428 263144 165148
rect 252544 157937 263144 158428
rect 207904 103999 263144 157937
rect 207904 102148 218504 103999
rect 207904 95428 217544 102148
rect 218344 95428 218504 102148
rect 207904 94937 218504 95428
rect 219304 94937 228944 103999
rect 229744 94937 229904 103999
rect 230704 94937 240344 103999
rect 241144 94937 241304 103999
rect 242104 94937 251744 103999
rect 252544 102148 263144 103999
rect 252544 95428 252704 102148
rect 253504 95428 263144 102148
rect 252544 94937 263144 95428
rect 207904 40999 263144 94937
rect 207904 39148 218504 40999
rect 207904 32508 217544 39148
rect 218344 32508 218504 39148
rect 207904 8128 218504 32508
rect 219304 32017 228944 40999
rect 229744 32017 229904 40999
rect 230704 32017 240344 40999
rect 241144 32017 241304 40999
rect 242104 32017 251744 40999
rect 219304 13031 251744 32017
rect 219304 8128 228944 13031
rect 229744 8128 229904 13031
rect 230704 8128 240344 13031
rect 241144 8128 241304 13031
rect 242104 8128 251744 13031
rect 252544 39148 263144 40999
rect 252544 32508 252704 39148
rect 253504 32508 263144 39148
rect 252544 8128 263144 32508
rect 263944 8128 264104 534448
rect 264904 533897 275504 534448
rect 276304 533897 285944 534448
rect 286744 533897 286904 534448
rect 287704 533897 297344 534448
rect 298144 533897 298304 534448
rect 299104 533897 308744 534448
rect 264904 483767 308744 533897
rect 264904 480148 275504 483767
rect 264904 473428 274544 480148
rect 275344 473428 275504 480148
rect 264904 472937 275504 473428
rect 276304 472937 285944 483767
rect 286744 472937 286904 483767
rect 287704 472937 297344 483767
rect 298144 472937 298304 483767
rect 299104 472937 308744 483767
rect 309544 480148 320144 534448
rect 309544 473428 309704 480148
rect 310504 473428 320144 480148
rect 309544 472937 320144 473428
rect 264904 418999 320144 472937
rect 264904 417148 275504 418999
rect 264904 410428 274544 417148
rect 275344 410428 275504 417148
rect 264904 409937 275504 410428
rect 276304 409937 285944 418999
rect 286744 409937 286904 418999
rect 287704 409937 297344 418999
rect 298144 409937 298304 418999
rect 299104 409937 308744 418999
rect 309544 417148 320144 418999
rect 309544 410428 309704 417148
rect 310504 410428 320144 417148
rect 309544 409937 320144 410428
rect 264904 355999 320144 409937
rect 264904 354148 275504 355999
rect 264904 347428 274544 354148
rect 275344 347428 275504 354148
rect 264904 346937 275504 347428
rect 276304 346937 285944 355999
rect 286744 346937 286904 355999
rect 287704 346937 297344 355999
rect 298144 346937 298304 355999
rect 299104 346937 308744 355999
rect 309544 354148 320144 355999
rect 309544 347428 309704 354148
rect 310504 347428 320144 354148
rect 309544 346937 320144 347428
rect 264904 292999 320144 346937
rect 264904 291148 275504 292999
rect 264904 284428 274544 291148
rect 275344 284428 275504 291148
rect 264904 283937 275504 284428
rect 276304 283937 285944 292999
rect 286744 283937 286904 292999
rect 287704 283937 297344 292999
rect 298144 283937 298304 292999
rect 299104 283937 308744 292999
rect 309544 291148 320144 292999
rect 309544 284428 309704 291148
rect 310504 284428 320144 291148
rect 309544 283937 320144 284428
rect 264904 229999 320144 283937
rect 264904 228148 275504 229999
rect 264904 221428 274544 228148
rect 275344 221428 275504 228148
rect 264904 220937 275504 221428
rect 276304 220937 285944 229999
rect 286744 220937 286904 229999
rect 287704 220937 297344 229999
rect 298144 220937 298304 229999
rect 299104 220937 308744 229999
rect 309544 228148 320144 229999
rect 309544 221428 309704 228148
rect 310504 221428 320144 228148
rect 309544 220937 320144 221428
rect 264904 166999 320144 220937
rect 264904 165148 275504 166999
rect 264904 158428 274544 165148
rect 275344 158428 275504 165148
rect 264904 157937 275504 158428
rect 276304 157937 285944 166999
rect 286744 157937 286904 166999
rect 287704 157937 297344 166999
rect 298144 157937 298304 166999
rect 299104 157937 308744 166999
rect 309544 165148 320144 166999
rect 309544 158428 309704 165148
rect 310504 158428 320144 165148
rect 309544 157937 320144 158428
rect 264904 103999 320144 157937
rect 264904 102148 275504 103999
rect 264904 95428 274544 102148
rect 275344 95428 275504 102148
rect 264904 94937 275504 95428
rect 276304 94937 285944 103999
rect 286744 94937 286904 103999
rect 287704 94937 297344 103999
rect 298144 94937 298304 103999
rect 299104 94937 308744 103999
rect 309544 102148 320144 103999
rect 309544 95428 309704 102148
rect 310504 95428 320144 102148
rect 309544 94937 320144 95428
rect 264904 40999 320144 94937
rect 264904 39148 275504 40999
rect 264904 32508 274544 39148
rect 275344 32508 275504 39148
rect 264904 8128 275504 32508
rect 276304 32017 285944 40999
rect 286744 32017 286904 40999
rect 287704 32017 297344 40999
rect 298144 32017 298304 40999
rect 299104 32017 308744 40999
rect 276304 13031 308744 32017
rect 276304 8128 285944 13031
rect 286744 8128 286904 13031
rect 287704 8128 297344 13031
rect 298144 8128 298304 13031
rect 299104 8128 308744 13031
rect 309544 39148 320144 40999
rect 309544 32508 309704 39148
rect 310504 32508 320144 39148
rect 309544 8128 320144 32508
rect 320944 8128 321104 534448
rect 321904 533897 332504 534448
rect 333304 533897 342944 534448
rect 343744 533897 343904 534448
rect 344704 533897 354344 534448
rect 355144 533897 355304 534448
rect 356104 533897 365744 534448
rect 321904 483767 365744 533897
rect 321904 480148 332504 483767
rect 321904 473428 331544 480148
rect 332344 473428 332504 480148
rect 321904 472937 332504 473428
rect 333304 472937 342944 483767
rect 343744 472937 343904 483767
rect 344704 472937 354344 483767
rect 355144 472937 355304 483767
rect 356104 472937 365744 483767
rect 366544 480148 377144 534448
rect 366544 473428 366704 480148
rect 367504 473428 377144 480148
rect 366544 472937 377144 473428
rect 321904 418999 377144 472937
rect 321904 417148 332504 418999
rect 321904 410428 331544 417148
rect 332344 410428 332504 417148
rect 321904 409937 332504 410428
rect 333304 409937 342944 418999
rect 343744 409937 343904 418999
rect 344704 409937 354344 418999
rect 355144 409937 355304 418999
rect 356104 409937 365744 418999
rect 366544 417148 377144 418999
rect 366544 410428 366704 417148
rect 367504 410428 377144 417148
rect 366544 409937 377144 410428
rect 321904 355999 377144 409937
rect 321904 354148 332504 355999
rect 321904 347428 331544 354148
rect 332344 347428 332504 354148
rect 321904 346937 332504 347428
rect 333304 346937 342944 355999
rect 343744 346937 343904 355999
rect 344704 346937 354344 355999
rect 355144 346937 355304 355999
rect 356104 346937 365744 355999
rect 366544 354148 377144 355999
rect 366544 347428 366704 354148
rect 367504 347428 377144 354148
rect 366544 346937 377144 347428
rect 321904 292999 377144 346937
rect 321904 291148 332504 292999
rect 321904 284428 331544 291148
rect 332344 284428 332504 291148
rect 321904 283937 332504 284428
rect 333304 283937 342944 292999
rect 343744 283937 343904 292999
rect 344704 283937 354344 292999
rect 355144 283937 355304 292999
rect 356104 283937 365744 292999
rect 366544 291148 377144 292999
rect 366544 284428 366704 291148
rect 367504 284428 377144 291148
rect 366544 283937 377144 284428
rect 321904 229999 377144 283937
rect 321904 228148 332504 229999
rect 321904 221428 331544 228148
rect 332344 221428 332504 228148
rect 321904 220937 332504 221428
rect 333304 220937 342944 229999
rect 343744 220937 343904 229999
rect 344704 220937 354344 229999
rect 355144 220937 355304 229999
rect 356104 220937 365744 229999
rect 366544 228148 377144 229999
rect 366544 221428 366704 228148
rect 367504 221428 377144 228148
rect 366544 220937 377144 221428
rect 321904 166999 377144 220937
rect 321904 165148 332504 166999
rect 321904 158428 331544 165148
rect 332344 158428 332504 165148
rect 321904 157937 332504 158428
rect 333304 157937 342944 166999
rect 343744 157937 343904 166999
rect 344704 157937 354344 166999
rect 355144 157937 355304 166999
rect 356104 157937 365744 166999
rect 366544 165148 377144 166999
rect 366544 158428 366704 165148
rect 367504 158428 377144 165148
rect 366544 157937 377144 158428
rect 321904 103999 377144 157937
rect 321904 102148 332504 103999
rect 321904 95428 331544 102148
rect 332344 95428 332504 102148
rect 321904 94937 332504 95428
rect 333304 94937 342944 103999
rect 343744 94937 343904 103999
rect 344704 94937 354344 103999
rect 355144 94937 355304 103999
rect 356104 94937 365744 103999
rect 366544 102148 377144 103999
rect 366544 95428 366704 102148
rect 367504 95428 377144 102148
rect 366544 94937 377144 95428
rect 321904 40999 377144 94937
rect 321904 39148 332504 40999
rect 321904 32508 331544 39148
rect 332344 32508 332504 39148
rect 321904 8128 332504 32508
rect 333304 32017 342944 40999
rect 343744 32017 343904 40999
rect 344704 32017 354344 40999
rect 355144 32017 355304 40999
rect 356104 32017 365744 40999
rect 333304 13031 365744 32017
rect 333304 8128 342944 13031
rect 343744 8128 343904 13031
rect 344704 8128 354344 13031
rect 355144 8128 355304 13031
rect 356104 8128 365744 13031
rect 366544 39148 377144 40999
rect 366544 32508 366704 39148
rect 367504 32508 377144 39148
rect 366544 8128 377144 32508
rect 377944 8128 378104 534448
rect 378904 533897 389504 534448
rect 390304 533897 399944 534448
rect 400744 533897 400904 534448
rect 401704 533897 411344 534448
rect 412144 533897 412304 534448
rect 413104 533897 422744 534448
rect 378904 483767 422744 533897
rect 378904 480148 389504 483767
rect 378904 473428 388544 480148
rect 389344 473428 389504 480148
rect 378904 472937 389504 473428
rect 390304 472937 399944 483767
rect 400744 472937 400904 483767
rect 401704 472937 411344 483767
rect 412144 472937 412304 483767
rect 413104 472937 422744 483767
rect 423544 480148 434144 534448
rect 423544 473428 423704 480148
rect 424504 473428 434144 480148
rect 423544 472937 434144 473428
rect 378904 418999 434144 472937
rect 378904 417148 389504 418999
rect 378904 410428 388544 417148
rect 389344 410428 389504 417148
rect 378904 409937 389504 410428
rect 390304 409937 399944 418999
rect 400744 409937 400904 418999
rect 401704 409937 411344 418999
rect 412144 409937 412304 418999
rect 413104 409937 422744 418999
rect 423544 417148 434144 418999
rect 423544 410428 423704 417148
rect 424504 410428 434144 417148
rect 423544 409937 434144 410428
rect 378904 355999 434144 409937
rect 378904 354148 389504 355999
rect 378904 347428 388544 354148
rect 389344 347428 389504 354148
rect 378904 346937 389504 347428
rect 390304 346937 399944 355999
rect 400744 346937 400904 355999
rect 401704 346937 411344 355999
rect 412144 346937 412304 355999
rect 413104 346937 422744 355999
rect 423544 354148 434144 355999
rect 423544 347428 423704 354148
rect 424504 347428 434144 354148
rect 423544 346937 434144 347428
rect 378904 292999 434144 346937
rect 378904 291148 389504 292999
rect 378904 284428 388544 291148
rect 389344 284428 389504 291148
rect 378904 283937 389504 284428
rect 390304 283937 399944 292999
rect 400744 283937 400904 292999
rect 401704 283937 411344 292999
rect 412144 283937 412304 292999
rect 413104 283937 422744 292999
rect 423544 291148 434144 292999
rect 423544 284428 423704 291148
rect 424504 284428 434144 291148
rect 423544 283937 434144 284428
rect 378904 229999 434144 283937
rect 378904 228148 389504 229999
rect 378904 221428 388544 228148
rect 389344 221428 389504 228148
rect 378904 220937 389504 221428
rect 390304 220937 399944 229999
rect 400744 220937 400904 229999
rect 401704 220937 411344 229999
rect 412144 220937 412304 229999
rect 413104 220937 422744 229999
rect 423544 228148 434144 229999
rect 423544 221428 423704 228148
rect 424504 221428 434144 228148
rect 423544 220937 434144 221428
rect 378904 166999 434144 220937
rect 378904 165148 389504 166999
rect 378904 158428 388544 165148
rect 389344 158428 389504 165148
rect 378904 157937 389504 158428
rect 390304 157937 399944 166999
rect 400744 157937 400904 166999
rect 401704 157937 411344 166999
rect 412144 157937 412304 166999
rect 413104 157937 422744 166999
rect 423544 165148 434144 166999
rect 423544 158428 423704 165148
rect 424504 158428 434144 165148
rect 423544 157937 434144 158428
rect 378904 103999 434144 157937
rect 378904 102148 389504 103999
rect 378904 95428 388544 102148
rect 389344 95428 389504 102148
rect 378904 94937 389504 95428
rect 390304 94937 399944 103999
rect 400744 94937 400904 103999
rect 401704 94937 411344 103999
rect 412144 94937 412304 103999
rect 413104 94937 422744 103999
rect 423544 102148 434144 103999
rect 423544 95428 423704 102148
rect 424504 95428 434144 102148
rect 423544 94937 434144 95428
rect 378904 40999 434144 94937
rect 378904 39148 389504 40999
rect 378904 32508 388544 39148
rect 389344 32508 389504 39148
rect 378904 8128 389504 32508
rect 390304 32017 399944 40999
rect 400744 32017 400904 40999
rect 401704 32017 411344 40999
rect 412144 32017 412304 40999
rect 413104 32017 422744 40999
rect 390304 13031 422744 32017
rect 390304 8128 399944 13031
rect 400744 8128 400904 13031
rect 401704 8128 411344 13031
rect 412144 8128 412304 13031
rect 413104 8128 422744 13031
rect 423544 39148 434144 40999
rect 423544 32508 423704 39148
rect 424504 32508 434144 39148
rect 423544 8128 434144 32508
rect 434944 8128 435104 534448
rect 435904 480367 486264 534448
rect 435904 480148 446504 480367
rect 435904 473428 445544 480148
rect 446344 473428 446504 480148
rect 435904 472937 446504 473428
rect 447304 472937 456944 480367
rect 457744 472937 457904 480367
rect 458704 472937 468344 480367
rect 469144 472937 469304 480367
rect 470104 472937 479744 480367
rect 480544 480148 486264 480367
rect 480544 473428 480704 480148
rect 481504 473428 486264 480148
rect 480544 472937 486264 473428
rect 435904 417367 486264 472937
rect 435904 417148 446504 417367
rect 435904 410428 445544 417148
rect 446344 410428 446504 417148
rect 435904 409937 446504 410428
rect 447304 409937 456944 417367
rect 457744 409937 457904 417367
rect 458704 409937 468344 417367
rect 469144 409937 469304 417367
rect 470104 409937 479744 417367
rect 480544 417148 486264 417367
rect 480544 410428 480704 417148
rect 481504 410428 486264 417148
rect 480544 409937 486264 410428
rect 435904 354367 486264 409937
rect 435904 354148 446504 354367
rect 435904 347428 445544 354148
rect 446344 347428 446504 354148
rect 435904 346937 446504 347428
rect 447304 346937 456944 354367
rect 457744 346937 457904 354367
rect 458704 346937 468344 354367
rect 469144 346937 469304 354367
rect 470104 346937 479744 354367
rect 480544 354148 486264 354367
rect 480544 347428 480704 354148
rect 481504 347428 486264 354148
rect 480544 346937 486264 347428
rect 435904 291367 486264 346937
rect 435904 291148 446504 291367
rect 435904 284428 445544 291148
rect 446344 284428 446504 291148
rect 435904 283937 446504 284428
rect 447304 283937 456944 291367
rect 457744 283937 457904 291367
rect 458704 283937 468344 291367
rect 469144 283937 469304 291367
rect 470104 283937 479744 291367
rect 480544 291148 486264 291367
rect 480544 284428 480704 291148
rect 481504 284428 486264 291148
rect 480544 283937 486264 284428
rect 435904 228367 486264 283937
rect 435904 228148 446504 228367
rect 435904 221428 445544 228148
rect 446344 221428 446504 228148
rect 435904 220937 446504 221428
rect 447304 220937 456944 228367
rect 457744 220937 457904 228367
rect 458704 220937 468344 228367
rect 469144 220937 469304 228367
rect 470104 220937 479744 228367
rect 480544 228148 486264 228367
rect 480544 221428 480704 228148
rect 481504 221428 486264 228148
rect 480544 220937 486264 221428
rect 435904 165367 486264 220937
rect 435904 165148 446504 165367
rect 435904 158428 445544 165148
rect 446344 158428 446504 165148
rect 435904 157937 446504 158428
rect 447304 157937 456944 165367
rect 457744 157937 457904 165367
rect 458704 157937 468344 165367
rect 469144 157937 469304 165367
rect 470104 157937 479744 165367
rect 480544 165148 486264 165367
rect 480544 158428 480704 165148
rect 481504 158428 486264 165148
rect 480544 157937 486264 158428
rect 435904 102367 486264 157937
rect 435904 102148 446504 102367
rect 435904 95428 445544 102148
rect 446344 95428 446504 102148
rect 435904 94937 446504 95428
rect 447304 94937 456944 102367
rect 457744 94937 457904 102367
rect 458704 94937 468344 102367
rect 469144 94937 469304 102367
rect 470104 94937 479744 102367
rect 480544 102148 486264 102367
rect 480544 95428 480704 102148
rect 481504 95428 486264 102148
rect 480544 94937 486264 95428
rect 435904 39367 486264 94937
rect 435904 39148 446504 39367
rect 435904 32508 445544 39148
rect 446344 32508 446504 39148
rect 435904 31609 446504 32508
rect 447304 31609 456944 39367
rect 457744 31609 457904 39367
rect 458704 31609 468344 39367
rect 435904 13167 468344 31609
rect 435904 8128 446504 13167
rect 447304 8128 456944 13167
rect 457744 8128 457904 13167
rect 458704 8128 468344 13167
rect 469144 8128 469304 39367
rect 470104 8128 479744 39367
rect 480544 39148 486264 39367
rect 480544 32508 480704 39148
rect 481504 32508 486264 39148
rect 480544 8128 486264 32508
<< metal5 >>
rect -2552 542696 497512 543656
rect -1192 541336 496152 542296
rect -2552 539356 497512 539996
rect -2552 530136 497512 530776
rect -2552 528856 497512 529496
rect -2552 519636 497512 520276
rect -2552 518356 497512 518996
rect -2552 509136 497512 509776
rect -2552 507856 497512 508496
rect -2552 498636 497512 499276
rect -2552 497356 497512 497996
rect -2552 488136 497512 488776
rect -2552 486856 497512 487496
rect -2552 477636 497512 478276
rect -2552 476356 497512 476996
rect -2552 467136 497512 467776
rect -2552 465856 497512 466496
rect -2552 456636 497512 457276
rect -2552 455356 497512 455996
rect -2552 446136 497512 446776
rect -2552 444856 497512 445496
rect -2552 435636 497512 436276
rect -2552 434356 497512 434996
rect -2552 425136 497512 425776
rect -2552 423856 497512 424496
rect -2552 414636 497512 415276
rect -2552 413356 497512 413996
rect -2552 404136 497512 404776
rect -2552 402856 497512 403496
rect -2552 393636 497512 394276
rect -2552 392356 497512 392996
rect -2552 383136 497512 383776
rect -2552 381856 497512 382496
rect -2552 372636 497512 373276
rect -2552 371356 497512 371996
rect -2552 362136 497512 362776
rect -2552 360856 497512 361496
rect -2552 351636 497512 352276
rect -2552 350356 497512 350996
rect -2552 341136 497512 341776
rect -2552 339856 497512 340496
rect -2552 330636 497512 331276
rect -2552 329356 497512 329996
rect -2552 320136 497512 320776
rect -2552 318856 497512 319496
rect -2552 309636 497512 310276
rect -2552 308356 497512 308996
rect -2552 299136 497512 299776
rect -2552 297856 497512 298496
rect -2552 288636 497512 289276
rect -2552 287356 497512 287996
rect -2552 278136 497512 278776
rect -2552 276856 497512 277496
rect -2552 267636 497512 268276
rect -2552 266356 497512 266996
rect -2552 257136 497512 257776
rect -2552 255856 497512 256496
rect -2552 246636 497512 247276
rect -2552 245356 497512 245996
rect -2552 236136 497512 236776
rect -2552 234856 497512 235496
rect -2552 225636 497512 226276
rect -2552 224356 497512 224996
rect -2552 215136 497512 215776
rect -2552 213856 497512 214496
rect -2552 204636 497512 205276
rect -2552 203356 497512 203996
rect -2552 194136 497512 194776
rect -2552 192856 497512 193496
rect -2552 183636 497512 184276
rect -2552 182356 497512 182996
rect -2552 173136 497512 173776
rect -2552 171856 497512 172496
rect -2552 162636 497512 163276
rect -2552 161356 497512 161996
rect -2552 152136 497512 152776
rect -2552 150856 497512 151496
rect -2552 141636 497512 142276
rect -2552 140356 497512 140996
rect -2552 131136 497512 131776
rect -2552 129856 497512 130496
rect -2552 120636 497512 121276
rect -2552 119356 497512 119996
rect -2552 110136 497512 110776
rect -2552 108856 497512 109496
rect -2552 99636 497512 100276
rect -2552 98356 497512 98996
rect -2552 89136 497512 89776
rect -2552 87856 497512 88496
rect -2552 78636 497512 79276
rect -2552 77356 497512 77996
rect -2552 68136 497512 68776
rect -2552 66856 497512 67496
rect -2552 57636 497512 58276
rect -2552 56356 497512 56996
rect -2552 47136 497512 47776
rect -2552 45856 497512 46496
rect -2552 36636 497512 37276
rect -2552 35356 497512 35996
rect -2552 26136 497512 26776
rect -2552 24856 497512 25496
rect -2552 15636 497512 16276
rect -2552 14356 497512 14996
rect -2552 5136 497512 5776
rect -2552 3856 497512 4496
rect -1192 616 496152 1576
rect -2552 -744 497512 216
<< labels >>
rlabel metal4 s -2552 -744 -1592 543656 4 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 -744 497512 216 8 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 542696 497512 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 496552 -744 497512 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 1984 -744 2624 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 13384 -744 14024 6068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 13384 34273 14024 39068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 13384 95508 14024 102068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 13384 158508 14024 165068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 13384 221508 14024 228068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 13384 284508 14024 291068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 13384 347508 14024 354068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 13384 410508 14024 417068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 13384 473508 14024 480068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 13384 536508 14024 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 24784 -744 25424 9415 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 24784 34273 25424 39559 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 24784 95017 25424 102559 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 24784 158017 25424 165559 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 24784 221017 25424 228559 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 24784 284017 25424 291559 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 24784 347017 25424 354559 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 24784 410017 25424 417559 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 24784 473017 25424 479743 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 24784 508001 25424 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 36184 -744 36824 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 47584 -744 48224 40919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 47584 95017 48224 103919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 47584 158017 48224 166919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 47584 221017 48224 229919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 47584 284017 48224 292919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 47584 347017 48224 355919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 47584 410017 48224 418919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 47584 473017 48224 483687 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 47584 533977 48224 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 58984 -744 59624 12951 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 58984 32097 59624 40919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 58984 95017 59624 103919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 58984 158017 59624 166919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 58984 221017 59624 229919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 58984 284017 59624 292919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 58984 347017 59624 355919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 58984 410017 59624 418919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 58984 473017 59624 483687 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 58984 533977 59624 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 70384 -744 71024 12951 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 70384 32097 71024 40919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 70384 95017 71024 103919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 70384 158017 71024 166919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 70384 221017 71024 229919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 70384 284017 71024 292919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 70384 347017 71024 355919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 70384 410017 71024 418919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 70384 473017 71024 483687 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 70384 533977 71024 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 81784 -744 82424 6068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 81784 32588 82424 39068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 81784 95508 82424 102068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 81784 158508 82424 165068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 81784 221508 82424 228068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 81784 284508 82424 291068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 81784 347508 82424 354068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 81784 410508 82424 417068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 81784 473508 82424 480068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 81784 536508 82424 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 93184 -744 93824 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 104584 -744 105224 40919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 104584 95017 105224 103919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 104584 158017 105224 166919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 104584 221017 105224 229919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 104584 284017 105224 292919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 104584 347017 105224 355919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 104584 410017 105224 418919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 104584 473017 105224 483687 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 104584 533977 105224 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 115984 -744 116624 12951 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 115984 32097 116624 40919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 115984 95017 116624 103919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 115984 158017 116624 166919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 115984 221017 116624 229919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 115984 284017 116624 292919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 115984 347017 116624 355919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 115984 410017 116624 418919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 115984 473017 116624 483687 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 115984 533977 116624 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 127384 -744 128024 12951 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 127384 32097 128024 40919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 127384 95017 128024 103919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 127384 158017 128024 166919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 127384 221017 128024 229919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 127384 284017 128024 292919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 127384 347017 128024 355919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 127384 410017 128024 418919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 127384 473017 128024 483687 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 127384 533977 128024 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 138784 -744 139424 6068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 138784 32588 139424 39068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 138784 95508 139424 102068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 138784 158508 139424 165068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 138784 221508 139424 228068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 138784 284508 139424 291068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 138784 347508 139424 354068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 138784 410508 139424 417068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 138784 473508 139424 480068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 138784 536508 139424 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 150184 -744 150824 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 161584 -744 162224 40919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 161584 95017 162224 103919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 161584 158017 162224 166919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 161584 221017 162224 229919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 161584 284017 162224 292919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 161584 347017 162224 355919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 161584 410017 162224 418919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 161584 473017 162224 483687 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 161584 533977 162224 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 172984 -744 173624 12951 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 172984 32097 173624 40919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 172984 95017 173624 103919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 172984 158017 173624 166919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 172984 221017 173624 229919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 172984 284017 173624 292919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 172984 347017 173624 355919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 172984 410017 173624 418919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 172984 473017 173624 483687 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 172984 533977 173624 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 184384 -744 185024 12951 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 184384 32097 185024 40919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 184384 95017 185024 103919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 184384 158017 185024 166919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 184384 221017 185024 229919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 184384 284017 185024 292919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 184384 347017 185024 355919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 184384 410017 185024 418919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 184384 473017 185024 483687 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 184384 533977 185024 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 195784 -744 196424 6068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 195784 32588 196424 39068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 195784 95508 196424 102068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 195784 158508 196424 165068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 195784 221508 196424 228068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 195784 284508 196424 291068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 195784 347508 196424 354068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 195784 410508 196424 417068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 195784 473508 196424 480068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 195784 536508 196424 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 207184 -744 207824 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 218584 -744 219224 40919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 218584 95017 219224 103919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 218584 158017 219224 166919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 218584 221017 219224 229919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 218584 284017 219224 292919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 218584 347017 219224 355919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 218584 410017 219224 418919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 218584 473017 219224 483687 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 218584 533977 219224 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 229984 -744 230624 12951 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 229984 32097 230624 40919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 229984 95017 230624 103919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 229984 158017 230624 166919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 229984 221017 230624 229919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 229984 284017 230624 292919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 229984 347017 230624 355919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 229984 410017 230624 418919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 229984 473017 230624 483687 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 229984 533977 230624 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 241384 -744 242024 12951 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 241384 32097 242024 40919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 241384 95017 242024 103919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 241384 158017 242024 166919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 241384 221017 242024 229919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 241384 284017 242024 292919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 241384 347017 242024 355919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 241384 410017 242024 418919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 241384 473017 242024 483687 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 241384 533977 242024 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 252784 -744 253424 6068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 252784 32588 253424 39068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 252784 95508 253424 102068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 252784 158508 253424 165068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 252784 221508 253424 228068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 252784 284508 253424 291068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 252784 347508 253424 354068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 252784 410508 253424 417068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 252784 473508 253424 480068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 252784 536508 253424 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 264184 -744 264824 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 275584 -744 276224 40919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 275584 95017 276224 103919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 275584 158017 276224 166919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 275584 221017 276224 229919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 275584 284017 276224 292919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 275584 347017 276224 355919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 275584 410017 276224 418919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 275584 473017 276224 483687 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 275584 533977 276224 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 286984 -744 287624 12951 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 286984 32097 287624 40919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 286984 95017 287624 103919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 286984 158017 287624 166919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 286984 221017 287624 229919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 286984 284017 287624 292919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 286984 347017 287624 355919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 286984 410017 287624 418919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 286984 473017 287624 483687 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 286984 533977 287624 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 298384 -744 299024 12951 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 298384 32097 299024 40919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 298384 95017 299024 103919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 298384 158017 299024 166919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 298384 221017 299024 229919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 298384 284017 299024 292919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 298384 347017 299024 355919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 298384 410017 299024 418919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 298384 473017 299024 483687 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 298384 533977 299024 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 309784 -744 310424 6068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 309784 32588 310424 39068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 309784 95508 310424 102068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 309784 158508 310424 165068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 309784 221508 310424 228068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 309784 284508 310424 291068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 309784 347508 310424 354068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 309784 410508 310424 417068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 309784 473508 310424 480068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 309784 536508 310424 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 321184 -744 321824 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 332584 -744 333224 40919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 332584 95017 333224 103919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 332584 158017 333224 166919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 332584 221017 333224 229919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 332584 284017 333224 292919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 332584 347017 333224 355919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 332584 410017 333224 418919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 332584 473017 333224 483687 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 332584 533977 333224 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 343984 -744 344624 12951 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 343984 32097 344624 40919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 343984 95017 344624 103919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 343984 158017 344624 166919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 343984 221017 344624 229919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 343984 284017 344624 292919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 343984 347017 344624 355919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 343984 410017 344624 418919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 343984 473017 344624 483687 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 343984 533977 344624 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 355384 -744 356024 12951 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 355384 32097 356024 40919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 355384 95017 356024 103919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 355384 158017 356024 166919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 355384 221017 356024 229919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 355384 284017 356024 292919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 355384 347017 356024 355919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 355384 410017 356024 418919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 355384 473017 356024 483687 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 355384 533977 356024 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 366784 -744 367424 6068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 366784 32588 367424 39068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 366784 95508 367424 102068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 366784 158508 367424 165068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 366784 221508 367424 228068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 366784 284508 367424 291068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 366784 347508 367424 354068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 366784 410508 367424 417068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 366784 473508 367424 480068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 366784 536508 367424 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 378184 -744 378824 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 389584 -744 390224 40919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 389584 95017 390224 103919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 389584 158017 390224 166919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 389584 221017 390224 229919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 389584 284017 390224 292919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 389584 347017 390224 355919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 389584 410017 390224 418919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 389584 473017 390224 483687 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 389584 533977 390224 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 400984 -744 401624 12951 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 400984 32097 401624 40919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 400984 95017 401624 103919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 400984 158017 401624 166919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 400984 221017 401624 229919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 400984 284017 401624 292919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 400984 347017 401624 355919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 400984 410017 401624 418919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 400984 473017 401624 483687 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 400984 533977 401624 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 412384 -744 413024 12951 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 412384 32097 413024 40919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 412384 95017 413024 103919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 412384 158017 413024 166919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 412384 221017 413024 229919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 412384 284017 413024 292919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 412384 347017 413024 355919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 412384 410017 413024 418919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 412384 473017 413024 483687 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 412384 533977 413024 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 423784 -744 424424 6068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 423784 32588 424424 39068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 423784 95508 424424 102068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 423784 158508 424424 165068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 423784 221508 424424 228068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 423784 284508 424424 291068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 423784 347508 424424 354068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 423784 410508 424424 417068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 423784 473508 424424 480068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 423784 536508 424424 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 435184 -744 435824 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 446584 -744 447224 13087 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 446584 31689 447224 39287 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 446584 95017 447224 102287 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 446584 158017 447224 165287 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 446584 221017 447224 228287 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 446584 284017 447224 291287 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 446584 347017 447224 354287 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 446584 410017 447224 417287 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 446584 473017 447224 480287 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 446584 536017 447224 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 457984 -744 458624 13087 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 457984 31689 458624 39287 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 457984 95017 458624 102287 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 457984 158017 458624 165287 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 457984 221017 458624 228287 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 457984 284017 458624 291287 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 457984 347017 458624 354287 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 457984 410017 458624 417287 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 457984 473017 458624 480287 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 457984 536017 458624 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 469384 -744 470024 39287 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 469384 95017 470024 102287 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 469384 158017 470024 165287 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 469384 221017 470024 228287 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 469384 284017 470024 291287 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 469384 347017 470024 354287 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 469384 410017 470024 417287 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 469384 473017 470024 480287 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 469384 536017 470024 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 480784 -744 481424 6068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 480784 32588 481424 39068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 480784 95508 481424 102068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 480784 158508 481424 165068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 480784 221508 481424 228068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 480784 284508 481424 291068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 480784 347508 481424 354068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 480784 410508 481424 417068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 480784 473508 481424 480068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 480784 536508 481424 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 492184 -744 492824 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 5136 497512 5776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 15636 497512 16276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 26136 497512 26776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 36636 497512 37276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 47136 497512 47776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 57636 497512 58276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 68136 497512 68776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 78636 497512 79276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 89136 497512 89776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 99636 497512 100276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 110136 497512 110776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 120636 497512 121276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 131136 497512 131776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 141636 497512 142276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 152136 497512 152776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 162636 497512 163276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 173136 497512 173776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 183636 497512 184276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 194136 497512 194776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 204636 497512 205276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 215136 497512 215776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 225636 497512 226276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 236136 497512 236776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 246636 497512 247276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 257136 497512 257776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 267636 497512 268276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 278136 497512 278776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 288636 497512 289276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 299136 497512 299776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 309636 497512 310276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 320136 497512 320776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 330636 497512 331276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 341136 497512 341776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 351636 497512 352276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 362136 497512 362776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 372636 497512 373276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 383136 497512 383776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 393636 497512 394276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 404136 497512 404776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 414636 497512 415276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 425136 497512 425776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 435636 497512 436276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 446136 497512 446776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 456636 497512 457276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 467136 497512 467776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 477636 497512 478276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 488136 497512 488776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 498636 497512 499276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 509136 497512 509776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 519636 497512 520276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 530136 497512 530776 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s -1192 616 -232 542296 4 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -1192 616 496152 1576 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -1192 541336 496152 542296 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 495192 616 496152 542296 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 1024 -744 1664 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 12424 -744 13064 9415 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 12424 34273 13064 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 23824 -744 24464 6068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 23824 34273 24464 39068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 23824 95508 24464 102068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 23824 158508 24464 165068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 23824 221508 24464 228068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 23824 284508 24464 291068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 23824 347508 24464 354068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 23824 410508 24464 417068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 23824 473508 24464 479743 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 23824 536508 24464 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 35224 -744 35864 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 46624 -744 47264 6068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 46624 32588 47264 39068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 46624 95508 47264 102068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 46624 158508 47264 165068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 46624 221508 47264 228068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 46624 284508 47264 291068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 46624 347508 47264 354068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 46624 410508 47264 417068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 46624 473508 47264 480068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 46624 536508 47264 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 58024 -744 58664 12951 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 58024 32097 58664 40919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 58024 95017 58664 103919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 58024 158017 58664 166919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 58024 221017 58664 229919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 58024 284017 58664 292919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 58024 347017 58664 355919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 58024 410017 58664 418919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 58024 473017 58664 483687 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 58024 533977 58664 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 69424 -744 70064 12951 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 69424 32097 70064 40919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 69424 95017 70064 103919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 69424 158017 70064 166919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 69424 221017 70064 229919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 69424 284017 70064 292919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 69424 347017 70064 355919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 69424 410017 70064 418919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 69424 473017 70064 483687 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 69424 533977 70064 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 80824 -744 81464 40919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 80824 95017 81464 103919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 80824 158017 81464 166919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 80824 221017 81464 229919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 80824 284017 81464 292919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 80824 347017 81464 355919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 80824 410017 81464 418919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 80824 473017 81464 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 92224 -744 92864 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 103624 -744 104264 6068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 103624 32588 104264 39068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 103624 95508 104264 102068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 103624 158508 104264 165068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 103624 221508 104264 228068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 103624 284508 104264 291068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 103624 347508 104264 354068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 103624 410508 104264 417068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 103624 473508 104264 480068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 103624 536508 104264 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 115024 -744 115664 12951 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 115024 32097 115664 40919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 115024 95017 115664 103919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 115024 158017 115664 166919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 115024 221017 115664 229919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 115024 284017 115664 292919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 115024 347017 115664 355919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 115024 410017 115664 418919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 115024 473017 115664 483687 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 115024 533977 115664 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 126424 -744 127064 12951 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 126424 32097 127064 40919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 126424 95017 127064 103919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 126424 158017 127064 166919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 126424 221017 127064 229919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 126424 284017 127064 292919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 126424 347017 127064 355919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 126424 410017 127064 418919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 126424 473017 127064 483687 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 126424 533977 127064 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 137824 -744 138464 40919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 137824 95017 138464 103919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 137824 158017 138464 166919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 137824 221017 138464 229919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 137824 284017 138464 292919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 137824 347017 138464 355919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 137824 410017 138464 418919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 137824 473017 138464 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 149224 -744 149864 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 160624 -744 161264 6068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 160624 32588 161264 39068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 160624 95508 161264 102068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 160624 158508 161264 165068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 160624 221508 161264 228068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 160624 284508 161264 291068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 160624 347508 161264 354068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 160624 410508 161264 417068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 160624 473508 161264 480068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 160624 536508 161264 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 172024 -744 172664 12951 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 172024 32097 172664 40919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 172024 95017 172664 103919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 172024 158017 172664 166919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 172024 221017 172664 229919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 172024 284017 172664 292919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 172024 347017 172664 355919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 172024 410017 172664 418919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 172024 473017 172664 483687 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 172024 533977 172664 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 183424 -744 184064 12951 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 183424 32097 184064 40919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 183424 95017 184064 103919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 183424 158017 184064 166919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 183424 221017 184064 229919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 183424 284017 184064 292919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 183424 347017 184064 355919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 183424 410017 184064 418919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 183424 473017 184064 483687 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 183424 533977 184064 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 194824 -744 195464 40919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 194824 95017 195464 103919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 194824 158017 195464 166919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 194824 221017 195464 229919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 194824 284017 195464 292919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 194824 347017 195464 355919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 194824 410017 195464 418919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 194824 473017 195464 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 206224 -744 206864 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 217624 -744 218264 6068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 217624 32588 218264 39068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 217624 95508 218264 102068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 217624 158508 218264 165068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 217624 221508 218264 228068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 217624 284508 218264 291068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 217624 347508 218264 354068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 217624 410508 218264 417068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 217624 473508 218264 480068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 217624 536508 218264 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 229024 -744 229664 12951 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 229024 32097 229664 40919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 229024 95017 229664 103919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 229024 158017 229664 166919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 229024 221017 229664 229919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 229024 284017 229664 292919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 229024 347017 229664 355919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 229024 410017 229664 418919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 229024 473017 229664 483687 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 229024 533977 229664 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 240424 -744 241064 12951 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 240424 32097 241064 40919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 240424 95017 241064 103919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 240424 158017 241064 166919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 240424 221017 241064 229919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 240424 284017 241064 292919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 240424 347017 241064 355919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 240424 410017 241064 418919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 240424 473017 241064 483687 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 240424 533977 241064 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 251824 -744 252464 40919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 251824 95017 252464 103919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 251824 158017 252464 166919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 251824 221017 252464 229919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 251824 284017 252464 292919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 251824 347017 252464 355919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 251824 410017 252464 418919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 251824 473017 252464 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 263224 -744 263864 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 274624 -744 275264 6068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 274624 32588 275264 39068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 274624 95508 275264 102068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 274624 158508 275264 165068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 274624 221508 275264 228068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 274624 284508 275264 291068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 274624 347508 275264 354068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 274624 410508 275264 417068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 274624 473508 275264 480068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 274624 536508 275264 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 286024 -744 286664 12951 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 286024 32097 286664 40919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 286024 95017 286664 103919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 286024 158017 286664 166919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 286024 221017 286664 229919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 286024 284017 286664 292919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 286024 347017 286664 355919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 286024 410017 286664 418919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 286024 473017 286664 483687 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 286024 533977 286664 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 297424 -744 298064 12951 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 297424 32097 298064 40919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 297424 95017 298064 103919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 297424 158017 298064 166919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 297424 221017 298064 229919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 297424 284017 298064 292919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 297424 347017 298064 355919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 297424 410017 298064 418919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 297424 473017 298064 483687 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 297424 533977 298064 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 308824 -744 309464 40919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 308824 95017 309464 103919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 308824 158017 309464 166919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 308824 221017 309464 229919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 308824 284017 309464 292919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 308824 347017 309464 355919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 308824 410017 309464 418919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 308824 473017 309464 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 320224 -744 320864 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 331624 -744 332264 6068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 331624 32588 332264 39068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 331624 95508 332264 102068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 331624 158508 332264 165068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 331624 221508 332264 228068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 331624 284508 332264 291068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 331624 347508 332264 354068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 331624 410508 332264 417068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 331624 473508 332264 480068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 331624 536508 332264 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 343024 -744 343664 12951 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 343024 32097 343664 40919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 343024 95017 343664 103919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 343024 158017 343664 166919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 343024 221017 343664 229919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 343024 284017 343664 292919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 343024 347017 343664 355919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 343024 410017 343664 418919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 343024 473017 343664 483687 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 343024 533977 343664 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 354424 -744 355064 12951 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 354424 32097 355064 40919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 354424 95017 355064 103919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 354424 158017 355064 166919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 354424 221017 355064 229919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 354424 284017 355064 292919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 354424 347017 355064 355919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 354424 410017 355064 418919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 354424 473017 355064 483687 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 354424 533977 355064 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 365824 -744 366464 40919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 365824 95017 366464 103919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 365824 158017 366464 166919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 365824 221017 366464 229919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 365824 284017 366464 292919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 365824 347017 366464 355919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 365824 410017 366464 418919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 365824 473017 366464 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 377224 -744 377864 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 388624 -744 389264 6068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 388624 32588 389264 39068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 388624 95508 389264 102068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 388624 158508 389264 165068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 388624 221508 389264 228068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 388624 284508 389264 291068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 388624 347508 389264 354068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 388624 410508 389264 417068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 388624 473508 389264 480068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 388624 536508 389264 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 400024 -744 400664 12951 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 400024 32097 400664 40919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 400024 95017 400664 103919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 400024 158017 400664 166919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 400024 221017 400664 229919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 400024 284017 400664 292919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 400024 347017 400664 355919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 400024 410017 400664 418919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 400024 473017 400664 483687 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 400024 533977 400664 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 411424 -744 412064 12951 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 411424 32097 412064 40919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 411424 95017 412064 103919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 411424 158017 412064 166919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 411424 221017 412064 229919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 411424 284017 412064 292919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 411424 347017 412064 355919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 411424 410017 412064 418919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 411424 473017 412064 483687 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 411424 533977 412064 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 422824 -744 423464 40919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 422824 95017 423464 103919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 422824 158017 423464 166919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 422824 221017 423464 229919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 422824 284017 423464 292919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 422824 347017 423464 355919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 422824 410017 423464 418919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 422824 473017 423464 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 434224 -744 434864 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 445624 -744 446264 6068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 445624 32588 446264 39068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 445624 95508 446264 102068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 445624 158508 446264 165068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 445624 221508 446264 228068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 445624 284508 446264 291068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 445624 347508 446264 354068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 445624 410508 446264 417068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 445624 473508 446264 480068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 445624 536508 446264 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 457024 -744 457664 13087 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 457024 31689 457664 39287 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 457024 95017 457664 102287 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 457024 158017 457664 165287 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 457024 221017 457664 228287 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 457024 284017 457664 291287 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 457024 347017 457664 354287 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 457024 410017 457664 417287 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 457024 473017 457664 480287 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 457024 536017 457664 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 468424 -744 469064 39287 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 468424 95017 469064 102287 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 468424 158017 469064 165287 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 468424 221017 469064 228287 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 468424 284017 469064 291287 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 468424 347017 469064 354287 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 468424 410017 469064 417287 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 468424 473017 469064 480287 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 468424 536017 469064 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 479824 -744 480464 39287 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 479824 95017 480464 102287 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 479824 158017 480464 165287 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 479824 221017 480464 228287 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 479824 284017 480464 291287 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 479824 347017 480464 354287 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 479824 410017 480464 417287 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 479824 473017 480464 480287 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 479824 536017 480464 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 491224 -744 491864 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 3856 497512 4496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 14356 497512 14996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 24856 497512 25496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 35356 497512 35996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 45856 497512 46496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 56356 497512 56996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 66856 497512 67496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 77356 497512 77996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 87856 497512 88496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 98356 497512 98996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 108856 497512 109496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 119356 497512 119996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 129856 497512 130496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 140356 497512 140996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 150856 497512 151496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 161356 497512 161996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 171856 497512 172496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 182356 497512 182996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 192856 497512 193496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 203356 497512 203996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 213856 497512 214496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 224356 497512 224996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 234856 497512 235496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 245356 497512 245996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 255856 497512 256496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 266356 497512 266996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 276856 497512 277496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 287356 497512 287996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 297856 497512 298496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 308356 497512 308996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 318856 497512 319496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 329356 497512 329996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 339856 497512 340496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 350356 497512 350996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 360856 497512 361496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 371356 497512 371996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 381856 497512 382496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 392356 497512 392996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 402856 497512 403496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 413356 497512 413996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 423856 497512 424496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 434356 497512 434996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 444856 497512 445496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 455356 497512 455996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 465856 497512 466496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 476356 497512 476996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 486856 497512 487496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 497356 497512 497996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 507856 497512 508496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 518356 497512 518996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 528856 497512 529496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 539356 497512 539996 6 VPWR
port 2 nsew power bidirectional
rlabel metal2 s 73526 0 73582 800 6 ccff_head
port 3 nsew signal input
rlabel metal2 s 59726 542200 59782 543000 6 ccff_tail
port 4 nsew signal output
rlabel metal3 s 0 10208 800 10328 6 clk
port 5 nsew signal input
rlabel metal2 s 15566 542200 15622 543000 6 gfpga_pad_io_soc_dir[0]
port 6 nsew signal output
rlabel metal3 s 0 91808 800 91928 6 gfpga_pad_io_soc_dir[100]
port 7 nsew signal output
rlabel metal3 s 0 108128 800 108248 6 gfpga_pad_io_soc_dir[101]
port 8 nsew signal output
rlabel metal3 s 0 124448 800 124568 6 gfpga_pad_io_soc_dir[102]
port 9 nsew signal output
rlabel metal3 s 0 140768 800 140888 6 gfpga_pad_io_soc_dir[103]
port 10 nsew signal output
rlabel metal3 s 0 157088 800 157208 6 gfpga_pad_io_soc_dir[104]
port 11 nsew signal output
rlabel metal3 s 0 173408 800 173528 6 gfpga_pad_io_soc_dir[105]
port 12 nsew signal output
rlabel metal3 s 0 189728 800 189848 6 gfpga_pad_io_soc_dir[106]
port 13 nsew signal output
rlabel metal3 s 0 206048 800 206168 6 gfpga_pad_io_soc_dir[107]
port 14 nsew signal output
rlabel metal3 s 0 222368 800 222488 6 gfpga_pad_io_soc_dir[108]
port 15 nsew signal output
rlabel metal3 s 0 238688 800 238808 6 gfpga_pad_io_soc_dir[109]
port 16 nsew signal output
rlabel metal2 s 156878 542200 156934 543000 6 gfpga_pad_io_soc_dir[10]
port 17 nsew signal output
rlabel metal3 s 0 255008 800 255128 6 gfpga_pad_io_soc_dir[110]
port 18 nsew signal output
rlabel metal3 s 0 276768 800 276888 6 gfpga_pad_io_soc_dir[111]
port 19 nsew signal output
rlabel metal3 s 0 293088 800 293208 6 gfpga_pad_io_soc_dir[112]
port 20 nsew signal output
rlabel metal3 s 0 309408 800 309528 6 gfpga_pad_io_soc_dir[113]
port 21 nsew signal output
rlabel metal3 s 0 325728 800 325848 6 gfpga_pad_io_soc_dir[114]
port 22 nsew signal output
rlabel metal3 s 0 342048 800 342168 6 gfpga_pad_io_soc_dir[115]
port 23 nsew signal output
rlabel metal3 s 0 358368 800 358488 6 gfpga_pad_io_soc_dir[116]
port 24 nsew signal output
rlabel metal3 s 0 374688 800 374808 6 gfpga_pad_io_soc_dir[117]
port 25 nsew signal output
rlabel metal3 s 0 391008 800 391128 6 gfpga_pad_io_soc_dir[118]
port 26 nsew signal output
rlabel metal3 s 0 407328 800 407448 6 gfpga_pad_io_soc_dir[119]
port 27 nsew signal output
rlabel metal2 s 170126 542200 170182 543000 6 gfpga_pad_io_soc_dir[11]
port 28 nsew signal output
rlabel metal3 s 0 423648 800 423768 6 gfpga_pad_io_soc_dir[120]
port 29 nsew signal output
rlabel metal3 s 0 439968 800 440088 6 gfpga_pad_io_soc_dir[121]
port 30 nsew signal output
rlabel metal3 s 0 456288 800 456408 6 gfpga_pad_io_soc_dir[122]
port 31 nsew signal output
rlabel metal3 s 0 472608 800 472728 6 gfpga_pad_io_soc_dir[123]
port 32 nsew signal output
rlabel metal3 s 0 488928 800 489048 6 gfpga_pad_io_soc_dir[124]
port 33 nsew signal output
rlabel metal3 s 0 505248 800 505368 6 gfpga_pad_io_soc_dir[125]
port 34 nsew signal output
rlabel metal3 s 0 521568 800 521688 6 gfpga_pad_io_soc_dir[126]
port 35 nsew signal output
rlabel metal3 s 0 537888 800 538008 6 gfpga_pad_io_soc_dir[127]
port 36 nsew signal output
rlabel metal2 s 183374 542200 183430 543000 6 gfpga_pad_io_soc_dir[12]
port 37 nsew signal output
rlabel metal2 s 196622 542200 196678 543000 6 gfpga_pad_io_soc_dir[13]
port 38 nsew signal output
rlabel metal2 s 209870 542200 209926 543000 6 gfpga_pad_io_soc_dir[14]
port 39 nsew signal output
rlabel metal2 s 223118 542200 223174 543000 6 gfpga_pad_io_soc_dir[15]
port 40 nsew signal output
rlabel metal2 s 236366 542200 236422 543000 6 gfpga_pad_io_soc_dir[16]
port 41 nsew signal output
rlabel metal2 s 249614 542200 249670 543000 6 gfpga_pad_io_soc_dir[17]
port 42 nsew signal output
rlabel metal2 s 262862 542200 262918 543000 6 gfpga_pad_io_soc_dir[18]
port 43 nsew signal output
rlabel metal2 s 276110 542200 276166 543000 6 gfpga_pad_io_soc_dir[19]
port 44 nsew signal output
rlabel metal2 s 28814 542200 28870 543000 6 gfpga_pad_io_soc_dir[1]
port 45 nsew signal output
rlabel metal2 s 289358 542200 289414 543000 6 gfpga_pad_io_soc_dir[20]
port 46 nsew signal output
rlabel metal2 s 302606 542200 302662 543000 6 gfpga_pad_io_soc_dir[21]
port 47 nsew signal output
rlabel metal2 s 315854 542200 315910 543000 6 gfpga_pad_io_soc_dir[22]
port 48 nsew signal output
rlabel metal2 s 329102 542200 329158 543000 6 gfpga_pad_io_soc_dir[23]
port 49 nsew signal output
rlabel metal2 s 342350 542200 342406 543000 6 gfpga_pad_io_soc_dir[24]
port 50 nsew signal output
rlabel metal2 s 355598 542200 355654 543000 6 gfpga_pad_io_soc_dir[25]
port 51 nsew signal output
rlabel metal2 s 368846 542200 368902 543000 6 gfpga_pad_io_soc_dir[26]
port 52 nsew signal output
rlabel metal2 s 382094 542200 382150 543000 6 gfpga_pad_io_soc_dir[27]
port 53 nsew signal output
rlabel metal2 s 395342 542200 395398 543000 6 gfpga_pad_io_soc_dir[28]
port 54 nsew signal output
rlabel metal2 s 408590 542200 408646 543000 6 gfpga_pad_io_soc_dir[29]
port 55 nsew signal output
rlabel metal2 s 42062 542200 42118 543000 6 gfpga_pad_io_soc_dir[2]
port 56 nsew signal output
rlabel metal2 s 421838 542200 421894 543000 6 gfpga_pad_io_soc_dir[30]
port 57 nsew signal output
rlabel metal2 s 435086 542200 435142 543000 6 gfpga_pad_io_soc_dir[31]
port 58 nsew signal output
rlabel metal2 s 448334 542200 448390 543000 6 gfpga_pad_io_soc_dir[32]
port 59 nsew signal output
rlabel metal2 s 461582 542200 461638 543000 6 gfpga_pad_io_soc_dir[33]
port 60 nsew signal output
rlabel metal2 s 474830 542200 474886 543000 6 gfpga_pad_io_soc_dir[34]
port 61 nsew signal output
rlabel metal2 s 488078 542200 488134 543000 6 gfpga_pad_io_soc_dir[35]
port 62 nsew signal output
rlabel metal3 s 494200 518032 495000 518152 6 gfpga_pad_io_soc_dir[36]
port 63 nsew signal output
rlabel metal3 s 494200 502120 495000 502240 6 gfpga_pad_io_soc_dir[37]
port 64 nsew signal output
rlabel metal3 s 494200 486208 495000 486328 6 gfpga_pad_io_soc_dir[38]
port 65 nsew signal output
rlabel metal3 s 494200 470296 495000 470416 6 gfpga_pad_io_soc_dir[39]
port 66 nsew signal output
rlabel metal2 s 55310 542200 55366 543000 6 gfpga_pad_io_soc_dir[3]
port 67 nsew signal output
rlabel metal3 s 494200 454384 495000 454504 6 gfpga_pad_io_soc_dir[40]
port 68 nsew signal output
rlabel metal3 s 494200 438472 495000 438592 6 gfpga_pad_io_soc_dir[41]
port 69 nsew signal output
rlabel metal3 s 494200 422560 495000 422680 6 gfpga_pad_io_soc_dir[42]
port 70 nsew signal output
rlabel metal3 s 494200 406648 495000 406768 6 gfpga_pad_io_soc_dir[43]
port 71 nsew signal output
rlabel metal3 s 494200 390736 495000 390856 6 gfpga_pad_io_soc_dir[44]
port 72 nsew signal output
rlabel metal3 s 494200 374824 495000 374944 6 gfpga_pad_io_soc_dir[45]
port 73 nsew signal output
rlabel metal3 s 494200 358912 495000 359032 6 gfpga_pad_io_soc_dir[46]
port 74 nsew signal output
rlabel metal3 s 494200 343000 495000 343120 6 gfpga_pad_io_soc_dir[47]
port 75 nsew signal output
rlabel metal3 s 494200 327088 495000 327208 6 gfpga_pad_io_soc_dir[48]
port 76 nsew signal output
rlabel metal3 s 494200 311176 495000 311296 6 gfpga_pad_io_soc_dir[49]
port 77 nsew signal output
rlabel metal2 s 77390 542200 77446 543000 6 gfpga_pad_io_soc_dir[4]
port 78 nsew signal output
rlabel metal3 s 494200 295264 495000 295384 6 gfpga_pad_io_soc_dir[50]
port 79 nsew signal output
rlabel metal3 s 494200 279352 495000 279472 6 gfpga_pad_io_soc_dir[51]
port 80 nsew signal output
rlabel metal3 s 494200 263440 495000 263560 6 gfpga_pad_io_soc_dir[52]
port 81 nsew signal output
rlabel metal3 s 494200 247528 495000 247648 6 gfpga_pad_io_soc_dir[53]
port 82 nsew signal output
rlabel metal3 s 494200 221008 495000 221128 6 gfpga_pad_io_soc_dir[54]
port 83 nsew signal output
rlabel metal3 s 494200 205096 495000 205216 6 gfpga_pad_io_soc_dir[55]
port 84 nsew signal output
rlabel metal3 s 494200 189184 495000 189304 6 gfpga_pad_io_soc_dir[56]
port 85 nsew signal output
rlabel metal3 s 494200 173272 495000 173392 6 gfpga_pad_io_soc_dir[57]
port 86 nsew signal output
rlabel metal3 s 494200 157360 495000 157480 6 gfpga_pad_io_soc_dir[58]
port 87 nsew signal output
rlabel metal3 s 494200 141448 495000 141568 6 gfpga_pad_io_soc_dir[59]
port 88 nsew signal output
rlabel metal2 s 90638 542200 90694 543000 6 gfpga_pad_io_soc_dir[5]
port 89 nsew signal output
rlabel metal3 s 494200 125536 495000 125656 6 gfpga_pad_io_soc_dir[60]
port 90 nsew signal output
rlabel metal3 s 494200 109624 495000 109744 6 gfpga_pad_io_soc_dir[61]
port 91 nsew signal output
rlabel metal3 s 494200 93712 495000 93832 6 gfpga_pad_io_soc_dir[62]
port 92 nsew signal output
rlabel metal3 s 494200 77800 495000 77920 6 gfpga_pad_io_soc_dir[63]
port 93 nsew signal output
rlabel metal3 s 494200 61888 495000 62008 6 gfpga_pad_io_soc_dir[64]
port 94 nsew signal output
rlabel metal3 s 494200 45976 495000 46096 6 gfpga_pad_io_soc_dir[65]
port 95 nsew signal output
rlabel metal3 s 494200 30064 495000 30184 6 gfpga_pad_io_soc_dir[66]
port 96 nsew signal output
rlabel metal3 s 494200 14152 495000 14272 6 gfpga_pad_io_soc_dir[67]
port 97 nsew signal output
rlabel metal2 s 479246 0 479302 800 6 gfpga_pad_io_soc_dir[68]
port 98 nsew signal output
rlabel metal2 s 461858 0 461914 800 6 gfpga_pad_io_soc_dir[69]
port 99 nsew signal output
rlabel metal2 s 103886 542200 103942 543000 6 gfpga_pad_io_soc_dir[6]
port 100 nsew signal output
rlabel metal2 s 444470 0 444526 800 6 gfpga_pad_io_soc_dir[70]
port 101 nsew signal output
rlabel metal2 s 427082 0 427138 800 6 gfpga_pad_io_soc_dir[71]
port 102 nsew signal output
rlabel metal2 s 409694 0 409750 800 6 gfpga_pad_io_soc_dir[72]
port 103 nsew signal output
rlabel metal2 s 392306 0 392362 800 6 gfpga_pad_io_soc_dir[73]
port 104 nsew signal output
rlabel metal2 s 374918 0 374974 800 6 gfpga_pad_io_soc_dir[74]
port 105 nsew signal output
rlabel metal2 s 357530 0 357586 800 6 gfpga_pad_io_soc_dir[75]
port 106 nsew signal output
rlabel metal2 s 340142 0 340198 800 6 gfpga_pad_io_soc_dir[76]
port 107 nsew signal output
rlabel metal2 s 322754 0 322810 800 6 gfpga_pad_io_soc_dir[77]
port 108 nsew signal output
rlabel metal2 s 305366 0 305422 800 6 gfpga_pad_io_soc_dir[78]
port 109 nsew signal output
rlabel metal2 s 287978 0 288034 800 6 gfpga_pad_io_soc_dir[79]
port 110 nsew signal output
rlabel metal2 s 117134 542200 117190 543000 6 gfpga_pad_io_soc_dir[7]
port 111 nsew signal output
rlabel metal2 s 270590 0 270646 800 6 gfpga_pad_io_soc_dir[80]
port 112 nsew signal output
rlabel metal2 s 253202 0 253258 800 6 gfpga_pad_io_soc_dir[81]
port 113 nsew signal output
rlabel metal2 s 235814 0 235870 800 6 gfpga_pad_io_soc_dir[82]
port 114 nsew signal output
rlabel metal2 s 218426 0 218482 800 6 gfpga_pad_io_soc_dir[83]
port 115 nsew signal output
rlabel metal2 s 201038 0 201094 800 6 gfpga_pad_io_soc_dir[84]
port 116 nsew signal output
rlabel metal2 s 183650 0 183706 800 6 gfpga_pad_io_soc_dir[85]
port 117 nsew signal output
rlabel metal2 s 166262 0 166318 800 6 gfpga_pad_io_soc_dir[86]
port 118 nsew signal output
rlabel metal2 s 148874 0 148930 800 6 gfpga_pad_io_soc_dir[87]
port 119 nsew signal output
rlabel metal2 s 131486 0 131542 800 6 gfpga_pad_io_soc_dir[88]
port 120 nsew signal output
rlabel metal2 s 114098 0 114154 800 6 gfpga_pad_io_soc_dir[89]
port 121 nsew signal output
rlabel metal2 s 130382 542200 130438 543000 6 gfpga_pad_io_soc_dir[8]
port 122 nsew signal output
rlabel metal2 s 96710 0 96766 800 6 gfpga_pad_io_soc_dir[90]
port 123 nsew signal output
rlabel metal2 s 79322 0 79378 800 6 gfpga_pad_io_soc_dir[91]
port 124 nsew signal output
rlabel metal2 s 56138 0 56194 800 6 gfpga_pad_io_soc_dir[92]
port 125 nsew signal output
rlabel metal2 s 38750 0 38806 800 6 gfpga_pad_io_soc_dir[93]
port 126 nsew signal output
rlabel metal2 s 21362 0 21418 800 6 gfpga_pad_io_soc_dir[94]
port 127 nsew signal output
rlabel metal2 s 3974 0 4030 800 6 gfpga_pad_io_soc_dir[95]
port 128 nsew signal output
rlabel metal3 s 0 26528 800 26648 6 gfpga_pad_io_soc_dir[96]
port 129 nsew signal output
rlabel metal3 s 0 42848 800 42968 6 gfpga_pad_io_soc_dir[97]
port 130 nsew signal output
rlabel metal3 s 0 59168 800 59288 6 gfpga_pad_io_soc_dir[98]
port 131 nsew signal output
rlabel metal3 s 0 75488 800 75608 6 gfpga_pad_io_soc_dir[99]
port 132 nsew signal output
rlabel metal2 s 143630 542200 143686 543000 6 gfpga_pad_io_soc_dir[9]
port 133 nsew signal output
rlabel metal2 s 6734 542200 6790 543000 6 gfpga_pad_io_soc_in[0]
port 134 nsew signal input
rlabel metal3 s 0 80928 800 81048 6 gfpga_pad_io_soc_in[100]
port 135 nsew signal input
rlabel metal3 s 0 97248 800 97368 6 gfpga_pad_io_soc_in[101]
port 136 nsew signal input
rlabel metal3 s 0 113568 800 113688 6 gfpga_pad_io_soc_in[102]
port 137 nsew signal input
rlabel metal3 s 0 129888 800 130008 6 gfpga_pad_io_soc_in[103]
port 138 nsew signal input
rlabel metal3 s 0 146208 800 146328 6 gfpga_pad_io_soc_in[104]
port 139 nsew signal input
rlabel metal3 s 0 162528 800 162648 6 gfpga_pad_io_soc_in[105]
port 140 nsew signal input
rlabel metal3 s 0 178848 800 178968 6 gfpga_pad_io_soc_in[106]
port 141 nsew signal input
rlabel metal3 s 0 195168 800 195288 6 gfpga_pad_io_soc_in[107]
port 142 nsew signal input
rlabel metal3 s 0 211488 800 211608 6 gfpga_pad_io_soc_in[108]
port 143 nsew signal input
rlabel metal3 s 0 227808 800 227928 6 gfpga_pad_io_soc_in[109]
port 144 nsew signal input
rlabel metal2 s 148046 542200 148102 543000 6 gfpga_pad_io_soc_in[10]
port 145 nsew signal input
rlabel metal3 s 0 244128 800 244248 6 gfpga_pad_io_soc_in[110]
port 146 nsew signal input
rlabel metal3 s 0 265888 800 266008 6 gfpga_pad_io_soc_in[111]
port 147 nsew signal input
rlabel metal3 s 0 282208 800 282328 6 gfpga_pad_io_soc_in[112]
port 148 nsew signal input
rlabel metal3 s 0 298528 800 298648 6 gfpga_pad_io_soc_in[113]
port 149 nsew signal input
rlabel metal3 s 0 314848 800 314968 6 gfpga_pad_io_soc_in[114]
port 150 nsew signal input
rlabel metal3 s 0 331168 800 331288 6 gfpga_pad_io_soc_in[115]
port 151 nsew signal input
rlabel metal3 s 0 347488 800 347608 6 gfpga_pad_io_soc_in[116]
port 152 nsew signal input
rlabel metal3 s 0 363808 800 363928 6 gfpga_pad_io_soc_in[117]
port 153 nsew signal input
rlabel metal3 s 0 380128 800 380248 6 gfpga_pad_io_soc_in[118]
port 154 nsew signal input
rlabel metal3 s 0 396448 800 396568 6 gfpga_pad_io_soc_in[119]
port 155 nsew signal input
rlabel metal2 s 161294 542200 161350 543000 6 gfpga_pad_io_soc_in[11]
port 156 nsew signal input
rlabel metal3 s 0 412768 800 412888 6 gfpga_pad_io_soc_in[120]
port 157 nsew signal input
rlabel metal3 s 0 429088 800 429208 6 gfpga_pad_io_soc_in[121]
port 158 nsew signal input
rlabel metal3 s 0 445408 800 445528 6 gfpga_pad_io_soc_in[122]
port 159 nsew signal input
rlabel metal3 s 0 461728 800 461848 6 gfpga_pad_io_soc_in[123]
port 160 nsew signal input
rlabel metal3 s 0 478048 800 478168 6 gfpga_pad_io_soc_in[124]
port 161 nsew signal input
rlabel metal3 s 0 494368 800 494488 6 gfpga_pad_io_soc_in[125]
port 162 nsew signal input
rlabel metal3 s 0 510688 800 510808 6 gfpga_pad_io_soc_in[126]
port 163 nsew signal input
rlabel metal3 s 0 527008 800 527128 6 gfpga_pad_io_soc_in[127]
port 164 nsew signal input
rlabel metal2 s 174542 542200 174598 543000 6 gfpga_pad_io_soc_in[12]
port 165 nsew signal input
rlabel metal2 s 187790 542200 187846 543000 6 gfpga_pad_io_soc_in[13]
port 166 nsew signal input
rlabel metal2 s 201038 542200 201094 543000 6 gfpga_pad_io_soc_in[14]
port 167 nsew signal input
rlabel metal2 s 214286 542200 214342 543000 6 gfpga_pad_io_soc_in[15]
port 168 nsew signal input
rlabel metal2 s 227534 542200 227590 543000 6 gfpga_pad_io_soc_in[16]
port 169 nsew signal input
rlabel metal2 s 240782 542200 240838 543000 6 gfpga_pad_io_soc_in[17]
port 170 nsew signal input
rlabel metal2 s 254030 542200 254086 543000 6 gfpga_pad_io_soc_in[18]
port 171 nsew signal input
rlabel metal2 s 267278 542200 267334 543000 6 gfpga_pad_io_soc_in[19]
port 172 nsew signal input
rlabel metal2 s 19982 542200 20038 543000 6 gfpga_pad_io_soc_in[1]
port 173 nsew signal input
rlabel metal2 s 280526 542200 280582 543000 6 gfpga_pad_io_soc_in[20]
port 174 nsew signal input
rlabel metal2 s 293774 542200 293830 543000 6 gfpga_pad_io_soc_in[21]
port 175 nsew signal input
rlabel metal2 s 307022 542200 307078 543000 6 gfpga_pad_io_soc_in[22]
port 176 nsew signal input
rlabel metal2 s 320270 542200 320326 543000 6 gfpga_pad_io_soc_in[23]
port 177 nsew signal input
rlabel metal2 s 333518 542200 333574 543000 6 gfpga_pad_io_soc_in[24]
port 178 nsew signal input
rlabel metal2 s 346766 542200 346822 543000 6 gfpga_pad_io_soc_in[25]
port 179 nsew signal input
rlabel metal2 s 360014 542200 360070 543000 6 gfpga_pad_io_soc_in[26]
port 180 nsew signal input
rlabel metal2 s 373262 542200 373318 543000 6 gfpga_pad_io_soc_in[27]
port 181 nsew signal input
rlabel metal2 s 386510 542200 386566 543000 6 gfpga_pad_io_soc_in[28]
port 182 nsew signal input
rlabel metal2 s 399758 542200 399814 543000 6 gfpga_pad_io_soc_in[29]
port 183 nsew signal input
rlabel metal2 s 33230 542200 33286 543000 6 gfpga_pad_io_soc_in[2]
port 184 nsew signal input
rlabel metal2 s 413006 542200 413062 543000 6 gfpga_pad_io_soc_in[30]
port 185 nsew signal input
rlabel metal2 s 426254 542200 426310 543000 6 gfpga_pad_io_soc_in[31]
port 186 nsew signal input
rlabel metal2 s 439502 542200 439558 543000 6 gfpga_pad_io_soc_in[32]
port 187 nsew signal input
rlabel metal2 s 452750 542200 452806 543000 6 gfpga_pad_io_soc_in[33]
port 188 nsew signal input
rlabel metal2 s 465998 542200 466054 543000 6 gfpga_pad_io_soc_in[34]
port 189 nsew signal input
rlabel metal2 s 479246 542200 479302 543000 6 gfpga_pad_io_soc_in[35]
port 190 nsew signal input
rlabel metal3 s 494200 528640 495000 528760 6 gfpga_pad_io_soc_in[36]
port 191 nsew signal input
rlabel metal3 s 494200 512728 495000 512848 6 gfpga_pad_io_soc_in[37]
port 192 nsew signal input
rlabel metal3 s 494200 496816 495000 496936 6 gfpga_pad_io_soc_in[38]
port 193 nsew signal input
rlabel metal3 s 494200 480904 495000 481024 6 gfpga_pad_io_soc_in[39]
port 194 nsew signal input
rlabel metal2 s 46478 542200 46534 543000 6 gfpga_pad_io_soc_in[3]
port 195 nsew signal input
rlabel metal3 s 494200 464992 495000 465112 6 gfpga_pad_io_soc_in[40]
port 196 nsew signal input
rlabel metal3 s 494200 449080 495000 449200 6 gfpga_pad_io_soc_in[41]
port 197 nsew signal input
rlabel metal3 s 494200 433168 495000 433288 6 gfpga_pad_io_soc_in[42]
port 198 nsew signal input
rlabel metal3 s 494200 417256 495000 417376 6 gfpga_pad_io_soc_in[43]
port 199 nsew signal input
rlabel metal3 s 494200 401344 495000 401464 6 gfpga_pad_io_soc_in[44]
port 200 nsew signal input
rlabel metal3 s 494200 385432 495000 385552 6 gfpga_pad_io_soc_in[45]
port 201 nsew signal input
rlabel metal3 s 494200 369520 495000 369640 6 gfpga_pad_io_soc_in[46]
port 202 nsew signal input
rlabel metal3 s 494200 353608 495000 353728 6 gfpga_pad_io_soc_in[47]
port 203 nsew signal input
rlabel metal3 s 494200 337696 495000 337816 6 gfpga_pad_io_soc_in[48]
port 204 nsew signal input
rlabel metal3 s 494200 321784 495000 321904 6 gfpga_pad_io_soc_in[49]
port 205 nsew signal input
rlabel metal2 s 68558 542200 68614 543000 6 gfpga_pad_io_soc_in[4]
port 206 nsew signal input
rlabel metal3 s 494200 305872 495000 305992 6 gfpga_pad_io_soc_in[50]
port 207 nsew signal input
rlabel metal3 s 494200 289960 495000 290080 6 gfpga_pad_io_soc_in[51]
port 208 nsew signal input
rlabel metal3 s 494200 274048 495000 274168 6 gfpga_pad_io_soc_in[52]
port 209 nsew signal input
rlabel metal3 s 494200 258136 495000 258256 6 gfpga_pad_io_soc_in[53]
port 210 nsew signal input
rlabel metal3 s 494200 231616 495000 231736 6 gfpga_pad_io_soc_in[54]
port 211 nsew signal input
rlabel metal3 s 494200 215704 495000 215824 6 gfpga_pad_io_soc_in[55]
port 212 nsew signal input
rlabel metal3 s 494200 199792 495000 199912 6 gfpga_pad_io_soc_in[56]
port 213 nsew signal input
rlabel metal3 s 494200 183880 495000 184000 6 gfpga_pad_io_soc_in[57]
port 214 nsew signal input
rlabel metal3 s 494200 167968 495000 168088 6 gfpga_pad_io_soc_in[58]
port 215 nsew signal input
rlabel metal3 s 494200 152056 495000 152176 6 gfpga_pad_io_soc_in[59]
port 216 nsew signal input
rlabel metal2 s 81806 542200 81862 543000 6 gfpga_pad_io_soc_in[5]
port 217 nsew signal input
rlabel metal3 s 494200 136144 495000 136264 6 gfpga_pad_io_soc_in[60]
port 218 nsew signal input
rlabel metal3 s 494200 120232 495000 120352 6 gfpga_pad_io_soc_in[61]
port 219 nsew signal input
rlabel metal3 s 494200 104320 495000 104440 6 gfpga_pad_io_soc_in[62]
port 220 nsew signal input
rlabel metal3 s 494200 88408 495000 88528 6 gfpga_pad_io_soc_in[63]
port 221 nsew signal input
rlabel metal3 s 494200 72496 495000 72616 6 gfpga_pad_io_soc_in[64]
port 222 nsew signal input
rlabel metal3 s 494200 56584 495000 56704 6 gfpga_pad_io_soc_in[65]
port 223 nsew signal input
rlabel metal3 s 494200 40672 495000 40792 6 gfpga_pad_io_soc_in[66]
port 224 nsew signal input
rlabel metal3 s 494200 24760 495000 24880 6 gfpga_pad_io_soc_in[67]
port 225 nsew signal input
rlabel metal2 s 490838 0 490894 800 6 gfpga_pad_io_soc_in[68]
port 226 nsew signal input
rlabel metal2 s 473450 0 473506 800 6 gfpga_pad_io_soc_in[69]
port 227 nsew signal input
rlabel metal2 s 95054 542200 95110 543000 6 gfpga_pad_io_soc_in[6]
port 228 nsew signal input
rlabel metal2 s 456062 0 456118 800 6 gfpga_pad_io_soc_in[70]
port 229 nsew signal input
rlabel metal2 s 438674 0 438730 800 6 gfpga_pad_io_soc_in[71]
port 230 nsew signal input
rlabel metal2 s 421286 0 421342 800 6 gfpga_pad_io_soc_in[72]
port 231 nsew signal input
rlabel metal2 s 403898 0 403954 800 6 gfpga_pad_io_soc_in[73]
port 232 nsew signal input
rlabel metal2 s 386510 0 386566 800 6 gfpga_pad_io_soc_in[74]
port 233 nsew signal input
rlabel metal2 s 369122 0 369178 800 6 gfpga_pad_io_soc_in[75]
port 234 nsew signal input
rlabel metal2 s 351734 0 351790 800 6 gfpga_pad_io_soc_in[76]
port 235 nsew signal input
rlabel metal2 s 334346 0 334402 800 6 gfpga_pad_io_soc_in[77]
port 236 nsew signal input
rlabel metal2 s 316958 0 317014 800 6 gfpga_pad_io_soc_in[78]
port 237 nsew signal input
rlabel metal2 s 299570 0 299626 800 6 gfpga_pad_io_soc_in[79]
port 238 nsew signal input
rlabel metal2 s 108302 542200 108358 543000 6 gfpga_pad_io_soc_in[7]
port 239 nsew signal input
rlabel metal2 s 282182 0 282238 800 6 gfpga_pad_io_soc_in[80]
port 240 nsew signal input
rlabel metal2 s 264794 0 264850 800 6 gfpga_pad_io_soc_in[81]
port 241 nsew signal input
rlabel metal2 s 247406 0 247462 800 6 gfpga_pad_io_soc_in[82]
port 242 nsew signal input
rlabel metal2 s 230018 0 230074 800 6 gfpga_pad_io_soc_in[83]
port 243 nsew signal input
rlabel metal2 s 212630 0 212686 800 6 gfpga_pad_io_soc_in[84]
port 244 nsew signal input
rlabel metal2 s 195242 0 195298 800 6 gfpga_pad_io_soc_in[85]
port 245 nsew signal input
rlabel metal2 s 177854 0 177910 800 6 gfpga_pad_io_soc_in[86]
port 246 nsew signal input
rlabel metal2 s 160466 0 160522 800 6 gfpga_pad_io_soc_in[87]
port 247 nsew signal input
rlabel metal2 s 143078 0 143134 800 6 gfpga_pad_io_soc_in[88]
port 248 nsew signal input
rlabel metal2 s 125690 0 125746 800 6 gfpga_pad_io_soc_in[89]
port 249 nsew signal input
rlabel metal2 s 121550 542200 121606 543000 6 gfpga_pad_io_soc_in[8]
port 250 nsew signal input
rlabel metal2 s 108302 0 108358 800 6 gfpga_pad_io_soc_in[90]
port 251 nsew signal input
rlabel metal2 s 90914 0 90970 800 6 gfpga_pad_io_soc_in[91]
port 252 nsew signal input
rlabel metal2 s 67730 0 67786 800 6 gfpga_pad_io_soc_in[92]
port 253 nsew signal input
rlabel metal2 s 50342 0 50398 800 6 gfpga_pad_io_soc_in[93]
port 254 nsew signal input
rlabel metal2 s 32954 0 33010 800 6 gfpga_pad_io_soc_in[94]
port 255 nsew signal input
rlabel metal2 s 15566 0 15622 800 6 gfpga_pad_io_soc_in[95]
port 256 nsew signal input
rlabel metal3 s 0 15648 800 15768 6 gfpga_pad_io_soc_in[96]
port 257 nsew signal input
rlabel metal3 s 0 31968 800 32088 6 gfpga_pad_io_soc_in[97]
port 258 nsew signal input
rlabel metal3 s 0 48288 800 48408 6 gfpga_pad_io_soc_in[98]
port 259 nsew signal input
rlabel metal3 s 0 64608 800 64728 6 gfpga_pad_io_soc_in[99]
port 260 nsew signal input
rlabel metal2 s 134798 542200 134854 543000 6 gfpga_pad_io_soc_in[9]
port 261 nsew signal input
rlabel metal2 s 11150 542200 11206 543000 6 gfpga_pad_io_soc_out[0]
port 262 nsew signal output
rlabel metal3 s 0 86368 800 86488 6 gfpga_pad_io_soc_out[100]
port 263 nsew signal output
rlabel metal3 s 0 102688 800 102808 6 gfpga_pad_io_soc_out[101]
port 264 nsew signal output
rlabel metal3 s 0 119008 800 119128 6 gfpga_pad_io_soc_out[102]
port 265 nsew signal output
rlabel metal3 s 0 135328 800 135448 6 gfpga_pad_io_soc_out[103]
port 266 nsew signal output
rlabel metal3 s 0 151648 800 151768 6 gfpga_pad_io_soc_out[104]
port 267 nsew signal output
rlabel metal3 s 0 167968 800 168088 6 gfpga_pad_io_soc_out[105]
port 268 nsew signal output
rlabel metal3 s 0 184288 800 184408 6 gfpga_pad_io_soc_out[106]
port 269 nsew signal output
rlabel metal3 s 0 200608 800 200728 6 gfpga_pad_io_soc_out[107]
port 270 nsew signal output
rlabel metal3 s 0 216928 800 217048 6 gfpga_pad_io_soc_out[108]
port 271 nsew signal output
rlabel metal3 s 0 233248 800 233368 6 gfpga_pad_io_soc_out[109]
port 272 nsew signal output
rlabel metal2 s 152462 542200 152518 543000 6 gfpga_pad_io_soc_out[10]
port 273 nsew signal output
rlabel metal3 s 0 249568 800 249688 6 gfpga_pad_io_soc_out[110]
port 274 nsew signal output
rlabel metal3 s 0 271328 800 271448 6 gfpga_pad_io_soc_out[111]
port 275 nsew signal output
rlabel metal3 s 0 287648 800 287768 6 gfpga_pad_io_soc_out[112]
port 276 nsew signal output
rlabel metal3 s 0 303968 800 304088 6 gfpga_pad_io_soc_out[113]
port 277 nsew signal output
rlabel metal3 s 0 320288 800 320408 6 gfpga_pad_io_soc_out[114]
port 278 nsew signal output
rlabel metal3 s 0 336608 800 336728 6 gfpga_pad_io_soc_out[115]
port 279 nsew signal output
rlabel metal3 s 0 352928 800 353048 6 gfpga_pad_io_soc_out[116]
port 280 nsew signal output
rlabel metal3 s 0 369248 800 369368 6 gfpga_pad_io_soc_out[117]
port 281 nsew signal output
rlabel metal3 s 0 385568 800 385688 6 gfpga_pad_io_soc_out[118]
port 282 nsew signal output
rlabel metal3 s 0 401888 800 402008 6 gfpga_pad_io_soc_out[119]
port 283 nsew signal output
rlabel metal2 s 165710 542200 165766 543000 6 gfpga_pad_io_soc_out[11]
port 284 nsew signal output
rlabel metal3 s 0 418208 800 418328 6 gfpga_pad_io_soc_out[120]
port 285 nsew signal output
rlabel metal3 s 0 434528 800 434648 6 gfpga_pad_io_soc_out[121]
port 286 nsew signal output
rlabel metal3 s 0 450848 800 450968 6 gfpga_pad_io_soc_out[122]
port 287 nsew signal output
rlabel metal3 s 0 467168 800 467288 6 gfpga_pad_io_soc_out[123]
port 288 nsew signal output
rlabel metal3 s 0 483488 800 483608 6 gfpga_pad_io_soc_out[124]
port 289 nsew signal output
rlabel metal3 s 0 499808 800 499928 6 gfpga_pad_io_soc_out[125]
port 290 nsew signal output
rlabel metal3 s 0 516128 800 516248 6 gfpga_pad_io_soc_out[126]
port 291 nsew signal output
rlabel metal3 s 0 532448 800 532568 6 gfpga_pad_io_soc_out[127]
port 292 nsew signal output
rlabel metal2 s 178958 542200 179014 543000 6 gfpga_pad_io_soc_out[12]
port 293 nsew signal output
rlabel metal2 s 192206 542200 192262 543000 6 gfpga_pad_io_soc_out[13]
port 294 nsew signal output
rlabel metal2 s 205454 542200 205510 543000 6 gfpga_pad_io_soc_out[14]
port 295 nsew signal output
rlabel metal2 s 218702 542200 218758 543000 6 gfpga_pad_io_soc_out[15]
port 296 nsew signal output
rlabel metal2 s 231950 542200 232006 543000 6 gfpga_pad_io_soc_out[16]
port 297 nsew signal output
rlabel metal2 s 245198 542200 245254 543000 6 gfpga_pad_io_soc_out[17]
port 298 nsew signal output
rlabel metal2 s 258446 542200 258502 543000 6 gfpga_pad_io_soc_out[18]
port 299 nsew signal output
rlabel metal2 s 271694 542200 271750 543000 6 gfpga_pad_io_soc_out[19]
port 300 nsew signal output
rlabel metal2 s 24398 542200 24454 543000 6 gfpga_pad_io_soc_out[1]
port 301 nsew signal output
rlabel metal2 s 284942 542200 284998 543000 6 gfpga_pad_io_soc_out[20]
port 302 nsew signal output
rlabel metal2 s 298190 542200 298246 543000 6 gfpga_pad_io_soc_out[21]
port 303 nsew signal output
rlabel metal2 s 311438 542200 311494 543000 6 gfpga_pad_io_soc_out[22]
port 304 nsew signal output
rlabel metal2 s 324686 542200 324742 543000 6 gfpga_pad_io_soc_out[23]
port 305 nsew signal output
rlabel metal2 s 337934 542200 337990 543000 6 gfpga_pad_io_soc_out[24]
port 306 nsew signal output
rlabel metal2 s 351182 542200 351238 543000 6 gfpga_pad_io_soc_out[25]
port 307 nsew signal output
rlabel metal2 s 364430 542200 364486 543000 6 gfpga_pad_io_soc_out[26]
port 308 nsew signal output
rlabel metal2 s 377678 542200 377734 543000 6 gfpga_pad_io_soc_out[27]
port 309 nsew signal output
rlabel metal2 s 390926 542200 390982 543000 6 gfpga_pad_io_soc_out[28]
port 310 nsew signal output
rlabel metal2 s 404174 542200 404230 543000 6 gfpga_pad_io_soc_out[29]
port 311 nsew signal output
rlabel metal2 s 37646 542200 37702 543000 6 gfpga_pad_io_soc_out[2]
port 312 nsew signal output
rlabel metal2 s 417422 542200 417478 543000 6 gfpga_pad_io_soc_out[30]
port 313 nsew signal output
rlabel metal2 s 430670 542200 430726 543000 6 gfpga_pad_io_soc_out[31]
port 314 nsew signal output
rlabel metal2 s 443918 542200 443974 543000 6 gfpga_pad_io_soc_out[32]
port 315 nsew signal output
rlabel metal2 s 457166 542200 457222 543000 6 gfpga_pad_io_soc_out[33]
port 316 nsew signal output
rlabel metal2 s 470414 542200 470470 543000 6 gfpga_pad_io_soc_out[34]
port 317 nsew signal output
rlabel metal2 s 483662 542200 483718 543000 6 gfpga_pad_io_soc_out[35]
port 318 nsew signal output
rlabel metal3 s 494200 523336 495000 523456 6 gfpga_pad_io_soc_out[36]
port 319 nsew signal output
rlabel metal3 s 494200 507424 495000 507544 6 gfpga_pad_io_soc_out[37]
port 320 nsew signal output
rlabel metal3 s 494200 491512 495000 491632 6 gfpga_pad_io_soc_out[38]
port 321 nsew signal output
rlabel metal3 s 494200 475600 495000 475720 6 gfpga_pad_io_soc_out[39]
port 322 nsew signal output
rlabel metal2 s 50894 542200 50950 543000 6 gfpga_pad_io_soc_out[3]
port 323 nsew signal output
rlabel metal3 s 494200 459688 495000 459808 6 gfpga_pad_io_soc_out[40]
port 324 nsew signal output
rlabel metal3 s 494200 443776 495000 443896 6 gfpga_pad_io_soc_out[41]
port 325 nsew signal output
rlabel metal3 s 494200 427864 495000 427984 6 gfpga_pad_io_soc_out[42]
port 326 nsew signal output
rlabel metal3 s 494200 411952 495000 412072 6 gfpga_pad_io_soc_out[43]
port 327 nsew signal output
rlabel metal3 s 494200 396040 495000 396160 6 gfpga_pad_io_soc_out[44]
port 328 nsew signal output
rlabel metal3 s 494200 380128 495000 380248 6 gfpga_pad_io_soc_out[45]
port 329 nsew signal output
rlabel metal3 s 494200 364216 495000 364336 6 gfpga_pad_io_soc_out[46]
port 330 nsew signal output
rlabel metal3 s 494200 348304 495000 348424 6 gfpga_pad_io_soc_out[47]
port 331 nsew signal output
rlabel metal3 s 494200 332392 495000 332512 6 gfpga_pad_io_soc_out[48]
port 332 nsew signal output
rlabel metal3 s 494200 316480 495000 316600 6 gfpga_pad_io_soc_out[49]
port 333 nsew signal output
rlabel metal2 s 72974 542200 73030 543000 6 gfpga_pad_io_soc_out[4]
port 334 nsew signal output
rlabel metal3 s 494200 300568 495000 300688 6 gfpga_pad_io_soc_out[50]
port 335 nsew signal output
rlabel metal3 s 494200 284656 495000 284776 6 gfpga_pad_io_soc_out[51]
port 336 nsew signal output
rlabel metal3 s 494200 268744 495000 268864 6 gfpga_pad_io_soc_out[52]
port 337 nsew signal output
rlabel metal3 s 494200 252832 495000 252952 6 gfpga_pad_io_soc_out[53]
port 338 nsew signal output
rlabel metal3 s 494200 226312 495000 226432 6 gfpga_pad_io_soc_out[54]
port 339 nsew signal output
rlabel metal3 s 494200 210400 495000 210520 6 gfpga_pad_io_soc_out[55]
port 340 nsew signal output
rlabel metal3 s 494200 194488 495000 194608 6 gfpga_pad_io_soc_out[56]
port 341 nsew signal output
rlabel metal3 s 494200 178576 495000 178696 6 gfpga_pad_io_soc_out[57]
port 342 nsew signal output
rlabel metal3 s 494200 162664 495000 162784 6 gfpga_pad_io_soc_out[58]
port 343 nsew signal output
rlabel metal3 s 494200 146752 495000 146872 6 gfpga_pad_io_soc_out[59]
port 344 nsew signal output
rlabel metal2 s 86222 542200 86278 543000 6 gfpga_pad_io_soc_out[5]
port 345 nsew signal output
rlabel metal3 s 494200 130840 495000 130960 6 gfpga_pad_io_soc_out[60]
port 346 nsew signal output
rlabel metal3 s 494200 114928 495000 115048 6 gfpga_pad_io_soc_out[61]
port 347 nsew signal output
rlabel metal3 s 494200 99016 495000 99136 6 gfpga_pad_io_soc_out[62]
port 348 nsew signal output
rlabel metal3 s 494200 83104 495000 83224 6 gfpga_pad_io_soc_out[63]
port 349 nsew signal output
rlabel metal3 s 494200 67192 495000 67312 6 gfpga_pad_io_soc_out[64]
port 350 nsew signal output
rlabel metal3 s 494200 51280 495000 51400 6 gfpga_pad_io_soc_out[65]
port 351 nsew signal output
rlabel metal3 s 494200 35368 495000 35488 6 gfpga_pad_io_soc_out[66]
port 352 nsew signal output
rlabel metal3 s 494200 19456 495000 19576 6 gfpga_pad_io_soc_out[67]
port 353 nsew signal output
rlabel metal2 s 485042 0 485098 800 6 gfpga_pad_io_soc_out[68]
port 354 nsew signal output
rlabel metal2 s 467654 0 467710 800 6 gfpga_pad_io_soc_out[69]
port 355 nsew signal output
rlabel metal2 s 99470 542200 99526 543000 6 gfpga_pad_io_soc_out[6]
port 356 nsew signal output
rlabel metal2 s 450266 0 450322 800 6 gfpga_pad_io_soc_out[70]
port 357 nsew signal output
rlabel metal2 s 432878 0 432934 800 6 gfpga_pad_io_soc_out[71]
port 358 nsew signal output
rlabel metal2 s 415490 0 415546 800 6 gfpga_pad_io_soc_out[72]
port 359 nsew signal output
rlabel metal2 s 398102 0 398158 800 6 gfpga_pad_io_soc_out[73]
port 360 nsew signal output
rlabel metal2 s 380714 0 380770 800 6 gfpga_pad_io_soc_out[74]
port 361 nsew signal output
rlabel metal2 s 363326 0 363382 800 6 gfpga_pad_io_soc_out[75]
port 362 nsew signal output
rlabel metal2 s 345938 0 345994 800 6 gfpga_pad_io_soc_out[76]
port 363 nsew signal output
rlabel metal2 s 328550 0 328606 800 6 gfpga_pad_io_soc_out[77]
port 364 nsew signal output
rlabel metal2 s 311162 0 311218 800 6 gfpga_pad_io_soc_out[78]
port 365 nsew signal output
rlabel metal2 s 293774 0 293830 800 6 gfpga_pad_io_soc_out[79]
port 366 nsew signal output
rlabel metal2 s 112718 542200 112774 543000 6 gfpga_pad_io_soc_out[7]
port 367 nsew signal output
rlabel metal2 s 276386 0 276442 800 6 gfpga_pad_io_soc_out[80]
port 368 nsew signal output
rlabel metal2 s 258998 0 259054 800 6 gfpga_pad_io_soc_out[81]
port 369 nsew signal output
rlabel metal2 s 241610 0 241666 800 6 gfpga_pad_io_soc_out[82]
port 370 nsew signal output
rlabel metal2 s 224222 0 224278 800 6 gfpga_pad_io_soc_out[83]
port 371 nsew signal output
rlabel metal2 s 206834 0 206890 800 6 gfpga_pad_io_soc_out[84]
port 372 nsew signal output
rlabel metal2 s 189446 0 189502 800 6 gfpga_pad_io_soc_out[85]
port 373 nsew signal output
rlabel metal2 s 172058 0 172114 800 6 gfpga_pad_io_soc_out[86]
port 374 nsew signal output
rlabel metal2 s 154670 0 154726 800 6 gfpga_pad_io_soc_out[87]
port 375 nsew signal output
rlabel metal2 s 137282 0 137338 800 6 gfpga_pad_io_soc_out[88]
port 376 nsew signal output
rlabel metal2 s 119894 0 119950 800 6 gfpga_pad_io_soc_out[89]
port 377 nsew signal output
rlabel metal2 s 125966 542200 126022 543000 6 gfpga_pad_io_soc_out[8]
port 378 nsew signal output
rlabel metal2 s 102506 0 102562 800 6 gfpga_pad_io_soc_out[90]
port 379 nsew signal output
rlabel metal2 s 85118 0 85174 800 6 gfpga_pad_io_soc_out[91]
port 380 nsew signal output
rlabel metal2 s 61934 0 61990 800 6 gfpga_pad_io_soc_out[92]
port 381 nsew signal output
rlabel metal2 s 44546 0 44602 800 6 gfpga_pad_io_soc_out[93]
port 382 nsew signal output
rlabel metal2 s 27158 0 27214 800 6 gfpga_pad_io_soc_out[94]
port 383 nsew signal output
rlabel metal2 s 9770 0 9826 800 6 gfpga_pad_io_soc_out[95]
port 384 nsew signal output
rlabel metal3 s 0 21088 800 21208 6 gfpga_pad_io_soc_out[96]
port 385 nsew signal output
rlabel metal3 s 0 37408 800 37528 6 gfpga_pad_io_soc_out[97]
port 386 nsew signal output
rlabel metal3 s 0 53728 800 53848 6 gfpga_pad_io_soc_out[98]
port 387 nsew signal output
rlabel metal3 s 0 70048 800 70168 6 gfpga_pad_io_soc_out[99]
port 388 nsew signal output
rlabel metal2 s 139214 542200 139270 543000 6 gfpga_pad_io_soc_out[9]
port 389 nsew signal output
rlabel metal3 s 494200 8848 495000 8968 6 isol_n
port 390 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 prog_clk
port 391 nsew signal input
rlabel metal3 s 0 260448 800 260568 6 prog_reset
port 392 nsew signal input
rlabel metal3 s 494200 236920 495000 237040 6 reset
port 393 nsew signal input
rlabel metal2 s 64142 542200 64198 543000 6 sc_head
port 394 nsew signal input
rlabel metal3 s 494200 533944 495000 534064 6 sc_tail
port 395 nsew signal output
rlabel metal3 s 494200 242224 495000 242344 6 test_enable
port 396 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 495000 543000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 77498306
string GDS_FILE /home/hosni/OpenFPGA/clear/openlane/fpga_core/runs/23_03_29_04_36/results/signoff/fpga_core.magic.gds
string GDS_START 41579182
<< end >>

