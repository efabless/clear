magic
tech sky130A
magscale 1 2
timestamp 1679357618
<< viali >>
rect 35909 24361 35943 24395
rect 39221 24361 39255 24395
rect 40049 24361 40083 24395
rect 40693 24361 40727 24395
rect 48329 24361 48363 24395
rect 17049 24293 17083 24327
rect 24593 24293 24627 24327
rect 32965 24293 32999 24327
rect 3249 24225 3283 24259
rect 5825 24225 5859 24259
rect 8217 24225 8251 24259
rect 10977 24225 11011 24259
rect 13553 24225 13587 24259
rect 16129 24225 16163 24259
rect 18705 24225 18739 24259
rect 20913 24225 20947 24259
rect 22477 24225 22511 24259
rect 25053 24225 25087 24259
rect 25145 24225 25179 24259
rect 26341 24225 26375 24259
rect 34069 24225 34103 24259
rect 34253 24225 34287 24259
rect 36553 24225 36587 24259
rect 37933 24225 37967 24259
rect 38117 24225 38151 24259
rect 48053 24225 48087 24259
rect 48513 24225 48547 24259
rect 2237 24157 2271 24191
rect 4169 24157 4203 24191
rect 4813 24157 4847 24191
rect 6745 24157 6779 24191
rect 7389 24157 7423 24191
rect 9321 24157 9355 24191
rect 9965 24157 9999 24191
rect 11897 24157 11931 24191
rect 12541 24157 12575 24191
rect 14473 24157 14507 24191
rect 15117 24157 15151 24191
rect 17601 24157 17635 24191
rect 19625 24157 19659 24191
rect 20085 24157 20119 24191
rect 22201 24157 22235 24191
rect 24041 24157 24075 24191
rect 26157 24157 26191 24191
rect 28089 24157 28123 24191
rect 28733 24157 28767 24191
rect 29929 24157 29963 24191
rect 30573 24157 30607 24191
rect 31217 24157 31251 24191
rect 32505 24157 32539 24191
rect 33149 24157 33183 24191
rect 35081 24157 35115 24191
rect 36369 24157 36403 24191
rect 40233 24157 40267 24191
rect 40877 24157 40911 24191
rect 41337 24157 41371 24191
rect 41705 24157 41739 24191
rect 42625 24157 42659 24191
rect 45293 24157 45327 24191
rect 45937 24157 45971 24191
rect 46765 24157 46799 24191
rect 48145 24157 48179 24191
rect 48789 24157 48823 24191
rect 24961 24089 24995 24123
rect 25789 24089 25823 24123
rect 27261 24089 27295 24123
rect 36277 24089 36311 24123
rect 45477 24089 45511 24123
rect 46949 24089 46983 24123
rect 3985 24021 4019 24055
rect 6561 24021 6595 24055
rect 9137 24021 9171 24055
rect 14289 24021 14323 24055
rect 19441 24021 19475 24055
rect 23857 24021 23891 24055
rect 27353 24021 27387 24055
rect 27905 24021 27939 24055
rect 28549 24021 28583 24055
rect 29745 24021 29779 24055
rect 30389 24021 30423 24055
rect 31033 24021 31067 24055
rect 32321 24021 32355 24055
rect 33609 24021 33643 24055
rect 33977 24021 34011 24055
rect 34897 24021 34931 24055
rect 37473 24021 37507 24055
rect 37841 24021 37875 24055
rect 41521 24021 41555 24055
rect 43913 24021 43947 24055
rect 46121 24021 46155 24055
rect 6561 23817 6595 23851
rect 23949 23817 23983 23851
rect 27905 23817 27939 23851
rect 32321 23817 32355 23851
rect 36093 23817 36127 23851
rect 39129 23817 39163 23851
rect 39865 23817 39899 23851
rect 44327 23817 44361 23851
rect 48973 23817 49007 23851
rect 3985 23749 4019 23783
rect 9137 23749 9171 23783
rect 10701 23749 10735 23783
rect 14381 23749 14415 23783
rect 16129 23749 16163 23783
rect 18153 23749 18187 23783
rect 19073 23749 19107 23783
rect 23857 23749 23891 23783
rect 32781 23749 32815 23783
rect 39037 23749 39071 23783
rect 46857 23749 46891 23783
rect 48145 23749 48179 23783
rect 2973 23681 3007 23715
rect 4629 23681 4663 23715
rect 6745 23681 6779 23715
rect 7481 23681 7515 23715
rect 8125 23681 8159 23715
rect 9965 23681 9999 23715
rect 11805 23681 11839 23715
rect 13461 23681 13495 23715
rect 15117 23681 15151 23715
rect 17141 23681 17175 23715
rect 18797 23681 18831 23715
rect 21465 23681 21499 23715
rect 22937 23681 22971 23715
rect 27261 23681 27295 23715
rect 27445 23681 27479 23715
rect 28089 23681 28123 23715
rect 28733 23681 28767 23715
rect 29377 23681 29411 23715
rect 32689 23681 32723 23715
rect 36461 23681 36495 23715
rect 37841 23681 37875 23715
rect 37933 23681 37967 23715
rect 45201 23681 45235 23715
rect 45477 23681 45511 23715
rect 48789 23681 48823 23715
rect 5457 23613 5491 23647
rect 12081 23613 12115 23647
rect 23029 23613 23063 23647
rect 23213 23613 23247 23647
rect 24869 23613 24903 23647
rect 25145 23613 25179 23647
rect 30021 23613 30055 23647
rect 30297 23613 30331 23647
rect 32965 23613 32999 23647
rect 33609 23613 33643 23647
rect 33885 23613 33919 23647
rect 36553 23613 36587 23647
rect 36737 23613 36771 23647
rect 38117 23613 38151 23647
rect 39221 23613 39255 23647
rect 39957 23613 39991 23647
rect 40049 23613 40083 23647
rect 41061 23613 41095 23647
rect 41337 23613 41371 23647
rect 43545 23613 43579 23647
rect 44097 23613 44131 23647
rect 13185 23545 13219 23579
rect 22569 23545 22603 23579
rect 38669 23545 38703 23579
rect 47041 23545 47075 23579
rect 7297 23477 7331 23511
rect 20545 23477 20579 23511
rect 21281 23477 21315 23511
rect 26617 23477 26651 23511
rect 28549 23477 28583 23511
rect 29193 23477 29227 23511
rect 31769 23477 31803 23511
rect 35357 23477 35391 23511
rect 37473 23477 37507 23511
rect 39497 23477 39531 23511
rect 42993 23477 43027 23511
rect 48237 23477 48271 23511
rect 19809 23273 19843 23307
rect 22661 23273 22695 23307
rect 27905 23273 27939 23307
rect 29745 23273 29779 23307
rect 33149 23273 33183 23307
rect 39037 23273 39071 23307
rect 40049 23273 40083 23307
rect 9873 23205 9907 23239
rect 24869 23205 24903 23239
rect 33701 23205 33735 23239
rect 47041 23205 47075 23239
rect 6101 23137 6135 23171
rect 7849 23137 7883 23171
rect 11253 23137 11287 23171
rect 13369 23137 13403 23171
rect 15761 23137 15795 23171
rect 20361 23137 20395 23171
rect 23765 23137 23799 23171
rect 23949 23137 23983 23171
rect 25973 23137 26007 23171
rect 28457 23137 28491 23171
rect 30205 23137 30239 23171
rect 30389 23137 30423 23171
rect 31677 23137 31711 23171
rect 35081 23137 35115 23171
rect 40601 23137 40635 23171
rect 41889 23137 41923 23171
rect 1777 23069 1811 23103
rect 4261 23069 4295 23103
rect 4913 23069 4947 23103
rect 5365 23069 5399 23103
rect 7389 23069 7423 23103
rect 9229 23069 9263 23103
rect 10057 23069 10091 23103
rect 10701 23069 10735 23103
rect 12541 23069 12575 23103
rect 14841 23069 14875 23103
rect 15485 23069 15519 23103
rect 17141 23069 17175 23103
rect 22845 23069 22879 23103
rect 25697 23069 25731 23103
rect 28273 23069 28307 23103
rect 31401 23069 31435 23103
rect 33885 23069 33919 23103
rect 37289 23069 37323 23103
rect 41613 23069 41647 23103
rect 43729 23069 43763 23103
rect 44005 23069 44039 23103
rect 45109 23069 45143 23103
rect 45569 23069 45603 23103
rect 46305 23069 46339 23103
rect 47225 23069 47259 23103
rect 47869 23069 47903 23103
rect 48329 23069 48363 23103
rect 49065 23069 49099 23103
rect 2789 23001 2823 23035
rect 17417 23001 17451 23035
rect 19717 23001 19751 23035
rect 20637 23001 20671 23035
rect 24685 23001 24719 23035
rect 35357 23001 35391 23035
rect 37565 23001 37599 23035
rect 40417 23001 40451 23035
rect 43637 23001 43671 23035
rect 4077 22933 4111 22967
rect 4721 22933 4755 22967
rect 9321 22933 9355 22967
rect 14657 22933 14691 22967
rect 18889 22933 18923 22967
rect 22109 22933 22143 22967
rect 23305 22933 23339 22967
rect 23673 22933 23707 22967
rect 27445 22933 27479 22967
rect 28365 22933 28399 22967
rect 30113 22933 30147 22967
rect 36829 22933 36863 22967
rect 40509 22933 40543 22967
rect 45201 22933 45235 22967
rect 45385 22933 45419 22967
rect 46121 22933 46155 22967
rect 47685 22933 47719 22967
rect 48513 22933 48547 22967
rect 49249 22933 49283 22967
rect 21189 22729 21223 22763
rect 30665 22729 30699 22763
rect 35909 22729 35943 22763
rect 39221 22729 39255 22763
rect 39681 22729 39715 22763
rect 40141 22729 40175 22763
rect 40877 22729 40911 22763
rect 47041 22729 47075 22763
rect 48513 22729 48547 22763
rect 2789 22661 2823 22695
rect 3985 22661 4019 22695
rect 19717 22661 19751 22695
rect 22293 22661 22327 22695
rect 25145 22661 25179 22695
rect 32689 22661 32723 22695
rect 1777 22593 1811 22627
rect 4813 22593 4847 22627
rect 6837 22593 6871 22627
rect 7481 22593 7515 22627
rect 9965 22593 9999 22627
rect 12173 22593 12207 22627
rect 12817 22593 12851 22627
rect 15117 22593 15151 22627
rect 16865 22593 16899 22627
rect 24869 22593 24903 22627
rect 27353 22593 27387 22627
rect 28089 22593 28123 22627
rect 31677 22593 31711 22627
rect 32781 22593 32815 22627
rect 33149 22593 33183 22627
rect 35449 22593 35483 22627
rect 36277 22593 36311 22627
rect 40049 22593 40083 22627
rect 41521 22593 41555 22627
rect 41797 22593 41831 22627
rect 42809 22593 42843 22627
rect 43269 22593 43303 22627
rect 44557 22593 44591 22627
rect 44925 22593 44959 22627
rect 47225 22593 47259 22627
rect 48329 22593 48363 22627
rect 49065 22593 49099 22627
rect 5089 22525 5123 22559
rect 7941 22525 7975 22559
rect 10241 22525 10275 22559
rect 13093 22525 13127 22559
rect 15393 22525 15427 22559
rect 17141 22525 17175 22559
rect 19441 22525 19475 22559
rect 22017 22525 22051 22559
rect 28365 22525 28399 22559
rect 30757 22525 30791 22559
rect 30849 22525 30883 22559
rect 32873 22525 32907 22559
rect 33425 22525 33459 22559
rect 34897 22525 34931 22559
rect 36369 22525 36403 22559
rect 36461 22525 36495 22559
rect 37473 22525 37507 22559
rect 37749 22525 37783 22559
rect 40233 22525 40267 22559
rect 40969 22525 41003 22559
rect 41061 22525 41095 22559
rect 43545 22525 43579 22559
rect 11989 22457 12023 22491
rect 27169 22457 27203 22491
rect 32321 22457 32355 22491
rect 40509 22457 40543 22491
rect 49249 22457 49283 22491
rect 4077 22389 4111 22423
rect 6653 22389 6687 22423
rect 18613 22389 18647 22423
rect 23765 22389 23799 22423
rect 26617 22389 26651 22423
rect 29837 22389 29871 22423
rect 30297 22389 30331 22423
rect 31493 22389 31527 22423
rect 41337 22389 41371 22423
rect 41613 22389 41647 22423
rect 42625 22389 42659 22423
rect 44741 22389 44775 22423
rect 7849 22185 7883 22219
rect 16957 22185 16991 22219
rect 28273 22185 28307 22219
rect 29745 22185 29779 22219
rect 41245 22185 41279 22219
rect 47777 22185 47811 22219
rect 2053 22049 2087 22083
rect 4445 22049 4479 22083
rect 6285 22049 6319 22083
rect 9597 22049 9631 22083
rect 11345 22049 11379 22083
rect 11805 22049 11839 22083
rect 17969 22049 18003 22083
rect 19901 22049 19935 22083
rect 22017 22049 22051 22083
rect 23213 22049 23247 22083
rect 25237 22049 25271 22083
rect 26433 22049 26467 22083
rect 26525 22049 26559 22083
rect 27629 22049 27663 22083
rect 28825 22049 28859 22083
rect 30849 22049 30883 22083
rect 32597 22049 32631 22083
rect 33701 22049 33735 22083
rect 35909 22049 35943 22083
rect 37565 22049 37599 22083
rect 40601 22049 40635 22083
rect 41797 22049 41831 22083
rect 1777 21981 1811 22015
rect 4077 21981 4111 22015
rect 6009 21981 6043 22015
rect 7757 21981 7791 22015
rect 8585 21981 8619 22015
rect 9137 21981 9171 22015
rect 12081 21981 12115 22015
rect 13369 21981 13403 22015
rect 15209 21981 15243 22015
rect 17601 21981 17635 22015
rect 19625 21981 19659 22015
rect 21833 21981 21867 22015
rect 27445 21981 27479 22015
rect 29929 21981 29963 22015
rect 36737 21981 36771 22015
rect 37289 21981 37323 22015
rect 40509 21981 40543 22015
rect 43453 21981 43487 22015
rect 47961 21981 47995 22015
rect 48605 21981 48639 22015
rect 11529 21913 11563 21947
rect 13185 21913 13219 21947
rect 14565 21913 14599 21947
rect 15485 21913 15519 21947
rect 21925 21913 21959 21947
rect 25053 21913 25087 21947
rect 28733 21913 28767 21947
rect 31125 21913 31159 21947
rect 33517 21913 33551 21947
rect 35725 21913 35759 21947
rect 41613 21913 41647 21947
rect 49157 21913 49191 21947
rect 8401 21845 8435 21879
rect 11621 21845 11655 21879
rect 14657 21845 14691 21879
rect 21465 21845 21499 21879
rect 22661 21845 22695 21879
rect 23029 21845 23063 21879
rect 23121 21845 23155 21879
rect 24593 21845 24627 21879
rect 24961 21845 24995 21879
rect 25881 21845 25915 21879
rect 25973 21845 26007 21879
rect 26341 21845 26375 21879
rect 27077 21845 27111 21879
rect 27537 21845 27571 21879
rect 28641 21845 28675 21879
rect 33057 21845 33091 21879
rect 33425 21845 33459 21879
rect 35357 21845 35391 21879
rect 35817 21845 35851 21879
rect 36553 21845 36587 21879
rect 39037 21845 39071 21879
rect 40049 21845 40083 21879
rect 40417 21845 40451 21879
rect 41705 21845 41739 21879
rect 43269 21845 43303 21879
rect 48421 21845 48455 21879
rect 49249 21845 49283 21879
rect 10333 21641 10367 21675
rect 10977 21641 11011 21675
rect 17417 21641 17451 21675
rect 17877 21641 17911 21675
rect 21005 21641 21039 21675
rect 24777 21641 24811 21675
rect 26433 21641 26467 21675
rect 27629 21641 27663 21675
rect 28365 21641 28399 21675
rect 34897 21641 34931 21675
rect 40233 21641 40267 21675
rect 12265 21573 12299 21607
rect 14841 21573 14875 21607
rect 18889 21573 18923 21607
rect 25237 21573 25271 21607
rect 27537 21573 27571 21607
rect 30021 21573 30055 21607
rect 36093 21573 36127 21607
rect 1777 21505 1811 21539
rect 3617 21505 3651 21539
rect 5917 21505 5951 21539
rect 6561 21505 6595 21539
rect 8401 21505 8435 21539
rect 10517 21505 10551 21539
rect 11161 21505 11195 21539
rect 13369 21505 13403 21539
rect 17785 21505 17819 21539
rect 20913 21505 20947 21539
rect 25145 21505 25179 21539
rect 26617 21505 26651 21539
rect 28733 21505 28767 21539
rect 29929 21505 29963 21539
rect 31125 21505 31159 21539
rect 32689 21505 32723 21539
rect 37473 21505 37507 21539
rect 40601 21505 40635 21539
rect 49065 21505 49099 21539
rect 2789 21437 2823 21471
rect 4169 21437 4203 21471
rect 7021 21437 7055 21471
rect 8861 21437 8895 21471
rect 13461 21437 13495 21471
rect 13645 21437 13679 21471
rect 14565 21437 14599 21471
rect 18061 21437 18095 21471
rect 18613 21437 18647 21471
rect 22477 21437 22511 21471
rect 22753 21437 22787 21471
rect 24225 21437 24259 21471
rect 25421 21437 25455 21471
rect 27721 21437 27755 21471
rect 28825 21437 28859 21471
rect 28917 21437 28951 21471
rect 30113 21437 30147 21471
rect 31217 21437 31251 21471
rect 31401 21437 31435 21471
rect 33149 21437 33183 21471
rect 33425 21437 33459 21471
rect 36185 21437 36219 21471
rect 36369 21437 36403 21471
rect 37749 21437 37783 21471
rect 40693 21437 40727 21471
rect 40785 21437 40819 21471
rect 5733 21369 5767 21403
rect 13001 21369 13035 21403
rect 27169 21369 27203 21403
rect 12357 21301 12391 21335
rect 16313 21301 16347 21335
rect 20361 21301 20395 21335
rect 29561 21301 29595 21335
rect 30757 21301 30791 21335
rect 35725 21301 35759 21335
rect 39221 21301 39255 21335
rect 39681 21301 39715 21335
rect 49249 21301 49283 21335
rect 9873 21097 9907 21131
rect 12909 21097 12943 21131
rect 13645 21097 13679 21131
rect 18889 21097 18923 21131
rect 21360 21097 21394 21131
rect 27905 21097 27939 21131
rect 28365 21097 28399 21131
rect 30849 21097 30883 21131
rect 33241 21097 33275 21131
rect 37289 21097 37323 21131
rect 40049 21097 40083 21131
rect 49249 21097 49283 21131
rect 7849 21029 7883 21063
rect 12081 21029 12115 21063
rect 19809 21029 19843 21063
rect 22845 21029 22879 21063
rect 29745 21029 29779 21063
rect 4445 20961 4479 20995
rect 6745 20961 6779 20995
rect 10517 20961 10551 20995
rect 17141 20961 17175 20995
rect 17417 20961 17451 20995
rect 20453 20961 20487 20995
rect 23857 20961 23891 20995
rect 25237 20961 25271 20995
rect 26433 20961 26467 20995
rect 28917 20961 28951 20995
rect 31309 20961 31343 20995
rect 31493 20961 31527 20995
rect 33793 20961 33827 20995
rect 34897 20961 34931 20995
rect 35173 20961 35207 20995
rect 36645 20961 36679 20995
rect 37749 20961 37783 20995
rect 38025 20961 38059 20995
rect 40509 20961 40543 20995
rect 40601 20961 40635 20995
rect 41797 20961 41831 20995
rect 1777 20893 1811 20927
rect 4077 20893 4111 20927
rect 6009 20893 6043 20927
rect 8033 20893 8067 20927
rect 11161 20893 11195 20927
rect 12817 20893 12851 20927
rect 14289 20893 14323 20927
rect 16681 20893 16715 20927
rect 20177 20893 20211 20927
rect 21097 20893 21131 20927
rect 23673 20893 23707 20927
rect 25053 20893 25087 20927
rect 27261 20893 27295 20927
rect 29929 20893 29963 20927
rect 32229 20893 32263 20927
rect 33609 20893 33643 20927
rect 41705 20893 41739 20927
rect 49065 20893 49099 20927
rect 2789 20825 2823 20859
rect 11897 20825 11931 20859
rect 13553 20825 13587 20859
rect 14565 20825 14599 20859
rect 23765 20825 23799 20859
rect 28825 20825 28859 20859
rect 41613 20825 41647 20859
rect 10977 20757 11011 20791
rect 16037 20757 16071 20791
rect 16497 20757 16531 20791
rect 20269 20757 20303 20791
rect 23305 20757 23339 20791
rect 24593 20757 24627 20791
rect 24961 20757 24995 20791
rect 25881 20757 25915 20791
rect 26249 20757 26283 20791
rect 26341 20757 26375 20791
rect 27077 20757 27111 20791
rect 28733 20757 28767 20791
rect 31217 20757 31251 20791
rect 32045 20757 32079 20791
rect 33701 20757 33735 20791
rect 39497 20757 39531 20791
rect 40417 20757 40451 20791
rect 41245 20757 41279 20791
rect 5273 20553 5307 20587
rect 8401 20553 8435 20587
rect 9965 20553 9999 20587
rect 10609 20553 10643 20587
rect 14105 20553 14139 20587
rect 16221 20553 16255 20587
rect 21465 20553 21499 20587
rect 29009 20553 29043 20587
rect 29837 20553 29871 20587
rect 31033 20553 31067 20587
rect 31125 20553 31159 20587
rect 34069 20553 34103 20587
rect 34529 20553 34563 20587
rect 40417 20553 40451 20587
rect 12725 20485 12759 20519
rect 15577 20485 15611 20519
rect 22477 20485 22511 20519
rect 27537 20485 27571 20519
rect 32597 20485 32631 20519
rect 38025 20485 38059 20519
rect 1777 20417 1811 20451
rect 3617 20417 3651 20451
rect 5457 20417 5491 20451
rect 6561 20417 6595 20451
rect 8585 20417 8619 20451
rect 9321 20417 9355 20451
rect 10149 20417 10183 20451
rect 10793 20417 10827 20451
rect 11805 20417 11839 20451
rect 12541 20417 12575 20451
rect 14197 20417 14231 20451
rect 15393 20417 15427 20451
rect 16129 20417 16163 20451
rect 17049 20417 17083 20451
rect 26249 20417 26283 20451
rect 34897 20417 34931 20451
rect 36461 20417 36495 20451
rect 36553 20417 36587 20451
rect 37749 20417 37783 20451
rect 40325 20417 40359 20451
rect 48605 20417 48639 20451
rect 49065 20417 49099 20451
rect 2789 20349 2823 20383
rect 3893 20349 3927 20383
rect 7021 20349 7055 20383
rect 14381 20349 14415 20383
rect 17325 20349 17359 20383
rect 19717 20349 19751 20383
rect 19993 20349 20027 20383
rect 22569 20349 22603 20383
rect 22661 20349 22695 20383
rect 23857 20349 23891 20383
rect 24133 20349 24167 20383
rect 27261 20349 27295 20383
rect 29929 20349 29963 20383
rect 30113 20349 30147 20383
rect 31217 20349 31251 20383
rect 32321 20349 32355 20383
rect 34989 20349 35023 20383
rect 35173 20349 35207 20383
rect 36737 20349 36771 20383
rect 40509 20349 40543 20383
rect 9137 20281 9171 20315
rect 13737 20281 13771 20315
rect 26065 20281 26099 20315
rect 36093 20281 36127 20315
rect 39497 20281 39531 20315
rect 49249 20281 49283 20315
rect 11897 20213 11931 20247
rect 18797 20213 18831 20247
rect 22109 20213 22143 20247
rect 25605 20213 25639 20247
rect 29469 20213 29503 20247
rect 30665 20213 30699 20247
rect 39957 20213 39991 20247
rect 48421 20213 48455 20247
rect 14749 20009 14783 20043
rect 16957 20009 16991 20043
rect 30389 20009 30423 20043
rect 33425 20009 33459 20043
rect 34897 20009 34931 20043
rect 40049 20009 40083 20043
rect 11529 19941 11563 19975
rect 16865 19941 16899 19975
rect 22293 19941 22327 19975
rect 24777 19941 24811 19975
rect 28089 19941 28123 19975
rect 31585 19941 31619 19975
rect 4905 19873 4939 19907
rect 6285 19873 6319 19907
rect 10793 19873 10827 19907
rect 17509 19873 17543 19907
rect 18613 19873 18647 19907
rect 18797 19873 18831 19907
rect 20821 19873 20855 19907
rect 23397 19873 23431 19907
rect 26157 19873 26191 19907
rect 26985 19873 27019 19907
rect 27905 19873 27939 19907
rect 28549 19873 28583 19907
rect 28641 19873 28675 19907
rect 31033 19873 31067 19907
rect 32137 19873 32171 19907
rect 33977 19873 34011 19907
rect 35357 19873 35391 19907
rect 35449 19873 35483 19907
rect 36737 19873 36771 19907
rect 38301 19873 38335 19907
rect 38485 19873 38519 19907
rect 40509 19873 40543 19907
rect 40601 19873 40635 19907
rect 41705 19873 41739 19907
rect 41797 19873 41831 19907
rect 49341 19873 49375 19907
rect 1777 19805 1811 19839
rect 4077 19805 4111 19839
rect 6009 19805 6043 19839
rect 7941 19805 7975 19839
rect 10057 19805 10091 19839
rect 11069 19805 11103 19839
rect 11345 19805 11379 19839
rect 11989 19805 12023 19839
rect 14933 19805 14967 19839
rect 15577 19805 15611 19839
rect 16497 19805 16531 19839
rect 19901 19805 19935 19839
rect 20545 19805 20579 19839
rect 26065 19805 26099 19839
rect 29929 19805 29963 19839
rect 31953 19805 31987 19839
rect 33793 19805 33827 19839
rect 33885 19805 33919 19839
rect 38209 19805 38243 19839
rect 39221 19805 39255 19839
rect 2789 19737 2823 19771
rect 12265 19737 12299 19771
rect 16681 19737 16715 19771
rect 17325 19737 17359 19771
rect 19717 19737 19751 19771
rect 25973 19737 26007 19771
rect 26801 19737 26835 19771
rect 27629 19737 27663 19771
rect 28457 19737 28491 19771
rect 35265 19737 35299 19771
rect 36461 19737 36495 19771
rect 40417 19737 40451 19771
rect 41613 19737 41647 19771
rect 49157 19737 49191 19771
rect 7757 19669 7791 19703
rect 9873 19669 9907 19703
rect 13737 19669 13771 19703
rect 17417 19669 17451 19703
rect 18153 19669 18187 19703
rect 18521 19669 18555 19703
rect 22753 19669 22787 19703
rect 23121 19669 23155 19703
rect 23213 19669 23247 19703
rect 25605 19669 25639 19703
rect 26433 19669 26467 19703
rect 26893 19669 26927 19703
rect 27261 19669 27295 19703
rect 27721 19669 27755 19703
rect 30757 19669 30791 19703
rect 30849 19669 30883 19703
rect 32045 19669 32079 19703
rect 36093 19669 36127 19703
rect 36553 19669 36587 19703
rect 37841 19669 37875 19703
rect 41245 19669 41279 19703
rect 10977 19465 11011 19499
rect 14473 19465 14507 19499
rect 15393 19465 15427 19499
rect 16865 19465 16899 19499
rect 17325 19465 17359 19499
rect 20729 19465 20763 19499
rect 21189 19465 21223 19499
rect 25145 19465 25179 19499
rect 28457 19465 28491 19499
rect 28825 19465 28859 19499
rect 29653 19465 29687 19499
rect 30113 19465 30147 19499
rect 32321 19465 32355 19499
rect 32689 19465 32723 19499
rect 32781 19465 32815 19499
rect 33517 19465 33551 19499
rect 33885 19465 33919 19499
rect 34713 19465 34747 19499
rect 40509 19465 40543 19499
rect 40601 19465 40635 19499
rect 4353 19397 4387 19431
rect 26157 19397 26191 19431
rect 27905 19397 27939 19431
rect 28917 19397 28951 19431
rect 31585 19397 31619 19431
rect 36277 19397 36311 19431
rect 1777 19329 1811 19363
rect 2789 19329 2823 19363
rect 3617 19329 3651 19363
rect 5365 19329 5399 19363
rect 11161 19329 11195 19363
rect 12081 19329 12115 19363
rect 12714 19329 12748 19363
rect 15577 19329 15611 19363
rect 16129 19329 16163 19363
rect 17233 19329 17267 19363
rect 18061 19329 18095 19363
rect 20085 19329 20119 19363
rect 21097 19329 21131 19363
rect 22017 19329 22051 19363
rect 22845 19329 22879 19363
rect 23397 19329 23431 19363
rect 30021 19329 30055 19363
rect 30849 19329 30883 19363
rect 35081 19329 35115 19363
rect 35173 19329 35207 19363
rect 36369 19329 36403 19363
rect 37933 19329 37967 19363
rect 49157 19329 49191 19363
rect 13001 19261 13035 19295
rect 17509 19261 17543 19295
rect 18337 19261 18371 19295
rect 21281 19261 21315 19295
rect 23673 19261 23707 19295
rect 26249 19261 26283 19295
rect 26433 19261 26467 19295
rect 29009 19261 29043 19295
rect 30297 19261 30331 19295
rect 32873 19261 32907 19295
rect 33977 19261 34011 19295
rect 34161 19261 34195 19295
rect 35357 19261 35391 19295
rect 36553 19261 36587 19295
rect 40693 19261 40727 19295
rect 35909 19193 35943 19227
rect 5457 19125 5491 19159
rect 9873 19125 9907 19159
rect 10517 19125 10551 19159
rect 12173 19125 12207 19159
rect 16221 19125 16255 19159
rect 25789 19125 25823 19159
rect 38196 19125 38230 19159
rect 39681 19125 39715 19159
rect 40141 19125 40175 19159
rect 49249 19125 49283 19159
rect 10885 18921 10919 18955
rect 11897 18921 11931 18955
rect 16037 18921 16071 18955
rect 16773 18921 16807 18955
rect 17969 18921 18003 18955
rect 19809 18921 19843 18955
rect 24593 18921 24627 18955
rect 29009 18921 29043 18955
rect 31493 18921 31527 18955
rect 32689 18921 32723 18955
rect 37013 18921 37047 18955
rect 41797 18921 41831 18955
rect 12541 18853 12575 18887
rect 27537 18853 27571 18887
rect 38025 18853 38059 18887
rect 4445 18785 4479 18819
rect 9137 18785 9171 18819
rect 9413 18785 9447 18819
rect 13001 18785 13035 18819
rect 13185 18785 13219 18819
rect 14289 18785 14323 18819
rect 14565 18785 14599 18819
rect 17233 18785 17267 18819
rect 17325 18785 17359 18819
rect 18613 18785 18647 18819
rect 20453 18785 20487 18819
rect 21557 18785 21591 18819
rect 21649 18785 21683 18819
rect 22569 18785 22603 18819
rect 25053 18785 25087 18819
rect 25237 18785 25271 18819
rect 25789 18785 25823 18819
rect 30205 18785 30239 18819
rect 30297 18785 30331 18819
rect 31953 18785 31987 18819
rect 32137 18785 32171 18819
rect 33149 18785 33183 18819
rect 33333 18785 33367 18819
rect 35265 18785 35299 18819
rect 38577 18785 38611 18819
rect 1777 18717 1811 18751
rect 4077 18717 4111 18751
rect 8217 18717 8251 18751
rect 12081 18717 12115 18751
rect 17141 18717 17175 18751
rect 20177 18717 20211 18751
rect 22293 18717 22327 18751
rect 29193 18717 29227 18751
rect 37473 18717 37507 18751
rect 38485 18717 38519 18751
rect 40049 18717 40083 18751
rect 48605 18717 48639 18751
rect 49065 18717 49099 18751
rect 2789 18649 2823 18683
rect 12909 18649 12943 18683
rect 26065 18649 26099 18683
rect 30113 18649 30147 18683
rect 35541 18649 35575 18683
rect 40325 18649 40359 18683
rect 8309 18581 8343 18615
rect 18337 18581 18371 18615
rect 18429 18581 18463 18615
rect 20269 18581 20303 18615
rect 21097 18581 21131 18615
rect 21465 18581 21499 18615
rect 24041 18581 24075 18615
rect 24961 18581 24995 18615
rect 29745 18581 29779 18615
rect 31861 18581 31895 18615
rect 33057 18581 33091 18615
rect 38393 18581 38427 18615
rect 48421 18581 48455 18615
rect 49249 18581 49283 18615
rect 7849 18377 7883 18411
rect 9781 18377 9815 18411
rect 10793 18377 10827 18411
rect 14289 18377 14323 18411
rect 15485 18377 15519 18411
rect 16129 18377 16163 18411
rect 16865 18377 16899 18411
rect 17233 18377 17267 18411
rect 18705 18377 18739 18411
rect 24685 18377 24719 18411
rect 25053 18377 25087 18411
rect 26249 18377 26283 18411
rect 27537 18377 27571 18411
rect 28917 18377 28951 18411
rect 30113 18377 30147 18411
rect 32321 18377 32355 18411
rect 36185 18377 36219 18411
rect 36277 18377 36311 18411
rect 39865 18377 39899 18411
rect 40417 18377 40451 18411
rect 40877 18377 40911 18411
rect 24133 18309 24167 18343
rect 29009 18309 29043 18343
rect 30573 18309 30607 18343
rect 40785 18309 40819 18343
rect 1777 18241 1811 18275
rect 4445 18241 4479 18275
rect 7757 18241 7791 18275
rect 9965 18241 9999 18275
rect 15669 18241 15703 18275
rect 16313 18241 16347 18275
rect 18613 18241 18647 18275
rect 19625 18241 19659 18275
rect 22385 18241 22419 18275
rect 23305 18241 23339 18275
rect 25145 18241 25179 18275
rect 26341 18241 26375 18275
rect 27629 18241 27663 18275
rect 30481 18241 30515 18275
rect 31493 18241 31527 18275
rect 32689 18241 32723 18275
rect 38117 18241 38151 18275
rect 49065 18241 49099 18275
rect 2789 18173 2823 18207
rect 4169 18173 4203 18207
rect 10885 18173 10919 18207
rect 10977 18173 11011 18207
rect 11713 18173 11747 18207
rect 11989 18173 12023 18207
rect 14381 18173 14415 18207
rect 14565 18173 14599 18207
rect 17325 18173 17359 18207
rect 17417 18173 17451 18207
rect 18889 18173 18923 18207
rect 19901 18173 19935 18207
rect 22477 18173 22511 18207
rect 22661 18173 22695 18207
rect 25329 18173 25363 18207
rect 26433 18173 26467 18207
rect 27721 18173 27755 18207
rect 29101 18173 29135 18207
rect 30757 18173 30791 18207
rect 32781 18173 32815 18207
rect 32965 18173 32999 18207
rect 33609 18173 33643 18207
rect 33885 18173 33919 18207
rect 35357 18173 35391 18207
rect 36369 18173 36403 18207
rect 38393 18173 38427 18207
rect 40969 18173 41003 18207
rect 10425 18105 10459 18139
rect 13921 18105 13955 18139
rect 18153 18105 18187 18139
rect 25881 18105 25915 18139
rect 28549 18105 28583 18139
rect 13461 18037 13495 18071
rect 18245 18037 18279 18071
rect 21373 18037 21407 18071
rect 22017 18037 22051 18071
rect 27169 18037 27203 18071
rect 28457 18037 28491 18071
rect 35817 18037 35851 18071
rect 49249 18037 49283 18071
rect 12357 17833 12391 17867
rect 12909 17833 12943 17867
rect 16037 17833 16071 17867
rect 16773 17833 16807 17867
rect 23305 17833 23339 17867
rect 25237 17833 25271 17867
rect 40509 17833 40543 17867
rect 13553 17765 13587 17799
rect 19441 17765 19475 17799
rect 24593 17765 24627 17799
rect 37565 17765 37599 17799
rect 38025 17765 38059 17799
rect 2053 17697 2087 17731
rect 14289 17697 14323 17731
rect 18705 17697 18739 17731
rect 20269 17697 20303 17731
rect 23857 17697 23891 17731
rect 25881 17697 25915 17731
rect 30941 17697 30975 17731
rect 32137 17697 32171 17731
rect 33241 17697 33275 17731
rect 33425 17697 33459 17731
rect 35817 17697 35851 17731
rect 36093 17697 36127 17731
rect 38485 17697 38519 17731
rect 38577 17697 38611 17731
rect 40969 17697 41003 17731
rect 41061 17697 41095 17731
rect 1777 17629 1811 17663
rect 10609 17629 10643 17663
rect 13093 17629 13127 17663
rect 13737 17629 13771 17663
rect 19625 17629 19659 17663
rect 22661 17629 22695 17663
rect 24777 17629 24811 17663
rect 27077 17629 27111 17663
rect 30205 17629 30239 17663
rect 35081 17629 35115 17663
rect 49065 17629 49099 17663
rect 10885 17561 10919 17595
rect 14565 17561 14599 17595
rect 17325 17561 17359 17595
rect 17969 17561 18003 17595
rect 20545 17561 20579 17595
rect 25697 17561 25731 17595
rect 27353 17561 27387 17595
rect 31953 17561 31987 17595
rect 32045 17561 32079 17595
rect 38393 17561 38427 17595
rect 40877 17561 40911 17595
rect 17417 17493 17451 17527
rect 22017 17493 22051 17527
rect 22477 17493 22511 17527
rect 23673 17493 23707 17527
rect 23765 17493 23799 17527
rect 25605 17493 25639 17527
rect 28825 17493 28859 17527
rect 31585 17493 31619 17527
rect 32781 17493 32815 17527
rect 33149 17493 33183 17527
rect 49249 17493 49283 17527
rect 10425 17289 10459 17323
rect 12725 17289 12759 17323
rect 15577 17289 15611 17323
rect 21005 17289 21039 17323
rect 24961 17289 24995 17323
rect 25421 17289 25455 17323
rect 27353 17289 27387 17323
rect 29101 17289 29135 17323
rect 29193 17289 29227 17323
rect 30205 17289 30239 17323
rect 36369 17289 36403 17323
rect 37473 17289 37507 17323
rect 48421 17289 48455 17323
rect 13185 17221 13219 17255
rect 14197 17221 14231 17255
rect 16957 17221 16991 17255
rect 30297 17221 30331 17255
rect 34621 17221 34655 17255
rect 37841 17221 37875 17255
rect 39221 17221 39255 17255
rect 49157 17221 49191 17255
rect 1777 17153 1811 17187
rect 10793 17153 10827 17187
rect 11805 17153 11839 17187
rect 13093 17153 13127 17187
rect 15393 17153 15427 17187
rect 15945 17153 15979 17187
rect 16037 17153 16071 17187
rect 17877 17153 17911 17187
rect 19257 17153 19291 17187
rect 22753 17153 22787 17187
rect 25329 17153 25363 17187
rect 27721 17153 27755 17187
rect 28549 17153 28583 17187
rect 31401 17153 31435 17187
rect 32321 17153 32355 17187
rect 37933 17153 37967 17187
rect 48605 17153 48639 17187
rect 2053 17085 2087 17119
rect 10885 17085 10919 17119
rect 10977 17085 11011 17119
rect 11989 17085 12023 17119
rect 13277 17085 13311 17119
rect 15117 17085 15151 17119
rect 16129 17085 16163 17119
rect 18705 17085 18739 17119
rect 19533 17085 19567 17119
rect 24501 17085 24535 17119
rect 25513 17085 25547 17119
rect 27813 17085 27847 17119
rect 27997 17085 28031 17119
rect 29285 17085 29319 17119
rect 30389 17085 30423 17119
rect 31493 17085 31527 17119
rect 31585 17085 31619 17119
rect 32597 17085 32631 17119
rect 35357 17085 35391 17119
rect 36461 17085 36495 17119
rect 36645 17085 36679 17119
rect 38025 17085 38059 17119
rect 38945 17085 38979 17119
rect 14381 17017 14415 17051
rect 36001 17017 36035 17051
rect 15209 16949 15243 16983
rect 17049 16949 17083 16983
rect 23016 16949 23050 16983
rect 28733 16949 28767 16983
rect 29837 16949 29871 16983
rect 31033 16949 31067 16983
rect 34069 16949 34103 16983
rect 40693 16949 40727 16983
rect 49249 16949 49283 16983
rect 10517 16745 10551 16779
rect 17404 16745 17438 16779
rect 24777 16745 24811 16779
rect 27353 16745 27387 16779
rect 15669 16677 15703 16711
rect 8217 16609 8251 16643
rect 8401 16609 8435 16643
rect 11621 16609 11655 16643
rect 13461 16609 13495 16643
rect 13645 16609 13679 16643
rect 14933 16609 14967 16643
rect 15117 16609 15151 16643
rect 16129 16609 16163 16643
rect 16313 16609 16347 16643
rect 17141 16609 17175 16643
rect 19625 16609 19659 16643
rect 21005 16609 21039 16643
rect 21281 16609 21315 16643
rect 23765 16609 23799 16643
rect 23857 16609 23891 16643
rect 25605 16609 25639 16643
rect 25881 16609 25915 16643
rect 30297 16609 30331 16643
rect 31401 16609 31435 16643
rect 31585 16609 31619 16643
rect 32321 16609 32355 16643
rect 32597 16609 32631 16643
rect 35725 16609 35759 16643
rect 36737 16609 36771 16643
rect 36829 16609 36863 16643
rect 38025 16609 38059 16643
rect 1777 16541 1811 16575
rect 8125 16541 8159 16575
rect 12541 16541 12575 16575
rect 16037 16541 16071 16575
rect 20269 16541 20303 16575
rect 34897 16541 34931 16575
rect 36645 16541 36679 16575
rect 37749 16541 37783 16575
rect 49065 16541 49099 16575
rect 2513 16473 2547 16507
rect 10425 16473 10459 16507
rect 11437 16473 11471 16507
rect 13369 16473 13403 16507
rect 23673 16473 23707 16507
rect 30113 16473 30147 16507
rect 30205 16473 30239 16507
rect 7757 16405 7791 16439
rect 11069 16405 11103 16439
rect 11529 16405 11563 16439
rect 12357 16405 12391 16439
rect 13001 16405 13035 16439
rect 14473 16405 14507 16439
rect 14841 16405 14875 16439
rect 18889 16405 18923 16439
rect 20085 16405 20119 16439
rect 22753 16405 22787 16439
rect 23305 16405 23339 16439
rect 29745 16405 29779 16439
rect 30941 16405 30975 16439
rect 31309 16405 31343 16439
rect 34069 16405 34103 16439
rect 36277 16405 36311 16439
rect 39497 16405 39531 16439
rect 49249 16405 49283 16439
rect 8309 16201 8343 16235
rect 9321 16201 9355 16235
rect 11069 16201 11103 16235
rect 11805 16201 11839 16235
rect 13001 16201 13035 16235
rect 15945 16201 15979 16235
rect 16037 16201 16071 16235
rect 23029 16201 23063 16235
rect 25881 16201 25915 16235
rect 26341 16201 26375 16235
rect 27629 16201 27663 16235
rect 30297 16201 30331 16235
rect 31033 16201 31067 16235
rect 31125 16201 31159 16235
rect 32781 16201 32815 16235
rect 33977 16201 34011 16235
rect 40509 16201 40543 16235
rect 40969 16201 41003 16235
rect 9229 16133 9263 16167
rect 13093 16133 13127 16167
rect 14749 16133 14783 16167
rect 17785 16133 17819 16167
rect 19441 16133 19475 16167
rect 24409 16133 24443 16167
rect 28825 16133 28859 16167
rect 38485 16133 38519 16167
rect 1777 16065 1811 16099
rect 10977 16065 11011 16099
rect 12173 16065 12207 16099
rect 23397 16065 23431 16099
rect 24133 16065 24167 16099
rect 27537 16065 27571 16099
rect 28365 16065 28399 16099
rect 28549 16065 28583 16099
rect 32689 16065 32723 16099
rect 33885 16065 33919 16099
rect 40877 16065 40911 16099
rect 49065 16065 49099 16099
rect 2053 15997 2087 16031
rect 8401 15997 8435 16031
rect 8585 15997 8619 16031
rect 12265 15997 12299 16031
rect 12449 15997 12483 16031
rect 13185 15997 13219 16031
rect 13921 15997 13955 16031
rect 14841 15997 14875 16031
rect 14933 15997 14967 16031
rect 16129 15997 16163 16031
rect 17877 15997 17911 16031
rect 18061 15997 18095 16031
rect 19165 15997 19199 16031
rect 23489 15997 23523 16031
rect 23673 15997 23707 16031
rect 27721 15997 27755 16031
rect 31217 15997 31251 16031
rect 32873 15997 32907 16031
rect 34069 15997 34103 16031
rect 35081 15997 35115 16031
rect 35357 15997 35391 16031
rect 38209 15997 38243 16031
rect 41061 15997 41095 16031
rect 15577 15929 15611 15963
rect 36829 15929 36863 15963
rect 7941 15861 7975 15895
rect 12633 15861 12667 15895
rect 14381 15861 14415 15895
rect 17417 15861 17451 15895
rect 20913 15861 20947 15895
rect 27169 15861 27203 15895
rect 30665 15861 30699 15895
rect 32321 15861 32355 15895
rect 33517 15861 33551 15895
rect 39957 15861 39991 15895
rect 49249 15861 49283 15895
rect 13185 15657 13219 15691
rect 15577 15657 15611 15691
rect 16773 15657 16807 15691
rect 18061 15657 18095 15691
rect 19901 15657 19935 15691
rect 21189 15657 21223 15691
rect 25881 15657 25915 15691
rect 29193 15657 29227 15691
rect 32229 15657 32263 15691
rect 35160 15657 35194 15691
rect 36645 15657 36679 15691
rect 39497 15657 39531 15691
rect 41797 15657 41831 15691
rect 49157 15657 49191 15691
rect 32689 15589 32723 15623
rect 2053 15521 2087 15555
rect 10793 15521 10827 15555
rect 13645 15521 13679 15555
rect 13737 15521 13771 15555
rect 16129 15521 16163 15555
rect 17325 15521 17359 15555
rect 20545 15521 20579 15555
rect 21741 15521 21775 15555
rect 23673 15521 23707 15555
rect 25329 15521 25363 15555
rect 26433 15521 26467 15555
rect 27997 15521 28031 15555
rect 30481 15521 30515 15555
rect 33149 15521 33183 15555
rect 33333 15521 33367 15555
rect 37289 15521 37323 15555
rect 40049 15521 40083 15555
rect 1777 15453 1811 15487
rect 13553 15453 13587 15487
rect 15945 15453 15979 15487
rect 17233 15453 17267 15487
rect 18613 15453 18647 15487
rect 23581 15453 23615 15487
rect 25145 15453 25179 15487
rect 26249 15453 26283 15487
rect 27813 15453 27847 15487
rect 30021 15453 30055 15487
rect 34069 15453 34103 15487
rect 34897 15453 34931 15487
rect 37749 15453 37783 15487
rect 49341 15453 49375 15487
rect 6561 15385 6595 15419
rect 11069 15385 11103 15419
rect 20361 15385 20395 15419
rect 23489 15385 23523 15419
rect 25053 15385 25087 15419
rect 26341 15385 26375 15419
rect 27905 15385 27939 15419
rect 30757 15385 30791 15419
rect 38025 15385 38059 15419
rect 40325 15385 40359 15419
rect 6653 15317 6687 15351
rect 12541 15317 12575 15351
rect 15117 15317 15151 15351
rect 16037 15317 16071 15351
rect 17141 15317 17175 15351
rect 18429 15317 18463 15351
rect 20269 15317 20303 15351
rect 21557 15317 21591 15351
rect 21649 15317 21683 15351
rect 23121 15317 23155 15351
rect 24685 15317 24719 15351
rect 27445 15317 27479 15351
rect 33057 15317 33091 15351
rect 9781 15113 9815 15147
rect 11069 15113 11103 15147
rect 11897 15113 11931 15147
rect 12265 15113 12299 15147
rect 15577 15113 15611 15147
rect 16037 15113 16071 15147
rect 19533 15113 19567 15147
rect 22937 15113 22971 15147
rect 24133 15113 24167 15147
rect 25145 15113 25179 15147
rect 26433 15113 26467 15147
rect 27629 15113 27663 15147
rect 30113 15113 30147 15147
rect 31401 15113 31435 15147
rect 32689 15113 32723 15147
rect 33517 15113 33551 15147
rect 33885 15113 33919 15147
rect 35081 15113 35115 15147
rect 39681 15113 39715 15147
rect 40141 15113 40175 15147
rect 9873 15045 9907 15079
rect 10977 15045 11011 15079
rect 15945 15045 15979 15079
rect 18705 15045 18739 15079
rect 19901 15045 19935 15079
rect 21097 15045 21131 15079
rect 25605 15045 25639 15079
rect 28825 15045 28859 15079
rect 31493 15045 31527 15079
rect 32781 15045 32815 15079
rect 36369 15045 36403 15079
rect 37749 15045 37783 15079
rect 1777 14977 1811 15011
rect 13185 14977 13219 15011
rect 13277 14977 13311 15011
rect 17233 14977 17267 15011
rect 18153 14977 18187 15011
rect 18797 14977 18831 15011
rect 19993 14977 20027 15011
rect 23305 14977 23339 15011
rect 24501 14977 24535 15011
rect 24593 14977 24627 15011
rect 25513 14977 25547 15011
rect 27537 14977 27571 15011
rect 28733 14977 28767 15011
rect 36277 14977 36311 15011
rect 40049 14977 40083 15011
rect 41061 14977 41095 15011
rect 49065 14977 49099 15011
rect 2053 14909 2087 14943
rect 10057 14909 10091 14943
rect 12357 14909 12391 14943
rect 12449 14909 12483 14943
rect 15025 14909 15059 14943
rect 16129 14909 16163 14943
rect 17325 14909 17359 14943
rect 17417 14909 17451 14943
rect 18889 14909 18923 14943
rect 20085 14909 20119 14943
rect 21189 14909 21223 14943
rect 21281 14909 21315 14943
rect 23397 14909 23431 14943
rect 23489 14909 23523 14943
rect 24685 14909 24719 14943
rect 25789 14909 25823 14943
rect 27721 14909 27755 14943
rect 28917 14909 28951 14943
rect 29561 14909 29595 14943
rect 30205 14909 30239 14943
rect 30297 14909 30331 14943
rect 31585 14909 31619 14943
rect 32873 14909 32907 14943
rect 33977 14909 34011 14943
rect 34161 14909 34195 14943
rect 35173 14909 35207 14943
rect 35357 14909 35391 14943
rect 36461 14909 36495 14943
rect 37473 14909 37507 14943
rect 39221 14909 39255 14943
rect 40233 14909 40267 14943
rect 20729 14841 20763 14875
rect 28365 14841 28399 14875
rect 29745 14841 29779 14875
rect 34713 14841 34747 14875
rect 49249 14841 49283 14875
rect 9413 14773 9447 14807
rect 13540 14773 13574 14807
rect 16865 14773 16899 14807
rect 18337 14773 18371 14807
rect 27169 14773 27203 14807
rect 31033 14773 31067 14807
rect 32321 14773 32355 14807
rect 35909 14773 35943 14807
rect 40877 14773 40911 14807
rect 10425 14569 10459 14603
rect 11805 14569 11839 14603
rect 14289 14569 14323 14603
rect 24041 14569 24075 14603
rect 27261 14569 27295 14603
rect 29745 14569 29779 14603
rect 33425 14569 33459 14603
rect 36645 14569 36679 14603
rect 13001 14501 13035 14535
rect 18153 14501 18187 14535
rect 22845 14501 22879 14535
rect 38853 14501 38887 14535
rect 2053 14433 2087 14467
rect 12357 14433 12391 14467
rect 13553 14433 13587 14467
rect 14749 14433 14783 14467
rect 14933 14433 14967 14467
rect 15761 14433 15795 14467
rect 16957 14433 16991 14467
rect 18705 14433 18739 14467
rect 20085 14433 20119 14467
rect 21097 14433 21131 14467
rect 21373 14433 21407 14467
rect 26801 14433 26835 14467
rect 28273 14433 28307 14467
rect 28457 14433 28491 14467
rect 30297 14433 30331 14467
rect 31585 14433 31619 14467
rect 32689 14433 32723 14467
rect 32873 14433 32907 14467
rect 33977 14433 34011 14467
rect 34897 14433 34931 14467
rect 37105 14433 37139 14467
rect 37381 14433 37415 14467
rect 1777 14365 1811 14399
rect 9781 14365 9815 14399
rect 13369 14365 13403 14399
rect 15485 14365 15519 14399
rect 16129 14365 16163 14399
rect 16773 14365 16807 14399
rect 19993 14365 20027 14399
rect 20821 14365 20855 14399
rect 24961 14365 24995 14399
rect 25053 14365 25087 14399
rect 28181 14365 28215 14399
rect 30113 14365 30147 14399
rect 33885 14365 33919 14399
rect 39497 14365 39531 14399
rect 49065 14365 49099 14399
rect 9597 14297 9631 14331
rect 10333 14297 10367 14331
rect 11161 14297 11195 14331
rect 12173 14297 12207 14331
rect 14657 14297 14691 14331
rect 18613 14297 18647 14331
rect 25329 14297 25363 14331
rect 30205 14297 30239 14331
rect 31401 14297 31435 14331
rect 32597 14297 32631 14331
rect 33793 14297 33827 14331
rect 35173 14297 35207 14331
rect 11253 14229 11287 14263
rect 12265 14229 12299 14263
rect 13461 14229 13495 14263
rect 15117 14229 15151 14263
rect 15577 14229 15611 14263
rect 16405 14229 16439 14263
rect 16865 14229 16899 14263
rect 17601 14229 17635 14263
rect 18521 14229 18555 14263
rect 19533 14229 19567 14263
rect 19901 14229 19935 14263
rect 27813 14229 27847 14263
rect 31033 14229 31067 14263
rect 31493 14229 31527 14263
rect 32229 14229 32263 14263
rect 39313 14229 39347 14263
rect 49249 14229 49283 14263
rect 3617 14025 3651 14059
rect 11713 14025 11747 14059
rect 14657 14025 14691 14059
rect 15577 14025 15611 14059
rect 15945 14025 15979 14059
rect 17141 14025 17175 14059
rect 17509 14025 17543 14059
rect 17601 14025 17635 14059
rect 18337 14025 18371 14059
rect 18705 14025 18739 14059
rect 21465 14025 21499 14059
rect 26617 14025 26651 14059
rect 31125 14025 31159 14059
rect 34069 14025 34103 14059
rect 34897 14025 34931 14059
rect 35725 14025 35759 14059
rect 37841 14025 37875 14059
rect 45661 14025 45695 14059
rect 48421 14025 48455 14059
rect 49249 14025 49283 14059
rect 16037 13957 16071 13991
rect 19993 13957 20027 13991
rect 25145 13957 25179 13991
rect 36093 13957 36127 13991
rect 37933 13957 37967 13991
rect 45017 13957 45051 13991
rect 49157 13957 49191 13991
rect 1777 13889 1811 13923
rect 3525 13889 3559 13923
rect 11161 13889 11195 13923
rect 12081 13889 12115 13923
rect 18797 13889 18831 13923
rect 24869 13889 24903 13923
rect 27169 13889 27203 13923
rect 29377 13889 29411 13923
rect 31769 13889 31803 13923
rect 45845 13889 45879 13923
rect 48605 13889 48639 13923
rect 2053 13821 2087 13855
rect 12173 13821 12207 13855
rect 12357 13821 12391 13855
rect 12909 13821 12943 13855
rect 13185 13821 13219 13855
rect 16129 13821 16163 13855
rect 17785 13821 17819 13855
rect 18889 13821 18923 13855
rect 19717 13821 19751 13855
rect 22017 13821 22051 13855
rect 22293 13821 22327 13855
rect 24409 13821 24443 13855
rect 28917 13821 28951 13855
rect 32321 13821 32355 13855
rect 32597 13821 32631 13855
rect 34989 13821 35023 13855
rect 35081 13821 35115 13855
rect 36185 13821 36219 13855
rect 36369 13821 36403 13855
rect 38025 13821 38059 13855
rect 45201 13821 45235 13855
rect 23765 13753 23799 13787
rect 34529 13753 34563 13787
rect 37473 13753 37507 13787
rect 29640 13685 29674 13719
rect 38853 13685 38887 13719
rect 13277 13481 13311 13515
rect 18153 13481 18187 13515
rect 20913 13481 20947 13515
rect 22109 13481 22143 13515
rect 23305 13481 23339 13515
rect 24869 13481 24903 13515
rect 29745 13481 29779 13515
rect 33333 13481 33367 13515
rect 34897 13481 34931 13515
rect 14565 13413 14599 13447
rect 15669 13345 15703 13379
rect 15853 13345 15887 13379
rect 16405 13345 16439 13379
rect 21465 13345 21499 13379
rect 22569 13345 22603 13379
rect 22753 13345 22787 13379
rect 23765 13345 23799 13379
rect 23949 13345 23983 13379
rect 25513 13345 25547 13379
rect 26801 13345 26835 13379
rect 27077 13345 27111 13379
rect 28825 13345 28859 13379
rect 30205 13345 30239 13379
rect 30297 13345 30331 13379
rect 31033 13345 31067 13379
rect 32781 13345 32815 13379
rect 33793 13345 33827 13379
rect 33885 13345 33919 13379
rect 35541 13345 35575 13379
rect 38117 13345 38151 13379
rect 1777 13277 1811 13311
rect 2789 13277 2823 13311
rect 10793 13277 10827 13311
rect 14381 13277 14415 13311
rect 18889 13277 18923 13311
rect 21281 13277 21315 13311
rect 25237 13277 25271 13311
rect 26249 13277 26283 13311
rect 30113 13277 30147 13311
rect 33701 13277 33735 13311
rect 35265 13277 35299 13311
rect 36369 13277 36403 13311
rect 41521 13277 41555 13311
rect 47961 13277 47995 13311
rect 49157 13277 49191 13311
rect 11069 13209 11103 13243
rect 15577 13209 15611 13243
rect 16681 13209 16715 13243
rect 21373 13209 21407 13243
rect 22477 13209 22511 13243
rect 31309 13209 31343 13243
rect 35357 13209 35391 13243
rect 36645 13209 36679 13243
rect 12541 13141 12575 13175
rect 15209 13141 15243 13175
rect 20361 13141 20395 13175
rect 23673 13141 23707 13175
rect 25329 13141 25363 13175
rect 41337 13141 41371 13175
rect 2881 12937 2915 12971
rect 12173 12937 12207 12971
rect 15945 12937 15979 12971
rect 18889 12937 18923 12971
rect 19717 12937 19751 12971
rect 20085 12937 20119 12971
rect 23121 12937 23155 12971
rect 23949 12937 23983 12971
rect 25789 12937 25823 12971
rect 30665 12937 30699 12971
rect 34069 12937 34103 12971
rect 36369 12937 36403 12971
rect 1685 12869 1719 12903
rect 1869 12869 1903 12903
rect 12081 12869 12115 12903
rect 18705 12869 18739 12903
rect 32597 12869 32631 12903
rect 34529 12869 34563 12903
rect 38669 12869 38703 12903
rect 3065 12801 3099 12835
rect 16037 12801 16071 12835
rect 17877 12801 17911 12835
rect 19257 12801 19291 12835
rect 19349 12801 19383 12835
rect 21097 12801 21131 12835
rect 23029 12801 23063 12835
rect 27997 12801 28031 12835
rect 30573 12801 30607 12835
rect 32321 12801 32355 12835
rect 36277 12801 36311 12835
rect 39497 12801 39531 12835
rect 40049 12801 40083 12835
rect 46121 12801 46155 12835
rect 47961 12801 47995 12835
rect 49157 12801 49191 12835
rect 12265 12733 12299 12767
rect 13001 12733 13035 12767
rect 13277 12733 13311 12767
rect 14749 12733 14783 12767
rect 16129 12733 16163 12767
rect 19533 12733 19567 12767
rect 20177 12733 20211 12767
rect 20269 12733 20303 12767
rect 21189 12733 21223 12767
rect 21281 12733 21315 12767
rect 23213 12733 23247 12767
rect 24041 12733 24075 12767
rect 24317 12733 24351 12767
rect 28273 12733 28307 12767
rect 30849 12733 30883 12767
rect 35265 12733 35299 12767
rect 36461 12733 36495 12767
rect 20729 12665 20763 12699
rect 30205 12665 30239 12699
rect 35909 12665 35943 12699
rect 11713 12597 11747 12631
rect 15577 12597 15611 12631
rect 17417 12597 17451 12631
rect 22201 12597 22235 12631
rect 22661 12597 22695 12631
rect 27537 12597 27571 12631
rect 29745 12597 29779 12631
rect 31585 12597 31619 12631
rect 40141 12597 40175 12631
rect 45937 12597 45971 12631
rect 13001 12393 13035 12427
rect 20821 12393 20855 12427
rect 22109 12393 22143 12427
rect 26341 12393 26375 12427
rect 31493 12393 31527 12427
rect 33885 12393 33919 12427
rect 19441 12325 19475 12359
rect 41245 12325 41279 12359
rect 1869 12257 1903 12291
rect 10517 12257 10551 12291
rect 10793 12257 10827 12291
rect 13461 12257 13495 12291
rect 13645 12257 13679 12291
rect 14289 12257 14323 12291
rect 17233 12257 17267 12291
rect 19993 12257 20027 12291
rect 21465 12257 21499 12291
rect 22661 12257 22695 12291
rect 23857 12257 23891 12291
rect 27537 12257 27571 12291
rect 30021 12257 30055 12291
rect 34897 12257 34931 12291
rect 37473 12257 37507 12291
rect 37749 12257 37783 12291
rect 49157 12257 49191 12291
rect 1593 12189 1627 12223
rect 17049 12189 17083 12223
rect 17877 12189 17911 12223
rect 19809 12189 19843 12223
rect 21189 12189 21223 12223
rect 23673 12189 23707 12223
rect 24593 12189 24627 12223
rect 29745 12189 29779 12223
rect 32137 12189 32171 12223
rect 39957 12189 39991 12223
rect 40417 12189 40451 12223
rect 41429 12189 41463 12223
rect 46121 12189 46155 12223
rect 47961 12189 47995 12223
rect 14565 12121 14599 12155
rect 18613 12121 18647 12155
rect 22477 12121 22511 12155
rect 24869 12121 24903 12155
rect 27445 12121 27479 12155
rect 28273 12121 28307 12155
rect 29009 12121 29043 12155
rect 32413 12121 32447 12155
rect 35173 12121 35207 12155
rect 39497 12121 39531 12155
rect 40141 12121 40175 12155
rect 12265 12053 12299 12087
rect 13369 12053 13403 12087
rect 16037 12053 16071 12087
rect 16681 12053 16715 12087
rect 17141 12053 17175 12087
rect 19901 12053 19935 12087
rect 21281 12053 21315 12087
rect 22569 12053 22603 12087
rect 23305 12053 23339 12087
rect 23765 12053 23799 12087
rect 26985 12053 27019 12087
rect 27353 12053 27387 12087
rect 36645 12053 36679 12087
rect 40233 12053 40267 12087
rect 45937 12053 45971 12087
rect 18613 11849 18647 11883
rect 19901 11849 19935 11883
rect 27169 11849 27203 11883
rect 37657 11849 37691 11883
rect 38117 11849 38151 11883
rect 22569 11781 22603 11815
rect 24225 11781 24259 11815
rect 27537 11781 27571 11815
rect 32689 11781 32723 11815
rect 33793 11781 33827 11815
rect 37749 11781 37783 11815
rect 39405 11781 39439 11815
rect 45109 11781 45143 11815
rect 49157 11781 49191 11815
rect 1593 11713 1627 11747
rect 2513 11713 2547 11747
rect 12081 11713 12115 11747
rect 14105 11713 14139 11747
rect 15485 11713 15519 11747
rect 15577 11713 15611 11747
rect 21097 11713 21131 11747
rect 21189 11713 21223 11747
rect 26617 11713 26651 11747
rect 28457 11713 28491 11747
rect 31125 11713 31159 11747
rect 31217 11713 31251 11747
rect 35173 11713 35207 11747
rect 38485 11713 38519 11747
rect 47961 11713 47995 11747
rect 12357 11645 12391 11679
rect 15761 11645 15795 11679
rect 16865 11645 16899 11679
rect 17141 11645 17175 11679
rect 19993 11645 20027 11679
rect 20085 11645 20119 11679
rect 21373 11645 21407 11679
rect 23397 11645 23431 11679
rect 23949 11645 23983 11679
rect 25697 11645 25731 11679
rect 27629 11645 27663 11679
rect 27813 11645 27847 11679
rect 28733 11645 28767 11679
rect 31401 11645 31435 11679
rect 32781 11645 32815 11679
rect 32873 11645 32907 11679
rect 34529 11645 34563 11679
rect 35449 11645 35483 11679
rect 37841 11645 37875 11679
rect 38577 11645 38611 11679
rect 38669 11645 38703 11679
rect 1777 11577 1811 11611
rect 32321 11577 32355 11611
rect 39589 11577 39623 11611
rect 45293 11577 45327 11611
rect 2329 11509 2363 11543
rect 15117 11509 15151 11543
rect 19533 11509 19567 11543
rect 20729 11509 20763 11543
rect 30205 11509 30239 11543
rect 30757 11509 30791 11543
rect 36921 11509 36955 11543
rect 37289 11509 37323 11543
rect 14381 11305 14415 11339
rect 16773 11305 16807 11339
rect 19993 11305 20027 11339
rect 22201 11305 22235 11339
rect 22753 11305 22787 11339
rect 26341 11305 26375 11339
rect 27156 11305 27190 11339
rect 29745 11305 29779 11339
rect 38301 11305 38335 11339
rect 1777 11237 1811 11271
rect 12725 11237 12759 11271
rect 15577 11237 15611 11271
rect 17969 11237 18003 11271
rect 32873 11237 32907 11271
rect 33333 11237 33367 11271
rect 40785 11237 40819 11271
rect 10977 11169 11011 11203
rect 14841 11169 14875 11203
rect 15025 11169 15059 11203
rect 16037 11169 16071 11203
rect 16221 11169 16255 11203
rect 17417 11169 17451 11203
rect 18613 11169 18647 11203
rect 20453 11169 20487 11203
rect 23213 11169 23247 11203
rect 23397 11169 23431 11203
rect 24593 11169 24627 11203
rect 24869 11169 24903 11203
rect 28641 11169 28675 11203
rect 30205 11169 30239 11203
rect 30297 11169 30331 11203
rect 33977 11169 34011 11203
rect 36093 11169 36127 11203
rect 49157 11169 49191 11203
rect 1593 11101 1627 11135
rect 14749 11101 14783 11135
rect 15945 11101 15979 11135
rect 17141 11101 17175 11135
rect 18337 11101 18371 11135
rect 26893 11101 26927 11135
rect 31125 11101 31159 11135
rect 35817 11101 35851 11135
rect 38485 11101 38519 11135
rect 40969 11101 41003 11135
rect 45661 11101 45695 11135
rect 47961 11101 47995 11135
rect 11253 11033 11287 11067
rect 17233 11033 17267 11067
rect 20729 11033 20763 11067
rect 23121 11033 23155 11067
rect 30113 11033 30147 11067
rect 31401 11033 31435 11067
rect 33701 11033 33735 11067
rect 33793 11033 33827 11067
rect 37841 11033 37875 11067
rect 40141 11033 40175 11067
rect 40325 11033 40359 11067
rect 45845 11033 45879 11067
rect 18429 10965 18463 10999
rect 1777 10761 1811 10795
rect 13185 10761 13219 10795
rect 15945 10761 15979 10795
rect 16037 10761 16071 10795
rect 17785 10761 17819 10795
rect 18245 10761 18279 10795
rect 18981 10761 19015 10795
rect 19441 10761 19475 10795
rect 20637 10761 20671 10795
rect 24225 10761 24259 10795
rect 27169 10761 27203 10795
rect 36093 10761 36127 10795
rect 13553 10693 13587 10727
rect 22293 10693 22327 10727
rect 28825 10693 28859 10727
rect 34069 10693 34103 10727
rect 37933 10693 37967 10727
rect 49157 10693 49191 10727
rect 1593 10625 1627 10659
rect 2329 10625 2363 10659
rect 13645 10625 13679 10659
rect 14749 10625 14783 10659
rect 14841 10625 14875 10659
rect 17325 10625 17359 10659
rect 18153 10625 18187 10659
rect 19349 10625 19383 10659
rect 20545 10625 20579 10659
rect 24593 10625 24627 10659
rect 25605 10625 25639 10659
rect 27537 10625 27571 10659
rect 30573 10625 30607 10659
rect 31585 10625 31619 10659
rect 32689 10625 32723 10659
rect 36461 10625 36495 10659
rect 36553 10625 36587 10659
rect 37841 10625 37875 10659
rect 39773 10625 39807 10659
rect 47961 10625 47995 10659
rect 13737 10557 13771 10591
rect 14933 10557 14967 10591
rect 16129 10557 16163 10591
rect 18337 10557 18371 10591
rect 19625 10557 19659 10591
rect 20729 10557 20763 10591
rect 22017 10557 22051 10591
rect 24685 10557 24719 10591
rect 24869 10557 24903 10591
rect 27629 10557 27663 10591
rect 27813 10557 27847 10591
rect 29653 10557 29687 10591
rect 30665 10557 30699 10591
rect 30757 10557 30791 10591
rect 32781 10557 32815 10591
rect 32965 10557 32999 10591
rect 33793 10557 33827 10591
rect 36645 10557 36679 10591
rect 38025 10557 38059 10591
rect 2513 10489 2547 10523
rect 14381 10489 14415 10523
rect 23765 10489 23799 10523
rect 28365 10489 28399 10523
rect 30205 10489 30239 10523
rect 32321 10489 32355 10523
rect 39957 10489 39991 10523
rect 15577 10421 15611 10455
rect 20177 10421 20211 10455
rect 35541 10421 35575 10455
rect 37473 10421 37507 10455
rect 12817 10217 12851 10251
rect 16037 10217 16071 10251
rect 19717 10217 19751 10251
rect 22017 10217 22051 10251
rect 24041 10217 24075 10251
rect 28733 10217 28767 10251
rect 32137 10217 32171 10251
rect 36645 10217 36679 10251
rect 37473 10217 37507 10251
rect 11621 10149 11655 10183
rect 16589 10149 16623 10183
rect 33977 10149 34011 10183
rect 1869 10081 1903 10115
rect 12081 10081 12115 10115
rect 12173 10081 12207 10115
rect 13369 10081 13403 10115
rect 17049 10081 17083 10115
rect 17141 10081 17175 10115
rect 18245 10081 18279 10115
rect 18337 10081 18371 10115
rect 20269 10081 20303 10115
rect 23213 10081 23247 10115
rect 24593 10081 24627 10115
rect 30389 10081 30423 10115
rect 33149 10081 33183 10115
rect 34897 10081 34931 10115
rect 37933 10081 37967 10115
rect 38025 10081 38059 10115
rect 40325 10081 40359 10115
rect 49157 10081 49191 10115
rect 1593 10013 1627 10047
rect 11989 10013 12023 10047
rect 13277 10013 13311 10047
rect 14289 10013 14323 10047
rect 18153 10013 18187 10047
rect 22477 10013 22511 10047
rect 26985 10013 27019 10047
rect 29929 10013 29963 10047
rect 33057 10013 33091 10047
rect 37841 10013 37875 10047
rect 38945 10013 38979 10047
rect 44373 10013 44407 10047
rect 46121 10013 46155 10047
rect 47961 10013 47995 10047
rect 13185 9945 13219 9979
rect 14565 9945 14599 9979
rect 20545 9945 20579 9979
rect 24869 9945 24903 9979
rect 27261 9945 27295 9979
rect 30665 9945 30699 9979
rect 35173 9945 35207 9979
rect 38761 9945 38795 9979
rect 40141 9945 40175 9979
rect 44557 9945 44591 9979
rect 47317 9945 47351 9979
rect 16957 9877 16991 9911
rect 17785 9877 17819 9911
rect 26341 9877 26375 9911
rect 32597 9877 32631 9911
rect 32965 9877 32999 9911
rect 25697 9673 25731 9707
rect 29285 9673 29319 9707
rect 12449 9605 12483 9639
rect 12541 9605 12575 9639
rect 15301 9605 15335 9639
rect 18889 9605 18923 9639
rect 19625 9605 19659 9639
rect 22753 9605 22787 9639
rect 23949 9605 23983 9639
rect 32965 9605 32999 9639
rect 49157 9605 49191 9639
rect 1593 9537 1627 9571
rect 13277 9537 13311 9571
rect 22661 9537 22695 9571
rect 23673 9537 23707 9571
rect 26065 9537 26099 9571
rect 26157 9537 26191 9571
rect 33057 9537 33091 9571
rect 33885 9537 33919 9571
rect 47961 9537 47995 9571
rect 12725 9469 12759 9503
rect 13553 9469 13587 9503
rect 16865 9469 16899 9503
rect 17141 9469 17175 9503
rect 19349 9469 19383 9503
rect 21097 9469 21131 9503
rect 22845 9469 22879 9503
rect 26341 9469 26375 9503
rect 27537 9469 27571 9503
rect 27813 9469 27847 9503
rect 29745 9469 29779 9503
rect 30021 9469 30055 9503
rect 33149 9469 33183 9503
rect 34161 9469 34195 9503
rect 1777 9401 1811 9435
rect 12081 9401 12115 9435
rect 35633 9401 35667 9435
rect 22293 9333 22327 9367
rect 23581 9333 23615 9367
rect 25421 9333 25455 9367
rect 31493 9333 31527 9367
rect 32597 9333 32631 9367
rect 1777 9129 1811 9163
rect 14381 9129 14415 9163
rect 18061 9129 18095 9163
rect 18889 9129 18923 9163
rect 24041 9129 24075 9163
rect 28181 9129 28215 9163
rect 33333 9129 33367 9163
rect 24593 9061 24627 9095
rect 36645 9061 36679 9095
rect 14841 8993 14875 9027
rect 15025 8993 15059 9027
rect 22293 8993 22327 9027
rect 22569 8993 22603 9027
rect 25145 8993 25179 9027
rect 28825 8993 28859 9027
rect 31033 8993 31067 9027
rect 33885 8993 33919 9027
rect 35357 8993 35391 9027
rect 35449 8993 35483 9027
rect 39497 8993 39531 9027
rect 49157 8993 49191 9027
rect 1593 8925 1627 8959
rect 2329 8925 2363 8959
rect 13737 8925 13771 8959
rect 16313 8925 16347 8959
rect 19441 8925 19475 8959
rect 21833 8925 21867 8959
rect 28549 8925 28583 8959
rect 29929 8925 29963 8959
rect 30757 8925 30791 8959
rect 33701 8925 33735 8959
rect 36829 8925 36863 8959
rect 37841 8925 37875 8959
rect 47961 8925 47995 8959
rect 16589 8857 16623 8891
rect 19717 8857 19751 8891
rect 25053 8857 25087 8891
rect 39313 8857 39347 8891
rect 2513 8789 2547 8823
rect 13553 8789 13587 8823
rect 14749 8789 14783 8823
rect 21189 8789 21223 8823
rect 24961 8789 24995 8823
rect 27629 8789 27663 8823
rect 28641 8789 28675 8823
rect 32505 8789 32539 8823
rect 33793 8789 33827 8823
rect 34897 8789 34931 8823
rect 35265 8789 35299 8823
rect 37657 8789 37691 8823
rect 15301 8585 15335 8619
rect 18613 8585 18647 8619
rect 21465 8585 21499 8619
rect 30573 8585 30607 8619
rect 31033 8585 31067 8619
rect 34069 8585 34103 8619
rect 37473 8585 37507 8619
rect 40417 8585 40451 8619
rect 22293 8517 22327 8551
rect 29101 8517 29135 8551
rect 32597 8517 32631 8551
rect 44281 8517 44315 8551
rect 49157 8517 49191 8551
rect 1869 8449 1903 8483
rect 13553 8449 13587 8483
rect 16865 8449 16899 8483
rect 19257 8449 19291 8483
rect 19717 8449 19751 8483
rect 22017 8449 22051 8483
rect 31401 8449 31435 8483
rect 32321 8449 32355 8483
rect 37657 8449 37691 8483
rect 39129 8449 39163 8483
rect 40325 8449 40359 8483
rect 45845 8449 45879 8483
rect 47961 8449 47995 8483
rect 1593 8381 1627 8415
rect 13829 8381 13863 8415
rect 17141 8381 17175 8415
rect 19993 8381 20027 8415
rect 28825 8381 28859 8415
rect 31493 8381 31527 8415
rect 31677 8381 31711 8415
rect 46857 8381 46891 8415
rect 23765 8313 23799 8347
rect 38945 8313 38979 8347
rect 44465 8313 44499 8347
rect 21189 8041 21223 8075
rect 22017 8041 22051 8075
rect 29929 8041 29963 8075
rect 30573 8041 30607 8075
rect 17693 7973 17727 8007
rect 32321 7973 32355 8007
rect 18153 7905 18187 7939
rect 18245 7905 18279 7939
rect 19441 7905 19475 7939
rect 22661 7905 22695 7939
rect 31217 7905 31251 7939
rect 32965 7905 32999 7939
rect 49157 7905 49191 7939
rect 1593 7837 1627 7871
rect 15853 7837 15887 7871
rect 18061 7837 18095 7871
rect 22385 7837 22419 7871
rect 30941 7837 30975 7871
rect 31033 7837 31067 7871
rect 31861 7837 31895 7871
rect 38761 7837 38795 7871
rect 47961 7837 47995 7871
rect 19717 7769 19751 7803
rect 38025 7769 38059 7803
rect 38945 7769 38979 7803
rect 1777 7701 1811 7735
rect 15669 7701 15703 7735
rect 22477 7701 22511 7735
rect 32689 7701 32723 7735
rect 32781 7701 32815 7735
rect 38117 7701 38151 7735
rect 1777 7497 1811 7531
rect 22017 7497 22051 7531
rect 22477 7497 22511 7531
rect 23305 7497 23339 7531
rect 37841 7429 37875 7463
rect 44925 7429 44959 7463
rect 49157 7429 49191 7463
rect 1593 7361 1627 7395
rect 17877 7361 17911 7395
rect 22385 7361 22419 7395
rect 31125 7361 31159 7395
rect 38577 7361 38611 7395
rect 47961 7361 47995 7395
rect 22661 7293 22695 7327
rect 38761 7225 38795 7259
rect 17693 7157 17727 7191
rect 37933 7157 37967 7191
rect 45017 7157 45051 7191
rect 49157 6817 49191 6851
rect 1685 6749 1719 6783
rect 2513 6749 2547 6783
rect 19901 6749 19935 6783
rect 46121 6749 46155 6783
rect 47961 6749 47995 6783
rect 1869 6681 1903 6715
rect 47317 6681 47351 6715
rect 2329 6613 2363 6647
rect 19717 6613 19751 6647
rect 37565 6341 37599 6375
rect 44005 6341 44039 6375
rect 49157 6341 49191 6375
rect 1593 6273 1627 6307
rect 18061 6273 18095 6307
rect 47961 6273 47995 6307
rect 18245 6205 18279 6239
rect 44189 6137 44223 6171
rect 1777 6069 1811 6103
rect 18705 6069 18739 6103
rect 37657 6069 37691 6103
rect 2513 5797 2547 5831
rect 49157 5729 49191 5763
rect 1593 5661 1627 5695
rect 2329 5661 2363 5695
rect 43729 5661 43763 5695
rect 47961 5661 47995 5695
rect 43913 5593 43947 5627
rect 1777 5525 1811 5559
rect 37749 5253 37783 5287
rect 38485 5253 38519 5287
rect 49157 5253 49191 5287
rect 18981 5185 19015 5219
rect 22728 5185 22762 5219
rect 45845 5185 45879 5219
rect 47961 5185 47995 5219
rect 1593 5117 1627 5151
rect 1869 5117 1903 5151
rect 19165 5117 19199 5151
rect 46857 5117 46891 5151
rect 38669 5049 38703 5083
rect 19625 4981 19659 5015
rect 22799 4981 22833 5015
rect 37841 4981 37875 5015
rect 46765 4709 46799 4743
rect 1869 4641 1903 4675
rect 20453 4641 20487 4675
rect 21925 4641 21959 4675
rect 25145 4641 25179 4675
rect 25605 4641 25639 4675
rect 47501 4641 47535 4675
rect 49157 4641 49191 4675
rect 20637 4573 20671 4607
rect 22109 4573 22143 4607
rect 23448 4573 23482 4607
rect 38025 4573 38059 4607
rect 47961 4573 47995 4607
rect 1685 4505 1719 4539
rect 23535 4505 23569 4539
rect 25329 4505 25363 4539
rect 37289 4505 37323 4539
rect 37473 4505 37507 4539
rect 46581 4505 46615 4539
rect 47317 4505 47351 4539
rect 21097 4437 21131 4471
rect 22569 4437 22603 4471
rect 38117 4437 38151 4471
rect 1685 4165 1719 4199
rect 27353 4165 27387 4199
rect 2329 4097 2363 4131
rect 22636 4097 22670 4131
rect 23524 4097 23558 4131
rect 27169 4097 27203 4131
rect 45845 4097 45879 4131
rect 47961 4097 47995 4131
rect 49157 4097 49191 4131
rect 1869 4029 1903 4063
rect 24133 4029 24167 4063
rect 24317 4029 24351 4063
rect 24593 4029 24627 4063
rect 27629 4029 27663 4063
rect 46673 4029 46707 4063
rect 23627 3961 23661 3995
rect 2513 3893 2547 3927
rect 22707 3893 22741 3927
rect 23857 3689 23891 3723
rect 36553 3689 36587 3723
rect 45569 3689 45603 3723
rect 24041 3553 24075 3587
rect 24593 3553 24627 3587
rect 24777 3553 24811 3587
rect 25053 3553 25087 3587
rect 49157 3553 49191 3587
rect 1593 3485 1627 3519
rect 1869 3485 1903 3519
rect 16497 3485 16531 3519
rect 20913 3485 20947 3519
rect 23581 3485 23615 3519
rect 45477 3485 45511 3519
rect 46121 3485 46155 3519
rect 47961 3485 47995 3519
rect 21189 3417 21223 3451
rect 36461 3417 36495 3451
rect 47317 3417 47351 3451
rect 16589 3349 16623 3383
rect 22661 3349 22695 3383
rect 21281 3145 21315 3179
rect 24409 3077 24443 3111
rect 49157 3077 49191 3111
rect 1593 3009 1627 3043
rect 14565 3009 14599 3043
rect 17601 3009 17635 3043
rect 18337 3009 18371 3043
rect 20177 3009 20211 3043
rect 20821 3009 20855 3043
rect 21465 3009 21499 3043
rect 22201 3009 22235 3043
rect 23213 3009 23247 3043
rect 26525 3009 26559 3043
rect 27445 3009 27479 3043
rect 28917 3009 28951 3043
rect 44005 3009 44039 3043
rect 45845 3009 45879 3043
rect 47961 3009 47995 3043
rect 14841 2941 14875 2975
rect 16313 2941 16347 2975
rect 18613 2941 18647 2975
rect 24133 2941 24167 2975
rect 25881 2941 25915 2975
rect 29193 2941 29227 2975
rect 45201 2941 45235 2975
rect 46857 2941 46891 2975
rect 1777 2873 1811 2907
rect 19993 2873 20027 2907
rect 20637 2873 20671 2907
rect 22661 2873 22695 2907
rect 17417 2805 17451 2839
rect 22293 2805 22327 2839
rect 23305 2805 23339 2839
rect 23673 2805 23707 2839
rect 26341 2805 26375 2839
rect 27721 2805 27755 2839
rect 27905 2805 27939 2839
rect 30665 2805 30699 2839
rect 2513 2601 2547 2635
rect 29009 2601 29043 2635
rect 35081 2601 35115 2635
rect 1777 2533 1811 2567
rect 3065 2533 3099 2567
rect 9689 2533 9723 2567
rect 19441 2533 19475 2567
rect 30849 2533 30883 2567
rect 12265 2465 12299 2499
rect 14749 2465 14783 2499
rect 17325 2465 17359 2499
rect 20545 2465 20579 2499
rect 22845 2465 22879 2499
rect 25053 2465 25087 2499
rect 27629 2465 27663 2499
rect 37749 2465 37783 2499
rect 41429 2465 41463 2499
rect 43821 2465 43855 2499
rect 49157 2465 49191 2499
rect 1593 2397 1627 2431
rect 3249 2397 3283 2431
rect 9873 2397 9907 2431
rect 11989 2397 12023 2431
rect 14473 2397 14507 2431
rect 17049 2397 17083 2431
rect 18889 2397 18923 2431
rect 19625 2397 19659 2431
rect 20085 2397 20119 2431
rect 22385 2397 22419 2431
rect 24593 2397 24627 2431
rect 27169 2397 27203 2431
rect 29193 2397 29227 2431
rect 31033 2397 31067 2431
rect 33149 2397 33183 2431
rect 35265 2397 35299 2431
rect 37473 2397 37507 2431
rect 40693 2397 40727 2431
rect 43545 2397 43579 2431
rect 45845 2397 45879 2431
rect 47961 2397 47995 2431
rect 2421 2329 2455 2363
rect 47041 2329 47075 2363
rect 18705 2261 18739 2295
rect 32965 2261 32999 2295
<< metal1 >>
rect 3418 25168 3424 25220
rect 3476 25208 3482 25220
rect 9214 25208 9220 25220
rect 3476 25180 9220 25208
rect 3476 25168 3482 25180
rect 9214 25168 9220 25180
rect 9272 25168 9278 25220
rect 3326 25032 3332 25084
rect 3384 25072 3390 25084
rect 8846 25072 8852 25084
rect 3384 25044 8852 25072
rect 3384 25032 3390 25044
rect 8846 25032 8852 25044
rect 8904 25032 8910 25084
rect 32122 24896 32128 24948
rect 32180 24936 32186 24948
rect 39206 24936 39212 24948
rect 32180 24908 39212 24936
rect 32180 24896 32186 24908
rect 39206 24896 39212 24908
rect 39264 24896 39270 24948
rect 28810 24828 28816 24880
rect 28868 24868 28874 24880
rect 48682 24868 48688 24880
rect 28868 24840 48688 24868
rect 28868 24828 28874 24840
rect 48682 24828 48688 24840
rect 48740 24828 48746 24880
rect 24026 24760 24032 24812
rect 24084 24800 24090 24812
rect 27798 24800 27804 24812
rect 24084 24772 27804 24800
rect 24084 24760 24090 24772
rect 27798 24760 27804 24772
rect 27856 24760 27862 24812
rect 32858 24760 32864 24812
rect 32916 24800 32922 24812
rect 36538 24800 36544 24812
rect 32916 24772 36544 24800
rect 32916 24760 32922 24772
rect 36538 24760 36544 24772
rect 36596 24760 36602 24812
rect 38930 24760 38936 24812
rect 38988 24800 38994 24812
rect 41782 24800 41788 24812
rect 38988 24772 41788 24800
rect 38988 24760 38994 24772
rect 41782 24760 41788 24772
rect 41840 24760 41846 24812
rect 19058 24692 19064 24744
rect 19116 24732 19122 24744
rect 22094 24732 22100 24744
rect 19116 24704 22100 24732
rect 19116 24692 19122 24704
rect 22094 24692 22100 24704
rect 22152 24692 22158 24744
rect 27430 24732 27436 24744
rect 24596 24704 27436 24732
rect 17586 24624 17592 24676
rect 17644 24664 17650 24676
rect 24596 24664 24624 24704
rect 27430 24692 27436 24704
rect 27488 24692 27494 24744
rect 36262 24692 36268 24744
rect 36320 24732 36326 24744
rect 40678 24732 40684 24744
rect 36320 24704 40684 24732
rect 36320 24692 36326 24704
rect 40678 24692 40684 24704
rect 40736 24692 40742 24744
rect 29086 24664 29092 24676
rect 17644 24636 24624 24664
rect 24688 24636 29092 24664
rect 17644 24624 17650 24636
rect 3142 24556 3148 24608
rect 3200 24596 3206 24608
rect 5718 24596 5724 24608
rect 3200 24568 5724 24596
rect 3200 24556 3206 24568
rect 5718 24556 5724 24568
rect 5776 24556 5782 24608
rect 17770 24556 17776 24608
rect 17828 24596 17834 24608
rect 20070 24596 20076 24608
rect 17828 24568 20076 24596
rect 17828 24556 17834 24568
rect 20070 24556 20076 24568
rect 20128 24556 20134 24608
rect 21450 24556 21456 24608
rect 21508 24596 21514 24608
rect 24688 24596 24716 24636
rect 29086 24624 29092 24636
rect 29144 24624 29150 24676
rect 29270 24624 29276 24676
rect 29328 24664 29334 24676
rect 35066 24664 35072 24676
rect 29328 24636 35072 24664
rect 29328 24624 29334 24636
rect 35066 24624 35072 24636
rect 35124 24624 35130 24676
rect 35710 24624 35716 24676
rect 35768 24664 35774 24676
rect 43530 24664 43536 24676
rect 35768 24636 43536 24664
rect 35768 24624 35774 24636
rect 43530 24624 43536 24636
rect 43588 24624 43594 24676
rect 21508 24568 24716 24596
rect 21508 24556 21514 24568
rect 24762 24556 24768 24608
rect 24820 24596 24826 24608
rect 31202 24596 31208 24608
rect 24820 24568 31208 24596
rect 24820 24556 24826 24568
rect 31202 24556 31208 24568
rect 31260 24556 31266 24608
rect 34974 24556 34980 24608
rect 35032 24596 35038 24608
rect 40034 24596 40040 24608
rect 35032 24568 40040 24596
rect 35032 24556 35038 24568
rect 40034 24556 40040 24568
rect 40092 24556 40098 24608
rect 1104 24506 49864 24528
rect 1104 24454 2950 24506
rect 3002 24454 3014 24506
rect 3066 24454 3078 24506
rect 3130 24454 3142 24506
rect 3194 24454 3206 24506
rect 3258 24454 12950 24506
rect 13002 24454 13014 24506
rect 13066 24454 13078 24506
rect 13130 24454 13142 24506
rect 13194 24454 13206 24506
rect 13258 24454 22950 24506
rect 23002 24454 23014 24506
rect 23066 24454 23078 24506
rect 23130 24454 23142 24506
rect 23194 24454 23206 24506
rect 23258 24454 32950 24506
rect 33002 24454 33014 24506
rect 33066 24454 33078 24506
rect 33130 24454 33142 24506
rect 33194 24454 33206 24506
rect 33258 24454 42950 24506
rect 43002 24454 43014 24506
rect 43066 24454 43078 24506
rect 43130 24454 43142 24506
rect 43194 24454 43206 24506
rect 43258 24454 49864 24506
rect 1104 24432 49864 24454
rect 2774 24352 2780 24404
rect 2832 24392 2838 24404
rect 6270 24392 6276 24404
rect 2832 24364 6276 24392
rect 2832 24352 2838 24364
rect 6270 24352 6276 24364
rect 6328 24352 6334 24404
rect 24026 24392 24032 24404
rect 19628 24364 24032 24392
rect 6730 24284 6736 24336
rect 6788 24284 6794 24336
rect 11882 24324 11888 24336
rect 10980 24296 11888 24324
rect 3237 24259 3295 24265
rect 3237 24225 3249 24259
rect 3283 24256 3295 24259
rect 3510 24256 3516 24268
rect 3283 24228 3516 24256
rect 3283 24225 3295 24228
rect 3237 24219 3295 24225
rect 3510 24216 3516 24228
rect 3568 24216 3574 24268
rect 5813 24259 5871 24265
rect 5813 24225 5825 24259
rect 5859 24256 5871 24259
rect 6748 24256 6776 24284
rect 5859 24228 6776 24256
rect 8205 24259 8263 24265
rect 5859 24225 5871 24228
rect 5813 24219 5871 24225
rect 8205 24225 8217 24259
rect 8251 24256 8263 24259
rect 8662 24256 8668 24268
rect 8251 24228 8668 24256
rect 8251 24225 8263 24228
rect 8205 24219 8263 24225
rect 8662 24216 8668 24228
rect 8720 24216 8726 24268
rect 10980 24265 11008 24296
rect 11882 24284 11888 24296
rect 11940 24284 11946 24336
rect 16022 24324 16028 24336
rect 12406 24296 16028 24324
rect 10965 24259 11023 24265
rect 10965 24225 10977 24259
rect 11011 24225 11023 24259
rect 12406 24256 12434 24296
rect 16022 24284 16028 24296
rect 16080 24284 16086 24336
rect 17037 24327 17095 24333
rect 17037 24293 17049 24327
rect 17083 24324 17095 24327
rect 19426 24324 19432 24336
rect 17083 24296 19432 24324
rect 17083 24293 17095 24296
rect 17037 24287 17095 24293
rect 19426 24284 19432 24296
rect 19484 24284 19490 24336
rect 10965 24219 11023 24225
rect 11900 24228 12434 24256
rect 13541 24259 13599 24265
rect 2225 24191 2283 24197
rect 2225 24157 2237 24191
rect 2271 24188 2283 24191
rect 2314 24188 2320 24200
rect 2271 24160 2320 24188
rect 2271 24157 2283 24160
rect 2225 24151 2283 24157
rect 2314 24148 2320 24160
rect 2372 24148 2378 24200
rect 4157 24191 4215 24197
rect 4157 24157 4169 24191
rect 4203 24188 4215 24191
rect 4706 24188 4712 24200
rect 4203 24160 4712 24188
rect 4203 24157 4215 24160
rect 4157 24151 4215 24157
rect 4706 24148 4712 24160
rect 4764 24148 4770 24200
rect 4801 24191 4859 24197
rect 4801 24157 4813 24191
rect 4847 24188 4859 24191
rect 6546 24188 6552 24200
rect 4847 24160 6552 24188
rect 4847 24157 4859 24160
rect 4801 24151 4859 24157
rect 6546 24148 6552 24160
rect 6604 24148 6610 24200
rect 6733 24191 6791 24197
rect 6733 24157 6745 24191
rect 6779 24188 6791 24191
rect 7377 24191 7435 24197
rect 6779 24160 6914 24188
rect 6779 24157 6791 24160
rect 6733 24151 6791 24157
rect 6886 24120 6914 24160
rect 7377 24157 7389 24191
rect 7423 24188 7435 24191
rect 7466 24188 7472 24200
rect 7423 24160 7472 24188
rect 7423 24157 7435 24160
rect 7377 24151 7435 24157
rect 7466 24148 7472 24160
rect 7524 24148 7530 24200
rect 9309 24191 9367 24197
rect 9309 24157 9321 24191
rect 9355 24188 9367 24191
rect 9674 24188 9680 24200
rect 9355 24160 9680 24188
rect 9355 24157 9367 24160
rect 9309 24151 9367 24157
rect 9674 24148 9680 24160
rect 9732 24148 9738 24200
rect 11900 24197 11928 24228
rect 13541 24225 13553 24259
rect 13587 24256 13599 24259
rect 13814 24256 13820 24268
rect 13587 24228 13820 24256
rect 13587 24225 13599 24228
rect 13541 24219 13599 24225
rect 13814 24216 13820 24228
rect 13872 24216 13878 24268
rect 16117 24259 16175 24265
rect 16117 24225 16129 24259
rect 16163 24256 16175 24259
rect 17678 24256 17684 24268
rect 16163 24228 17684 24256
rect 16163 24225 16175 24228
rect 16117 24219 16175 24225
rect 17678 24216 17684 24228
rect 17736 24216 17742 24268
rect 18693 24259 18751 24265
rect 18693 24225 18705 24259
rect 18739 24256 18751 24259
rect 19518 24256 19524 24268
rect 18739 24228 19524 24256
rect 18739 24225 18751 24228
rect 18693 24219 18751 24225
rect 19518 24216 19524 24228
rect 19576 24216 19582 24268
rect 9953 24191 10011 24197
rect 9953 24157 9965 24191
rect 9999 24188 10011 24191
rect 11885 24191 11943 24197
rect 9999 24160 11744 24188
rect 9999 24157 10011 24160
rect 9953 24151 10011 24157
rect 10318 24120 10324 24132
rect 6886 24092 10324 24120
rect 10318 24080 10324 24092
rect 10376 24080 10382 24132
rect 11716 24120 11744 24160
rect 11885 24157 11897 24191
rect 11931 24157 11943 24191
rect 11885 24151 11943 24157
rect 12529 24191 12587 24197
rect 12529 24157 12541 24191
rect 12575 24188 12587 24191
rect 12618 24188 12624 24200
rect 12575 24160 12624 24188
rect 12575 24157 12587 24160
rect 12529 24151 12587 24157
rect 12618 24148 12624 24160
rect 12676 24148 12682 24200
rect 14458 24148 14464 24200
rect 14516 24148 14522 24200
rect 15105 24191 15163 24197
rect 15105 24157 15117 24191
rect 15151 24188 15163 24191
rect 16574 24188 16580 24200
rect 15151 24160 16580 24188
rect 15151 24157 15163 24160
rect 15105 24151 15163 24157
rect 16574 24148 16580 24160
rect 16632 24148 16638 24200
rect 17586 24148 17592 24200
rect 17644 24148 17650 24200
rect 19628 24197 19656 24364
rect 24026 24352 24032 24364
rect 24084 24352 24090 24404
rect 24118 24352 24124 24404
rect 24176 24392 24182 24404
rect 24176 24364 31432 24392
rect 24176 24352 24182 24364
rect 20530 24284 20536 24336
rect 20588 24324 20594 24336
rect 20588 24296 22094 24324
rect 20588 24284 20594 24296
rect 19720 24228 20208 24256
rect 19613 24191 19671 24197
rect 19613 24157 19625 24191
rect 19659 24157 19671 24191
rect 19613 24151 19671 24157
rect 13630 24120 13636 24132
rect 11716 24092 13636 24120
rect 13630 24080 13636 24092
rect 13688 24080 13694 24132
rect 13722 24080 13728 24132
rect 13780 24120 13786 24132
rect 19720 24120 19748 24228
rect 20073 24191 20131 24197
rect 20073 24157 20085 24191
rect 20119 24157 20131 24191
rect 20073 24151 20131 24157
rect 13780 24092 19748 24120
rect 13780 24080 13786 24092
rect 3973 24055 4031 24061
rect 3973 24021 3985 24055
rect 4019 24052 4031 24055
rect 4614 24052 4620 24064
rect 4019 24024 4620 24052
rect 4019 24021 4031 24024
rect 3973 24015 4031 24021
rect 4614 24012 4620 24024
rect 4672 24012 4678 24064
rect 6549 24055 6607 24061
rect 6549 24021 6561 24055
rect 6595 24052 6607 24055
rect 7466 24052 7472 24064
rect 6595 24024 7472 24052
rect 6595 24021 6607 24024
rect 6549 24015 6607 24021
rect 7466 24012 7472 24024
rect 7524 24012 7530 24064
rect 9122 24012 9128 24064
rect 9180 24012 9186 24064
rect 13446 24012 13452 24064
rect 13504 24052 13510 24064
rect 14277 24055 14335 24061
rect 14277 24052 14289 24055
rect 13504 24024 14289 24052
rect 13504 24012 13510 24024
rect 14277 24021 14289 24024
rect 14323 24021 14335 24055
rect 14277 24015 14335 24021
rect 19429 24055 19487 24061
rect 19429 24021 19441 24055
rect 19475 24052 19487 24055
rect 20088 24052 20116 24151
rect 19475 24024 20116 24052
rect 20180 24052 20208 24228
rect 20898 24216 20904 24268
rect 20956 24216 20962 24268
rect 22066 24256 22094 24296
rect 23566 24284 23572 24336
rect 23624 24324 23630 24336
rect 24581 24327 24639 24333
rect 24581 24324 24593 24327
rect 23624 24296 24593 24324
rect 23624 24284 23630 24296
rect 24581 24293 24593 24296
rect 24627 24293 24639 24327
rect 24581 24287 24639 24293
rect 24946 24284 24952 24336
rect 25004 24324 25010 24336
rect 25004 24296 25084 24324
rect 25004 24284 25010 24296
rect 25056 24265 25084 24296
rect 26142 24284 26148 24336
rect 26200 24324 26206 24336
rect 28718 24324 28724 24336
rect 26200 24296 28724 24324
rect 26200 24284 26206 24296
rect 28718 24284 28724 24296
rect 28776 24284 28782 24336
rect 28902 24284 28908 24336
rect 28960 24324 28966 24336
rect 28960 24296 31340 24324
rect 28960 24284 28966 24296
rect 22465 24259 22523 24265
rect 22465 24256 22477 24259
rect 22066 24228 22477 24256
rect 22465 24225 22477 24228
rect 22511 24225 22523 24259
rect 22465 24219 22523 24225
rect 25041 24259 25099 24265
rect 25041 24225 25053 24259
rect 25087 24225 25099 24259
rect 25041 24219 25099 24225
rect 25130 24216 25136 24268
rect 25188 24216 25194 24268
rect 26326 24216 26332 24268
rect 26384 24216 26390 24268
rect 27982 24216 27988 24268
rect 28040 24256 28046 24268
rect 28040 24228 29960 24256
rect 28040 24216 28046 24228
rect 22186 24148 22192 24200
rect 22244 24148 22250 24200
rect 24029 24191 24087 24197
rect 24029 24157 24041 24191
rect 24075 24188 24087 24191
rect 25406 24188 25412 24200
rect 24075 24160 25412 24188
rect 24075 24157 24087 24160
rect 24029 24151 24087 24157
rect 25406 24148 25412 24160
rect 25464 24148 25470 24200
rect 26050 24148 26056 24200
rect 26108 24188 26114 24200
rect 26145 24191 26203 24197
rect 26145 24188 26157 24191
rect 26108 24160 26157 24188
rect 26108 24148 26114 24160
rect 26145 24157 26157 24160
rect 26191 24157 26203 24191
rect 26145 24151 26203 24157
rect 26694 24148 26700 24200
rect 26752 24188 26758 24200
rect 28077 24191 28135 24197
rect 28077 24188 28089 24191
rect 26752 24160 28089 24188
rect 26752 24148 26758 24160
rect 28077 24157 28089 24160
rect 28123 24157 28135 24191
rect 28077 24151 28135 24157
rect 28718 24148 28724 24200
rect 28776 24148 28782 24200
rect 29932 24197 29960 24228
rect 29917 24191 29975 24197
rect 29917 24157 29929 24191
rect 29963 24157 29975 24191
rect 29917 24151 29975 24157
rect 30561 24191 30619 24197
rect 30561 24157 30573 24191
rect 30607 24157 30619 24191
rect 30561 24151 30619 24157
rect 24949 24123 25007 24129
rect 24949 24120 24961 24123
rect 22066 24092 24961 24120
rect 22066 24052 22094 24092
rect 24949 24089 24961 24092
rect 24995 24120 25007 24123
rect 25777 24123 25835 24129
rect 25777 24120 25789 24123
rect 24995 24092 25789 24120
rect 24995 24089 25007 24092
rect 24949 24083 25007 24089
rect 25777 24089 25789 24092
rect 25823 24089 25835 24123
rect 26418 24120 26424 24132
rect 25777 24083 25835 24089
rect 26160 24092 26424 24120
rect 20180 24024 22094 24052
rect 23845 24055 23903 24061
rect 19475 24021 19487 24024
rect 19429 24015 19487 24021
rect 23845 24021 23857 24055
rect 23891 24052 23903 24055
rect 26160 24052 26188 24092
rect 26418 24080 26424 24092
rect 26476 24080 26482 24132
rect 27246 24080 27252 24132
rect 27304 24080 27310 24132
rect 29086 24080 29092 24132
rect 29144 24120 29150 24132
rect 30576 24120 30604 24151
rect 31202 24148 31208 24200
rect 31260 24148 31266 24200
rect 31312 24188 31340 24296
rect 31404 24256 31432 24364
rect 31478 24352 31484 24404
rect 31536 24392 31542 24404
rect 35897 24395 35955 24401
rect 35897 24392 35909 24395
rect 31536 24364 35909 24392
rect 31536 24352 31542 24364
rect 35897 24361 35909 24364
rect 35943 24361 35955 24395
rect 35897 24355 35955 24361
rect 36004 24364 36584 24392
rect 31846 24284 31852 24336
rect 31904 24324 31910 24336
rect 32953 24327 33011 24333
rect 32953 24324 32965 24327
rect 31904 24296 32965 24324
rect 31904 24284 31910 24296
rect 32953 24293 32965 24296
rect 32999 24293 33011 24327
rect 36004 24324 36032 24364
rect 32953 24287 33011 24293
rect 34072 24296 36032 24324
rect 36556 24324 36584 24364
rect 37550 24352 37556 24404
rect 37608 24392 37614 24404
rect 38562 24392 38568 24404
rect 37608 24364 38568 24392
rect 37608 24352 37614 24364
rect 38562 24352 38568 24364
rect 38620 24352 38626 24404
rect 39206 24352 39212 24404
rect 39264 24352 39270 24404
rect 40034 24352 40040 24404
rect 40092 24352 40098 24404
rect 40678 24352 40684 24404
rect 40736 24352 40742 24404
rect 48314 24352 48320 24404
rect 48372 24352 48378 24404
rect 39666 24324 39672 24336
rect 36556 24296 39672 24324
rect 34072 24265 34100 24296
rect 39666 24284 39672 24296
rect 39724 24284 39730 24336
rect 39942 24284 39948 24336
rect 40000 24324 40006 24336
rect 40954 24324 40960 24336
rect 40000 24296 40960 24324
rect 40000 24284 40006 24296
rect 40954 24284 40960 24296
rect 41012 24284 41018 24336
rect 34057 24259 34115 24265
rect 31404 24228 33180 24256
rect 33152 24197 33180 24228
rect 34057 24225 34069 24259
rect 34103 24225 34115 24259
rect 34057 24219 34115 24225
rect 34241 24259 34299 24265
rect 34241 24225 34253 24259
rect 34287 24256 34299 24259
rect 34287 24228 36492 24256
rect 34287 24225 34299 24228
rect 34241 24219 34299 24225
rect 32493 24191 32551 24197
rect 32493 24188 32505 24191
rect 31312 24160 32505 24188
rect 32493 24157 32505 24160
rect 32539 24157 32551 24191
rect 32493 24151 32551 24157
rect 33137 24191 33195 24197
rect 33137 24157 33149 24191
rect 33183 24157 33195 24191
rect 33137 24151 33195 24157
rect 35066 24148 35072 24200
rect 35124 24148 35130 24200
rect 36354 24148 36360 24200
rect 36412 24148 36418 24200
rect 36464 24188 36492 24228
rect 36538 24216 36544 24268
rect 36596 24216 36602 24268
rect 37550 24256 37556 24268
rect 37200 24228 37556 24256
rect 37200 24188 37228 24228
rect 37550 24216 37556 24228
rect 37608 24216 37614 24268
rect 37918 24216 37924 24268
rect 37976 24216 37982 24268
rect 38105 24259 38163 24265
rect 38105 24225 38117 24259
rect 38151 24256 38163 24259
rect 38378 24256 38384 24268
rect 38151 24228 38384 24256
rect 38151 24225 38163 24228
rect 38105 24219 38163 24225
rect 38378 24216 38384 24228
rect 38436 24216 38442 24268
rect 38654 24216 38660 24268
rect 38712 24256 38718 24268
rect 48041 24259 48099 24265
rect 38712 24228 41736 24256
rect 38712 24216 38718 24228
rect 39114 24188 39120 24200
rect 36464 24160 37228 24188
rect 37292 24160 39120 24188
rect 36265 24123 36323 24129
rect 29144 24092 30420 24120
rect 30576 24092 33640 24120
rect 29144 24080 29150 24092
rect 23891 24024 26188 24052
rect 23891 24021 23903 24024
rect 23845 24015 23903 24021
rect 26234 24012 26240 24064
rect 26292 24052 26298 24064
rect 27341 24055 27399 24061
rect 27341 24052 27353 24055
rect 26292 24024 27353 24052
rect 26292 24012 26298 24024
rect 27341 24021 27353 24024
rect 27387 24021 27399 24055
rect 27341 24015 27399 24021
rect 27706 24012 27712 24064
rect 27764 24052 27770 24064
rect 27893 24055 27951 24061
rect 27893 24052 27905 24055
rect 27764 24024 27905 24052
rect 27764 24012 27770 24024
rect 27893 24021 27905 24024
rect 27939 24021 27951 24055
rect 27893 24015 27951 24021
rect 28442 24012 28448 24064
rect 28500 24052 28506 24064
rect 28537 24055 28595 24061
rect 28537 24052 28549 24055
rect 28500 24024 28549 24052
rect 28500 24012 28506 24024
rect 28537 24021 28549 24024
rect 28583 24021 28595 24055
rect 28537 24015 28595 24021
rect 29178 24012 29184 24064
rect 29236 24052 29242 24064
rect 30392 24061 30420 24092
rect 29733 24055 29791 24061
rect 29733 24052 29745 24055
rect 29236 24024 29745 24052
rect 29236 24012 29242 24024
rect 29733 24021 29745 24024
rect 29779 24021 29791 24055
rect 29733 24015 29791 24021
rect 30377 24055 30435 24061
rect 30377 24021 30389 24055
rect 30423 24021 30435 24055
rect 30377 24015 30435 24021
rect 30466 24012 30472 24064
rect 30524 24052 30530 24064
rect 31021 24055 31079 24061
rect 31021 24052 31033 24055
rect 30524 24024 31033 24052
rect 30524 24012 30530 24024
rect 31021 24021 31033 24024
rect 31067 24021 31079 24055
rect 31021 24015 31079 24021
rect 31938 24012 31944 24064
rect 31996 24052 32002 24064
rect 33612 24061 33640 24092
rect 36265 24089 36277 24123
rect 36311 24120 36323 24123
rect 37292 24120 37320 24160
rect 39114 24148 39120 24160
rect 39172 24148 39178 24200
rect 39206 24148 39212 24200
rect 39264 24188 39270 24200
rect 41708 24197 41736 24228
rect 48041 24225 48053 24259
rect 48087 24256 48099 24259
rect 48222 24256 48228 24268
rect 48087 24228 48228 24256
rect 48087 24225 48099 24228
rect 48041 24219 48099 24225
rect 48222 24216 48228 24228
rect 48280 24256 48286 24268
rect 48501 24259 48559 24265
rect 48501 24256 48513 24259
rect 48280 24228 48513 24256
rect 48280 24216 48286 24228
rect 48501 24225 48513 24228
rect 48547 24225 48559 24259
rect 48501 24219 48559 24225
rect 40221 24191 40279 24197
rect 40221 24188 40233 24191
rect 39264 24160 40233 24188
rect 39264 24148 39270 24160
rect 40221 24157 40233 24160
rect 40267 24157 40279 24191
rect 40221 24151 40279 24157
rect 40865 24191 40923 24197
rect 40865 24157 40877 24191
rect 40911 24188 40923 24191
rect 41325 24191 41383 24197
rect 41325 24188 41337 24191
rect 40911 24160 41337 24188
rect 40911 24157 40923 24160
rect 40865 24151 40923 24157
rect 41325 24157 41337 24160
rect 41371 24157 41383 24191
rect 41325 24151 41383 24157
rect 41693 24191 41751 24197
rect 41693 24157 41705 24191
rect 41739 24157 41751 24191
rect 41693 24151 41751 24157
rect 36311 24092 37320 24120
rect 37384 24092 37688 24120
rect 36311 24089 36323 24092
rect 36265 24083 36323 24089
rect 32309 24055 32367 24061
rect 32309 24052 32321 24055
rect 31996 24024 32321 24052
rect 31996 24012 32002 24024
rect 32309 24021 32321 24024
rect 32355 24021 32367 24055
rect 32309 24015 32367 24021
rect 33597 24055 33655 24061
rect 33597 24021 33609 24055
rect 33643 24021 33655 24055
rect 33597 24015 33655 24021
rect 33962 24012 33968 24064
rect 34020 24012 34026 24064
rect 34882 24012 34888 24064
rect 34940 24012 34946 24064
rect 35618 24012 35624 24064
rect 35676 24052 35682 24064
rect 37384 24052 37412 24092
rect 35676 24024 37412 24052
rect 35676 24012 35682 24024
rect 37458 24012 37464 24064
rect 37516 24012 37522 24064
rect 37660 24052 37688 24092
rect 37734 24080 37740 24132
rect 37792 24120 37798 24132
rect 40880 24120 40908 24151
rect 42150 24148 42156 24200
rect 42208 24188 42214 24200
rect 42613 24191 42671 24197
rect 42613 24188 42625 24191
rect 42208 24160 42625 24188
rect 42208 24148 42214 24160
rect 42613 24157 42625 24160
rect 42659 24157 42671 24191
rect 42613 24151 42671 24157
rect 44726 24148 44732 24200
rect 44784 24188 44790 24200
rect 45281 24191 45339 24197
rect 45281 24188 45293 24191
rect 44784 24160 45293 24188
rect 44784 24148 44790 24160
rect 45281 24157 45293 24160
rect 45327 24157 45339 24191
rect 45281 24151 45339 24157
rect 45554 24148 45560 24200
rect 45612 24188 45618 24200
rect 45925 24191 45983 24197
rect 45925 24188 45937 24191
rect 45612 24160 45937 24188
rect 45612 24148 45618 24160
rect 45925 24157 45937 24160
rect 45971 24157 45983 24191
rect 45925 24151 45983 24157
rect 46014 24148 46020 24200
rect 46072 24188 46078 24200
rect 46753 24191 46811 24197
rect 46753 24188 46765 24191
rect 46072 24160 46765 24188
rect 46072 24148 46078 24160
rect 46753 24157 46765 24160
rect 46799 24157 46811 24191
rect 46753 24151 46811 24157
rect 47302 24148 47308 24200
rect 47360 24188 47366 24200
rect 48133 24191 48191 24197
rect 48133 24188 48145 24191
rect 47360 24160 48145 24188
rect 47360 24148 47366 24160
rect 48133 24157 48145 24160
rect 48179 24157 48191 24191
rect 48133 24151 48191 24157
rect 48590 24148 48596 24200
rect 48648 24188 48654 24200
rect 48777 24191 48835 24197
rect 48777 24188 48789 24191
rect 48648 24160 48789 24188
rect 48648 24148 48654 24160
rect 48777 24157 48789 24160
rect 48823 24157 48835 24191
rect 48777 24151 48835 24157
rect 37792 24092 40908 24120
rect 37792 24080 37798 24092
rect 40954 24080 40960 24132
rect 41012 24120 41018 24132
rect 41138 24120 41144 24132
rect 41012 24092 41144 24120
rect 41012 24080 41018 24092
rect 41138 24080 41144 24092
rect 41196 24120 41202 24132
rect 45465 24123 45523 24129
rect 45465 24120 45477 24123
rect 41196 24092 45477 24120
rect 41196 24080 41202 24092
rect 45465 24089 45477 24092
rect 45511 24089 45523 24123
rect 45465 24083 45523 24089
rect 46934 24080 46940 24132
rect 46992 24080 46998 24132
rect 37829 24055 37887 24061
rect 37829 24052 37841 24055
rect 37660 24024 37841 24052
rect 37829 24021 37841 24024
rect 37875 24052 37887 24055
rect 39850 24052 39856 24064
rect 37875 24024 39856 24052
rect 37875 24021 37887 24024
rect 37829 24015 37887 24021
rect 39850 24012 39856 24024
rect 39908 24012 39914 24064
rect 40770 24012 40776 24064
rect 40828 24052 40834 24064
rect 41509 24055 41567 24061
rect 41509 24052 41521 24055
rect 40828 24024 41521 24052
rect 40828 24012 40834 24024
rect 41509 24021 41521 24024
rect 41555 24021 41567 24055
rect 41509 24015 41567 24021
rect 43346 24012 43352 24064
rect 43404 24052 43410 24064
rect 43901 24055 43959 24061
rect 43901 24052 43913 24055
rect 43404 24024 43913 24052
rect 43404 24012 43410 24024
rect 43901 24021 43913 24024
rect 43947 24021 43959 24055
rect 43901 24015 43959 24021
rect 46106 24012 46112 24064
rect 46164 24012 46170 24064
rect 1104 23962 49864 23984
rect 1104 23910 7950 23962
rect 8002 23910 8014 23962
rect 8066 23910 8078 23962
rect 8130 23910 8142 23962
rect 8194 23910 8206 23962
rect 8258 23910 17950 23962
rect 18002 23910 18014 23962
rect 18066 23910 18078 23962
rect 18130 23910 18142 23962
rect 18194 23910 18206 23962
rect 18258 23910 27950 23962
rect 28002 23910 28014 23962
rect 28066 23910 28078 23962
rect 28130 23910 28142 23962
rect 28194 23910 28206 23962
rect 28258 23910 37950 23962
rect 38002 23910 38014 23962
rect 38066 23910 38078 23962
rect 38130 23910 38142 23962
rect 38194 23910 38206 23962
rect 38258 23910 47950 23962
rect 48002 23910 48014 23962
rect 48066 23910 48078 23962
rect 48130 23910 48142 23962
rect 48194 23910 48206 23962
rect 48258 23910 49864 23962
rect 1104 23888 49864 23910
rect 6546 23808 6552 23860
rect 6604 23808 6610 23860
rect 12710 23848 12716 23860
rect 8128 23820 12716 23848
rect 3973 23783 4031 23789
rect 3973 23749 3985 23783
rect 4019 23780 4031 23783
rect 4154 23780 4160 23792
rect 4019 23752 4160 23780
rect 4019 23749 4031 23752
rect 3973 23743 4031 23749
rect 4154 23740 4160 23752
rect 4212 23740 4218 23792
rect 2961 23715 3019 23721
rect 2961 23681 2973 23715
rect 3007 23712 3019 23715
rect 3510 23712 3516 23724
rect 3007 23684 3516 23712
rect 3007 23681 3019 23684
rect 2961 23675 3019 23681
rect 3510 23672 3516 23684
rect 3568 23672 3574 23724
rect 4614 23672 4620 23724
rect 4672 23672 4678 23724
rect 6733 23715 6791 23721
rect 6733 23681 6745 23715
rect 6779 23712 6791 23715
rect 7282 23712 7288 23724
rect 6779 23684 7288 23712
rect 6779 23681 6791 23684
rect 6733 23675 6791 23681
rect 7282 23672 7288 23684
rect 7340 23672 7346 23724
rect 8128 23721 8156 23820
rect 12710 23808 12716 23820
rect 12768 23808 12774 23860
rect 18708 23820 20392 23848
rect 9125 23783 9183 23789
rect 9125 23749 9137 23783
rect 9171 23780 9183 23783
rect 9306 23780 9312 23792
rect 9171 23752 9312 23780
rect 9171 23749 9183 23752
rect 9125 23743 9183 23749
rect 9306 23740 9312 23752
rect 9364 23740 9370 23792
rect 10594 23740 10600 23792
rect 10652 23780 10658 23792
rect 10689 23783 10747 23789
rect 10689 23780 10701 23783
rect 10652 23752 10701 23780
rect 10652 23740 10658 23752
rect 10689 23749 10701 23752
rect 10735 23749 10747 23783
rect 10689 23743 10747 23749
rect 14366 23740 14372 23792
rect 14424 23740 14430 23792
rect 16114 23740 16120 23792
rect 16172 23740 16178 23792
rect 18141 23783 18199 23789
rect 18141 23749 18153 23783
rect 18187 23780 18199 23783
rect 18322 23780 18328 23792
rect 18187 23752 18328 23780
rect 18187 23749 18199 23752
rect 18141 23743 18199 23749
rect 18322 23740 18328 23752
rect 18380 23740 18386 23792
rect 7469 23715 7527 23721
rect 7469 23681 7481 23715
rect 7515 23681 7527 23715
rect 7469 23675 7527 23681
rect 8113 23715 8171 23721
rect 8113 23681 8125 23715
rect 8159 23681 8171 23715
rect 8113 23675 8171 23681
rect 9953 23715 10011 23721
rect 9953 23681 9965 23715
rect 9999 23712 10011 23715
rect 11793 23715 11851 23721
rect 9999 23684 11560 23712
rect 9999 23681 10011 23684
rect 9953 23675 10011 23681
rect 5442 23604 5448 23656
rect 5500 23604 5506 23656
rect 7484 23644 7512 23675
rect 9582 23644 9588 23656
rect 7484 23616 9588 23644
rect 9582 23604 9588 23616
rect 9640 23604 9646 23656
rect 3418 23536 3424 23588
rect 3476 23576 3482 23588
rect 5534 23576 5540 23588
rect 3476 23548 5540 23576
rect 3476 23536 3482 23548
rect 5534 23536 5540 23548
rect 5592 23536 5598 23588
rect 11532 23576 11560 23684
rect 11793 23681 11805 23715
rect 11839 23712 11851 23715
rect 11839 23684 13216 23712
rect 11839 23681 11851 23684
rect 11793 23675 11851 23681
rect 12066 23604 12072 23656
rect 12124 23604 12130 23656
rect 12434 23576 12440 23588
rect 11532 23548 12440 23576
rect 12434 23536 12440 23548
rect 12492 23536 12498 23588
rect 13188 23585 13216 23684
rect 13446 23672 13452 23724
rect 13504 23672 13510 23724
rect 15105 23715 15163 23721
rect 15105 23681 15117 23715
rect 15151 23681 15163 23715
rect 15105 23675 15163 23681
rect 17129 23715 17187 23721
rect 17129 23681 17141 23715
rect 17175 23712 17187 23715
rect 18708 23712 18736 23820
rect 19058 23740 19064 23792
rect 19116 23740 19122 23792
rect 20364 23780 20392 23820
rect 20438 23808 20444 23860
rect 20496 23848 20502 23860
rect 23474 23848 23480 23860
rect 20496 23820 23480 23848
rect 20496 23808 20502 23820
rect 23474 23808 23480 23820
rect 23532 23808 23538 23860
rect 23937 23851 23995 23857
rect 23937 23848 23949 23851
rect 23584 23820 23949 23848
rect 20364 23752 20484 23780
rect 17175 23684 18736 23712
rect 17175 23681 17187 23684
rect 17129 23675 17187 23681
rect 15120 23644 15148 23675
rect 18782 23672 18788 23724
rect 18840 23672 18846 23724
rect 20162 23672 20168 23724
rect 20220 23672 20226 23724
rect 17954 23644 17960 23656
rect 15120 23616 17960 23644
rect 17954 23604 17960 23616
rect 18012 23604 18018 23656
rect 20254 23644 20260 23656
rect 18892 23616 20260 23644
rect 13173 23579 13231 23585
rect 13173 23545 13185 23579
rect 13219 23576 13231 23579
rect 18892 23576 18920 23616
rect 20254 23604 20260 23616
rect 20312 23604 20318 23656
rect 20456 23644 20484 23752
rect 20530 23740 20536 23792
rect 20588 23780 20594 23792
rect 23584 23780 23612 23820
rect 23937 23817 23949 23820
rect 23983 23817 23995 23851
rect 23937 23811 23995 23817
rect 27798 23808 27804 23860
rect 27856 23848 27862 23860
rect 27893 23851 27951 23857
rect 27893 23848 27905 23851
rect 27856 23820 27905 23848
rect 27856 23808 27862 23820
rect 27893 23817 27905 23820
rect 27939 23817 27951 23851
rect 32309 23851 32367 23857
rect 32309 23848 32321 23851
rect 27893 23811 27951 23817
rect 29380 23820 32321 23848
rect 20588 23752 23612 23780
rect 23845 23783 23903 23789
rect 20588 23740 20594 23752
rect 23845 23749 23857 23783
rect 23891 23780 23903 23783
rect 25222 23780 25228 23792
rect 23891 23752 25228 23780
rect 23891 23749 23903 23752
rect 23845 23743 23903 23749
rect 25222 23740 25228 23752
rect 25280 23740 25286 23792
rect 26418 23780 26424 23792
rect 26358 23752 26424 23780
rect 26418 23740 26424 23752
rect 26476 23740 26482 23792
rect 27338 23740 27344 23792
rect 27396 23780 27402 23792
rect 27396 23752 28764 23780
rect 27396 23740 27402 23752
rect 21450 23672 21456 23724
rect 21508 23672 21514 23724
rect 22925 23715 22983 23721
rect 22925 23681 22937 23715
rect 22971 23712 22983 23715
rect 23474 23712 23480 23724
rect 22971 23684 23480 23712
rect 22971 23681 22983 23684
rect 22925 23675 22983 23681
rect 23474 23672 23480 23684
rect 23532 23672 23538 23724
rect 27154 23672 27160 23724
rect 27212 23712 27218 23724
rect 27249 23715 27307 23721
rect 27249 23712 27261 23715
rect 27212 23684 27261 23712
rect 27212 23672 27218 23684
rect 27249 23681 27261 23684
rect 27295 23681 27307 23715
rect 27249 23675 27307 23681
rect 27430 23672 27436 23724
rect 27488 23672 27494 23724
rect 28736 23721 28764 23752
rect 29380 23721 29408 23820
rect 32309 23817 32321 23820
rect 32355 23817 32367 23851
rect 32309 23811 32367 23817
rect 33962 23808 33968 23860
rect 34020 23848 34026 23860
rect 36081 23851 36139 23857
rect 36081 23848 36093 23851
rect 34020 23820 36093 23848
rect 34020 23808 34026 23820
rect 36081 23817 36093 23820
rect 36127 23817 36139 23851
rect 36081 23811 36139 23817
rect 37458 23808 37464 23860
rect 37516 23848 37522 23860
rect 39117 23851 39175 23857
rect 39117 23848 39129 23851
rect 37516 23820 39129 23848
rect 37516 23808 37522 23820
rect 39117 23817 39129 23820
rect 39163 23817 39175 23851
rect 39117 23811 39175 23817
rect 39850 23808 39856 23860
rect 39908 23848 39914 23860
rect 39908 23820 41184 23848
rect 39908 23808 39914 23820
rect 30742 23740 30748 23792
rect 30800 23740 30806 23792
rect 32769 23783 32827 23789
rect 32769 23749 32781 23783
rect 32815 23780 32827 23783
rect 34146 23780 34152 23792
rect 32815 23752 34152 23780
rect 32815 23749 32827 23752
rect 32769 23743 32827 23749
rect 34146 23740 34152 23752
rect 34204 23740 34210 23792
rect 34330 23740 34336 23792
rect 34388 23740 34394 23792
rect 35250 23740 35256 23792
rect 35308 23780 35314 23792
rect 39025 23783 39083 23789
rect 35308 23752 38884 23780
rect 35308 23740 35314 23752
rect 28077 23715 28135 23721
rect 28077 23681 28089 23715
rect 28123 23681 28135 23715
rect 28077 23675 28135 23681
rect 28721 23715 28779 23721
rect 28721 23681 28733 23715
rect 28767 23681 28779 23715
rect 28721 23675 28779 23681
rect 29365 23715 29423 23721
rect 29365 23681 29377 23715
rect 29411 23681 29423 23715
rect 29365 23675 29423 23681
rect 23017 23647 23075 23653
rect 20456 23616 22876 23644
rect 13219 23548 18920 23576
rect 13219 23545 13231 23548
rect 13173 23539 13231 23545
rect 20070 23536 20076 23588
rect 20128 23576 20134 23588
rect 22557 23579 22615 23585
rect 22557 23576 22569 23579
rect 20128 23548 22569 23576
rect 20128 23536 20134 23548
rect 22557 23545 22569 23548
rect 22603 23545 22615 23579
rect 22557 23539 22615 23545
rect 4798 23468 4804 23520
rect 4856 23508 4862 23520
rect 7285 23511 7343 23517
rect 7285 23508 7297 23511
rect 4856 23480 7297 23508
rect 4856 23468 4862 23480
rect 7285 23477 7297 23480
rect 7331 23477 7343 23511
rect 7285 23471 7343 23477
rect 9674 23468 9680 23520
rect 9732 23508 9738 23520
rect 16574 23508 16580 23520
rect 9732 23480 16580 23508
rect 9732 23468 9738 23480
rect 16574 23468 16580 23480
rect 16632 23468 16638 23520
rect 18782 23468 18788 23520
rect 18840 23508 18846 23520
rect 20346 23508 20352 23520
rect 18840 23480 20352 23508
rect 18840 23468 18846 23480
rect 20346 23468 20352 23480
rect 20404 23468 20410 23520
rect 20530 23468 20536 23520
rect 20588 23468 20594 23520
rect 21266 23468 21272 23520
rect 21324 23468 21330 23520
rect 22848 23508 22876 23616
rect 23017 23613 23029 23647
rect 23063 23613 23075 23647
rect 23017 23607 23075 23613
rect 23201 23647 23259 23653
rect 23201 23613 23213 23647
rect 23247 23644 23259 23647
rect 23290 23644 23296 23656
rect 23247 23616 23296 23644
rect 23247 23613 23259 23616
rect 23201 23607 23259 23613
rect 23032 23576 23060 23607
rect 23290 23604 23296 23616
rect 23348 23604 23354 23656
rect 24854 23604 24860 23656
rect 24912 23604 24918 23656
rect 25133 23647 25191 23653
rect 25133 23613 25145 23647
rect 25179 23644 25191 23647
rect 27614 23644 27620 23656
rect 25179 23616 27620 23644
rect 25179 23613 25191 23616
rect 25133 23607 25191 23613
rect 27614 23604 27620 23616
rect 27672 23604 27678 23656
rect 28092 23644 28120 23675
rect 32674 23672 32680 23724
rect 32732 23672 32738 23724
rect 36449 23715 36507 23721
rect 36449 23681 36461 23715
rect 36495 23712 36507 23715
rect 37366 23712 37372 23724
rect 36495 23684 37372 23712
rect 36495 23681 36507 23684
rect 36449 23675 36507 23681
rect 37366 23672 37372 23684
rect 37424 23672 37430 23724
rect 37826 23672 37832 23724
rect 37884 23672 37890 23724
rect 37921 23715 37979 23721
rect 37921 23681 37933 23715
rect 37967 23712 37979 23715
rect 38746 23712 38752 23724
rect 37967 23684 38752 23712
rect 37967 23681 37979 23684
rect 37921 23675 37979 23681
rect 38746 23672 38752 23684
rect 38804 23672 38810 23724
rect 29730 23644 29736 23656
rect 28092 23616 29736 23644
rect 29730 23604 29736 23616
rect 29788 23604 29794 23656
rect 30006 23604 30012 23656
rect 30064 23604 30070 23656
rect 30285 23647 30343 23653
rect 30285 23644 30297 23647
rect 30116 23616 30297 23644
rect 24762 23576 24768 23588
rect 23032 23548 24768 23576
rect 24762 23536 24768 23548
rect 24820 23536 24826 23588
rect 29270 23576 29276 23588
rect 26436 23548 29276 23576
rect 25130 23508 25136 23520
rect 22848 23480 25136 23508
rect 25130 23468 25136 23480
rect 25188 23468 25194 23520
rect 25222 23468 25228 23520
rect 25280 23508 25286 23520
rect 26436 23508 26464 23548
rect 29270 23536 29276 23548
rect 29328 23536 29334 23588
rect 29362 23536 29368 23588
rect 29420 23576 29426 23588
rect 30116 23576 30144 23616
rect 30285 23613 30297 23616
rect 30331 23644 30343 23647
rect 32398 23644 32404 23656
rect 30331 23616 32404 23644
rect 30331 23613 30343 23616
rect 30285 23607 30343 23613
rect 32398 23604 32404 23616
rect 32456 23644 32462 23656
rect 32858 23644 32864 23656
rect 32456 23616 32864 23644
rect 32456 23604 32462 23616
rect 32858 23604 32864 23616
rect 32916 23604 32922 23656
rect 32953 23647 33011 23653
rect 32953 23613 32965 23647
rect 32999 23613 33011 23647
rect 32953 23607 33011 23613
rect 29420 23548 30144 23576
rect 29420 23536 29426 23548
rect 25280 23480 26464 23508
rect 25280 23468 25286 23480
rect 26602 23468 26608 23520
rect 26660 23468 26666 23520
rect 28537 23511 28595 23517
rect 28537 23477 28549 23511
rect 28583 23508 28595 23511
rect 28626 23508 28632 23520
rect 28583 23480 28632 23508
rect 28583 23477 28595 23480
rect 28537 23471 28595 23477
rect 28626 23468 28632 23480
rect 28684 23468 28690 23520
rect 28994 23468 29000 23520
rect 29052 23508 29058 23520
rect 29181 23511 29239 23517
rect 29181 23508 29193 23511
rect 29052 23480 29193 23508
rect 29052 23468 29058 23480
rect 29181 23477 29193 23480
rect 29227 23477 29239 23511
rect 29181 23471 29239 23477
rect 30282 23468 30288 23520
rect 30340 23508 30346 23520
rect 31478 23508 31484 23520
rect 30340 23480 31484 23508
rect 30340 23468 30346 23480
rect 31478 23468 31484 23480
rect 31536 23468 31542 23520
rect 31662 23468 31668 23520
rect 31720 23508 31726 23520
rect 31757 23511 31815 23517
rect 31757 23508 31769 23511
rect 31720 23480 31769 23508
rect 31720 23468 31726 23480
rect 31757 23477 31769 23480
rect 31803 23477 31815 23511
rect 32968 23508 32996 23607
rect 33318 23604 33324 23656
rect 33376 23644 33382 23656
rect 33597 23647 33655 23653
rect 33597 23644 33609 23647
rect 33376 23616 33609 23644
rect 33376 23604 33382 23616
rect 33597 23613 33609 23616
rect 33643 23613 33655 23647
rect 33597 23607 33655 23613
rect 33870 23604 33876 23656
rect 33928 23604 33934 23656
rect 34238 23604 34244 23656
rect 34296 23644 34302 23656
rect 34296 23616 35756 23644
rect 34296 23604 34302 23616
rect 34882 23536 34888 23588
rect 34940 23576 34946 23588
rect 35618 23576 35624 23588
rect 34940 23548 35624 23576
rect 34940 23536 34946 23548
rect 35618 23536 35624 23548
rect 35676 23536 35682 23588
rect 35728 23576 35756 23616
rect 36538 23604 36544 23656
rect 36596 23604 36602 23656
rect 36722 23604 36728 23656
rect 36780 23604 36786 23656
rect 38105 23647 38163 23653
rect 38105 23613 38117 23647
rect 38151 23644 38163 23647
rect 38286 23644 38292 23656
rect 38151 23616 38292 23644
rect 38151 23613 38163 23616
rect 38105 23607 38163 23613
rect 38286 23604 38292 23616
rect 38344 23604 38350 23656
rect 38856 23644 38884 23752
rect 39025 23749 39037 23783
rect 39071 23780 39083 23783
rect 40034 23780 40040 23792
rect 39071 23752 40040 23780
rect 39071 23749 39083 23752
rect 39025 23743 39083 23749
rect 40034 23740 40040 23752
rect 40092 23740 40098 23792
rect 39316 23684 41092 23712
rect 39209 23647 39267 23653
rect 39209 23644 39221 23647
rect 38856 23616 39221 23644
rect 39209 23613 39221 23616
rect 39255 23613 39267 23647
rect 39209 23607 39267 23613
rect 38657 23579 38715 23585
rect 38657 23576 38669 23579
rect 35728 23548 38669 23576
rect 38657 23545 38669 23548
rect 38703 23545 38715 23579
rect 38657 23539 38715 23545
rect 35342 23508 35348 23520
rect 32968 23480 35348 23508
rect 31757 23471 31815 23477
rect 35342 23468 35348 23480
rect 35400 23468 35406 23520
rect 35434 23468 35440 23520
rect 35492 23508 35498 23520
rect 37461 23511 37519 23517
rect 37461 23508 37473 23511
rect 35492 23480 37473 23508
rect 35492 23468 35498 23480
rect 37461 23477 37473 23480
rect 37507 23477 37519 23511
rect 37461 23471 37519 23477
rect 38562 23468 38568 23520
rect 38620 23508 38626 23520
rect 39316 23508 39344 23684
rect 39942 23604 39948 23656
rect 40000 23604 40006 23656
rect 41064 23653 41092 23684
rect 40037 23647 40095 23653
rect 40037 23613 40049 23647
rect 40083 23613 40095 23647
rect 40037 23607 40095 23613
rect 41049 23647 41107 23653
rect 41049 23613 41061 23647
rect 41095 23613 41107 23647
rect 41049 23607 41107 23613
rect 39758 23536 39764 23588
rect 39816 23576 39822 23588
rect 40052 23576 40080 23607
rect 39816 23548 40080 23576
rect 41156 23576 41184 23820
rect 41230 23808 41236 23860
rect 41288 23848 41294 23860
rect 44315 23851 44373 23857
rect 44315 23848 44327 23851
rect 41288 23820 44327 23848
rect 41288 23808 41294 23820
rect 44315 23817 44327 23820
rect 44361 23817 44373 23851
rect 48961 23851 49019 23857
rect 48961 23848 48973 23851
rect 44315 23811 44373 23817
rect 44560 23820 48973 23848
rect 41322 23740 41328 23792
rect 41380 23740 41386 23792
rect 41414 23740 41420 23792
rect 41472 23780 41478 23792
rect 44560 23780 44588 23820
rect 48961 23817 48973 23820
rect 49007 23817 49019 23851
rect 48961 23811 49019 23817
rect 41472 23752 44588 23780
rect 41472 23740 41478 23752
rect 46842 23740 46848 23792
rect 46900 23740 46906 23792
rect 47854 23740 47860 23792
rect 47912 23780 47918 23792
rect 48133 23783 48191 23789
rect 48133 23780 48145 23783
rect 47912 23752 48145 23780
rect 47912 23740 47918 23752
rect 48133 23749 48145 23752
rect 48179 23749 48191 23783
rect 48133 23743 48191 23749
rect 41340 23712 41368 23740
rect 45189 23715 45247 23721
rect 45189 23712 45201 23715
rect 41340 23684 45201 23712
rect 45189 23681 45201 23684
rect 45235 23681 45247 23715
rect 45189 23675 45247 23681
rect 45462 23672 45468 23724
rect 45520 23672 45526 23724
rect 48774 23672 48780 23724
rect 48832 23672 48838 23724
rect 41230 23604 41236 23656
rect 41288 23644 41294 23656
rect 41325 23647 41383 23653
rect 41325 23644 41337 23647
rect 41288 23616 41337 23644
rect 41288 23604 41294 23616
rect 41325 23613 41337 23616
rect 41371 23613 41383 23647
rect 41325 23607 41383 23613
rect 43530 23604 43536 23656
rect 43588 23644 43594 23656
rect 44085 23647 44143 23653
rect 44085 23644 44097 23647
rect 43588 23616 44097 23644
rect 43588 23604 43594 23616
rect 44085 23613 44097 23616
rect 44131 23613 44143 23647
rect 44085 23607 44143 23613
rect 47029 23579 47087 23585
rect 47029 23576 47041 23579
rect 41156 23548 47041 23576
rect 39816 23536 39822 23548
rect 47029 23545 47041 23548
rect 47075 23545 47087 23579
rect 47029 23539 47087 23545
rect 38620 23480 39344 23508
rect 39485 23511 39543 23517
rect 38620 23468 38626 23480
rect 39485 23477 39497 23511
rect 39531 23508 39543 23511
rect 40494 23508 40500 23520
rect 39531 23480 40500 23508
rect 39531 23477 39543 23480
rect 39485 23471 39543 23477
rect 40494 23468 40500 23480
rect 40552 23468 40558 23520
rect 42794 23468 42800 23520
rect 42852 23508 42858 23520
rect 42981 23511 43039 23517
rect 42981 23508 42993 23511
rect 42852 23480 42993 23508
rect 42852 23468 42858 23480
rect 42981 23477 42993 23480
rect 43027 23477 43039 23511
rect 42981 23471 43039 23477
rect 47118 23468 47124 23520
rect 47176 23508 47182 23520
rect 48225 23511 48283 23517
rect 48225 23508 48237 23511
rect 47176 23480 48237 23508
rect 47176 23468 47182 23480
rect 48225 23477 48237 23480
rect 48271 23477 48283 23511
rect 48225 23471 48283 23477
rect 1104 23418 49864 23440
rect 1104 23366 2950 23418
rect 3002 23366 3014 23418
rect 3066 23366 3078 23418
rect 3130 23366 3142 23418
rect 3194 23366 3206 23418
rect 3258 23366 12950 23418
rect 13002 23366 13014 23418
rect 13066 23366 13078 23418
rect 13130 23366 13142 23418
rect 13194 23366 13206 23418
rect 13258 23366 22950 23418
rect 23002 23366 23014 23418
rect 23066 23366 23078 23418
rect 23130 23366 23142 23418
rect 23194 23366 23206 23418
rect 23258 23366 32950 23418
rect 33002 23366 33014 23418
rect 33066 23366 33078 23418
rect 33130 23366 33142 23418
rect 33194 23366 33206 23418
rect 33258 23366 42950 23418
rect 43002 23366 43014 23418
rect 43066 23366 43078 23418
rect 43130 23366 43142 23418
rect 43194 23366 43206 23418
rect 43258 23366 49864 23418
rect 1104 23344 49864 23366
rect 17586 23304 17592 23316
rect 10060 23276 17592 23304
rect 1578 23196 1584 23248
rect 1636 23236 1642 23248
rect 4338 23236 4344 23248
rect 1636 23208 4344 23236
rect 1636 23196 1642 23208
rect 4338 23196 4344 23208
rect 4396 23196 4402 23248
rect 7742 23196 7748 23248
rect 7800 23236 7806 23248
rect 9861 23239 9919 23245
rect 9861 23236 9873 23239
rect 7800 23208 9873 23236
rect 7800 23196 7806 23208
rect 9861 23205 9873 23208
rect 9907 23205 9919 23239
rect 9861 23199 9919 23205
rect 1780 23140 5488 23168
rect 1780 23109 1808 23140
rect 1765 23103 1823 23109
rect 1765 23069 1777 23103
rect 1811 23069 1823 23103
rect 1765 23063 1823 23069
rect 4249 23103 4307 23109
rect 4249 23069 4261 23103
rect 4295 23100 4307 23103
rect 4430 23100 4436 23112
rect 4295 23072 4436 23100
rect 4295 23069 4307 23072
rect 4249 23063 4307 23069
rect 4430 23060 4436 23072
rect 4488 23060 4494 23112
rect 4901 23103 4959 23109
rect 4901 23069 4913 23103
rect 4947 23100 4959 23103
rect 5258 23100 5264 23112
rect 4947 23072 5264 23100
rect 4947 23069 4959 23072
rect 4901 23063 4959 23069
rect 5258 23060 5264 23072
rect 5316 23060 5322 23112
rect 5353 23103 5411 23109
rect 5353 23069 5365 23103
rect 5399 23069 5411 23103
rect 5460 23100 5488 23140
rect 6086 23128 6092 23180
rect 6144 23128 6150 23180
rect 7834 23128 7840 23180
rect 7892 23128 7898 23180
rect 7098 23100 7104 23112
rect 5460 23072 7104 23100
rect 5353 23063 5411 23069
rect 2774 22992 2780 23044
rect 2832 22992 2838 23044
rect 2866 22992 2872 23044
rect 2924 23032 2930 23044
rect 4154 23032 4160 23044
rect 2924 23004 4160 23032
rect 2924 22992 2930 23004
rect 4154 22992 4160 23004
rect 4212 22992 4218 23044
rect 3602 22924 3608 22976
rect 3660 22964 3666 22976
rect 4065 22967 4123 22973
rect 4065 22964 4077 22967
rect 3660 22936 4077 22964
rect 3660 22924 3666 22936
rect 4065 22933 4077 22936
rect 4111 22933 4123 22967
rect 4065 22927 4123 22933
rect 4709 22967 4767 22973
rect 4709 22933 4721 22967
rect 4755 22964 4767 22967
rect 5368 22964 5396 23063
rect 7098 23060 7104 23072
rect 7156 23060 7162 23112
rect 7377 23103 7435 23109
rect 7377 23069 7389 23103
rect 7423 23100 7435 23103
rect 8294 23100 8300 23112
rect 7423 23072 8300 23100
rect 7423 23069 7435 23072
rect 7377 23063 7435 23069
rect 8294 23060 8300 23072
rect 8352 23060 8358 23112
rect 9122 23060 9128 23112
rect 9180 23100 9186 23112
rect 10060 23109 10088 23276
rect 17586 23264 17592 23276
rect 17644 23264 17650 23316
rect 17954 23264 17960 23316
rect 18012 23304 18018 23316
rect 19797 23307 19855 23313
rect 19797 23304 19809 23307
rect 18012 23276 19809 23304
rect 18012 23264 18018 23276
rect 19797 23273 19809 23276
rect 19843 23273 19855 23307
rect 22002 23304 22008 23316
rect 19797 23267 19855 23273
rect 19904 23276 22008 23304
rect 13814 23196 13820 23248
rect 13872 23236 13878 23248
rect 13872 23208 15884 23236
rect 13872 23196 13878 23208
rect 11238 23128 11244 23180
rect 11296 23128 11302 23180
rect 13354 23128 13360 23180
rect 13412 23128 13418 23180
rect 15746 23128 15752 23180
rect 15804 23128 15810 23180
rect 15856 23168 15884 23208
rect 19904 23168 19932 23276
rect 22002 23264 22008 23276
rect 22060 23264 22066 23316
rect 22186 23264 22192 23316
rect 22244 23304 22250 23316
rect 22649 23307 22707 23313
rect 22649 23304 22661 23307
rect 22244 23276 22661 23304
rect 22244 23264 22250 23276
rect 22649 23273 22661 23276
rect 22695 23273 22707 23307
rect 22649 23267 22707 23273
rect 22830 23264 22836 23316
rect 22888 23304 22894 23316
rect 23382 23304 23388 23316
rect 22888 23276 23388 23304
rect 22888 23264 22894 23276
rect 23382 23264 23388 23276
rect 23440 23264 23446 23316
rect 27798 23304 27804 23316
rect 23768 23276 27804 23304
rect 22094 23196 22100 23248
rect 22152 23236 22158 23248
rect 23290 23236 23296 23248
rect 22152 23208 23296 23236
rect 22152 23196 22158 23208
rect 23290 23196 23296 23208
rect 23348 23196 23354 23248
rect 15856 23140 19932 23168
rect 20346 23128 20352 23180
rect 20404 23168 20410 23180
rect 20714 23168 20720 23180
rect 20404 23140 20720 23168
rect 20404 23128 20410 23140
rect 20714 23128 20720 23140
rect 20772 23128 20778 23180
rect 22738 23168 22744 23180
rect 21744 23140 22744 23168
rect 9217 23103 9275 23109
rect 9217 23100 9229 23103
rect 9180 23072 9229 23100
rect 9180 23060 9186 23072
rect 9217 23069 9229 23072
rect 9263 23069 9275 23103
rect 9217 23063 9275 23069
rect 10045 23103 10103 23109
rect 10045 23069 10057 23103
rect 10091 23069 10103 23103
rect 10045 23063 10103 23069
rect 10686 23060 10692 23112
rect 10744 23060 10750 23112
rect 12529 23103 12587 23109
rect 12529 23069 12541 23103
rect 12575 23100 12587 23103
rect 14366 23100 14372 23112
rect 12575 23072 14372 23100
rect 12575 23069 12587 23072
rect 12529 23063 12587 23069
rect 14366 23060 14372 23072
rect 14424 23060 14430 23112
rect 14829 23103 14887 23109
rect 14829 23069 14841 23103
rect 14875 23100 14887 23103
rect 15102 23100 15108 23112
rect 14875 23072 15108 23100
rect 14875 23069 14887 23072
rect 14829 23063 14887 23069
rect 15102 23060 15108 23072
rect 15160 23060 15166 23112
rect 15473 23103 15531 23109
rect 15473 23069 15485 23103
rect 15519 23069 15531 23103
rect 15473 23063 15531 23069
rect 5442 22992 5448 23044
rect 5500 23032 5506 23044
rect 7650 23032 7656 23044
rect 5500 23004 7656 23032
rect 5500 22992 5506 23004
rect 7650 22992 7656 23004
rect 7708 22992 7714 23044
rect 15488 23032 15516 23063
rect 17034 23060 17040 23112
rect 17092 23100 17098 23112
rect 17129 23103 17187 23109
rect 17129 23100 17141 23103
rect 17092 23072 17141 23100
rect 17092 23060 17098 23072
rect 17129 23069 17141 23072
rect 17175 23069 17187 23103
rect 21744 23086 21772 23140
rect 22738 23128 22744 23140
rect 22796 23128 22802 23180
rect 23768 23177 23796 23276
rect 27798 23264 27804 23276
rect 27856 23264 27862 23316
rect 27890 23264 27896 23316
rect 27948 23264 27954 23316
rect 29730 23264 29736 23316
rect 29788 23264 29794 23316
rect 30558 23264 30564 23316
rect 30616 23304 30622 23316
rect 30616 23276 32904 23304
rect 30616 23264 30622 23276
rect 24857 23239 24915 23245
rect 24857 23205 24869 23239
rect 24903 23236 24915 23239
rect 25130 23236 25136 23248
rect 24903 23208 25136 23236
rect 24903 23205 24915 23208
rect 24857 23199 24915 23205
rect 25130 23196 25136 23208
rect 25188 23196 25194 23248
rect 30650 23236 30656 23248
rect 29932 23208 30656 23236
rect 23753 23171 23811 23177
rect 23753 23137 23765 23171
rect 23799 23137 23811 23171
rect 23753 23131 23811 23137
rect 23937 23171 23995 23177
rect 23937 23137 23949 23171
rect 23983 23168 23995 23171
rect 25961 23171 26019 23177
rect 25961 23168 25973 23171
rect 23983 23140 25973 23168
rect 23983 23137 23995 23140
rect 23937 23131 23995 23137
rect 25961 23137 25973 23140
rect 26007 23168 26019 23171
rect 26602 23168 26608 23180
rect 26007 23140 26608 23168
rect 26007 23137 26019 23140
rect 25961 23131 26019 23137
rect 26602 23128 26608 23140
rect 26660 23128 26666 23180
rect 26970 23128 26976 23180
rect 27028 23168 27034 23180
rect 28445 23171 28503 23177
rect 28445 23168 28457 23171
rect 27028 23140 28457 23168
rect 27028 23128 27034 23140
rect 28445 23137 28457 23140
rect 28491 23137 28503 23171
rect 28445 23131 28503 23137
rect 17129 23063 17187 23069
rect 21910 23060 21916 23112
rect 21968 23100 21974 23112
rect 22833 23103 22891 23109
rect 21968 23072 22784 23100
rect 21968 23060 21974 23072
rect 17310 23032 17316 23044
rect 15488 23004 17316 23032
rect 17310 22992 17316 23004
rect 17368 22992 17374 23044
rect 17405 23035 17463 23041
rect 17405 23001 17417 23035
rect 17451 23032 17463 23035
rect 17494 23032 17500 23044
rect 17451 23004 17500 23032
rect 17451 23001 17463 23004
rect 17405 22995 17463 23001
rect 17494 22992 17500 23004
rect 17552 22992 17558 23044
rect 18690 23032 18696 23044
rect 18630 23004 18696 23032
rect 18690 22992 18696 23004
rect 18748 22992 18754 23044
rect 19705 23035 19763 23041
rect 19705 23001 19717 23035
rect 19751 23001 19763 23035
rect 19705 22995 19763 23001
rect 4755 22936 5396 22964
rect 4755 22933 4767 22936
rect 4709 22927 4767 22933
rect 9306 22924 9312 22976
rect 9364 22924 9370 22976
rect 12802 22924 12808 22976
rect 12860 22964 12866 22976
rect 14645 22967 14703 22973
rect 14645 22964 14657 22967
rect 12860 22936 14657 22964
rect 12860 22924 12866 22936
rect 14645 22933 14657 22936
rect 14691 22933 14703 22967
rect 14645 22927 14703 22933
rect 18877 22967 18935 22973
rect 18877 22933 18889 22967
rect 18923 22964 18935 22967
rect 19058 22964 19064 22976
rect 18923 22936 19064 22964
rect 18923 22933 18935 22936
rect 18877 22927 18935 22933
rect 19058 22924 19064 22936
rect 19116 22924 19122 22976
rect 19720 22964 19748 22995
rect 20622 22992 20628 23044
rect 20680 22992 20686 23044
rect 22002 22992 22008 23044
rect 22060 23032 22066 23044
rect 22278 23032 22284 23044
rect 22060 23004 22284 23032
rect 22060 22992 22066 23004
rect 22278 22992 22284 23004
rect 22336 22992 22342 23044
rect 22756 23032 22784 23072
rect 22833 23069 22845 23103
rect 22879 23100 22891 23103
rect 24946 23100 24952 23112
rect 22879 23072 24952 23100
rect 22879 23069 22891 23072
rect 22833 23063 22891 23069
rect 24946 23060 24952 23072
rect 25004 23060 25010 23112
rect 25682 23060 25688 23112
rect 25740 23060 25746 23112
rect 28261 23103 28319 23109
rect 28261 23069 28273 23103
rect 28307 23100 28319 23103
rect 29932 23100 29960 23208
rect 30650 23196 30656 23208
rect 30708 23196 30714 23248
rect 30193 23171 30251 23177
rect 30193 23137 30205 23171
rect 30239 23168 30251 23171
rect 30282 23168 30288 23180
rect 30239 23140 30288 23168
rect 30239 23137 30251 23140
rect 30193 23131 30251 23137
rect 30282 23128 30288 23140
rect 30340 23128 30346 23180
rect 30377 23171 30435 23177
rect 30377 23137 30389 23171
rect 30423 23168 30435 23171
rect 31662 23168 31668 23180
rect 30423 23140 31668 23168
rect 30423 23137 30435 23140
rect 30377 23131 30435 23137
rect 31662 23128 31668 23140
rect 31720 23128 31726 23180
rect 28307 23072 29960 23100
rect 28307 23069 28319 23072
rect 28261 23063 28319 23069
rect 30006 23060 30012 23112
rect 30064 23100 30070 23112
rect 31389 23103 31447 23109
rect 31389 23100 31401 23103
rect 30064 23072 31401 23100
rect 30064 23060 30070 23072
rect 31389 23069 31401 23072
rect 31435 23069 31447 23103
rect 32876 23100 32904 23276
rect 33042 23264 33048 23316
rect 33100 23304 33106 23316
rect 33137 23307 33195 23313
rect 33137 23304 33149 23307
rect 33100 23276 33149 23304
rect 33100 23264 33106 23276
rect 33137 23273 33149 23276
rect 33183 23304 33195 23307
rect 34698 23304 34704 23316
rect 33183 23276 34704 23304
rect 33183 23273 33195 23276
rect 33137 23267 33195 23273
rect 34698 23264 34704 23276
rect 34756 23264 34762 23316
rect 35158 23264 35164 23316
rect 35216 23304 35222 23316
rect 38562 23304 38568 23316
rect 35216 23276 38568 23304
rect 35216 23264 35222 23276
rect 38562 23264 38568 23276
rect 38620 23264 38626 23316
rect 38654 23264 38660 23316
rect 38712 23304 38718 23316
rect 39025 23307 39083 23313
rect 39025 23304 39037 23307
rect 38712 23276 39037 23304
rect 38712 23264 38718 23276
rect 39025 23273 39037 23276
rect 39071 23273 39083 23307
rect 39025 23267 39083 23273
rect 40034 23264 40040 23316
rect 40092 23264 40098 23316
rect 40218 23264 40224 23316
rect 40276 23304 40282 23316
rect 41598 23304 41604 23316
rect 40276 23276 41604 23304
rect 40276 23264 40282 23276
rect 41598 23264 41604 23276
rect 41656 23264 41662 23316
rect 43346 23304 43352 23316
rect 41708 23276 43352 23304
rect 32950 23196 32956 23248
rect 33008 23236 33014 23248
rect 33689 23239 33747 23245
rect 33689 23236 33701 23239
rect 33008 23208 33701 23236
rect 33008 23196 33014 23208
rect 33689 23205 33701 23208
rect 33735 23205 33747 23239
rect 33689 23199 33747 23205
rect 38838 23196 38844 23248
rect 38896 23236 38902 23248
rect 41708 23236 41736 23276
rect 43346 23264 43352 23276
rect 43404 23264 43410 23316
rect 38896 23208 41736 23236
rect 47029 23239 47087 23245
rect 38896 23196 38902 23208
rect 47029 23205 47041 23239
rect 47075 23205 47087 23239
rect 47029 23199 47087 23205
rect 33318 23128 33324 23180
rect 33376 23168 33382 23180
rect 34606 23168 34612 23180
rect 33376 23140 34612 23168
rect 33376 23128 33382 23140
rect 34606 23128 34612 23140
rect 34664 23168 34670 23180
rect 35069 23171 35127 23177
rect 35069 23168 35081 23171
rect 34664 23140 35081 23168
rect 34664 23128 34670 23140
rect 35069 23137 35081 23140
rect 35115 23168 35127 23171
rect 35115 23140 38792 23168
rect 35115 23137 35127 23140
rect 35069 23131 35127 23137
rect 37292 23112 37320 23140
rect 33873 23103 33931 23109
rect 33873 23100 33885 23103
rect 32876 23072 33885 23100
rect 31389 23063 31447 23069
rect 33873 23069 33885 23072
rect 33919 23069 33931 23103
rect 33873 23063 33931 23069
rect 22756 23004 23796 23032
rect 21910 22964 21916 22976
rect 19720 22936 21916 22964
rect 21910 22924 21916 22936
rect 21968 22924 21974 22976
rect 22094 22924 22100 22976
rect 22152 22924 22158 22976
rect 22186 22924 22192 22976
rect 22244 22964 22250 22976
rect 23293 22967 23351 22973
rect 23293 22964 23305 22967
rect 22244 22936 23305 22964
rect 22244 22924 22250 22936
rect 23293 22933 23305 22936
rect 23339 22933 23351 22967
rect 23293 22927 23351 22933
rect 23658 22924 23664 22976
rect 23716 22924 23722 22976
rect 23768 22964 23796 23004
rect 24670 22992 24676 23044
rect 24728 22992 24734 23044
rect 25314 23032 25320 23044
rect 24780 23004 25320 23032
rect 24780 22964 24808 23004
rect 25314 22992 25320 23004
rect 25372 22992 25378 23044
rect 26418 22992 26424 23044
rect 26476 22992 26482 23044
rect 30834 23032 30840 23044
rect 27448 23004 30840 23032
rect 23768 22936 24808 22964
rect 25130 22924 25136 22976
rect 25188 22964 25194 22976
rect 27448 22973 27476 23004
rect 30834 22992 30840 23004
rect 30892 22992 30898 23044
rect 31404 23032 31432 23063
rect 37274 23060 37280 23112
rect 37332 23060 37338 23112
rect 38764 23100 38792 23140
rect 40586 23128 40592 23180
rect 40644 23128 40650 23180
rect 41877 23171 41935 23177
rect 41877 23137 41889 23171
rect 41923 23168 41935 23171
rect 47044 23168 47072 23199
rect 49234 23168 49240 23180
rect 41923 23140 47072 23168
rect 47228 23140 49240 23168
rect 41923 23137 41935 23140
rect 41877 23131 41935 23137
rect 41601 23103 41659 23109
rect 41601 23100 41613 23103
rect 38764 23072 41613 23100
rect 41601 23069 41613 23072
rect 41647 23069 41659 23103
rect 41601 23063 41659 23069
rect 43717 23103 43775 23109
rect 43717 23069 43729 23103
rect 43763 23069 43775 23103
rect 43717 23063 43775 23069
rect 31570 23032 31576 23044
rect 31404 23004 31576 23032
rect 31570 22992 31576 23004
rect 31628 22992 31634 23044
rect 32122 23032 32128 23044
rect 31680 23004 32128 23032
rect 27433 22967 27491 22973
rect 27433 22964 27445 22967
rect 25188 22936 27445 22964
rect 25188 22924 25194 22936
rect 27433 22933 27445 22936
rect 27479 22933 27491 22967
rect 27433 22927 27491 22933
rect 28350 22924 28356 22976
rect 28408 22924 28414 22976
rect 30098 22924 30104 22976
rect 30156 22924 30162 22976
rect 30742 22924 30748 22976
rect 30800 22964 30806 22976
rect 31202 22964 31208 22976
rect 30800 22936 31208 22964
rect 30800 22924 30806 22936
rect 31202 22924 31208 22936
rect 31260 22964 31266 22976
rect 31680 22964 31708 23004
rect 32122 22992 32128 23004
rect 32180 22992 32186 23044
rect 35342 22992 35348 23044
rect 35400 22992 35406 23044
rect 35802 22992 35808 23044
rect 35860 22992 35866 23044
rect 36722 22992 36728 23044
rect 36780 23032 36786 23044
rect 37182 23032 37188 23044
rect 36780 23004 37188 23032
rect 36780 22992 36786 23004
rect 37182 22992 37188 23004
rect 37240 23032 37246 23044
rect 37553 23035 37611 23041
rect 37553 23032 37565 23035
rect 37240 23004 37565 23032
rect 37240 22992 37246 23004
rect 37553 23001 37565 23004
rect 37599 23001 37611 23035
rect 38838 23032 38844 23044
rect 38778 23004 38844 23032
rect 37553 22995 37611 23001
rect 38838 22992 38844 23004
rect 38896 22992 38902 23044
rect 39574 22992 39580 23044
rect 39632 23032 39638 23044
rect 40310 23032 40316 23044
rect 39632 23004 40316 23032
rect 39632 22992 39638 23004
rect 40310 22992 40316 23004
rect 40368 22992 40374 23044
rect 40405 23035 40463 23041
rect 40405 23001 40417 23035
rect 40451 23032 40463 23035
rect 42150 23032 42156 23044
rect 40451 23004 42156 23032
rect 40451 23001 40463 23004
rect 40405 22995 40463 23001
rect 42150 22992 42156 23004
rect 42208 22992 42214 23044
rect 43346 23032 43352 23044
rect 43102 23004 43352 23032
rect 43346 22992 43352 23004
rect 43404 22992 43410 23044
rect 43622 22992 43628 23044
rect 43680 22992 43686 23044
rect 31260 22936 31708 22964
rect 31260 22924 31266 22936
rect 31754 22924 31760 22976
rect 31812 22964 31818 22976
rect 33042 22964 33048 22976
rect 31812 22936 33048 22964
rect 31812 22924 31818 22936
rect 33042 22924 33048 22936
rect 33100 22924 33106 22976
rect 33318 22924 33324 22976
rect 33376 22964 33382 22976
rect 35066 22964 35072 22976
rect 33376 22936 35072 22964
rect 33376 22924 33382 22936
rect 35066 22924 35072 22936
rect 35124 22924 35130 22976
rect 35158 22924 35164 22976
rect 35216 22964 35222 22976
rect 36817 22967 36875 22973
rect 36817 22964 36829 22967
rect 35216 22936 36829 22964
rect 35216 22924 35222 22936
rect 36817 22933 36829 22936
rect 36863 22964 36875 22967
rect 38562 22964 38568 22976
rect 36863 22936 38568 22964
rect 36863 22933 36875 22936
rect 36817 22927 36875 22933
rect 38562 22924 38568 22936
rect 38620 22924 38626 22976
rect 40218 22924 40224 22976
rect 40276 22964 40282 22976
rect 40497 22967 40555 22973
rect 40497 22964 40509 22967
rect 40276 22936 40509 22964
rect 40276 22924 40282 22936
rect 40497 22933 40509 22936
rect 40543 22964 40555 22967
rect 41414 22964 41420 22976
rect 40543 22936 41420 22964
rect 40543 22933 40555 22936
rect 40497 22927 40555 22933
rect 41414 22924 41420 22936
rect 41472 22924 41478 22976
rect 41598 22924 41604 22976
rect 41656 22964 41662 22976
rect 42610 22964 42616 22976
rect 41656 22936 42616 22964
rect 41656 22924 41662 22936
rect 42610 22924 42616 22936
rect 42668 22924 42674 22976
rect 42794 22924 42800 22976
rect 42852 22964 42858 22976
rect 43732 22964 43760 23063
rect 43990 23060 43996 23112
rect 44048 23060 44054 23112
rect 44082 23060 44088 23112
rect 44140 23100 44146 23112
rect 45097 23103 45155 23109
rect 45097 23100 45109 23103
rect 44140 23072 45109 23100
rect 44140 23060 44146 23072
rect 45097 23069 45109 23072
rect 45143 23069 45155 23103
rect 45097 23063 45155 23069
rect 45557 23103 45615 23109
rect 45557 23069 45569 23103
rect 45603 23069 45615 23103
rect 45557 23063 45615 23069
rect 43806 22992 43812 23044
rect 43864 23032 43870 23044
rect 45572 23032 45600 23063
rect 46290 23060 46296 23112
rect 46348 23060 46354 23112
rect 47228 23109 47256 23140
rect 49234 23128 49240 23140
rect 49292 23128 49298 23180
rect 47213 23103 47271 23109
rect 47213 23069 47225 23103
rect 47259 23069 47271 23103
rect 47213 23063 47271 23069
rect 47854 23060 47860 23112
rect 47912 23060 47918 23112
rect 48314 23060 48320 23112
rect 48372 23060 48378 23112
rect 49053 23103 49111 23109
rect 49053 23069 49065 23103
rect 49099 23100 49111 23103
rect 49142 23100 49148 23112
rect 49099 23072 49148 23100
rect 49099 23069 49111 23072
rect 49053 23063 49111 23069
rect 49142 23060 49148 23072
rect 49200 23060 49206 23112
rect 43864 23004 45600 23032
rect 43864 22992 43870 23004
rect 46842 22992 46848 23044
rect 46900 23032 46906 23044
rect 46900 23004 49280 23032
rect 46900 22992 46906 23004
rect 42852 22936 43760 22964
rect 42852 22924 42858 22936
rect 45186 22924 45192 22976
rect 45244 22924 45250 22976
rect 45370 22924 45376 22976
rect 45428 22924 45434 22976
rect 45462 22924 45468 22976
rect 45520 22964 45526 22976
rect 46109 22967 46167 22973
rect 46109 22964 46121 22967
rect 45520 22936 46121 22964
rect 45520 22924 45526 22936
rect 46109 22933 46121 22936
rect 46155 22933 46167 22967
rect 46109 22927 46167 22933
rect 47670 22924 47676 22976
rect 47728 22924 47734 22976
rect 48498 22924 48504 22976
rect 48556 22924 48562 22976
rect 49252 22973 49280 23004
rect 49237 22967 49295 22973
rect 49237 22933 49249 22967
rect 49283 22933 49295 22967
rect 49237 22927 49295 22933
rect 1104 22874 49864 22896
rect 1104 22822 7950 22874
rect 8002 22822 8014 22874
rect 8066 22822 8078 22874
rect 8130 22822 8142 22874
rect 8194 22822 8206 22874
rect 8258 22822 17950 22874
rect 18002 22822 18014 22874
rect 18066 22822 18078 22874
rect 18130 22822 18142 22874
rect 18194 22822 18206 22874
rect 18258 22822 27950 22874
rect 28002 22822 28014 22874
rect 28066 22822 28078 22874
rect 28130 22822 28142 22874
rect 28194 22822 28206 22874
rect 28258 22822 37950 22874
rect 38002 22822 38014 22874
rect 38066 22822 38078 22874
rect 38130 22822 38142 22874
rect 38194 22822 38206 22874
rect 38258 22822 47950 22874
rect 48002 22822 48014 22874
rect 48066 22822 48078 22874
rect 48130 22822 48142 22874
rect 48194 22822 48206 22874
rect 48258 22822 49864 22874
rect 1104 22800 49864 22822
rect 3326 22720 3332 22772
rect 3384 22760 3390 22772
rect 6730 22760 6736 22772
rect 3384 22732 6736 22760
rect 3384 22720 3390 22732
rect 6730 22720 6736 22732
rect 6788 22720 6794 22772
rect 13354 22760 13360 22772
rect 6886 22732 13360 22760
rect 2777 22695 2835 22701
rect 2777 22661 2789 22695
rect 2823 22692 2835 22695
rect 2866 22692 2872 22704
rect 2823 22664 2872 22692
rect 2823 22661 2835 22664
rect 2777 22655 2835 22661
rect 2866 22652 2872 22664
rect 2924 22652 2930 22704
rect 3973 22695 4031 22701
rect 3973 22661 3985 22695
rect 4019 22692 4031 22695
rect 6886 22692 6914 22732
rect 13354 22720 13360 22732
rect 13412 22720 13418 22772
rect 17402 22760 17408 22772
rect 15120 22732 17408 22760
rect 7558 22692 7564 22704
rect 4019 22664 5764 22692
rect 4019 22661 4031 22664
rect 3973 22655 4031 22661
rect 1765 22627 1823 22633
rect 1765 22593 1777 22627
rect 1811 22624 1823 22627
rect 1811 22596 2820 22624
rect 1811 22593 1823 22596
rect 1765 22587 1823 22593
rect 2792 22488 2820 22596
rect 4798 22584 4804 22636
rect 4856 22584 4862 22636
rect 5074 22516 5080 22568
rect 5132 22516 5138 22568
rect 5736 22556 5764 22664
rect 6840 22664 6914 22692
rect 7300 22664 7564 22692
rect 6840 22633 6868 22664
rect 6825 22627 6883 22633
rect 6825 22593 6837 22627
rect 6871 22593 6883 22627
rect 6825 22587 6883 22593
rect 7300 22556 7328 22664
rect 7558 22652 7564 22664
rect 7616 22652 7622 22704
rect 7466 22584 7472 22636
rect 7524 22584 7530 22636
rect 9953 22627 10011 22633
rect 9953 22593 9965 22627
rect 9999 22593 10011 22627
rect 9953 22587 10011 22593
rect 12161 22627 12219 22633
rect 12161 22593 12173 22627
rect 12207 22593 12219 22627
rect 12161 22587 12219 22593
rect 5736 22528 7328 22556
rect 7374 22516 7380 22568
rect 7432 22556 7438 22568
rect 7929 22559 7987 22565
rect 7929 22556 7941 22559
rect 7432 22528 7941 22556
rect 7432 22516 7438 22528
rect 7929 22525 7941 22528
rect 7975 22525 7987 22559
rect 7929 22519 7987 22525
rect 9968 22488 9996 22587
rect 10042 22516 10048 22568
rect 10100 22556 10106 22568
rect 10229 22559 10287 22565
rect 10229 22556 10241 22559
rect 10100 22528 10241 22556
rect 10100 22516 10106 22528
rect 10229 22525 10241 22528
rect 10275 22525 10287 22559
rect 10229 22519 10287 22525
rect 11977 22491 12035 22497
rect 11977 22488 11989 22491
rect 2792 22460 9904 22488
rect 9968 22460 11989 22488
rect 4065 22423 4123 22429
rect 4065 22389 4077 22423
rect 4111 22420 4123 22423
rect 6454 22420 6460 22432
rect 4111 22392 6460 22420
rect 4111 22389 4123 22392
rect 4065 22383 4123 22389
rect 6454 22380 6460 22392
rect 6512 22380 6518 22432
rect 6641 22423 6699 22429
rect 6641 22389 6653 22423
rect 6687 22420 6699 22423
rect 9122 22420 9128 22432
rect 6687 22392 9128 22420
rect 6687 22389 6699 22392
rect 6641 22383 6699 22389
rect 9122 22380 9128 22392
rect 9180 22380 9186 22432
rect 9876 22420 9904 22460
rect 11977 22457 11989 22460
rect 12023 22457 12035 22491
rect 12176 22488 12204 22587
rect 12802 22584 12808 22636
rect 12860 22584 12866 22636
rect 15120 22633 15148 22732
rect 17402 22720 17408 22732
rect 17460 22720 17466 22772
rect 20622 22720 20628 22772
rect 20680 22760 20686 22772
rect 21177 22763 21235 22769
rect 21177 22760 21189 22763
rect 20680 22732 21189 22760
rect 20680 22720 20686 22732
rect 21177 22729 21189 22732
rect 21223 22760 21235 22763
rect 22646 22760 22652 22772
rect 21223 22732 22652 22760
rect 21223 22729 21235 22732
rect 21177 22723 21235 22729
rect 22646 22720 22652 22732
rect 22704 22760 22710 22772
rect 24762 22760 24768 22772
rect 22704 22732 24768 22760
rect 22704 22720 22710 22732
rect 24762 22720 24768 22732
rect 24820 22720 24826 22772
rect 24854 22720 24860 22772
rect 24912 22760 24918 22772
rect 30006 22760 30012 22772
rect 24912 22732 30012 22760
rect 24912 22720 24918 22732
rect 17034 22692 17040 22704
rect 16868 22664 17040 22692
rect 16868 22633 16896 22664
rect 17034 22652 17040 22664
rect 17092 22652 17098 22704
rect 18690 22692 18696 22704
rect 18354 22664 18696 22692
rect 18690 22652 18696 22664
rect 18748 22652 18754 22704
rect 18874 22652 18880 22704
rect 18932 22692 18938 22704
rect 19705 22695 19763 22701
rect 19705 22692 19717 22695
rect 18932 22664 19717 22692
rect 18932 22652 18938 22664
rect 19705 22661 19717 22664
rect 19751 22661 19763 22695
rect 19705 22655 19763 22661
rect 20162 22652 20168 22704
rect 20220 22652 20226 22704
rect 22278 22652 22284 22704
rect 22336 22652 22342 22704
rect 22738 22652 22744 22704
rect 22796 22652 22802 22704
rect 25038 22692 25044 22704
rect 23584 22664 25044 22692
rect 15105 22627 15163 22633
rect 15105 22593 15117 22627
rect 15151 22593 15163 22627
rect 15105 22587 15163 22593
rect 16853 22627 16911 22633
rect 16853 22593 16865 22627
rect 16899 22593 16911 22627
rect 23584 22624 23612 22664
rect 25038 22652 25044 22664
rect 25096 22652 25102 22704
rect 25130 22652 25136 22704
rect 25188 22652 25194 22704
rect 26418 22692 26424 22704
rect 26358 22664 26424 22692
rect 26418 22652 26424 22664
rect 26476 22692 26482 22704
rect 27430 22692 27436 22704
rect 26476 22664 27436 22692
rect 26476 22652 26482 22664
rect 27430 22652 27436 22664
rect 27488 22652 27494 22704
rect 27614 22652 27620 22704
rect 27672 22692 27678 22704
rect 27890 22692 27896 22704
rect 27672 22664 27896 22692
rect 27672 22652 27678 22664
rect 27890 22652 27896 22664
rect 27948 22652 27954 22704
rect 16853 22587 16911 22593
rect 23492 22596 23612 22624
rect 12526 22516 12532 22568
rect 12584 22556 12590 22568
rect 13081 22559 13139 22565
rect 13081 22556 13093 22559
rect 12584 22528 13093 22556
rect 12584 22516 12590 22528
rect 13081 22525 13093 22528
rect 13127 22525 13139 22559
rect 13081 22519 13139 22525
rect 15010 22516 15016 22568
rect 15068 22556 15074 22568
rect 15381 22559 15439 22565
rect 15381 22556 15393 22559
rect 15068 22528 15393 22556
rect 15068 22516 15074 22528
rect 15381 22525 15393 22528
rect 15427 22525 15439 22559
rect 15381 22519 15439 22525
rect 17126 22516 17132 22568
rect 17184 22516 17190 22568
rect 18598 22516 18604 22568
rect 18656 22556 18662 22568
rect 19429 22559 19487 22565
rect 19429 22556 19441 22559
rect 18656 22528 19441 22556
rect 18656 22516 18662 22528
rect 19429 22525 19441 22528
rect 19475 22525 19487 22559
rect 19429 22519 19487 22525
rect 22002 22516 22008 22568
rect 22060 22516 22066 22568
rect 14734 22488 14740 22500
rect 12176 22460 14740 22488
rect 11977 22451 12035 22457
rect 14734 22448 14740 22460
rect 14792 22448 14798 22500
rect 15654 22420 15660 22432
rect 9876 22392 15660 22420
rect 15654 22380 15660 22392
rect 15712 22380 15718 22432
rect 17494 22380 17500 22432
rect 17552 22420 17558 22432
rect 18601 22423 18659 22429
rect 18601 22420 18613 22423
rect 17552 22392 18613 22420
rect 17552 22380 17558 22392
rect 18601 22389 18613 22392
rect 18647 22420 18659 22423
rect 23492 22420 23520 22596
rect 24854 22584 24860 22636
rect 24912 22584 24918 22636
rect 27338 22584 27344 22636
rect 27396 22584 27402 22636
rect 28092 22633 28120 22732
rect 30006 22720 30012 22732
rect 30064 22720 30070 22772
rect 30653 22763 30711 22769
rect 30653 22729 30665 22763
rect 30699 22760 30711 22763
rect 30699 22732 32444 22760
rect 30699 22729 30711 22732
rect 30653 22723 30711 22729
rect 30742 22692 30748 22704
rect 29578 22664 30748 22692
rect 30742 22652 30748 22664
rect 30800 22652 30806 22704
rect 32416 22692 32444 22732
rect 32490 22720 32496 22772
rect 32548 22760 32554 22772
rect 35897 22763 35955 22769
rect 32548 22732 35848 22760
rect 32548 22720 32554 22732
rect 32582 22692 32588 22704
rect 32416 22664 32588 22692
rect 32582 22652 32588 22664
rect 32640 22652 32646 22704
rect 32677 22695 32735 22701
rect 32677 22661 32689 22695
rect 32723 22692 32735 22695
rect 33318 22692 33324 22704
rect 32723 22664 33324 22692
rect 32723 22661 32735 22664
rect 32677 22655 32735 22661
rect 33318 22652 33324 22664
rect 33376 22652 33382 22704
rect 33686 22652 33692 22704
rect 33744 22692 33750 22704
rect 35820 22692 35848 22732
rect 35897 22729 35909 22763
rect 35943 22760 35955 22763
rect 36354 22760 36360 22772
rect 35943 22732 36360 22760
rect 35943 22729 35955 22732
rect 35897 22723 35955 22729
rect 36354 22720 36360 22732
rect 36412 22720 36418 22772
rect 37182 22720 37188 22772
rect 37240 22760 37246 22772
rect 39209 22763 39267 22769
rect 39209 22760 39221 22763
rect 37240 22732 39221 22760
rect 37240 22720 37246 22732
rect 39209 22729 39221 22732
rect 39255 22729 39267 22763
rect 39209 22723 39267 22729
rect 37734 22692 37740 22704
rect 33744 22664 33902 22692
rect 35820 22664 37740 22692
rect 33744 22652 33750 22664
rect 37734 22652 37740 22664
rect 37792 22652 37798 22704
rect 28077 22627 28135 22633
rect 28077 22593 28089 22627
rect 28123 22593 28135 22627
rect 28077 22587 28135 22593
rect 29564 22596 30972 22624
rect 23658 22516 23664 22568
rect 23716 22556 23722 22568
rect 27614 22556 27620 22568
rect 23716 22528 27620 22556
rect 23716 22516 23722 22528
rect 27614 22516 27620 22528
rect 27672 22516 27678 22568
rect 28353 22559 28411 22565
rect 28353 22525 28365 22559
rect 28399 22556 28411 22559
rect 28994 22556 29000 22568
rect 28399 22528 29000 22556
rect 28399 22525 28411 22528
rect 28353 22519 28411 22525
rect 28994 22516 29000 22528
rect 29052 22556 29058 22568
rect 29564 22556 29592 22596
rect 29052 22528 29592 22556
rect 29052 22516 29058 22528
rect 30742 22516 30748 22568
rect 30800 22516 30806 22568
rect 30834 22516 30840 22568
rect 30892 22516 30898 22568
rect 30944 22556 30972 22596
rect 31662 22584 31668 22636
rect 31720 22584 31726 22636
rect 32769 22627 32827 22633
rect 32769 22593 32781 22627
rect 32815 22624 32827 22627
rect 32815 22596 32996 22624
rect 32815 22593 32827 22596
rect 32769 22587 32827 22593
rect 32861 22559 32919 22565
rect 30944 22528 32444 22556
rect 26142 22448 26148 22500
rect 26200 22488 26206 22500
rect 26970 22488 26976 22500
rect 26200 22460 26976 22488
rect 26200 22448 26206 22460
rect 26970 22448 26976 22460
rect 27028 22448 27034 22500
rect 27154 22448 27160 22500
rect 27212 22448 27218 22500
rect 30374 22448 30380 22500
rect 30432 22488 30438 22500
rect 32309 22491 32367 22497
rect 32309 22488 32321 22491
rect 30432 22460 32321 22488
rect 30432 22448 30438 22460
rect 32309 22457 32321 22460
rect 32355 22457 32367 22491
rect 32416 22488 32444 22528
rect 32861 22525 32873 22559
rect 32907 22525 32919 22559
rect 32861 22519 32919 22525
rect 32876 22488 32904 22519
rect 32416 22460 32904 22488
rect 32309 22451 32367 22457
rect 18647 22392 23520 22420
rect 18647 22389 18659 22392
rect 18601 22383 18659 22389
rect 23658 22380 23664 22432
rect 23716 22420 23722 22432
rect 23753 22423 23811 22429
rect 23753 22420 23765 22423
rect 23716 22392 23765 22420
rect 23716 22380 23722 22392
rect 23753 22389 23765 22392
rect 23799 22389 23811 22423
rect 23753 22383 23811 22389
rect 26602 22380 26608 22432
rect 26660 22380 26666 22432
rect 28902 22380 28908 22432
rect 28960 22420 28966 22432
rect 29825 22423 29883 22429
rect 29825 22420 29837 22423
rect 28960 22392 29837 22420
rect 28960 22380 28966 22392
rect 29825 22389 29837 22392
rect 29871 22389 29883 22423
rect 29825 22383 29883 22389
rect 30282 22380 30288 22432
rect 30340 22380 30346 22432
rect 31478 22380 31484 22432
rect 31536 22380 31542 22432
rect 32968 22420 32996 22596
rect 33134 22584 33140 22636
rect 33192 22584 33198 22636
rect 35437 22627 35495 22633
rect 35437 22593 35449 22627
rect 35483 22624 35495 22627
rect 36078 22624 36084 22636
rect 35483 22596 36084 22624
rect 35483 22593 35495 22596
rect 35437 22587 35495 22593
rect 36078 22584 36084 22596
rect 36136 22624 36142 22636
rect 36265 22627 36323 22633
rect 36265 22624 36277 22627
rect 36136 22596 36277 22624
rect 36136 22584 36142 22596
rect 36265 22593 36277 22596
rect 36311 22593 36323 22627
rect 36265 22587 36323 22593
rect 38838 22584 38844 22636
rect 38896 22584 38902 22636
rect 33042 22516 33048 22568
rect 33100 22556 33106 22568
rect 33413 22559 33471 22565
rect 33413 22556 33425 22559
rect 33100 22528 33425 22556
rect 33100 22516 33106 22528
rect 33413 22525 33425 22528
rect 33459 22525 33471 22559
rect 33413 22519 33471 22525
rect 33870 22516 33876 22568
rect 33928 22556 33934 22568
rect 34885 22559 34943 22565
rect 34885 22556 34897 22559
rect 33928 22528 34897 22556
rect 33928 22516 33934 22528
rect 34885 22525 34897 22528
rect 34931 22556 34943 22559
rect 35250 22556 35256 22568
rect 34931 22528 35256 22556
rect 34931 22525 34943 22528
rect 34885 22519 34943 22525
rect 35250 22516 35256 22528
rect 35308 22516 35314 22568
rect 36170 22516 36176 22568
rect 36228 22556 36234 22568
rect 36357 22559 36415 22565
rect 36357 22556 36369 22559
rect 36228 22528 36369 22556
rect 36228 22516 36234 22528
rect 36357 22525 36369 22528
rect 36403 22525 36415 22559
rect 36357 22519 36415 22525
rect 36446 22516 36452 22568
rect 36504 22516 36510 22568
rect 37274 22516 37280 22568
rect 37332 22556 37338 22568
rect 37461 22559 37519 22565
rect 37461 22556 37473 22559
rect 37332 22528 37473 22556
rect 37332 22516 37338 22528
rect 37461 22525 37473 22528
rect 37507 22525 37519 22559
rect 37461 22519 37519 22525
rect 37734 22516 37740 22568
rect 37792 22516 37798 22568
rect 39224 22556 39252 22723
rect 39666 22720 39672 22772
rect 39724 22720 39730 22772
rect 40126 22720 40132 22772
rect 40184 22720 40190 22772
rect 40865 22763 40923 22769
rect 40865 22729 40877 22763
rect 40911 22760 40923 22763
rect 47029 22763 47087 22769
rect 47029 22760 47041 22763
rect 40911 22732 47041 22760
rect 40911 22729 40923 22732
rect 40865 22723 40923 22729
rect 47029 22729 47041 22732
rect 47075 22729 47087 22763
rect 47029 22723 47087 22729
rect 48501 22763 48559 22769
rect 48501 22729 48513 22763
rect 48547 22760 48559 22763
rect 48682 22760 48688 22772
rect 48547 22732 48688 22760
rect 48547 22729 48559 22732
rect 48501 22723 48559 22729
rect 48682 22720 48688 22732
rect 48740 22720 48746 22772
rect 40310 22652 40316 22704
rect 40368 22692 40374 22704
rect 40368 22664 44956 22692
rect 40368 22652 40374 22664
rect 40034 22584 40040 22636
rect 40092 22584 40098 22636
rect 41506 22584 41512 22636
rect 41564 22584 41570 22636
rect 41782 22584 41788 22636
rect 41840 22584 41846 22636
rect 41874 22584 41880 22636
rect 41932 22624 41938 22636
rect 42797 22627 42855 22633
rect 42797 22624 42809 22627
rect 41932 22596 42809 22624
rect 41932 22584 41938 22596
rect 42797 22593 42809 22596
rect 42843 22593 42855 22627
rect 42797 22587 42855 22593
rect 43257 22627 43315 22633
rect 43257 22593 43269 22627
rect 43303 22624 43315 22627
rect 43438 22624 43444 22636
rect 43303 22596 43444 22624
rect 43303 22593 43315 22596
rect 43257 22587 43315 22593
rect 43438 22584 43444 22596
rect 43496 22624 43502 22636
rect 44928 22633 44956 22664
rect 44545 22627 44603 22633
rect 44545 22624 44557 22627
rect 43496 22596 44557 22624
rect 43496 22584 43502 22596
rect 44545 22593 44557 22596
rect 44591 22593 44603 22627
rect 44545 22587 44603 22593
rect 44913 22627 44971 22633
rect 44913 22593 44925 22627
rect 44959 22593 44971 22627
rect 44913 22587 44971 22593
rect 46750 22584 46756 22636
rect 46808 22624 46814 22636
rect 47213 22627 47271 22633
rect 47213 22624 47225 22627
rect 46808 22596 47225 22624
rect 46808 22584 46814 22596
rect 47213 22593 47225 22596
rect 47259 22593 47271 22627
rect 47213 22587 47271 22593
rect 48317 22627 48375 22633
rect 48317 22593 48329 22627
rect 48363 22624 48375 22627
rect 48406 22624 48412 22636
rect 48363 22596 48412 22624
rect 48363 22593 48375 22596
rect 48317 22587 48375 22593
rect 48406 22584 48412 22596
rect 48464 22584 48470 22636
rect 49050 22584 49056 22636
rect 49108 22584 49114 22636
rect 40221 22559 40279 22565
rect 40221 22556 40233 22559
rect 39224 22528 40233 22556
rect 40221 22525 40233 22528
rect 40267 22525 40279 22559
rect 40221 22519 40279 22525
rect 40954 22516 40960 22568
rect 41012 22516 41018 22568
rect 41046 22516 41052 22568
rect 41104 22516 41110 22568
rect 43530 22516 43536 22568
rect 43588 22516 43594 22568
rect 39022 22488 39028 22500
rect 38856 22460 39028 22488
rect 35250 22420 35256 22432
rect 32968 22392 35256 22420
rect 35250 22380 35256 22392
rect 35308 22380 35314 22432
rect 36998 22380 37004 22432
rect 37056 22420 37062 22432
rect 38856 22420 38884 22460
rect 39022 22448 39028 22460
rect 39080 22448 39086 22500
rect 39114 22448 39120 22500
rect 39172 22488 39178 22500
rect 40497 22491 40555 22497
rect 40497 22488 40509 22491
rect 39172 22460 40509 22488
rect 39172 22448 39178 22460
rect 40497 22457 40509 22460
rect 40543 22457 40555 22491
rect 40497 22451 40555 22457
rect 47302 22448 47308 22500
rect 47360 22488 47366 22500
rect 49237 22491 49295 22497
rect 49237 22488 49249 22491
rect 47360 22460 49249 22488
rect 47360 22448 47366 22460
rect 49237 22457 49249 22460
rect 49283 22457 49295 22491
rect 49237 22451 49295 22457
rect 37056 22392 38884 22420
rect 37056 22380 37062 22392
rect 41322 22380 41328 22432
rect 41380 22380 41386 22432
rect 41598 22380 41604 22432
rect 41656 22380 41662 22432
rect 41690 22380 41696 22432
rect 41748 22420 41754 22432
rect 42613 22423 42671 22429
rect 42613 22420 42625 22423
rect 41748 22392 42625 22420
rect 41748 22380 41754 22392
rect 42613 22389 42625 22392
rect 42659 22389 42671 22423
rect 42613 22383 42671 22389
rect 44726 22380 44732 22432
rect 44784 22380 44790 22432
rect 1104 22330 49864 22352
rect 1104 22278 2950 22330
rect 3002 22278 3014 22330
rect 3066 22278 3078 22330
rect 3130 22278 3142 22330
rect 3194 22278 3206 22330
rect 3258 22278 12950 22330
rect 13002 22278 13014 22330
rect 13066 22278 13078 22330
rect 13130 22278 13142 22330
rect 13194 22278 13206 22330
rect 13258 22278 22950 22330
rect 23002 22278 23014 22330
rect 23066 22278 23078 22330
rect 23130 22278 23142 22330
rect 23194 22278 23206 22330
rect 23258 22278 32950 22330
rect 33002 22278 33014 22330
rect 33066 22278 33078 22330
rect 33130 22278 33142 22330
rect 33194 22278 33206 22330
rect 33258 22278 42950 22330
rect 43002 22278 43014 22330
rect 43066 22278 43078 22330
rect 43130 22278 43142 22330
rect 43194 22278 43206 22330
rect 43258 22278 49864 22330
rect 1104 22256 49864 22278
rect 2222 22176 2228 22228
rect 2280 22216 2286 22228
rect 4890 22216 4896 22228
rect 2280 22188 4896 22216
rect 2280 22176 2286 22188
rect 4890 22176 4896 22188
rect 4948 22176 4954 22228
rect 7098 22176 7104 22228
rect 7156 22216 7162 22228
rect 7837 22219 7895 22225
rect 7837 22216 7849 22219
rect 7156 22188 7849 22216
rect 7156 22176 7162 22188
rect 7837 22185 7849 22188
rect 7883 22185 7895 22219
rect 7837 22179 7895 22185
rect 16945 22219 17003 22225
rect 16945 22185 16957 22219
rect 16991 22216 17003 22219
rect 17126 22216 17132 22228
rect 16991 22188 17132 22216
rect 16991 22185 17003 22188
rect 16945 22179 17003 22185
rect 17126 22176 17132 22188
rect 17184 22176 17190 22228
rect 17402 22176 17408 22228
rect 17460 22216 17466 22228
rect 20990 22216 20996 22228
rect 17460 22188 20996 22216
rect 17460 22176 17466 22188
rect 20990 22176 20996 22188
rect 21048 22176 21054 22228
rect 22370 22176 22376 22228
rect 22428 22216 22434 22228
rect 23198 22216 23204 22228
rect 22428 22188 23204 22216
rect 22428 22176 22434 22188
rect 23198 22176 23204 22188
rect 23256 22216 23262 22228
rect 23256 22188 26556 22216
rect 23256 22176 23262 22188
rect 3418 22108 3424 22160
rect 3476 22148 3482 22160
rect 3476 22120 5672 22148
rect 3476 22108 3482 22120
rect 1302 22040 1308 22092
rect 1360 22080 1366 22092
rect 2041 22083 2099 22089
rect 2041 22080 2053 22083
rect 1360 22052 2053 22080
rect 1360 22040 1366 22052
rect 2041 22049 2053 22052
rect 2087 22049 2099 22083
rect 2041 22043 2099 22049
rect 3786 22040 3792 22092
rect 3844 22080 3850 22092
rect 4433 22083 4491 22089
rect 4433 22080 4445 22083
rect 3844 22052 4445 22080
rect 3844 22040 3850 22052
rect 4433 22049 4445 22052
rect 4479 22049 4491 22083
rect 5644 22080 5672 22120
rect 10502 22108 10508 22160
rect 10560 22148 10566 22160
rect 13722 22148 13728 22160
rect 10560 22120 13728 22148
rect 10560 22108 10566 22120
rect 13722 22108 13728 22120
rect 13780 22108 13786 22160
rect 17218 22108 17224 22160
rect 17276 22148 17282 22160
rect 17276 22120 18000 22148
rect 17276 22108 17282 22120
rect 6273 22083 6331 22089
rect 6273 22080 6285 22083
rect 5644 22052 6285 22080
rect 4433 22043 4491 22049
rect 6273 22049 6285 22052
rect 6319 22049 6331 22083
rect 6273 22043 6331 22049
rect 9214 22040 9220 22092
rect 9272 22080 9278 22092
rect 9585 22083 9643 22089
rect 9585 22080 9597 22083
rect 9272 22052 9597 22080
rect 9272 22040 9278 22052
rect 9585 22049 9597 22052
rect 9631 22049 9643 22083
rect 9585 22043 9643 22049
rect 11333 22083 11391 22089
rect 11333 22049 11345 22083
rect 11379 22080 11391 22083
rect 11793 22083 11851 22089
rect 11793 22080 11805 22083
rect 11379 22052 11805 22080
rect 11379 22049 11391 22052
rect 11333 22043 11391 22049
rect 11793 22049 11805 22052
rect 11839 22080 11851 22083
rect 13814 22080 13820 22092
rect 11839 22052 13820 22080
rect 11839 22049 11851 22052
rect 11793 22043 11851 22049
rect 13814 22040 13820 22052
rect 13872 22040 13878 22092
rect 17972 22089 18000 22120
rect 18966 22108 18972 22160
rect 19024 22148 19030 22160
rect 19024 22120 19932 22148
rect 19024 22108 19030 22120
rect 19904 22089 19932 22120
rect 21726 22108 21732 22160
rect 21784 22148 21790 22160
rect 21784 22120 22048 22148
rect 21784 22108 21790 22120
rect 22020 22089 22048 22120
rect 23124 22120 23336 22148
rect 17957 22083 18015 22089
rect 17957 22049 17969 22083
rect 18003 22049 18015 22083
rect 17957 22043 18015 22049
rect 19889 22083 19947 22089
rect 19889 22049 19901 22083
rect 19935 22049 19947 22083
rect 19889 22043 19947 22049
rect 22005 22083 22063 22089
rect 22005 22049 22017 22083
rect 22051 22049 22063 22083
rect 22005 22043 22063 22049
rect 1765 22015 1823 22021
rect 1765 21981 1777 22015
rect 1811 21981 1823 22015
rect 1765 21975 1823 21981
rect 1780 21876 1808 21975
rect 4062 21972 4068 22024
rect 4120 21972 4126 22024
rect 5994 21972 6000 22024
rect 6052 21972 6058 22024
rect 7742 21972 7748 22024
rect 7800 21972 7806 22024
rect 8573 22015 8631 22021
rect 8573 21981 8585 22015
rect 8619 21981 8631 22015
rect 8573 21975 8631 21981
rect 8588 21944 8616 21975
rect 9122 21972 9128 22024
rect 9180 21972 9186 22024
rect 11974 22012 11980 22024
rect 11440 21984 11980 22012
rect 11440 21944 11468 21984
rect 11974 21972 11980 21984
rect 12032 21972 12038 22024
rect 12066 21972 12072 22024
rect 12124 21972 12130 22024
rect 12434 21972 12440 22024
rect 12492 22012 12498 22024
rect 13357 22015 13415 22021
rect 13357 22012 13369 22015
rect 12492 21984 13369 22012
rect 12492 21972 12498 21984
rect 13357 21981 13369 21984
rect 13403 21981 13415 22015
rect 13357 21975 13415 21981
rect 13998 21972 14004 22024
rect 14056 22012 14062 22024
rect 15197 22015 15255 22021
rect 15197 22012 15209 22015
rect 14056 21984 15209 22012
rect 14056 21972 14062 21984
rect 15197 21981 15209 21984
rect 15243 21981 15255 22015
rect 15197 21975 15255 21981
rect 17589 22015 17647 22021
rect 17589 21981 17601 22015
rect 17635 21981 17647 22015
rect 17589 21975 17647 21981
rect 19613 22015 19671 22021
rect 19613 21981 19625 22015
rect 19659 22012 19671 22015
rect 21266 22012 21272 22024
rect 19659 21984 21272 22012
rect 19659 21981 19671 21984
rect 19613 21975 19671 21981
rect 2746 21916 8524 21944
rect 8588 21916 11468 21944
rect 11517 21947 11575 21953
rect 2746 21876 2774 21916
rect 1780 21848 2774 21876
rect 4706 21836 4712 21888
rect 4764 21876 4770 21888
rect 8389 21879 8447 21885
rect 8389 21876 8401 21879
rect 4764 21848 8401 21876
rect 4764 21836 4770 21848
rect 8389 21845 8401 21848
rect 8435 21845 8447 21879
rect 8496 21876 8524 21916
rect 11517 21913 11529 21947
rect 11563 21944 11575 21947
rect 11563 21916 12434 21944
rect 11563 21913 11575 21916
rect 11517 21907 11575 21913
rect 12406 21888 12434 21916
rect 12802 21904 12808 21956
rect 12860 21944 12866 21956
rect 13173 21947 13231 21953
rect 13173 21944 13185 21947
rect 12860 21916 13185 21944
rect 12860 21904 12866 21916
rect 13173 21913 13185 21916
rect 13219 21913 13231 21947
rect 13173 21907 13231 21913
rect 14553 21947 14611 21953
rect 14553 21913 14565 21947
rect 14599 21944 14611 21947
rect 14918 21944 14924 21956
rect 14599 21916 14924 21944
rect 14599 21913 14611 21916
rect 14553 21907 14611 21913
rect 14918 21904 14924 21916
rect 14976 21904 14982 21956
rect 15473 21947 15531 21953
rect 15473 21913 15485 21947
rect 15519 21913 15531 21947
rect 17604 21944 17632 21975
rect 21266 21972 21272 21984
rect 21324 21972 21330 22024
rect 21821 22015 21879 22021
rect 21821 21981 21833 22015
rect 21867 22012 21879 22015
rect 23124 22012 23152 22120
rect 23198 22040 23204 22092
rect 23256 22040 23262 22092
rect 23308 22080 23336 22120
rect 23382 22108 23388 22160
rect 23440 22148 23446 22160
rect 25498 22148 25504 22160
rect 23440 22120 25504 22148
rect 23440 22108 23446 22120
rect 25498 22108 25504 22120
rect 25556 22108 25562 22160
rect 26528 22148 26556 22188
rect 27798 22176 27804 22228
rect 27856 22216 27862 22228
rect 28261 22219 28319 22225
rect 28261 22216 28273 22219
rect 27856 22188 28273 22216
rect 27856 22176 27862 22188
rect 28261 22185 28273 22188
rect 28307 22185 28319 22219
rect 28261 22179 28319 22185
rect 29270 22176 29276 22228
rect 29328 22216 29334 22228
rect 29733 22219 29791 22225
rect 29733 22216 29745 22219
rect 29328 22188 29745 22216
rect 29328 22176 29334 22188
rect 29733 22185 29745 22188
rect 29779 22185 29791 22219
rect 29733 22179 29791 22185
rect 31294 22176 31300 22228
rect 31352 22216 31358 22228
rect 32214 22216 32220 22228
rect 31352 22188 32220 22216
rect 31352 22176 31358 22188
rect 32214 22176 32220 22188
rect 32272 22176 32278 22228
rect 35802 22176 35808 22228
rect 35860 22216 35866 22228
rect 38838 22216 38844 22228
rect 35860 22188 38844 22216
rect 35860 22176 35866 22188
rect 38838 22176 38844 22188
rect 38896 22176 38902 22228
rect 40034 22176 40040 22228
rect 40092 22216 40098 22228
rect 41233 22219 41291 22225
rect 41233 22216 41245 22219
rect 40092 22188 41245 22216
rect 40092 22176 40098 22188
rect 41233 22185 41245 22188
rect 41279 22185 41291 22219
rect 41233 22179 41291 22185
rect 42150 22176 42156 22228
rect 42208 22216 42214 22228
rect 47765 22219 47823 22225
rect 47765 22216 47777 22219
rect 42208 22188 47777 22216
rect 42208 22176 42214 22188
rect 47765 22185 47777 22188
rect 47811 22185 47823 22219
rect 47765 22179 47823 22185
rect 26602 22148 26608 22160
rect 26528 22120 26608 22148
rect 24578 22080 24584 22092
rect 23308 22052 24584 22080
rect 24578 22040 24584 22052
rect 24636 22040 24642 22092
rect 24762 22040 24768 22092
rect 24820 22080 24826 22092
rect 25225 22083 25283 22089
rect 25225 22080 25237 22083
rect 24820 22052 25237 22080
rect 24820 22040 24826 22052
rect 25225 22049 25237 22052
rect 25271 22080 25283 22083
rect 26142 22080 26148 22092
rect 25271 22052 26148 22080
rect 25271 22049 25283 22052
rect 25225 22043 25283 22049
rect 26142 22040 26148 22052
rect 26200 22040 26206 22092
rect 26418 22040 26424 22092
rect 26476 22040 26482 22092
rect 26528 22089 26556 22120
rect 26602 22108 26608 22120
rect 26660 22108 26666 22160
rect 33870 22148 33876 22160
rect 33704 22120 33876 22148
rect 26513 22083 26571 22089
rect 26513 22049 26525 22083
rect 26559 22080 26571 22083
rect 26559 22052 26593 22080
rect 26559 22049 26571 22052
rect 26513 22043 26571 22049
rect 27062 22040 27068 22092
rect 27120 22080 27126 22092
rect 27617 22083 27675 22089
rect 27617 22080 27629 22083
rect 27120 22052 27629 22080
rect 27120 22040 27126 22052
rect 27617 22049 27629 22052
rect 27663 22049 27675 22083
rect 27617 22043 27675 22049
rect 27890 22040 27896 22092
rect 27948 22080 27954 22092
rect 28813 22083 28871 22089
rect 28813 22080 28825 22083
rect 27948 22052 28825 22080
rect 27948 22040 27954 22052
rect 28813 22049 28825 22052
rect 28859 22080 28871 22083
rect 28902 22080 28908 22092
rect 28859 22052 28908 22080
rect 28859 22049 28871 22052
rect 28813 22043 28871 22049
rect 28902 22040 28908 22052
rect 28960 22040 28966 22092
rect 29546 22040 29552 22092
rect 29604 22080 29610 22092
rect 30466 22080 30472 22092
rect 29604 22052 30472 22080
rect 29604 22040 29610 22052
rect 30466 22040 30472 22052
rect 30524 22040 30530 22092
rect 30837 22083 30895 22089
rect 30837 22049 30849 22083
rect 30883 22080 30895 22083
rect 31570 22080 31576 22092
rect 30883 22052 31576 22080
rect 30883 22049 30895 22052
rect 30837 22043 30895 22049
rect 31570 22040 31576 22052
rect 31628 22040 31634 22092
rect 32398 22040 32404 22092
rect 32456 22080 32462 22092
rect 33704 22089 33732 22120
rect 33870 22108 33876 22120
rect 33928 22108 33934 22160
rect 38562 22108 38568 22160
rect 38620 22148 38626 22160
rect 38620 22120 40632 22148
rect 38620 22108 38626 22120
rect 32585 22083 32643 22089
rect 32585 22080 32597 22083
rect 32456 22052 32597 22080
rect 32456 22040 32462 22052
rect 32585 22049 32597 22052
rect 32631 22049 32643 22083
rect 32585 22043 32643 22049
rect 33689 22083 33747 22089
rect 33689 22049 33701 22083
rect 33735 22080 33747 22083
rect 33735 22052 33769 22080
rect 33735 22049 33747 22052
rect 33689 22043 33747 22049
rect 35894 22040 35900 22092
rect 35952 22040 35958 22092
rect 37550 22040 37556 22092
rect 37608 22040 37614 22092
rect 37642 22040 37648 22092
rect 37700 22080 37706 22092
rect 40604 22089 40632 22120
rect 40770 22108 40776 22160
rect 40828 22148 40834 22160
rect 40828 22120 41828 22148
rect 40828 22108 40834 22120
rect 41800 22089 41828 22120
rect 42536 22120 43024 22148
rect 40589 22083 40647 22089
rect 37700 22052 40172 22080
rect 37700 22040 37706 22052
rect 21867 21984 23152 22012
rect 21867 21981 21879 21984
rect 21821 21975 21879 21981
rect 23934 21972 23940 22024
rect 23992 22012 23998 22024
rect 27433 22015 27491 22021
rect 23992 21984 26004 22012
rect 23992 21972 23998 21984
rect 20438 21944 20444 21956
rect 16698 21916 17540 21944
rect 17604 21916 20444 21944
rect 15473 21907 15531 21913
rect 11422 21876 11428 21888
rect 8496 21848 11428 21876
rect 8389 21839 8447 21845
rect 11422 21836 11428 21848
rect 11480 21836 11486 21888
rect 11606 21836 11612 21888
rect 11664 21836 11670 21888
rect 12406 21848 12440 21888
rect 12434 21836 12440 21848
rect 12492 21836 12498 21888
rect 12618 21836 12624 21888
rect 12676 21876 12682 21888
rect 14645 21879 14703 21885
rect 14645 21876 14657 21879
rect 12676 21848 14657 21876
rect 12676 21836 12682 21848
rect 14645 21845 14657 21848
rect 14691 21845 14703 21879
rect 15488 21876 15516 21907
rect 16298 21876 16304 21888
rect 15488 21848 16304 21876
rect 14645 21839 14703 21845
rect 16298 21836 16304 21848
rect 16356 21836 16362 21888
rect 16482 21836 16488 21888
rect 16540 21876 16546 21888
rect 16776 21876 16804 21916
rect 16540 21848 16804 21876
rect 17512 21876 17540 21916
rect 20438 21904 20444 21916
rect 20496 21904 20502 21956
rect 21913 21947 21971 21953
rect 21913 21913 21925 21947
rect 21959 21944 21971 21947
rect 22278 21944 22284 21956
rect 21959 21916 22284 21944
rect 21959 21913 21971 21916
rect 21913 21907 21971 21913
rect 22278 21904 22284 21916
rect 22336 21904 22342 21956
rect 25041 21947 25099 21953
rect 25041 21913 25053 21947
rect 25087 21944 25099 21947
rect 25222 21944 25228 21956
rect 25087 21916 25228 21944
rect 25087 21913 25099 21916
rect 25041 21907 25099 21913
rect 25222 21904 25228 21916
rect 25280 21904 25286 21956
rect 18690 21876 18696 21888
rect 17512 21848 18696 21876
rect 16540 21836 16546 21848
rect 18690 21836 18696 21848
rect 18748 21836 18754 21888
rect 19242 21836 19248 21888
rect 19300 21876 19306 21888
rect 21453 21879 21511 21885
rect 21453 21876 21465 21879
rect 19300 21848 21465 21876
rect 19300 21836 19306 21848
rect 21453 21845 21465 21848
rect 21499 21845 21511 21879
rect 21453 21839 21511 21845
rect 21542 21836 21548 21888
rect 21600 21876 21606 21888
rect 22649 21879 22707 21885
rect 22649 21876 22661 21879
rect 21600 21848 22661 21876
rect 21600 21836 21606 21848
rect 22649 21845 22661 21848
rect 22695 21845 22707 21879
rect 22649 21839 22707 21845
rect 22830 21836 22836 21888
rect 22888 21876 22894 21888
rect 23017 21879 23075 21885
rect 23017 21876 23029 21879
rect 22888 21848 23029 21876
rect 22888 21836 22894 21848
rect 23017 21845 23029 21848
rect 23063 21845 23075 21879
rect 23017 21839 23075 21845
rect 23106 21836 23112 21888
rect 23164 21836 23170 21888
rect 23474 21836 23480 21888
rect 23532 21876 23538 21888
rect 24581 21879 24639 21885
rect 24581 21876 24593 21879
rect 23532 21848 24593 21876
rect 23532 21836 23538 21848
rect 24581 21845 24593 21848
rect 24627 21845 24639 21879
rect 24581 21839 24639 21845
rect 24946 21836 24952 21888
rect 25004 21836 25010 21888
rect 25130 21836 25136 21888
rect 25188 21876 25194 21888
rect 25866 21876 25872 21888
rect 25188 21848 25872 21876
rect 25188 21836 25194 21848
rect 25866 21836 25872 21848
rect 25924 21836 25930 21888
rect 25976 21885 26004 21984
rect 27433 21981 27445 22015
rect 27479 22012 27491 22015
rect 27706 22012 27712 22024
rect 27479 21984 27712 22012
rect 27479 21981 27491 21984
rect 27433 21975 27491 21981
rect 27706 21972 27712 21984
rect 27764 22012 27770 22024
rect 29822 22012 29828 22024
rect 27764 21984 29828 22012
rect 27764 21972 27770 21984
rect 29822 21972 29828 21984
rect 29880 21972 29886 22024
rect 29917 22015 29975 22021
rect 29917 21981 29929 22015
rect 29963 22012 29975 22015
rect 29963 21984 30880 22012
rect 29963 21981 29975 21984
rect 29917 21975 29975 21981
rect 28721 21947 28779 21953
rect 28721 21913 28733 21947
rect 28767 21944 28779 21947
rect 30374 21944 30380 21956
rect 28767 21916 30380 21944
rect 28767 21913 28779 21916
rect 28721 21907 28779 21913
rect 30374 21904 30380 21916
rect 30432 21904 30438 21956
rect 25961 21879 26019 21885
rect 25961 21845 25973 21879
rect 26007 21845 26019 21879
rect 25961 21839 26019 21845
rect 26234 21836 26240 21888
rect 26292 21876 26298 21888
rect 26329 21879 26387 21885
rect 26329 21876 26341 21879
rect 26292 21848 26341 21876
rect 26292 21836 26298 21848
rect 26329 21845 26341 21848
rect 26375 21876 26387 21879
rect 26510 21876 26516 21888
rect 26375 21848 26516 21876
rect 26375 21845 26387 21848
rect 26329 21839 26387 21845
rect 26510 21836 26516 21848
rect 26568 21836 26574 21888
rect 26602 21836 26608 21888
rect 26660 21876 26666 21888
rect 27065 21879 27123 21885
rect 27065 21876 27077 21879
rect 26660 21848 27077 21876
rect 26660 21836 26666 21848
rect 27065 21845 27077 21848
rect 27111 21845 27123 21879
rect 27065 21839 27123 21845
rect 27154 21836 27160 21888
rect 27212 21876 27218 21888
rect 27430 21876 27436 21888
rect 27212 21848 27436 21876
rect 27212 21836 27218 21848
rect 27430 21836 27436 21848
rect 27488 21836 27494 21888
rect 27525 21879 27583 21885
rect 27525 21845 27537 21879
rect 27571 21876 27583 21879
rect 28534 21876 28540 21888
rect 27571 21848 28540 21876
rect 27571 21845 27583 21848
rect 27525 21839 27583 21845
rect 28534 21836 28540 21848
rect 28592 21836 28598 21888
rect 28629 21879 28687 21885
rect 28629 21845 28641 21879
rect 28675 21876 28687 21879
rect 29546 21876 29552 21888
rect 28675 21848 29552 21876
rect 28675 21845 28687 21848
rect 28629 21839 28687 21845
rect 29546 21836 29552 21848
rect 29604 21836 29610 21888
rect 30852 21876 30880 21984
rect 34146 21972 34152 22024
rect 34204 22012 34210 22024
rect 36725 22015 36783 22021
rect 36725 22012 36737 22015
rect 34204 21984 36737 22012
rect 34204 21972 34210 21984
rect 36725 21981 36737 21984
rect 36771 21981 36783 22015
rect 36725 21975 36783 21981
rect 37274 21972 37280 22024
rect 37332 21972 37338 22024
rect 38838 22012 38844 22024
rect 38686 21984 38844 22012
rect 38838 21972 38844 21984
rect 38896 22012 38902 22024
rect 39022 22012 39028 22024
rect 38896 21984 39028 22012
rect 38896 21972 38902 21984
rect 39022 21972 39028 21984
rect 39080 21972 39086 22024
rect 31110 21904 31116 21956
rect 31168 21904 31174 21956
rect 31202 21904 31208 21956
rect 31260 21944 31266 21956
rect 33505 21947 33563 21953
rect 33505 21944 33517 21947
rect 31260 21916 31602 21944
rect 32600 21916 33517 21944
rect 31260 21904 31266 21916
rect 31294 21876 31300 21888
rect 30852 21848 31300 21876
rect 31294 21836 31300 21848
rect 31352 21836 31358 21888
rect 31386 21836 31392 21888
rect 31444 21876 31450 21888
rect 32600 21876 32628 21916
rect 33505 21913 33517 21916
rect 33551 21913 33563 21947
rect 33505 21907 33563 21913
rect 35713 21947 35771 21953
rect 35713 21913 35725 21947
rect 35759 21944 35771 21947
rect 40144 21944 40172 22052
rect 40589 22049 40601 22083
rect 40635 22049 40647 22083
rect 40589 22043 40647 22049
rect 41785 22083 41843 22089
rect 41785 22049 41797 22083
rect 41831 22049 41843 22083
rect 41785 22043 41843 22049
rect 40497 22015 40555 22021
rect 40497 21981 40509 22015
rect 40543 22012 40555 22015
rect 42536 22012 42564 22120
rect 42610 22040 42616 22092
rect 42668 22080 42674 22092
rect 42996 22080 43024 22120
rect 45462 22080 45468 22092
rect 42668 22052 42932 22080
rect 42996 22052 45468 22080
rect 42668 22040 42674 22052
rect 40543 21984 42564 22012
rect 42904 22012 42932 22052
rect 45462 22040 45468 22052
rect 45520 22040 45526 22092
rect 43441 22015 43499 22021
rect 43441 22012 43453 22015
rect 42904 21984 43453 22012
rect 40543 21981 40555 21984
rect 40497 21975 40555 21981
rect 43441 21981 43453 21984
rect 43487 21981 43499 22015
rect 43441 21975 43499 21981
rect 46750 21972 46756 22024
rect 46808 22012 46814 22024
rect 47949 22015 48007 22021
rect 47949 22012 47961 22015
rect 46808 21984 47961 22012
rect 46808 21972 46814 21984
rect 47949 21981 47961 21984
rect 47995 21981 48007 22015
rect 47949 21975 48007 21981
rect 48590 21972 48596 22024
rect 48648 21972 48654 22024
rect 41506 21944 41512 21956
rect 35759 21916 37964 21944
rect 35759 21913 35771 21916
rect 35713 21907 35771 21913
rect 31444 21848 32628 21876
rect 31444 21836 31450 21848
rect 32674 21836 32680 21888
rect 32732 21876 32738 21888
rect 33045 21879 33103 21885
rect 33045 21876 33057 21879
rect 32732 21848 33057 21876
rect 32732 21836 32738 21848
rect 33045 21845 33057 21848
rect 33091 21845 33103 21879
rect 33045 21839 33103 21845
rect 33410 21836 33416 21888
rect 33468 21836 33474 21888
rect 34790 21836 34796 21888
rect 34848 21876 34854 21888
rect 35345 21879 35403 21885
rect 35345 21876 35357 21879
rect 34848 21848 35357 21876
rect 34848 21836 34854 21848
rect 35345 21845 35357 21848
rect 35391 21845 35403 21879
rect 35345 21839 35403 21845
rect 35802 21836 35808 21888
rect 35860 21836 35866 21888
rect 36538 21836 36544 21888
rect 36596 21836 36602 21888
rect 37936 21876 37964 21916
rect 38948 21916 40080 21944
rect 40144 21916 41512 21944
rect 38948 21876 38976 21916
rect 37936 21848 38976 21876
rect 39025 21879 39083 21885
rect 39025 21845 39037 21879
rect 39071 21876 39083 21879
rect 39114 21876 39120 21888
rect 39071 21848 39120 21876
rect 39071 21845 39083 21848
rect 39025 21839 39083 21845
rect 39114 21836 39120 21848
rect 39172 21876 39178 21888
rect 39758 21876 39764 21888
rect 39172 21848 39764 21876
rect 39172 21836 39178 21848
rect 39758 21836 39764 21848
rect 39816 21836 39822 21888
rect 40052 21885 40080 21916
rect 41506 21904 41512 21916
rect 41564 21904 41570 21956
rect 41601 21947 41659 21953
rect 41601 21913 41613 21947
rect 41647 21944 41659 21947
rect 47670 21944 47676 21956
rect 41647 21916 47676 21944
rect 41647 21913 41659 21916
rect 41601 21907 41659 21913
rect 47670 21904 47676 21916
rect 47728 21904 47734 21956
rect 49142 21904 49148 21956
rect 49200 21904 49206 21956
rect 40037 21879 40095 21885
rect 40037 21845 40049 21879
rect 40083 21845 40095 21879
rect 40037 21839 40095 21845
rect 40405 21879 40463 21885
rect 40405 21845 40417 21879
rect 40451 21876 40463 21879
rect 40586 21876 40592 21888
rect 40451 21848 40592 21876
rect 40451 21845 40463 21848
rect 40405 21839 40463 21845
rect 40586 21836 40592 21848
rect 40644 21836 40650 21888
rect 40954 21836 40960 21888
rect 41012 21876 41018 21888
rect 41138 21876 41144 21888
rect 41012 21848 41144 21876
rect 41012 21836 41018 21848
rect 41138 21836 41144 21848
rect 41196 21876 41202 21888
rect 41693 21879 41751 21885
rect 41693 21876 41705 21879
rect 41196 21848 41705 21876
rect 41196 21836 41202 21848
rect 41693 21845 41705 21848
rect 41739 21845 41751 21879
rect 41693 21839 41751 21845
rect 43254 21836 43260 21888
rect 43312 21836 43318 21888
rect 48406 21836 48412 21888
rect 48464 21836 48470 21888
rect 48682 21836 48688 21888
rect 48740 21876 48746 21888
rect 49237 21879 49295 21885
rect 49237 21876 49249 21879
rect 48740 21848 49249 21876
rect 48740 21836 48746 21848
rect 49237 21845 49249 21848
rect 49283 21845 49295 21879
rect 49237 21839 49295 21845
rect 1104 21786 49864 21808
rect 1104 21734 7950 21786
rect 8002 21734 8014 21786
rect 8066 21734 8078 21786
rect 8130 21734 8142 21786
rect 8194 21734 8206 21786
rect 8258 21734 17950 21786
rect 18002 21734 18014 21786
rect 18066 21734 18078 21786
rect 18130 21734 18142 21786
rect 18194 21734 18206 21786
rect 18258 21734 27950 21786
rect 28002 21734 28014 21786
rect 28066 21734 28078 21786
rect 28130 21734 28142 21786
rect 28194 21734 28206 21786
rect 28258 21734 37950 21786
rect 38002 21734 38014 21786
rect 38066 21734 38078 21786
rect 38130 21734 38142 21786
rect 38194 21734 38206 21786
rect 38258 21734 47950 21786
rect 48002 21734 48014 21786
rect 48066 21734 48078 21786
rect 48130 21734 48142 21786
rect 48194 21734 48206 21786
rect 48258 21734 49864 21786
rect 1104 21712 49864 21734
rect 4062 21632 4068 21684
rect 4120 21672 4126 21684
rect 9674 21672 9680 21684
rect 4120 21644 9680 21672
rect 4120 21632 4126 21644
rect 9674 21632 9680 21644
rect 9732 21632 9738 21684
rect 10318 21632 10324 21684
rect 10376 21632 10382 21684
rect 10686 21632 10692 21684
rect 10744 21672 10750 21684
rect 10965 21675 11023 21681
rect 10965 21672 10977 21675
rect 10744 21644 10977 21672
rect 10744 21632 10750 21644
rect 10965 21641 10977 21644
rect 11011 21641 11023 21675
rect 13722 21672 13728 21684
rect 10965 21635 11023 21641
rect 12268 21644 13728 21672
rect 5626 21604 5632 21616
rect 1780 21576 5632 21604
rect 1780 21545 1808 21576
rect 5626 21564 5632 21576
rect 5684 21564 5690 21616
rect 10410 21604 10416 21616
rect 5920 21576 10416 21604
rect 1765 21539 1823 21545
rect 1765 21505 1777 21539
rect 1811 21505 1823 21539
rect 1765 21499 1823 21505
rect 3602 21496 3608 21548
rect 3660 21496 3666 21548
rect 5920 21545 5948 21576
rect 10410 21564 10416 21576
rect 10468 21564 10474 21616
rect 12158 21604 12164 21616
rect 10520 21576 12164 21604
rect 5905 21539 5963 21545
rect 5905 21505 5917 21539
rect 5951 21505 5963 21539
rect 5905 21499 5963 21505
rect 6546 21496 6552 21548
rect 6604 21496 6610 21548
rect 10520 21545 10548 21576
rect 12158 21564 12164 21576
rect 12216 21564 12222 21616
rect 12268 21613 12296 21644
rect 13722 21632 13728 21644
rect 13780 21632 13786 21684
rect 17126 21672 17132 21684
rect 13832 21644 17132 21672
rect 12253 21607 12311 21613
rect 12253 21573 12265 21607
rect 12299 21573 12311 21607
rect 12253 21567 12311 21573
rect 12342 21564 12348 21616
rect 12400 21604 12406 21616
rect 13446 21604 13452 21616
rect 12400 21576 13452 21604
rect 12400 21564 12406 21576
rect 13446 21564 13452 21576
rect 13504 21564 13510 21616
rect 8389 21539 8447 21545
rect 8389 21505 8401 21539
rect 8435 21505 8447 21539
rect 8389 21499 8447 21505
rect 10505 21539 10563 21545
rect 10505 21505 10517 21539
rect 10551 21505 10563 21539
rect 10505 21499 10563 21505
rect 11149 21539 11207 21545
rect 11149 21505 11161 21539
rect 11195 21536 11207 21539
rect 11195 21508 12434 21536
rect 11195 21505 11207 21508
rect 11149 21499 11207 21505
rect 2777 21471 2835 21477
rect 2777 21437 2789 21471
rect 2823 21468 2835 21471
rect 3326 21468 3332 21480
rect 2823 21440 3332 21468
rect 2823 21437 2835 21440
rect 2777 21431 2835 21437
rect 3326 21428 3332 21440
rect 3384 21428 3390 21480
rect 4154 21428 4160 21480
rect 4212 21428 4218 21480
rect 5534 21428 5540 21480
rect 5592 21468 5598 21480
rect 7009 21471 7067 21477
rect 7009 21468 7021 21471
rect 5592 21440 7021 21468
rect 5592 21428 5598 21440
rect 7009 21437 7021 21440
rect 7055 21437 7067 21471
rect 7009 21431 7067 21437
rect 5721 21403 5779 21409
rect 5721 21369 5733 21403
rect 5767 21400 5779 21403
rect 8404 21400 8432 21499
rect 8846 21428 8852 21480
rect 8904 21428 8910 21480
rect 9858 21428 9864 21480
rect 9916 21468 9922 21480
rect 11606 21468 11612 21480
rect 9916 21440 11612 21468
rect 9916 21428 9922 21440
rect 11606 21428 11612 21440
rect 11664 21428 11670 21480
rect 12406 21468 12434 21508
rect 12618 21496 12624 21548
rect 12676 21536 12682 21548
rect 13357 21539 13415 21545
rect 13357 21536 13369 21539
rect 12676 21508 13369 21536
rect 12676 21496 12682 21508
rect 13357 21505 13369 21508
rect 13403 21505 13415 21539
rect 13832 21536 13860 21644
rect 17126 21632 17132 21644
rect 17184 21632 17190 21684
rect 17402 21632 17408 21684
rect 17460 21632 17466 21684
rect 17770 21632 17776 21684
rect 17828 21672 17834 21684
rect 17865 21675 17923 21681
rect 17865 21672 17877 21675
rect 17828 21644 17877 21672
rect 17828 21632 17834 21644
rect 17865 21641 17877 21644
rect 17911 21641 17923 21675
rect 20530 21672 20536 21684
rect 17865 21635 17923 21641
rect 18064 21644 20536 21672
rect 14826 21564 14832 21616
rect 14884 21564 14890 21616
rect 16114 21604 16120 21616
rect 16054 21576 16120 21604
rect 16114 21564 16120 21576
rect 16172 21604 16178 21616
rect 16482 21604 16488 21616
rect 16172 21576 16488 21604
rect 16172 21564 16178 21576
rect 16482 21564 16488 21576
rect 16540 21564 16546 21616
rect 13357 21499 13415 21505
rect 13648 21508 13860 21536
rect 12526 21468 12532 21480
rect 12406 21440 12532 21468
rect 12526 21428 12532 21440
rect 12584 21428 12590 21480
rect 13648 21477 13676 21508
rect 17770 21496 17776 21548
rect 17828 21496 17834 21548
rect 13449 21471 13507 21477
rect 13449 21437 13461 21471
rect 13495 21437 13507 21471
rect 13449 21431 13507 21437
rect 13633 21471 13691 21477
rect 13633 21437 13645 21471
rect 13679 21437 13691 21471
rect 13633 21431 13691 21437
rect 5767 21372 8432 21400
rect 5767 21369 5779 21372
rect 5721 21363 5779 21369
rect 11238 21360 11244 21412
rect 11296 21400 11302 21412
rect 12989 21403 13047 21409
rect 12989 21400 13001 21403
rect 11296 21372 13001 21400
rect 11296 21360 11302 21372
rect 12989 21369 13001 21372
rect 13035 21369 13047 21403
rect 13464 21400 13492 21431
rect 13722 21428 13728 21480
rect 13780 21468 13786 21480
rect 14550 21468 14556 21480
rect 13780 21440 14556 21468
rect 13780 21428 13786 21440
rect 14550 21428 14556 21440
rect 14608 21428 14614 21480
rect 16390 21468 16396 21480
rect 14660 21440 16396 21468
rect 14660 21400 14688 21440
rect 16390 21428 16396 21440
rect 16448 21428 16454 21480
rect 18064 21477 18092 21644
rect 20530 21632 20536 21644
rect 20588 21632 20594 21684
rect 20990 21632 20996 21684
rect 21048 21632 21054 21684
rect 22554 21632 22560 21684
rect 22612 21672 22618 21684
rect 23106 21672 23112 21684
rect 22612 21644 23112 21672
rect 22612 21632 22618 21644
rect 23106 21632 23112 21644
rect 23164 21632 23170 21684
rect 24762 21632 24768 21684
rect 24820 21632 24826 21684
rect 26421 21675 26479 21681
rect 26421 21641 26433 21675
rect 26467 21672 26479 21675
rect 27246 21672 27252 21684
rect 26467 21644 27252 21672
rect 26467 21641 26479 21644
rect 26421 21635 26479 21641
rect 27246 21632 27252 21644
rect 27304 21632 27310 21684
rect 27617 21675 27675 21681
rect 27617 21641 27629 21675
rect 27663 21672 27675 21675
rect 27706 21672 27712 21684
rect 27663 21644 27712 21672
rect 27663 21641 27675 21644
rect 27617 21635 27675 21641
rect 27706 21632 27712 21644
rect 27764 21632 27770 21684
rect 27798 21632 27804 21684
rect 27856 21672 27862 21684
rect 28353 21675 28411 21681
rect 28353 21672 28365 21675
rect 27856 21644 28365 21672
rect 27856 21632 27862 21644
rect 28353 21641 28365 21644
rect 28399 21641 28411 21675
rect 28353 21635 28411 21641
rect 28442 21632 28448 21684
rect 28500 21672 28506 21684
rect 31110 21672 31116 21684
rect 28500 21644 31116 21672
rect 28500 21632 28506 21644
rect 31110 21632 31116 21644
rect 31168 21632 31174 21684
rect 32600 21644 34744 21672
rect 18782 21564 18788 21616
rect 18840 21604 18846 21616
rect 18877 21607 18935 21613
rect 18877 21604 18889 21607
rect 18840 21576 18889 21604
rect 18840 21564 18846 21576
rect 18877 21573 18889 21576
rect 18923 21573 18935 21607
rect 20346 21604 20352 21616
rect 20102 21576 20352 21604
rect 18877 21567 18935 21573
rect 20346 21564 20352 21576
rect 20404 21604 20410 21616
rect 22278 21604 22284 21616
rect 20404 21576 22284 21604
rect 20404 21564 20410 21576
rect 22278 21564 22284 21576
rect 22336 21604 22342 21616
rect 22738 21604 22744 21616
rect 22336 21576 22744 21604
rect 22336 21564 22342 21576
rect 22738 21564 22744 21576
rect 22796 21604 22802 21616
rect 25225 21607 25283 21613
rect 25225 21604 25237 21607
rect 22796 21576 23230 21604
rect 24872 21576 25237 21604
rect 22796 21564 22802 21576
rect 20901 21539 20959 21545
rect 20901 21505 20913 21539
rect 20947 21536 20959 21539
rect 21634 21536 21640 21548
rect 20947 21508 21640 21536
rect 20947 21505 20959 21508
rect 20901 21499 20959 21505
rect 21634 21496 21640 21508
rect 21692 21496 21698 21548
rect 24872 21536 24900 21576
rect 25225 21573 25237 21576
rect 25271 21604 25283 21607
rect 27430 21604 27436 21616
rect 25271 21576 27436 21604
rect 25271 21573 25283 21576
rect 25225 21567 25283 21573
rect 27430 21564 27436 21576
rect 27488 21564 27494 21616
rect 27525 21607 27583 21613
rect 27525 21573 27537 21607
rect 27571 21604 27583 21607
rect 29086 21604 29092 21616
rect 27571 21576 29092 21604
rect 27571 21573 27583 21576
rect 27525 21567 27583 21573
rect 29086 21564 29092 21576
rect 29144 21564 29150 21616
rect 30009 21607 30067 21613
rect 30009 21573 30021 21607
rect 30055 21604 30067 21607
rect 32490 21604 32496 21616
rect 30055 21576 32496 21604
rect 30055 21573 30067 21576
rect 30009 21567 30067 21573
rect 32490 21564 32496 21576
rect 32548 21564 32554 21616
rect 23952 21508 24900 21536
rect 18049 21471 18107 21477
rect 18049 21437 18061 21471
rect 18095 21437 18107 21471
rect 18049 21431 18107 21437
rect 18598 21428 18604 21480
rect 18656 21428 18662 21480
rect 20714 21428 20720 21480
rect 20772 21468 20778 21480
rect 22002 21468 22008 21480
rect 20772 21440 22008 21468
rect 20772 21428 20778 21440
rect 22002 21428 22008 21440
rect 22060 21468 22066 21480
rect 22465 21471 22523 21477
rect 22465 21468 22477 21471
rect 22060 21440 22477 21468
rect 22060 21428 22066 21440
rect 22465 21437 22477 21440
rect 22511 21437 22523 21471
rect 22741 21471 22799 21477
rect 22741 21468 22753 21471
rect 22465 21431 22523 21437
rect 22572 21440 22753 21468
rect 13464 21372 14688 21400
rect 12989 21363 13047 21369
rect 17034 21360 17040 21412
rect 17092 21400 17098 21412
rect 18616 21400 18644 21428
rect 22572 21400 22600 21440
rect 22741 21437 22753 21440
rect 22787 21437 22799 21471
rect 22741 21431 22799 21437
rect 23382 21428 23388 21480
rect 23440 21468 23446 21480
rect 23952 21468 23980 21508
rect 25130 21496 25136 21548
rect 25188 21496 25194 21548
rect 26605 21539 26663 21545
rect 26605 21505 26617 21539
rect 26651 21536 26663 21539
rect 26651 21508 27844 21536
rect 26651 21505 26663 21508
rect 26605 21499 26663 21505
rect 23440 21440 23980 21468
rect 23440 21428 23446 21440
rect 24210 21428 24216 21480
rect 24268 21428 24274 21480
rect 25406 21428 25412 21480
rect 25464 21468 25470 21480
rect 27709 21471 27767 21477
rect 25464 21440 27568 21468
rect 25464 21428 25470 21440
rect 17092 21372 18644 21400
rect 19904 21372 22600 21400
rect 17092 21360 17098 21372
rect 4062 21292 4068 21344
rect 4120 21332 4126 21344
rect 12345 21335 12403 21341
rect 12345 21332 12357 21335
rect 4120 21304 12357 21332
rect 4120 21292 4126 21304
rect 12345 21301 12357 21304
rect 12391 21301 12403 21335
rect 12345 21295 12403 21301
rect 13538 21292 13544 21344
rect 13596 21332 13602 21344
rect 15470 21332 15476 21344
rect 13596 21304 15476 21332
rect 13596 21292 13602 21304
rect 15470 21292 15476 21304
rect 15528 21292 15534 21344
rect 16298 21292 16304 21344
rect 16356 21292 16362 21344
rect 19058 21292 19064 21344
rect 19116 21332 19122 21344
rect 19904 21332 19932 21372
rect 23750 21360 23756 21412
rect 23808 21400 23814 21412
rect 27157 21403 27215 21409
rect 27157 21400 27169 21403
rect 23808 21372 27169 21400
rect 23808 21360 23814 21372
rect 27157 21369 27169 21372
rect 27203 21369 27215 21403
rect 27540 21400 27568 21440
rect 27709 21437 27721 21471
rect 27755 21437 27767 21471
rect 27709 21431 27767 21437
rect 27724 21400 27752 21431
rect 27540 21372 27752 21400
rect 27816 21400 27844 21508
rect 27890 21496 27896 21548
rect 27948 21536 27954 21548
rect 28721 21539 28779 21545
rect 28721 21536 28733 21539
rect 27948 21508 28733 21536
rect 27948 21496 27954 21508
rect 28721 21505 28733 21508
rect 28767 21505 28779 21539
rect 28721 21499 28779 21505
rect 29917 21539 29975 21545
rect 29917 21505 29929 21539
rect 29963 21505 29975 21539
rect 29917 21499 29975 21505
rect 28258 21428 28264 21480
rect 28316 21468 28322 21480
rect 28813 21471 28871 21477
rect 28813 21468 28825 21471
rect 28316 21440 28825 21468
rect 28316 21428 28322 21440
rect 28813 21437 28825 21440
rect 28859 21437 28871 21471
rect 28813 21431 28871 21437
rect 28902 21428 28908 21480
rect 28960 21428 28966 21480
rect 29730 21400 29736 21412
rect 27816 21372 29736 21400
rect 27157 21363 27215 21369
rect 29730 21360 29736 21372
rect 29788 21360 29794 21412
rect 29932 21400 29960 21499
rect 30466 21496 30472 21548
rect 30524 21536 30530 21548
rect 31018 21536 31024 21548
rect 30524 21508 31024 21536
rect 30524 21496 30530 21508
rect 31018 21496 31024 21508
rect 31076 21496 31082 21548
rect 31113 21539 31171 21545
rect 31113 21505 31125 21539
rect 31159 21536 31171 21539
rect 32600 21536 32628 21644
rect 33410 21604 33416 21616
rect 32692 21576 33416 21604
rect 32692 21545 32720 21576
rect 33410 21564 33416 21576
rect 33468 21564 33474 21616
rect 33686 21564 33692 21616
rect 33744 21604 33750 21616
rect 33870 21604 33876 21616
rect 33744 21576 33876 21604
rect 33744 21564 33750 21576
rect 33870 21564 33876 21576
rect 33928 21564 33934 21616
rect 34716 21548 34744 21644
rect 34882 21632 34888 21684
rect 34940 21672 34946 21684
rect 37734 21672 37740 21684
rect 34940 21644 37740 21672
rect 34940 21632 34946 21644
rect 37734 21632 37740 21644
rect 37792 21632 37798 21684
rect 40126 21632 40132 21684
rect 40184 21672 40190 21684
rect 40221 21675 40279 21681
rect 40221 21672 40233 21675
rect 40184 21644 40233 21672
rect 40184 21632 40190 21644
rect 40221 21641 40233 21644
rect 40267 21641 40279 21675
rect 40221 21635 40279 21641
rect 40586 21632 40592 21684
rect 40644 21672 40650 21684
rect 46842 21672 46848 21684
rect 40644 21644 46848 21672
rect 40644 21632 40650 21644
rect 46842 21632 46848 21644
rect 46900 21632 46906 21684
rect 36081 21607 36139 21613
rect 36081 21573 36093 21607
rect 36127 21604 36139 21607
rect 36262 21604 36268 21616
rect 36127 21576 36268 21604
rect 36127 21573 36139 21576
rect 36081 21567 36139 21573
rect 36262 21564 36268 21576
rect 36320 21564 36326 21616
rect 39022 21604 39028 21616
rect 38962 21576 39028 21604
rect 39022 21564 39028 21576
rect 39080 21604 39086 21616
rect 39482 21604 39488 21616
rect 39080 21576 39488 21604
rect 39080 21564 39086 21576
rect 39482 21564 39488 21576
rect 39540 21564 39546 21616
rect 41138 21564 41144 21616
rect 41196 21604 41202 21616
rect 41322 21604 41328 21616
rect 41196 21576 41328 21604
rect 41196 21564 41202 21576
rect 41322 21564 41328 21576
rect 41380 21604 41386 21616
rect 47118 21604 47124 21616
rect 41380 21576 47124 21604
rect 41380 21564 41386 21576
rect 47118 21564 47124 21576
rect 47176 21564 47182 21616
rect 31159 21508 32628 21536
rect 32677 21539 32735 21545
rect 31159 21505 31171 21508
rect 31113 21499 31171 21505
rect 32677 21505 32689 21539
rect 32723 21505 32735 21539
rect 32677 21499 32735 21505
rect 34698 21496 34704 21548
rect 34756 21536 34762 21548
rect 37090 21536 37096 21548
rect 34756 21508 37096 21536
rect 34756 21496 34762 21508
rect 37090 21496 37096 21508
rect 37148 21496 37154 21548
rect 37274 21496 37280 21548
rect 37332 21536 37338 21548
rect 37461 21539 37519 21545
rect 37461 21536 37473 21539
rect 37332 21508 37473 21536
rect 37332 21496 37338 21508
rect 37461 21505 37473 21508
rect 37507 21505 37519 21539
rect 37461 21499 37519 21505
rect 39666 21496 39672 21548
rect 39724 21536 39730 21548
rect 40589 21539 40647 21545
rect 40589 21536 40601 21539
rect 39724 21508 40601 21536
rect 39724 21496 39730 21508
rect 40589 21505 40601 21508
rect 40635 21536 40647 21539
rect 46934 21536 46940 21548
rect 40635 21508 46940 21536
rect 40635 21505 40647 21508
rect 40589 21499 40647 21505
rect 46934 21496 46940 21508
rect 46992 21496 46998 21548
rect 49050 21496 49056 21548
rect 49108 21496 49114 21548
rect 30006 21428 30012 21480
rect 30064 21468 30070 21480
rect 30101 21471 30159 21477
rect 30101 21468 30113 21471
rect 30064 21440 30113 21468
rect 30064 21428 30070 21440
rect 30101 21437 30113 21440
rect 30147 21437 30159 21471
rect 30101 21431 30159 21437
rect 31202 21428 31208 21480
rect 31260 21428 31266 21480
rect 31389 21471 31447 21477
rect 31389 21437 31401 21471
rect 31435 21468 31447 21471
rect 31478 21468 31484 21480
rect 31435 21440 31484 21468
rect 31435 21437 31447 21440
rect 31389 21431 31447 21437
rect 31478 21428 31484 21440
rect 31536 21428 31542 21480
rect 31570 21428 31576 21480
rect 31628 21468 31634 21480
rect 33137 21471 33195 21477
rect 33137 21468 33149 21471
rect 31628 21440 33149 21468
rect 31628 21428 31634 21440
rect 33137 21437 33149 21440
rect 33183 21437 33195 21471
rect 33137 21431 33195 21437
rect 33410 21428 33416 21480
rect 33468 21428 33474 21480
rect 36170 21428 36176 21480
rect 36228 21428 36234 21480
rect 36357 21471 36415 21477
rect 36357 21437 36369 21471
rect 36403 21468 36415 21471
rect 36906 21468 36912 21480
rect 36403 21440 36912 21468
rect 36403 21437 36415 21440
rect 36357 21431 36415 21437
rect 36906 21428 36912 21440
rect 36964 21428 36970 21480
rect 37737 21471 37795 21477
rect 37737 21468 37749 21471
rect 37568 21440 37749 21468
rect 32674 21400 32680 21412
rect 29932 21372 32680 21400
rect 32674 21360 32680 21372
rect 32732 21400 32738 21412
rect 32858 21400 32864 21412
rect 32732 21372 32864 21400
rect 32732 21360 32738 21372
rect 32858 21360 32864 21372
rect 32916 21360 32922 21412
rect 36538 21400 36544 21412
rect 34808 21372 36544 21400
rect 19116 21304 19932 21332
rect 19116 21292 19122 21304
rect 20254 21292 20260 21344
rect 20312 21332 20318 21344
rect 20349 21335 20407 21341
rect 20349 21332 20361 21335
rect 20312 21304 20361 21332
rect 20312 21292 20318 21304
rect 20349 21301 20361 21304
rect 20395 21301 20407 21335
rect 20349 21295 20407 21301
rect 21910 21292 21916 21344
rect 21968 21332 21974 21344
rect 26142 21332 26148 21344
rect 21968 21304 26148 21332
rect 21968 21292 21974 21304
rect 26142 21292 26148 21304
rect 26200 21292 26206 21344
rect 26234 21292 26240 21344
rect 26292 21332 26298 21344
rect 28626 21332 28632 21344
rect 26292 21304 28632 21332
rect 26292 21292 26298 21304
rect 28626 21292 28632 21304
rect 28684 21332 28690 21344
rect 28902 21332 28908 21344
rect 28684 21304 28908 21332
rect 28684 21292 28690 21304
rect 28902 21292 28908 21304
rect 28960 21292 28966 21344
rect 29086 21292 29092 21344
rect 29144 21332 29150 21344
rect 29270 21332 29276 21344
rect 29144 21304 29276 21332
rect 29144 21292 29150 21304
rect 29270 21292 29276 21304
rect 29328 21292 29334 21344
rect 29546 21292 29552 21344
rect 29604 21292 29610 21344
rect 30374 21292 30380 21344
rect 30432 21332 30438 21344
rect 30745 21335 30803 21341
rect 30745 21332 30757 21335
rect 30432 21304 30757 21332
rect 30432 21292 30438 21304
rect 30745 21301 30757 21304
rect 30791 21301 30803 21335
rect 30745 21295 30803 21301
rect 30834 21292 30840 21344
rect 30892 21332 30898 21344
rect 34808 21332 34836 21372
rect 36538 21360 36544 21372
rect 36596 21360 36602 21412
rect 37568 21400 37596 21440
rect 37737 21437 37749 21440
rect 37783 21468 37795 21471
rect 39114 21468 39120 21480
rect 37783 21440 39120 21468
rect 37783 21437 37795 21440
rect 37737 21431 37795 21437
rect 39114 21428 39120 21440
rect 39172 21428 39178 21480
rect 40402 21428 40408 21480
rect 40460 21468 40466 21480
rect 40678 21468 40684 21480
rect 40460 21440 40684 21468
rect 40460 21428 40466 21440
rect 40678 21428 40684 21440
rect 40736 21428 40742 21480
rect 40770 21428 40776 21480
rect 40828 21428 40834 21480
rect 43254 21400 43260 21412
rect 37384 21372 37596 21400
rect 38764 21372 43260 21400
rect 30892 21304 34836 21332
rect 30892 21292 30898 21304
rect 35618 21292 35624 21344
rect 35676 21332 35682 21344
rect 35713 21335 35771 21341
rect 35713 21332 35725 21335
rect 35676 21304 35725 21332
rect 35676 21292 35682 21304
rect 35713 21301 35725 21304
rect 35759 21301 35771 21335
rect 35713 21295 35771 21301
rect 36170 21292 36176 21344
rect 36228 21332 36234 21344
rect 37384 21332 37412 21372
rect 36228 21304 37412 21332
rect 36228 21292 36234 21304
rect 37918 21292 37924 21344
rect 37976 21332 37982 21344
rect 38764 21332 38792 21372
rect 43254 21360 43260 21372
rect 43312 21360 43318 21412
rect 43622 21360 43628 21412
rect 43680 21400 43686 21412
rect 48958 21400 48964 21412
rect 43680 21372 48964 21400
rect 43680 21360 43686 21372
rect 48958 21360 48964 21372
rect 49016 21360 49022 21412
rect 37976 21304 38792 21332
rect 37976 21292 37982 21304
rect 39206 21292 39212 21344
rect 39264 21292 39270 21344
rect 39666 21292 39672 21344
rect 39724 21292 39730 21344
rect 41598 21292 41604 21344
rect 41656 21332 41662 21344
rect 49237 21335 49295 21341
rect 49237 21332 49249 21335
rect 41656 21304 49249 21332
rect 41656 21292 41662 21304
rect 49237 21301 49249 21304
rect 49283 21301 49295 21335
rect 49237 21295 49295 21301
rect 1104 21242 49864 21264
rect 1104 21190 2950 21242
rect 3002 21190 3014 21242
rect 3066 21190 3078 21242
rect 3130 21190 3142 21242
rect 3194 21190 3206 21242
rect 3258 21190 12950 21242
rect 13002 21190 13014 21242
rect 13066 21190 13078 21242
rect 13130 21190 13142 21242
rect 13194 21190 13206 21242
rect 13258 21190 22950 21242
rect 23002 21190 23014 21242
rect 23066 21190 23078 21242
rect 23130 21190 23142 21242
rect 23194 21190 23206 21242
rect 23258 21190 32950 21242
rect 33002 21190 33014 21242
rect 33066 21190 33078 21242
rect 33130 21190 33142 21242
rect 33194 21190 33206 21242
rect 33258 21190 42950 21242
rect 43002 21190 43014 21242
rect 43066 21190 43078 21242
rect 43130 21190 43142 21242
rect 43194 21190 43206 21242
rect 43258 21190 49864 21242
rect 1104 21168 49864 21190
rect 5994 21088 6000 21140
rect 6052 21128 6058 21140
rect 9861 21131 9919 21137
rect 6052 21100 7972 21128
rect 6052 21088 6058 21100
rect 7837 21063 7895 21069
rect 7837 21060 7849 21063
rect 6012 21032 7849 21060
rect 4246 20952 4252 21004
rect 4304 20992 4310 21004
rect 4433 20995 4491 21001
rect 4433 20992 4445 20995
rect 4304 20964 4445 20992
rect 4304 20952 4310 20964
rect 4433 20961 4445 20964
rect 4479 20961 4491 20995
rect 4433 20955 4491 20961
rect 1765 20927 1823 20933
rect 1765 20893 1777 20927
rect 1811 20924 1823 20927
rect 1811 20896 4016 20924
rect 1811 20893 1823 20896
rect 1765 20887 1823 20893
rect 2774 20816 2780 20868
rect 2832 20816 2838 20868
rect 3988 20856 4016 20896
rect 4062 20884 4068 20936
rect 4120 20884 4126 20936
rect 6012 20933 6040 21032
rect 7837 21029 7849 21032
rect 7883 21029 7895 21063
rect 7944 21060 7972 21100
rect 9861 21097 9873 21131
rect 9907 21128 9919 21131
rect 12618 21128 12624 21140
rect 9907 21100 12624 21128
rect 9907 21097 9919 21100
rect 9861 21091 9919 21097
rect 12618 21088 12624 21100
rect 12676 21088 12682 21140
rect 12710 21088 12716 21140
rect 12768 21128 12774 21140
rect 12897 21131 12955 21137
rect 12897 21128 12909 21131
rect 12768 21100 12909 21128
rect 12768 21088 12774 21100
rect 12897 21097 12909 21100
rect 12943 21097 12955 21131
rect 12897 21091 12955 21097
rect 13630 21088 13636 21140
rect 13688 21088 13694 21140
rect 15286 21128 15292 21140
rect 13740 21100 15292 21128
rect 12069 21063 12127 21069
rect 12069 21060 12081 21063
rect 7944 21032 12081 21060
rect 7837 21023 7895 21029
rect 12069 21029 12081 21032
rect 12115 21029 12127 21063
rect 12069 21023 12127 21029
rect 6730 20952 6736 21004
rect 6788 20952 6794 21004
rect 10505 20995 10563 21001
rect 10505 20961 10517 20995
rect 10551 20992 10563 20995
rect 13630 20992 13636 21004
rect 10551 20964 13636 20992
rect 10551 20961 10563 20964
rect 10505 20955 10563 20961
rect 13630 20952 13636 20964
rect 13688 20952 13694 21004
rect 5997 20927 6055 20933
rect 5997 20893 6009 20927
rect 6043 20893 6055 20927
rect 5997 20887 6055 20893
rect 8021 20927 8079 20933
rect 8021 20893 8033 20927
rect 8067 20924 8079 20927
rect 10962 20924 10968 20936
rect 8067 20896 10968 20924
rect 8067 20893 8079 20896
rect 8021 20887 8079 20893
rect 10962 20884 10968 20896
rect 11020 20884 11026 20936
rect 11146 20884 11152 20936
rect 11204 20884 11210 20936
rect 12805 20927 12863 20933
rect 12805 20893 12817 20927
rect 12851 20924 12863 20927
rect 13740 20924 13768 21100
rect 15286 21088 15292 21100
rect 15344 21088 15350 21140
rect 17770 21088 17776 21140
rect 17828 21128 17834 21140
rect 17828 21100 18828 21128
rect 17828 21088 17834 21100
rect 13906 21020 13912 21072
rect 13964 21060 13970 21072
rect 14182 21060 14188 21072
rect 13964 21032 14188 21060
rect 13964 21020 13970 21032
rect 14182 21020 14188 21032
rect 14240 21020 14246 21072
rect 18800 21060 18828 21100
rect 18874 21088 18880 21140
rect 18932 21088 18938 21140
rect 21348 21131 21406 21137
rect 21348 21097 21360 21131
rect 21394 21128 21406 21131
rect 22370 21128 22376 21140
rect 21394 21100 22376 21128
rect 21394 21097 21406 21100
rect 21348 21091 21406 21097
rect 22370 21088 22376 21100
rect 22428 21088 22434 21140
rect 27798 21128 27804 21140
rect 25240 21100 27804 21128
rect 19797 21063 19855 21069
rect 19797 21060 19809 21063
rect 18800 21032 19809 21060
rect 19797 21029 19809 21032
rect 19843 21029 19855 21063
rect 20990 21060 20996 21072
rect 19797 21023 19855 21029
rect 20364 21032 20996 21060
rect 14550 20952 14556 21004
rect 14608 20992 14614 21004
rect 17034 20992 17040 21004
rect 14608 20964 17040 20992
rect 14608 20952 14614 20964
rect 17034 20952 17040 20964
rect 17092 20992 17098 21004
rect 17129 20995 17187 21001
rect 17129 20992 17141 20995
rect 17092 20964 17141 20992
rect 17092 20952 17098 20964
rect 17129 20961 17141 20964
rect 17175 20961 17187 20995
rect 17129 20955 17187 20961
rect 17405 20995 17463 21001
rect 17405 20961 17417 20995
rect 17451 20992 17463 20995
rect 20364 20992 20392 21032
rect 20990 21020 20996 21032
rect 21048 21020 21054 21072
rect 22462 21020 22468 21072
rect 22520 21060 22526 21072
rect 22833 21063 22891 21069
rect 22833 21060 22845 21063
rect 22520 21032 22845 21060
rect 22520 21020 22526 21032
rect 22833 21029 22845 21032
rect 22879 21029 22891 21063
rect 22833 21023 22891 21029
rect 17451 20964 20392 20992
rect 20441 20995 20499 21001
rect 17451 20961 17463 20964
rect 17405 20955 17463 20961
rect 20441 20961 20453 20995
rect 20487 20992 20499 20995
rect 22094 20992 22100 21004
rect 20487 20964 22100 20992
rect 20487 20961 20499 20964
rect 20441 20955 20499 20961
rect 22094 20952 22100 20964
rect 22152 20952 22158 21004
rect 22370 20952 22376 21004
rect 22428 20992 22434 21004
rect 22554 20992 22560 21004
rect 22428 20964 22560 20992
rect 22428 20952 22434 20964
rect 22554 20952 22560 20964
rect 22612 20952 22618 21004
rect 25240 21001 25268 21100
rect 27798 21088 27804 21100
rect 27856 21088 27862 21140
rect 27890 21088 27896 21140
rect 27948 21088 27954 21140
rect 28353 21131 28411 21137
rect 28353 21097 28365 21131
rect 28399 21128 28411 21131
rect 30098 21128 30104 21140
rect 28399 21100 30104 21128
rect 28399 21097 28411 21100
rect 28353 21091 28411 21097
rect 30098 21088 30104 21100
rect 30156 21088 30162 21140
rect 30282 21088 30288 21140
rect 30340 21128 30346 21140
rect 30837 21131 30895 21137
rect 30837 21128 30849 21131
rect 30340 21100 30849 21128
rect 30340 21088 30346 21100
rect 30837 21097 30849 21100
rect 30883 21097 30895 21131
rect 30837 21091 30895 21097
rect 31202 21088 31208 21140
rect 31260 21128 31266 21140
rect 33134 21128 33140 21140
rect 31260 21100 33140 21128
rect 31260 21088 31266 21100
rect 33134 21088 33140 21100
rect 33192 21088 33198 21140
rect 33229 21131 33287 21137
rect 33229 21097 33241 21131
rect 33275 21128 33287 21131
rect 36262 21128 36268 21140
rect 33275 21100 36268 21128
rect 33275 21097 33287 21100
rect 33229 21091 33287 21097
rect 36262 21088 36268 21100
rect 36320 21088 36326 21140
rect 37277 21131 37335 21137
rect 37277 21097 37289 21131
rect 37323 21128 37335 21131
rect 37366 21128 37372 21140
rect 37323 21100 37372 21128
rect 37323 21097 37335 21100
rect 37277 21091 37335 21097
rect 37366 21088 37372 21100
rect 37424 21088 37430 21140
rect 38746 21088 38752 21140
rect 38804 21128 38810 21140
rect 40037 21131 40095 21137
rect 40037 21128 40049 21131
rect 38804 21100 40049 21128
rect 38804 21088 38810 21100
rect 40037 21097 40049 21100
rect 40083 21097 40095 21131
rect 40037 21091 40095 21097
rect 40310 21088 40316 21140
rect 40368 21128 40374 21140
rect 43622 21128 43628 21140
rect 40368 21100 43628 21128
rect 40368 21088 40374 21100
rect 43622 21088 43628 21100
rect 43680 21088 43686 21140
rect 48958 21088 48964 21140
rect 49016 21128 49022 21140
rect 49237 21131 49295 21137
rect 49237 21128 49249 21131
rect 49016 21100 49249 21128
rect 49016 21088 49022 21100
rect 49237 21097 49249 21100
rect 49283 21097 49295 21131
rect 49237 21091 49295 21097
rect 26142 21020 26148 21072
rect 26200 21060 26206 21072
rect 29733 21063 29791 21069
rect 29733 21060 29745 21063
rect 26200 21032 29745 21060
rect 26200 21020 26206 21032
rect 29733 21029 29745 21032
rect 29779 21029 29791 21063
rect 34790 21060 34796 21072
rect 29733 21023 29791 21029
rect 31312 21032 34796 21060
rect 23845 20995 23903 21001
rect 23845 20992 23857 20995
rect 22664 20964 23857 20992
rect 12851 20896 13768 20924
rect 12851 20893 12863 20896
rect 12805 20887 12863 20893
rect 13998 20884 14004 20936
rect 14056 20924 14062 20936
rect 14277 20927 14335 20933
rect 14277 20924 14289 20927
rect 14056 20896 14289 20924
rect 14056 20884 14062 20896
rect 14277 20893 14289 20896
rect 14323 20893 14335 20927
rect 14277 20887 14335 20893
rect 16669 20927 16727 20933
rect 16669 20893 16681 20927
rect 16715 20893 16727 20927
rect 16669 20887 16727 20893
rect 11514 20856 11520 20868
rect 3988 20828 11520 20856
rect 11514 20816 11520 20828
rect 11572 20816 11578 20868
rect 11885 20859 11943 20865
rect 11885 20825 11897 20859
rect 11931 20856 11943 20859
rect 11931 20828 12434 20856
rect 11931 20825 11943 20828
rect 11885 20819 11943 20825
rect 7834 20748 7840 20800
rect 7892 20788 7898 20800
rect 10965 20791 11023 20797
rect 10965 20788 10977 20791
rect 7892 20760 10977 20788
rect 7892 20748 7898 20760
rect 10965 20757 10977 20760
rect 11011 20757 11023 20791
rect 12406 20788 12434 20828
rect 13538 20816 13544 20868
rect 13596 20816 13602 20868
rect 13906 20816 13912 20868
rect 13964 20856 13970 20868
rect 14553 20859 14611 20865
rect 14553 20856 14565 20859
rect 13964 20828 14565 20856
rect 13964 20816 13970 20828
rect 14553 20825 14565 20828
rect 14599 20825 14611 20859
rect 15838 20856 15844 20868
rect 15778 20828 15844 20856
rect 14553 20819 14611 20825
rect 15838 20816 15844 20828
rect 15896 20856 15902 20868
rect 16114 20856 16120 20868
rect 15896 20828 16120 20856
rect 15896 20816 15902 20828
rect 16114 20816 16120 20828
rect 16172 20816 16178 20868
rect 14642 20788 14648 20800
rect 12406 20760 14648 20788
rect 10965 20751 11023 20757
rect 14642 20748 14648 20760
rect 14700 20748 14706 20800
rect 14826 20748 14832 20800
rect 14884 20788 14890 20800
rect 16025 20791 16083 20797
rect 16025 20788 16037 20791
rect 14884 20760 16037 20788
rect 14884 20748 14890 20760
rect 16025 20757 16037 20760
rect 16071 20757 16083 20791
rect 16025 20751 16083 20757
rect 16482 20748 16488 20800
rect 16540 20748 16546 20800
rect 16684 20788 16712 20887
rect 19518 20884 19524 20936
rect 19576 20924 19582 20936
rect 20165 20927 20223 20933
rect 20165 20924 20177 20927
rect 19576 20896 20177 20924
rect 19576 20884 19582 20896
rect 20165 20893 20177 20896
rect 20211 20893 20223 20927
rect 20165 20887 20223 20893
rect 20714 20884 20720 20936
rect 20772 20924 20778 20936
rect 21085 20927 21143 20933
rect 21085 20924 21097 20927
rect 20772 20896 21097 20924
rect 20772 20884 20778 20896
rect 21085 20893 21097 20896
rect 21131 20893 21143 20927
rect 21085 20887 21143 20893
rect 18690 20856 18696 20868
rect 18630 20828 18696 20856
rect 18690 20816 18696 20828
rect 18748 20816 18754 20868
rect 20806 20856 20812 20868
rect 20180 20828 20812 20856
rect 20180 20788 20208 20828
rect 20806 20816 20812 20828
rect 20864 20816 20870 20868
rect 21818 20816 21824 20868
rect 21876 20816 21882 20868
rect 16684 20760 20208 20788
rect 20257 20791 20315 20797
rect 20257 20757 20269 20791
rect 20303 20788 20315 20791
rect 22002 20788 22008 20800
rect 20303 20760 22008 20788
rect 20303 20757 20315 20760
rect 20257 20751 20315 20757
rect 22002 20748 22008 20760
rect 22060 20748 22066 20800
rect 22094 20748 22100 20800
rect 22152 20788 22158 20800
rect 22664 20788 22692 20964
rect 23845 20961 23857 20964
rect 23891 20961 23903 20995
rect 23845 20955 23903 20961
rect 25225 20995 25283 21001
rect 25225 20961 25237 20995
rect 25271 20961 25283 20995
rect 25225 20955 25283 20961
rect 26326 20952 26332 21004
rect 26384 20992 26390 21004
rect 26421 20995 26479 21001
rect 26421 20992 26433 20995
rect 26384 20964 26433 20992
rect 26384 20952 26390 20964
rect 26421 20961 26433 20964
rect 26467 20961 26479 20995
rect 26421 20955 26479 20961
rect 27798 20952 27804 21004
rect 27856 20992 27862 21004
rect 28442 20992 28448 21004
rect 27856 20964 28448 20992
rect 27856 20952 27862 20964
rect 28442 20952 28448 20964
rect 28500 20952 28506 21004
rect 28905 20995 28963 21001
rect 28905 20961 28917 20995
rect 28951 20992 28963 20995
rect 29362 20992 29368 21004
rect 28951 20964 29368 20992
rect 28951 20961 28963 20964
rect 28905 20955 28963 20961
rect 29362 20952 29368 20964
rect 29420 20952 29426 21004
rect 31312 21001 31340 21032
rect 34790 21020 34796 21032
rect 34848 21020 34854 21072
rect 39224 21032 40632 21060
rect 39224 21004 39252 21032
rect 40604 21004 40632 21032
rect 40696 21032 41828 21060
rect 31297 20995 31355 21001
rect 31297 20961 31309 20995
rect 31343 20961 31355 20995
rect 31297 20955 31355 20961
rect 31481 20995 31539 21001
rect 31481 20961 31493 20995
rect 31527 20992 31539 20995
rect 33410 20992 33416 21004
rect 31527 20964 33416 20992
rect 31527 20961 31539 20964
rect 31481 20955 31539 20961
rect 33410 20952 33416 20964
rect 33468 20952 33474 21004
rect 33686 20952 33692 21004
rect 33744 20992 33750 21004
rect 33781 20995 33839 21001
rect 33781 20992 33793 20995
rect 33744 20964 33793 20992
rect 33744 20952 33750 20964
rect 33781 20961 33793 20964
rect 33827 20961 33839 20995
rect 33781 20955 33839 20961
rect 34606 20952 34612 21004
rect 34664 20992 34670 21004
rect 34885 20995 34943 21001
rect 34885 20992 34897 20995
rect 34664 20964 34897 20992
rect 34664 20952 34670 20964
rect 34885 20961 34897 20964
rect 34931 20961 34943 20995
rect 34885 20955 34943 20961
rect 35158 20952 35164 21004
rect 35216 20952 35222 21004
rect 35894 20952 35900 21004
rect 35952 20992 35958 21004
rect 36633 20995 36691 21001
rect 36633 20992 36645 20995
rect 35952 20964 36645 20992
rect 35952 20952 35958 20964
rect 36633 20961 36645 20964
rect 36679 20961 36691 20995
rect 36633 20955 36691 20961
rect 37274 20952 37280 21004
rect 37332 20992 37338 21004
rect 37734 20992 37740 21004
rect 37332 20964 37740 20992
rect 37332 20952 37338 20964
rect 37734 20952 37740 20964
rect 37792 20952 37798 21004
rect 38013 20995 38071 21001
rect 38013 20961 38025 20995
rect 38059 20992 38071 20995
rect 39206 20992 39212 21004
rect 38059 20964 39212 20992
rect 38059 20961 38071 20964
rect 38013 20955 38071 20961
rect 39206 20952 39212 20964
rect 39264 20952 39270 21004
rect 40494 20952 40500 21004
rect 40552 20952 40558 21004
rect 40586 20952 40592 21004
rect 40644 20952 40650 21004
rect 23661 20927 23719 20933
rect 23661 20893 23673 20927
rect 23707 20924 23719 20927
rect 24762 20924 24768 20936
rect 23707 20896 24768 20924
rect 23707 20893 23719 20896
rect 23661 20887 23719 20893
rect 24762 20884 24768 20896
rect 24820 20884 24826 20936
rect 25038 20884 25044 20936
rect 25096 20884 25102 20936
rect 25314 20884 25320 20936
rect 25372 20924 25378 20936
rect 27249 20927 27307 20933
rect 27249 20924 27261 20927
rect 25372 20896 27261 20924
rect 25372 20884 25378 20896
rect 27249 20893 27261 20896
rect 27295 20893 27307 20927
rect 27249 20887 27307 20893
rect 29917 20927 29975 20933
rect 29917 20893 29929 20927
rect 29963 20924 29975 20927
rect 30282 20924 30288 20936
rect 29963 20896 30288 20924
rect 29963 20893 29975 20896
rect 29917 20887 29975 20893
rect 30282 20884 30288 20896
rect 30340 20884 30346 20936
rect 32214 20884 32220 20936
rect 32272 20884 32278 20936
rect 33597 20927 33655 20933
rect 33597 20893 33609 20927
rect 33643 20924 33655 20927
rect 34698 20924 34704 20936
rect 33643 20896 34704 20924
rect 33643 20893 33655 20896
rect 33597 20887 33655 20893
rect 34698 20884 34704 20896
rect 34756 20884 34762 20936
rect 39482 20924 39488 20936
rect 39146 20896 39488 20924
rect 39482 20884 39488 20896
rect 39540 20884 39546 20936
rect 39758 20884 39764 20936
rect 39816 20924 39822 20936
rect 40696 20924 40724 21032
rect 41800 21001 41828 21032
rect 41785 20995 41843 21001
rect 41785 20961 41797 20995
rect 41831 20961 41843 20995
rect 41785 20955 41843 20961
rect 41693 20927 41751 20933
rect 41693 20924 41705 20927
rect 39816 20896 40724 20924
rect 41386 20896 41705 20924
rect 39816 20884 39822 20896
rect 23750 20816 23756 20868
rect 23808 20816 23814 20868
rect 28813 20859 28871 20865
rect 28813 20856 28825 20859
rect 24596 20828 28825 20856
rect 22152 20760 22692 20788
rect 22152 20748 22158 20760
rect 23290 20748 23296 20800
rect 23348 20748 23354 20800
rect 24596 20797 24624 20828
rect 28813 20825 28825 20828
rect 28859 20825 28871 20859
rect 28813 20819 28871 20825
rect 29362 20816 29368 20868
rect 29420 20856 29426 20868
rect 31478 20856 31484 20868
rect 29420 20828 31484 20856
rect 29420 20816 29426 20828
rect 31478 20816 31484 20828
rect 31536 20816 31542 20868
rect 33134 20816 33140 20868
rect 33192 20856 33198 20868
rect 33192 20828 33732 20856
rect 33192 20816 33198 20828
rect 24581 20791 24639 20797
rect 24581 20757 24593 20791
rect 24627 20757 24639 20791
rect 24581 20751 24639 20757
rect 24946 20748 24952 20800
rect 25004 20748 25010 20800
rect 25314 20748 25320 20800
rect 25372 20788 25378 20800
rect 25869 20791 25927 20797
rect 25869 20788 25881 20791
rect 25372 20760 25881 20788
rect 25372 20748 25378 20760
rect 25869 20757 25881 20760
rect 25915 20757 25927 20791
rect 25869 20751 25927 20757
rect 26234 20748 26240 20800
rect 26292 20748 26298 20800
rect 26329 20791 26387 20797
rect 26329 20757 26341 20791
rect 26375 20788 26387 20791
rect 26418 20788 26424 20800
rect 26375 20760 26424 20788
rect 26375 20757 26387 20760
rect 26329 20751 26387 20757
rect 26418 20748 26424 20760
rect 26476 20748 26482 20800
rect 26878 20748 26884 20800
rect 26936 20788 26942 20800
rect 27065 20791 27123 20797
rect 27065 20788 27077 20791
rect 26936 20760 27077 20788
rect 26936 20748 26942 20760
rect 27065 20757 27077 20760
rect 27111 20757 27123 20791
rect 27065 20751 27123 20757
rect 27614 20748 27620 20800
rect 27672 20788 27678 20800
rect 28626 20788 28632 20800
rect 27672 20760 28632 20788
rect 27672 20748 27678 20760
rect 28626 20748 28632 20760
rect 28684 20748 28690 20800
rect 28718 20748 28724 20800
rect 28776 20748 28782 20800
rect 31202 20748 31208 20800
rect 31260 20748 31266 20800
rect 32030 20748 32036 20800
rect 32088 20748 32094 20800
rect 32490 20748 32496 20800
rect 32548 20788 32554 20800
rect 32858 20788 32864 20800
rect 32548 20760 32864 20788
rect 32548 20748 32554 20760
rect 32858 20748 32864 20760
rect 32916 20748 32922 20800
rect 33704 20797 33732 20828
rect 34422 20816 34428 20868
rect 34480 20856 34486 20868
rect 37918 20856 37924 20868
rect 34480 20828 35650 20856
rect 36464 20828 37924 20856
rect 34480 20816 34486 20828
rect 33689 20791 33747 20797
rect 33689 20757 33701 20791
rect 33735 20788 33747 20791
rect 36464 20788 36492 20828
rect 37918 20816 37924 20828
rect 37976 20816 37982 20868
rect 39942 20816 39948 20868
rect 40000 20856 40006 20868
rect 41386 20856 41414 20896
rect 41693 20893 41705 20896
rect 41739 20893 41751 20927
rect 41693 20887 41751 20893
rect 49050 20884 49056 20936
rect 49108 20884 49114 20936
rect 40000 20828 41414 20856
rect 41601 20859 41659 20865
rect 40000 20816 40006 20828
rect 41601 20825 41613 20859
rect 41647 20856 41659 20859
rect 48406 20856 48412 20868
rect 41647 20828 48412 20856
rect 41647 20825 41659 20828
rect 41601 20819 41659 20825
rect 48406 20816 48412 20828
rect 48464 20816 48470 20868
rect 33735 20760 36492 20788
rect 33735 20757 33747 20760
rect 33689 20751 33747 20757
rect 38286 20748 38292 20800
rect 38344 20788 38350 20800
rect 39485 20791 39543 20797
rect 39485 20788 39497 20791
rect 38344 20760 39497 20788
rect 38344 20748 38350 20760
rect 39485 20757 39497 20760
rect 39531 20757 39543 20791
rect 39485 20751 39543 20757
rect 40405 20791 40463 20797
rect 40405 20757 40417 20791
rect 40451 20788 40463 20791
rect 41233 20791 41291 20797
rect 41233 20788 41245 20791
rect 40451 20760 41245 20788
rect 40451 20757 40463 20760
rect 40405 20751 40463 20757
rect 41233 20757 41245 20760
rect 41279 20757 41291 20791
rect 41233 20751 41291 20757
rect 1104 20698 49864 20720
rect 1104 20646 7950 20698
rect 8002 20646 8014 20698
rect 8066 20646 8078 20698
rect 8130 20646 8142 20698
rect 8194 20646 8206 20698
rect 8258 20646 17950 20698
rect 18002 20646 18014 20698
rect 18066 20646 18078 20698
rect 18130 20646 18142 20698
rect 18194 20646 18206 20698
rect 18258 20646 27950 20698
rect 28002 20646 28014 20698
rect 28066 20646 28078 20698
rect 28130 20646 28142 20698
rect 28194 20646 28206 20698
rect 28258 20646 37950 20698
rect 38002 20646 38014 20698
rect 38066 20646 38078 20698
rect 38130 20646 38142 20698
rect 38194 20646 38206 20698
rect 38258 20646 47950 20698
rect 48002 20646 48014 20698
rect 48066 20646 48078 20698
rect 48130 20646 48142 20698
rect 48194 20646 48206 20698
rect 48258 20646 49864 20698
rect 1104 20624 49864 20646
rect 5261 20587 5319 20593
rect 5261 20553 5273 20587
rect 5307 20584 5319 20587
rect 6546 20584 6552 20596
rect 5307 20556 6552 20584
rect 5307 20553 5319 20556
rect 5261 20547 5319 20553
rect 6546 20544 6552 20556
rect 6604 20544 6610 20596
rect 8294 20544 8300 20596
rect 8352 20584 8358 20596
rect 8389 20587 8447 20593
rect 8389 20584 8401 20587
rect 8352 20556 8401 20584
rect 8352 20544 8358 20556
rect 8389 20553 8401 20556
rect 8435 20553 8447 20587
rect 8389 20547 8447 20553
rect 9582 20544 9588 20596
rect 9640 20584 9646 20596
rect 9953 20587 10011 20593
rect 9953 20584 9965 20587
rect 9640 20556 9965 20584
rect 9640 20544 9646 20556
rect 9953 20553 9965 20556
rect 9999 20553 10011 20587
rect 9953 20547 10011 20553
rect 10410 20544 10416 20596
rect 10468 20584 10474 20596
rect 10597 20587 10655 20593
rect 10597 20584 10609 20587
rect 10468 20556 10609 20584
rect 10468 20544 10474 20556
rect 10597 20553 10609 20556
rect 10643 20584 10655 20587
rect 10686 20584 10692 20596
rect 10643 20556 10692 20584
rect 10643 20553 10655 20556
rect 10597 20547 10655 20553
rect 10686 20544 10692 20556
rect 10744 20544 10750 20596
rect 11330 20544 11336 20596
rect 11388 20584 11394 20596
rect 11388 20556 12848 20584
rect 11388 20544 11394 20556
rect 11238 20516 11244 20528
rect 10152 20488 11244 20516
rect 1762 20408 1768 20460
rect 1820 20408 1826 20460
rect 3602 20408 3608 20460
rect 3660 20408 3666 20460
rect 5445 20451 5503 20457
rect 5445 20417 5457 20451
rect 5491 20448 5503 20451
rect 6362 20448 6368 20460
rect 5491 20420 6368 20448
rect 5491 20417 5503 20420
rect 5445 20411 5503 20417
rect 6362 20408 6368 20420
rect 6420 20408 6426 20460
rect 6454 20408 6460 20460
rect 6512 20448 6518 20460
rect 6549 20451 6607 20457
rect 6549 20448 6561 20451
rect 6512 20420 6561 20448
rect 6512 20408 6518 20420
rect 6549 20417 6561 20420
rect 6595 20417 6607 20451
rect 6549 20411 6607 20417
rect 8573 20451 8631 20457
rect 8573 20417 8585 20451
rect 8619 20417 8631 20451
rect 8573 20411 8631 20417
rect 9309 20451 9367 20457
rect 9309 20417 9321 20451
rect 9355 20448 9367 20451
rect 10042 20448 10048 20460
rect 9355 20420 10048 20448
rect 9355 20417 9367 20420
rect 9309 20411 9367 20417
rect 2777 20383 2835 20389
rect 2777 20349 2789 20383
rect 2823 20380 2835 20383
rect 2866 20380 2872 20392
rect 2823 20352 2872 20380
rect 2823 20349 2835 20352
rect 2777 20343 2835 20349
rect 2866 20340 2872 20352
rect 2924 20340 2930 20392
rect 3878 20340 3884 20392
rect 3936 20340 3942 20392
rect 5718 20340 5724 20392
rect 5776 20380 5782 20392
rect 7009 20383 7067 20389
rect 7009 20380 7021 20383
rect 5776 20352 7021 20380
rect 5776 20340 5782 20352
rect 7009 20349 7021 20352
rect 7055 20349 7067 20383
rect 8588 20380 8616 20411
rect 10042 20408 10048 20420
rect 10100 20408 10106 20460
rect 10152 20457 10180 20488
rect 11238 20476 11244 20488
rect 11296 20476 11302 20528
rect 11422 20476 11428 20528
rect 11480 20516 11486 20528
rect 12713 20519 12771 20525
rect 12713 20516 12725 20519
rect 11480 20488 12725 20516
rect 11480 20476 11486 20488
rect 12713 20485 12725 20488
rect 12759 20485 12771 20519
rect 12820 20516 12848 20556
rect 13630 20544 13636 20596
rect 13688 20584 13694 20596
rect 14093 20587 14151 20593
rect 14093 20584 14105 20587
rect 13688 20556 14105 20584
rect 13688 20544 13694 20556
rect 14093 20553 14105 20556
rect 14139 20553 14151 20587
rect 14093 20547 14151 20553
rect 14366 20544 14372 20596
rect 14424 20584 14430 20596
rect 16209 20587 16267 20593
rect 16209 20584 16221 20587
rect 14424 20556 16221 20584
rect 14424 20544 14430 20556
rect 16209 20553 16221 20556
rect 16255 20553 16267 20587
rect 19150 20584 19156 20596
rect 16209 20547 16267 20553
rect 16316 20556 19156 20584
rect 15565 20519 15623 20525
rect 12820 20488 15516 20516
rect 12713 20479 12771 20485
rect 10137 20451 10195 20457
rect 10137 20417 10149 20451
rect 10183 20417 10195 20451
rect 10137 20411 10195 20417
rect 10781 20451 10839 20457
rect 10781 20417 10793 20451
rect 10827 20417 10839 20451
rect 10781 20411 10839 20417
rect 11793 20451 11851 20457
rect 11793 20417 11805 20451
rect 11839 20448 11851 20451
rect 11882 20448 11888 20460
rect 11839 20420 11888 20448
rect 11839 20417 11851 20420
rect 11793 20411 11851 20417
rect 9766 20380 9772 20392
rect 8588 20352 9772 20380
rect 7009 20343 7067 20349
rect 9766 20340 9772 20352
rect 9824 20340 9830 20392
rect 7650 20272 7656 20324
rect 7708 20312 7714 20324
rect 9125 20315 9183 20321
rect 9125 20312 9137 20315
rect 7708 20284 9137 20312
rect 7708 20272 7714 20284
rect 9125 20281 9137 20284
rect 9171 20281 9183 20315
rect 10796 20312 10824 20411
rect 11882 20408 11888 20420
rect 11940 20408 11946 20460
rect 12529 20451 12587 20457
rect 12529 20417 12541 20451
rect 12575 20448 12587 20451
rect 13630 20448 13636 20460
rect 12575 20420 13636 20448
rect 12575 20417 12587 20420
rect 12529 20411 12587 20417
rect 13630 20408 13636 20420
rect 13688 20408 13694 20460
rect 14185 20451 14243 20457
rect 14185 20417 14197 20451
rect 14231 20448 14243 20451
rect 14231 20420 15332 20448
rect 14231 20417 14243 20420
rect 14185 20411 14243 20417
rect 14369 20383 14427 20389
rect 12544 20352 14320 20380
rect 12544 20312 12572 20352
rect 13725 20315 13783 20321
rect 13725 20312 13737 20315
rect 10796 20284 12572 20312
rect 12636 20284 13737 20312
rect 9125 20275 9183 20281
rect 9674 20204 9680 20256
rect 9732 20244 9738 20256
rect 11885 20247 11943 20253
rect 11885 20244 11897 20247
rect 9732 20216 11897 20244
rect 9732 20204 9738 20216
rect 11885 20213 11897 20216
rect 11931 20213 11943 20247
rect 11885 20207 11943 20213
rect 11974 20204 11980 20256
rect 12032 20244 12038 20256
rect 12636 20244 12664 20284
rect 13725 20281 13737 20284
rect 13771 20281 13783 20315
rect 14292 20312 14320 20352
rect 14369 20349 14381 20383
rect 14415 20380 14427 20383
rect 14826 20380 14832 20392
rect 14415 20352 14832 20380
rect 14415 20349 14427 20352
rect 14369 20343 14427 20349
rect 14826 20340 14832 20352
rect 14884 20340 14890 20392
rect 15304 20380 15332 20420
rect 15378 20408 15384 20460
rect 15436 20408 15442 20460
rect 15488 20448 15516 20488
rect 15565 20485 15577 20519
rect 15611 20516 15623 20519
rect 15654 20516 15660 20528
rect 15611 20488 15660 20516
rect 15611 20485 15623 20488
rect 15565 20479 15623 20485
rect 15654 20476 15660 20488
rect 15712 20476 15718 20528
rect 16316 20516 16344 20556
rect 19150 20544 19156 20556
rect 19208 20544 19214 20596
rect 20622 20584 20628 20596
rect 19720 20556 20628 20584
rect 18690 20516 18696 20528
rect 15764 20488 16344 20516
rect 18538 20488 18696 20516
rect 15764 20448 15792 20488
rect 18690 20476 18696 20488
rect 18748 20516 18754 20528
rect 19426 20516 19432 20528
rect 18748 20488 19432 20516
rect 18748 20476 18754 20488
rect 19426 20476 19432 20488
rect 19484 20476 19490 20528
rect 15488 20420 15792 20448
rect 16114 20408 16120 20460
rect 16172 20408 16178 20460
rect 17034 20408 17040 20460
rect 17092 20408 17098 20460
rect 16758 20380 16764 20392
rect 15304 20352 16764 20380
rect 16758 20340 16764 20352
rect 16816 20340 16822 20392
rect 17313 20383 17371 20389
rect 17313 20349 17325 20383
rect 17359 20380 17371 20383
rect 17359 20352 19012 20380
rect 17359 20349 17371 20352
rect 17313 20343 17371 20349
rect 16850 20312 16856 20324
rect 14292 20284 16856 20312
rect 13725 20275 13783 20281
rect 16850 20272 16856 20284
rect 16908 20272 16914 20324
rect 18984 20256 19012 20352
rect 19610 20340 19616 20392
rect 19668 20380 19674 20392
rect 19720 20389 19748 20556
rect 20622 20544 20628 20556
rect 20680 20544 20686 20596
rect 20990 20544 20996 20596
rect 21048 20584 21054 20596
rect 21453 20587 21511 20593
rect 21453 20584 21465 20587
rect 21048 20556 21465 20584
rect 21048 20544 21054 20556
rect 21453 20553 21465 20556
rect 21499 20584 21511 20587
rect 22094 20584 22100 20596
rect 21499 20556 22100 20584
rect 21499 20553 21511 20556
rect 21453 20547 21511 20553
rect 22094 20544 22100 20556
rect 22152 20544 22158 20596
rect 25406 20584 25412 20596
rect 22388 20556 25412 20584
rect 21266 20516 21272 20528
rect 21206 20488 21272 20516
rect 21266 20476 21272 20488
rect 21324 20516 21330 20528
rect 21818 20516 21824 20528
rect 21324 20488 21824 20516
rect 21324 20476 21330 20488
rect 21818 20476 21824 20488
rect 21876 20476 21882 20528
rect 22388 20448 22416 20556
rect 25406 20544 25412 20556
rect 25464 20544 25470 20596
rect 26602 20544 26608 20596
rect 26660 20584 26666 20596
rect 27154 20584 27160 20596
rect 26660 20556 27160 20584
rect 26660 20544 26666 20556
rect 27154 20544 27160 20556
rect 27212 20584 27218 20596
rect 27212 20556 27660 20584
rect 27212 20544 27218 20556
rect 22465 20519 22523 20525
rect 22465 20485 22477 20519
rect 22511 20516 22523 20519
rect 22554 20516 22560 20528
rect 22511 20488 22560 20516
rect 22511 20485 22523 20488
rect 22465 20479 22523 20485
rect 22554 20476 22560 20488
rect 22612 20476 22618 20528
rect 23658 20476 23664 20528
rect 23716 20516 23722 20528
rect 24118 20516 24124 20528
rect 23716 20488 24124 20516
rect 23716 20476 23722 20488
rect 24118 20476 24124 20488
rect 24176 20476 24182 20528
rect 26620 20516 26648 20544
rect 25346 20488 26648 20516
rect 27430 20476 27436 20528
rect 27488 20516 27494 20528
rect 27525 20519 27583 20525
rect 27525 20516 27537 20519
rect 27488 20488 27537 20516
rect 27488 20476 27494 20488
rect 27525 20485 27537 20488
rect 27571 20485 27583 20519
rect 27632 20516 27660 20556
rect 27706 20544 27712 20596
rect 27764 20584 27770 20596
rect 28534 20584 28540 20596
rect 27764 20556 28540 20584
rect 27764 20544 27770 20556
rect 28534 20544 28540 20556
rect 28592 20584 28598 20596
rect 28592 20556 28856 20584
rect 28592 20544 28598 20556
rect 27632 20488 28014 20516
rect 27525 20479 27583 20485
rect 23750 20448 23756 20460
rect 22066 20420 22416 20448
rect 22572 20420 23756 20448
rect 19705 20383 19763 20389
rect 19705 20380 19717 20383
rect 19668 20352 19717 20380
rect 19668 20340 19674 20352
rect 19705 20349 19717 20352
rect 19751 20349 19763 20383
rect 19705 20343 19763 20349
rect 19981 20383 20039 20389
rect 19981 20349 19993 20383
rect 20027 20380 20039 20383
rect 21358 20380 21364 20392
rect 20027 20352 21364 20380
rect 20027 20349 20039 20352
rect 19981 20343 20039 20349
rect 21358 20340 21364 20352
rect 21416 20380 21422 20392
rect 22066 20380 22094 20420
rect 22572 20389 22600 20420
rect 23750 20408 23756 20420
rect 23808 20408 23814 20460
rect 25498 20408 25504 20460
rect 25556 20448 25562 20460
rect 26237 20451 26295 20457
rect 26237 20448 26249 20451
rect 25556 20420 26249 20448
rect 25556 20408 25562 20420
rect 26237 20417 26249 20420
rect 26283 20417 26295 20451
rect 28828 20448 28856 20556
rect 28994 20544 29000 20596
rect 29052 20544 29058 20596
rect 29825 20587 29883 20593
rect 29825 20553 29837 20587
rect 29871 20553 29883 20587
rect 29825 20547 29883 20553
rect 29840 20460 29868 20547
rect 30834 20544 30840 20596
rect 30892 20584 30898 20596
rect 31021 20587 31079 20593
rect 31021 20584 31033 20587
rect 30892 20556 31033 20584
rect 30892 20544 30898 20556
rect 31021 20553 31033 20556
rect 31067 20553 31079 20587
rect 31021 20547 31079 20553
rect 31110 20544 31116 20596
rect 31168 20544 31174 20596
rect 33410 20544 33416 20596
rect 33468 20584 33474 20596
rect 34057 20587 34115 20593
rect 34057 20584 34069 20587
rect 33468 20556 34069 20584
rect 33468 20544 33474 20556
rect 34057 20553 34069 20556
rect 34103 20553 34115 20587
rect 34057 20547 34115 20553
rect 34517 20587 34575 20593
rect 34517 20553 34529 20587
rect 34563 20584 34575 20587
rect 35802 20584 35808 20596
rect 34563 20556 35808 20584
rect 34563 20553 34575 20556
rect 34517 20547 34575 20553
rect 35802 20544 35808 20556
rect 35860 20544 35866 20596
rect 40402 20544 40408 20596
rect 40460 20544 40466 20596
rect 32490 20476 32496 20528
rect 32548 20516 32554 20528
rect 32585 20519 32643 20525
rect 32585 20516 32597 20519
rect 32548 20488 32597 20516
rect 32548 20476 32554 20488
rect 32585 20485 32597 20488
rect 32631 20485 32643 20519
rect 33870 20516 33876 20528
rect 33810 20488 33876 20516
rect 32585 20479 32643 20485
rect 33870 20476 33876 20488
rect 33928 20516 33934 20528
rect 34422 20516 34428 20528
rect 33928 20488 34428 20516
rect 33928 20476 33934 20488
rect 34422 20476 34428 20488
rect 34480 20476 34486 20528
rect 34606 20476 34612 20528
rect 34664 20516 34670 20528
rect 35894 20516 35900 20528
rect 34664 20488 35900 20516
rect 34664 20476 34670 20488
rect 35894 20476 35900 20488
rect 35952 20476 35958 20528
rect 37918 20516 37924 20528
rect 36004 20488 37924 20516
rect 29638 20448 29644 20460
rect 28828 20420 29644 20448
rect 26237 20411 26295 20417
rect 29638 20408 29644 20420
rect 29696 20408 29702 20460
rect 29822 20408 29828 20460
rect 29880 20408 29886 20460
rect 34514 20408 34520 20460
rect 34572 20448 34578 20460
rect 34885 20452 34943 20457
rect 34808 20451 34943 20452
rect 34808 20448 34897 20451
rect 34572 20424 34897 20448
rect 34572 20420 34836 20424
rect 34572 20408 34578 20420
rect 34885 20417 34897 20424
rect 34931 20417 34943 20451
rect 34885 20411 34943 20417
rect 34992 20448 35296 20452
rect 35342 20448 35348 20460
rect 34992 20424 35348 20448
rect 21416 20352 22094 20380
rect 22557 20383 22615 20389
rect 21416 20340 21422 20352
rect 22557 20349 22569 20383
rect 22603 20349 22615 20383
rect 22557 20343 22615 20349
rect 22649 20383 22707 20389
rect 22649 20349 22661 20383
rect 22695 20349 22707 20383
rect 22649 20343 22707 20349
rect 22370 20272 22376 20324
rect 22428 20312 22434 20324
rect 22664 20312 22692 20343
rect 23382 20340 23388 20392
rect 23440 20380 23446 20392
rect 23845 20383 23903 20389
rect 23845 20380 23857 20383
rect 23440 20352 23857 20380
rect 23440 20340 23446 20352
rect 23845 20349 23857 20352
rect 23891 20349 23903 20383
rect 23845 20343 23903 20349
rect 24118 20340 24124 20392
rect 24176 20340 24182 20392
rect 25590 20340 25596 20392
rect 25648 20380 25654 20392
rect 26970 20380 26976 20392
rect 25648 20352 26976 20380
rect 25648 20340 25654 20352
rect 26970 20340 26976 20352
rect 27028 20340 27034 20392
rect 27249 20383 27307 20389
rect 27249 20349 27261 20383
rect 27295 20349 27307 20383
rect 27249 20343 27307 20349
rect 22428 20284 22692 20312
rect 22428 20272 22434 20284
rect 25222 20272 25228 20324
rect 25280 20312 25286 20324
rect 26050 20312 26056 20324
rect 25280 20284 26056 20312
rect 25280 20272 25286 20284
rect 26050 20272 26056 20284
rect 26108 20272 26114 20324
rect 12032 20216 12664 20244
rect 12032 20204 12038 20216
rect 12710 20204 12716 20256
rect 12768 20244 12774 20256
rect 18414 20244 18420 20256
rect 12768 20216 18420 20244
rect 12768 20204 12774 20216
rect 18414 20204 18420 20216
rect 18472 20204 18478 20256
rect 18782 20204 18788 20256
rect 18840 20204 18846 20256
rect 18966 20204 18972 20256
rect 19024 20244 19030 20256
rect 21726 20244 21732 20256
rect 19024 20216 21732 20244
rect 19024 20204 19030 20216
rect 21726 20204 21732 20216
rect 21784 20204 21790 20256
rect 21910 20204 21916 20256
rect 21968 20244 21974 20256
rect 22097 20247 22155 20253
rect 22097 20244 22109 20247
rect 21968 20216 22109 20244
rect 21968 20204 21974 20216
rect 22097 20213 22109 20216
rect 22143 20213 22155 20247
rect 22097 20207 22155 20213
rect 23658 20204 23664 20256
rect 23716 20244 23722 20256
rect 25590 20244 25596 20256
rect 23716 20216 25596 20244
rect 23716 20204 23722 20216
rect 25590 20204 25596 20216
rect 25648 20204 25654 20256
rect 27264 20244 27292 20343
rect 27890 20340 27896 20392
rect 27948 20380 27954 20392
rect 29362 20380 29368 20392
rect 27948 20352 29368 20380
rect 27948 20340 27954 20352
rect 29362 20340 29368 20352
rect 29420 20340 29426 20392
rect 29914 20340 29920 20392
rect 29972 20340 29978 20392
rect 30098 20340 30104 20392
rect 30156 20340 30162 20392
rect 30190 20340 30196 20392
rect 30248 20380 30254 20392
rect 31205 20383 31263 20389
rect 31205 20380 31217 20383
rect 30248 20352 31217 20380
rect 30248 20340 30254 20352
rect 31205 20349 31217 20352
rect 31251 20349 31263 20383
rect 31570 20380 31576 20392
rect 31205 20343 31263 20349
rect 31312 20352 31576 20380
rect 31312 20312 31340 20352
rect 31570 20340 31576 20352
rect 31628 20380 31634 20392
rect 32309 20383 32367 20389
rect 32309 20380 32321 20383
rect 31628 20352 32321 20380
rect 31628 20340 31634 20352
rect 32309 20349 32321 20352
rect 32355 20349 32367 20383
rect 32309 20343 32367 20349
rect 32582 20340 32588 20392
rect 32640 20380 32646 20392
rect 33594 20380 33600 20392
rect 32640 20352 33600 20380
rect 32640 20340 32646 20352
rect 33594 20340 33600 20352
rect 33652 20340 33658 20392
rect 34992 20389 35020 20424
rect 35268 20420 35348 20424
rect 35342 20408 35348 20420
rect 35400 20448 35406 20460
rect 36004 20448 36032 20488
rect 37918 20476 37924 20488
rect 37976 20476 37982 20528
rect 38013 20519 38071 20525
rect 38013 20485 38025 20519
rect 38059 20516 38071 20519
rect 38286 20516 38292 20528
rect 38059 20488 38292 20516
rect 38059 20485 38071 20488
rect 38013 20479 38071 20485
rect 38286 20476 38292 20488
rect 38344 20476 38350 20528
rect 39482 20516 39488 20528
rect 39238 20488 39488 20516
rect 39482 20476 39488 20488
rect 39540 20476 39546 20528
rect 35400 20420 36032 20448
rect 35400 20408 35406 20420
rect 36078 20408 36084 20460
rect 36136 20448 36142 20460
rect 36449 20451 36507 20457
rect 36449 20448 36461 20451
rect 36136 20420 36461 20448
rect 36136 20408 36142 20420
rect 36449 20417 36461 20420
rect 36495 20417 36507 20451
rect 36449 20411 36507 20417
rect 36541 20451 36599 20457
rect 36541 20417 36553 20451
rect 36587 20448 36599 20451
rect 37550 20448 37556 20460
rect 36587 20420 37556 20448
rect 36587 20417 36599 20420
rect 36541 20411 36599 20417
rect 37550 20408 37556 20420
rect 37608 20408 37614 20460
rect 37734 20408 37740 20460
rect 37792 20408 37798 20460
rect 40310 20408 40316 20460
rect 40368 20408 40374 20460
rect 45370 20448 45376 20460
rect 40420 20420 45376 20448
rect 34977 20383 35035 20389
rect 34977 20349 34989 20383
rect 35023 20349 35035 20383
rect 34977 20343 35035 20349
rect 35158 20340 35164 20392
rect 35216 20340 35222 20392
rect 36725 20383 36783 20389
rect 36725 20349 36737 20383
rect 36771 20380 36783 20383
rect 37642 20380 37648 20392
rect 36771 20352 37648 20380
rect 36771 20349 36783 20352
rect 36725 20343 36783 20349
rect 37642 20340 37648 20352
rect 37700 20340 37706 20392
rect 40420 20380 40448 20420
rect 45370 20408 45376 20420
rect 45428 20408 45434 20460
rect 48590 20408 48596 20460
rect 48648 20408 48654 20460
rect 49050 20408 49056 20460
rect 49108 20408 49114 20460
rect 37844 20352 40448 20380
rect 36081 20315 36139 20321
rect 36081 20312 36093 20315
rect 29380 20284 31340 20312
rect 33888 20284 36093 20312
rect 29380 20244 29408 20284
rect 27264 20216 29408 20244
rect 29457 20247 29515 20253
rect 29457 20213 29469 20247
rect 29503 20244 29515 20247
rect 30558 20244 30564 20256
rect 29503 20216 30564 20244
rect 29503 20213 29515 20216
rect 29457 20207 29515 20213
rect 30558 20204 30564 20216
rect 30616 20204 30622 20256
rect 30653 20247 30711 20253
rect 30653 20213 30665 20247
rect 30699 20244 30711 20247
rect 31110 20244 31116 20256
rect 30699 20216 31116 20244
rect 30699 20213 30711 20216
rect 30653 20207 30711 20213
rect 31110 20204 31116 20216
rect 31168 20204 31174 20256
rect 31294 20204 31300 20256
rect 31352 20244 31358 20256
rect 33888 20244 33916 20284
rect 36081 20281 36093 20284
rect 36127 20281 36139 20315
rect 36081 20275 36139 20281
rect 31352 20216 33916 20244
rect 31352 20204 31358 20216
rect 34054 20204 34060 20256
rect 34112 20244 34118 20256
rect 37844 20244 37872 20352
rect 40494 20340 40500 20392
rect 40552 20340 40558 20392
rect 41386 20352 45554 20380
rect 39485 20315 39543 20321
rect 39485 20281 39497 20315
rect 39531 20312 39543 20315
rect 40126 20312 40132 20324
rect 39531 20284 40132 20312
rect 39531 20281 39543 20284
rect 39485 20275 39543 20281
rect 34112 20216 37872 20244
rect 34112 20204 34118 20216
rect 38654 20204 38660 20256
rect 38712 20244 38718 20256
rect 39500 20244 39528 20275
rect 40126 20272 40132 20284
rect 40184 20272 40190 20324
rect 40402 20272 40408 20324
rect 40460 20312 40466 20324
rect 41386 20312 41414 20352
rect 40460 20284 41414 20312
rect 45526 20312 45554 20352
rect 49237 20315 49295 20321
rect 49237 20312 49249 20315
rect 45526 20284 49249 20312
rect 40460 20272 40466 20284
rect 49237 20281 49249 20284
rect 49283 20281 49295 20315
rect 49237 20275 49295 20281
rect 38712 20216 39528 20244
rect 39945 20247 40003 20253
rect 38712 20204 38718 20216
rect 39945 20213 39957 20247
rect 39991 20244 40003 20247
rect 40862 20244 40868 20256
rect 39991 20216 40868 20244
rect 39991 20213 40003 20216
rect 39945 20207 40003 20213
rect 40862 20204 40868 20216
rect 40920 20204 40926 20256
rect 48406 20204 48412 20256
rect 48464 20204 48470 20256
rect 1104 20154 49864 20176
rect 1104 20102 2950 20154
rect 3002 20102 3014 20154
rect 3066 20102 3078 20154
rect 3130 20102 3142 20154
rect 3194 20102 3206 20154
rect 3258 20102 12950 20154
rect 13002 20102 13014 20154
rect 13066 20102 13078 20154
rect 13130 20102 13142 20154
rect 13194 20102 13206 20154
rect 13258 20102 22950 20154
rect 23002 20102 23014 20154
rect 23066 20102 23078 20154
rect 23130 20102 23142 20154
rect 23194 20102 23206 20154
rect 23258 20102 32950 20154
rect 33002 20102 33014 20154
rect 33066 20102 33078 20154
rect 33130 20102 33142 20154
rect 33194 20102 33206 20154
rect 33258 20102 42950 20154
rect 43002 20102 43014 20154
rect 43066 20102 43078 20154
rect 43130 20102 43142 20154
rect 43194 20102 43206 20154
rect 43258 20102 49864 20154
rect 1104 20080 49864 20102
rect 2746 20012 14596 20040
rect 1765 19839 1823 19845
rect 1765 19805 1777 19839
rect 1811 19836 1823 19839
rect 2746 19836 2774 20012
rect 3602 19932 3608 19984
rect 3660 19972 3666 19984
rect 11517 19975 11575 19981
rect 11517 19972 11529 19975
rect 3660 19944 11529 19972
rect 3660 19932 3666 19944
rect 11517 19941 11529 19944
rect 11563 19941 11575 19975
rect 11517 19935 11575 19941
rect 13354 19932 13360 19984
rect 13412 19972 13418 19984
rect 13538 19972 13544 19984
rect 13412 19944 13544 19972
rect 13412 19932 13418 19944
rect 13538 19932 13544 19944
rect 13596 19932 13602 19984
rect 14568 19972 14596 20012
rect 14734 20000 14740 20052
rect 14792 20000 14798 20052
rect 16390 20000 16396 20052
rect 16448 20040 16454 20052
rect 16945 20043 17003 20049
rect 16945 20040 16957 20043
rect 16448 20012 16957 20040
rect 16448 20000 16454 20012
rect 16945 20009 16957 20012
rect 16991 20009 17003 20043
rect 23290 20040 23296 20052
rect 16945 20003 17003 20009
rect 18616 20012 23296 20040
rect 16853 19975 16911 19981
rect 16853 19972 16865 19975
rect 14568 19944 16865 19972
rect 16853 19941 16865 19944
rect 16899 19941 16911 19975
rect 16853 19935 16911 19941
rect 17310 19932 17316 19984
rect 17368 19972 17374 19984
rect 17368 19944 17632 19972
rect 17368 19932 17374 19944
rect 4890 19864 4896 19916
rect 4948 19864 4954 19916
rect 5920 19876 6132 19904
rect 1811 19808 2774 19836
rect 4065 19839 4123 19845
rect 1811 19805 1823 19808
rect 1765 19799 1823 19805
rect 4065 19805 4077 19839
rect 4111 19836 4123 19839
rect 5920 19836 5948 19876
rect 4111 19808 5948 19836
rect 5997 19839 6055 19845
rect 4111 19805 4123 19808
rect 4065 19799 4123 19805
rect 5997 19805 6009 19839
rect 6043 19805 6055 19839
rect 6104 19836 6132 19876
rect 6270 19864 6276 19916
rect 6328 19864 6334 19916
rect 9306 19904 9312 19916
rect 6656 19876 9312 19904
rect 6656 19836 6684 19876
rect 9306 19864 9312 19876
rect 9364 19864 9370 19916
rect 10781 19907 10839 19913
rect 10781 19873 10793 19907
rect 10827 19904 10839 19907
rect 10827 19876 11376 19904
rect 10827 19873 10839 19876
rect 10781 19867 10839 19873
rect 11348 19848 11376 19876
rect 16298 19864 16304 19916
rect 16356 19904 16362 19916
rect 17497 19907 17555 19913
rect 17497 19904 17509 19907
rect 16356 19876 17509 19904
rect 16356 19864 16362 19876
rect 17497 19873 17509 19876
rect 17543 19873 17555 19907
rect 17497 19867 17555 19873
rect 6104 19808 6684 19836
rect 7929 19839 7987 19845
rect 5997 19799 6055 19805
rect 7929 19805 7941 19839
rect 7975 19836 7987 19839
rect 9490 19836 9496 19848
rect 7975 19808 9496 19836
rect 7975 19805 7987 19808
rect 7929 19799 7987 19805
rect 2774 19728 2780 19780
rect 2832 19728 2838 19780
rect 6012 19700 6040 19799
rect 9490 19796 9496 19808
rect 9548 19796 9554 19848
rect 10045 19839 10103 19845
rect 10045 19805 10057 19839
rect 10091 19805 10103 19839
rect 10045 19799 10103 19805
rect 7282 19728 7288 19780
rect 7340 19768 7346 19780
rect 10060 19768 10088 19799
rect 11054 19796 11060 19848
rect 11112 19796 11118 19848
rect 11330 19796 11336 19848
rect 11388 19796 11394 19848
rect 11974 19796 11980 19848
rect 12032 19796 12038 19848
rect 14274 19836 14280 19848
rect 13386 19808 14280 19836
rect 14274 19796 14280 19808
rect 14332 19796 14338 19848
rect 14642 19796 14648 19848
rect 14700 19836 14706 19848
rect 14921 19839 14979 19845
rect 14921 19836 14933 19839
rect 14700 19808 14933 19836
rect 14700 19796 14706 19808
rect 14921 19805 14933 19808
rect 14967 19805 14979 19839
rect 14921 19799 14979 19805
rect 15565 19839 15623 19845
rect 15565 19805 15577 19839
rect 15611 19805 15623 19839
rect 15565 19799 15623 19805
rect 16485 19839 16543 19845
rect 16485 19805 16497 19839
rect 16531 19836 16543 19839
rect 17604 19836 17632 19944
rect 18616 19913 18644 20012
rect 23290 20000 23296 20012
rect 23348 20000 23354 20052
rect 24118 20000 24124 20052
rect 24176 20040 24182 20052
rect 30006 20040 30012 20052
rect 24176 20012 30012 20040
rect 24176 20000 24182 20012
rect 21818 19932 21824 19984
rect 21876 19972 21882 19984
rect 22281 19975 22339 19981
rect 22281 19972 22293 19975
rect 21876 19944 22293 19972
rect 21876 19932 21882 19944
rect 22281 19941 22293 19944
rect 22327 19941 22339 19975
rect 22281 19935 22339 19941
rect 22830 19932 22836 19984
rect 22888 19972 22894 19984
rect 24765 19975 24823 19981
rect 24765 19972 24777 19975
rect 22888 19944 24777 19972
rect 22888 19932 22894 19944
rect 24765 19941 24777 19944
rect 24811 19941 24823 19975
rect 24765 19935 24823 19941
rect 18601 19907 18659 19913
rect 18601 19873 18613 19907
rect 18647 19873 18659 19907
rect 18601 19867 18659 19873
rect 18785 19907 18843 19913
rect 18785 19873 18797 19907
rect 18831 19904 18843 19907
rect 18874 19904 18880 19916
rect 18831 19876 18880 19904
rect 18831 19873 18843 19876
rect 18785 19867 18843 19873
rect 18874 19864 18880 19876
rect 18932 19864 18938 19916
rect 20809 19907 20867 19913
rect 20809 19873 20821 19907
rect 20855 19904 20867 19907
rect 23385 19907 23443 19913
rect 20855 19876 22094 19904
rect 20855 19873 20867 19876
rect 20809 19867 20867 19873
rect 19889 19839 19947 19845
rect 19889 19836 19901 19839
rect 16531 19808 17448 19836
rect 17604 19808 19901 19836
rect 16531 19805 16543 19808
rect 16485 19799 16543 19805
rect 12158 19768 12164 19780
rect 7340 19740 9904 19768
rect 10060 19740 12164 19768
rect 7340 19728 7346 19740
rect 9876 19709 9904 19740
rect 12158 19728 12164 19740
rect 12216 19728 12222 19780
rect 12250 19728 12256 19780
rect 12308 19728 12314 19780
rect 14734 19768 14740 19780
rect 13648 19740 14740 19768
rect 7745 19703 7803 19709
rect 7745 19700 7757 19703
rect 6012 19672 7757 19700
rect 7745 19669 7757 19672
rect 7791 19669 7803 19703
rect 7745 19663 7803 19669
rect 9861 19703 9919 19709
rect 9861 19669 9873 19703
rect 9907 19669 9919 19703
rect 9861 19663 9919 19669
rect 12066 19660 12072 19712
rect 12124 19700 12130 19712
rect 12618 19700 12624 19712
rect 12124 19672 12624 19700
rect 12124 19660 12130 19672
rect 12618 19660 12624 19672
rect 12676 19660 12682 19712
rect 13262 19660 13268 19712
rect 13320 19700 13326 19712
rect 13648 19700 13676 19740
rect 14734 19728 14740 19740
rect 14792 19728 14798 19780
rect 13320 19672 13676 19700
rect 13725 19703 13783 19709
rect 13320 19660 13326 19672
rect 13725 19669 13737 19703
rect 13771 19700 13783 19703
rect 13814 19700 13820 19712
rect 13771 19672 13820 19700
rect 13771 19669 13783 19672
rect 13725 19663 13783 19669
rect 13814 19660 13820 19672
rect 13872 19660 13878 19712
rect 15580 19700 15608 19799
rect 16666 19728 16672 19780
rect 16724 19728 16730 19780
rect 16942 19728 16948 19780
rect 17000 19768 17006 19780
rect 17313 19771 17371 19777
rect 17313 19768 17325 19771
rect 17000 19740 17325 19768
rect 17000 19728 17006 19740
rect 17313 19737 17325 19740
rect 17359 19737 17371 19771
rect 17313 19731 17371 19737
rect 17420 19712 17448 19808
rect 19889 19805 19901 19808
rect 19935 19805 19947 19839
rect 19889 19799 19947 19805
rect 20530 19796 20536 19848
rect 20588 19796 20594 19848
rect 22066 19836 22094 19876
rect 23385 19873 23397 19907
rect 23431 19904 23443 19907
rect 25130 19904 25136 19916
rect 23431 19876 25136 19904
rect 23431 19873 23443 19876
rect 23385 19867 23443 19873
rect 25130 19864 25136 19876
rect 25188 19864 25194 19916
rect 25590 19864 25596 19916
rect 25648 19904 25654 19916
rect 26988 19913 27016 20012
rect 30006 20000 30012 20012
rect 30064 20000 30070 20052
rect 30377 20043 30435 20049
rect 30377 20009 30389 20043
rect 30423 20040 30435 20043
rect 31386 20040 31392 20052
rect 30423 20012 31392 20040
rect 30423 20009 30435 20012
rect 30377 20003 30435 20009
rect 31386 20000 31392 20012
rect 31444 20000 31450 20052
rect 33413 20043 33471 20049
rect 33413 20009 33425 20043
rect 33459 20040 33471 20043
rect 34698 20040 34704 20052
rect 33459 20012 34704 20040
rect 33459 20009 33471 20012
rect 33413 20003 33471 20009
rect 34698 20000 34704 20012
rect 34756 20000 34762 20052
rect 34885 20043 34943 20049
rect 34885 20009 34897 20043
rect 34931 20040 34943 20043
rect 36722 20040 36728 20052
rect 34931 20012 36728 20040
rect 34931 20009 34943 20012
rect 34885 20003 34943 20009
rect 36722 20000 36728 20012
rect 36780 20000 36786 20052
rect 37826 20000 37832 20052
rect 37884 20040 37890 20052
rect 40037 20043 40095 20049
rect 40037 20040 40049 20043
rect 37884 20012 40049 20040
rect 37884 20000 37890 20012
rect 40037 20009 40049 20012
rect 40083 20009 40095 20043
rect 40037 20003 40095 20009
rect 40126 20000 40132 20052
rect 40184 20040 40190 20052
rect 40184 20012 41828 20040
rect 40184 20000 40190 20012
rect 27154 19932 27160 19984
rect 27212 19972 27218 19984
rect 28077 19975 28135 19981
rect 28077 19972 28089 19975
rect 27212 19944 28089 19972
rect 27212 19932 27218 19944
rect 28077 19941 28089 19944
rect 28123 19941 28135 19975
rect 28077 19935 28135 19941
rect 28994 19932 29000 19984
rect 29052 19972 29058 19984
rect 31573 19975 31631 19981
rect 31573 19972 31585 19975
rect 29052 19944 31585 19972
rect 29052 19932 29058 19944
rect 31573 19941 31585 19944
rect 31619 19941 31631 19975
rect 31573 19935 31631 19941
rect 33502 19932 33508 19984
rect 33560 19972 33566 19984
rect 33560 19944 40540 19972
rect 33560 19932 33566 19944
rect 26145 19907 26203 19913
rect 26145 19904 26157 19907
rect 25648 19876 26157 19904
rect 25648 19864 25654 19876
rect 26145 19873 26157 19876
rect 26191 19873 26203 19907
rect 26145 19867 26203 19873
rect 26973 19907 27031 19913
rect 26973 19873 26985 19907
rect 27019 19873 27031 19907
rect 26973 19867 27031 19873
rect 27522 19864 27528 19916
rect 27580 19904 27586 19916
rect 27890 19904 27896 19916
rect 27580 19876 27896 19904
rect 27580 19864 27586 19876
rect 27890 19864 27896 19876
rect 27948 19864 27954 19916
rect 28534 19864 28540 19916
rect 28592 19864 28598 19916
rect 28626 19864 28632 19916
rect 28684 19864 28690 19916
rect 29546 19904 29552 19916
rect 28736 19876 29552 19904
rect 23842 19836 23848 19848
rect 22066 19808 23848 19836
rect 23842 19796 23848 19808
rect 23900 19796 23906 19848
rect 26053 19839 26111 19845
rect 26053 19805 26065 19839
rect 26099 19836 26111 19839
rect 28736 19836 28764 19876
rect 29546 19864 29552 19876
rect 29604 19864 29610 19916
rect 31021 19907 31079 19913
rect 31021 19873 31033 19907
rect 31067 19904 31079 19907
rect 31754 19904 31760 19916
rect 31067 19876 31760 19904
rect 31067 19873 31079 19876
rect 31021 19867 31079 19873
rect 31754 19864 31760 19876
rect 31812 19864 31818 19916
rect 32122 19864 32128 19916
rect 32180 19864 32186 19916
rect 33410 19864 33416 19916
rect 33468 19904 33474 19916
rect 33965 19907 34023 19913
rect 33965 19904 33977 19907
rect 33468 19876 33977 19904
rect 33468 19864 33474 19876
rect 33965 19873 33977 19876
rect 34011 19873 34023 19907
rect 33965 19867 34023 19873
rect 35250 19864 35256 19916
rect 35308 19904 35314 19916
rect 35345 19907 35403 19913
rect 35345 19904 35357 19907
rect 35308 19876 35357 19904
rect 35308 19864 35314 19876
rect 35345 19873 35357 19876
rect 35391 19873 35403 19907
rect 35345 19867 35403 19873
rect 35434 19864 35440 19916
rect 35492 19864 35498 19916
rect 36725 19907 36783 19913
rect 36725 19873 36737 19907
rect 36771 19904 36783 19907
rect 37274 19904 37280 19916
rect 36771 19876 37280 19904
rect 36771 19873 36783 19876
rect 36725 19867 36783 19873
rect 37274 19864 37280 19876
rect 37332 19864 37338 19916
rect 37918 19864 37924 19916
rect 37976 19904 37982 19916
rect 38289 19907 38347 19913
rect 38289 19904 38301 19907
rect 37976 19876 38301 19904
rect 37976 19864 37982 19876
rect 38289 19873 38301 19876
rect 38335 19904 38347 19907
rect 38378 19904 38384 19916
rect 38335 19876 38384 19904
rect 38335 19873 38347 19876
rect 38289 19867 38347 19873
rect 38378 19864 38384 19876
rect 38436 19864 38442 19916
rect 38473 19907 38531 19913
rect 38473 19873 38485 19907
rect 38519 19904 38531 19907
rect 38562 19904 38568 19916
rect 38519 19876 38568 19904
rect 38519 19873 38531 19876
rect 38473 19867 38531 19873
rect 38562 19864 38568 19876
rect 38620 19864 38626 19916
rect 40512 19913 40540 19944
rect 40497 19907 40555 19913
rect 40497 19873 40509 19907
rect 40543 19873 40555 19907
rect 40497 19867 40555 19873
rect 40586 19864 40592 19916
rect 40644 19864 40650 19916
rect 41598 19864 41604 19916
rect 41656 19904 41662 19916
rect 41800 19913 41828 20012
rect 41693 19907 41751 19913
rect 41693 19904 41705 19907
rect 41656 19876 41705 19904
rect 41656 19864 41662 19876
rect 41693 19873 41705 19876
rect 41739 19873 41751 19907
rect 41693 19867 41751 19873
rect 41785 19907 41843 19913
rect 41785 19873 41797 19907
rect 41831 19873 41843 19907
rect 41785 19867 41843 19873
rect 41874 19864 41880 19916
rect 41932 19904 41938 19916
rect 49329 19907 49387 19913
rect 49329 19904 49341 19907
rect 41932 19876 49341 19904
rect 41932 19864 41938 19876
rect 49329 19873 49341 19876
rect 49375 19873 49387 19907
rect 49329 19867 49387 19873
rect 26099 19808 28764 19836
rect 26099 19805 26111 19808
rect 26053 19799 26111 19805
rect 28810 19796 28816 19848
rect 28868 19836 28874 19848
rect 29917 19839 29975 19845
rect 29917 19836 29929 19839
rect 28868 19808 29929 19836
rect 28868 19796 28874 19808
rect 29917 19805 29929 19808
rect 29963 19805 29975 19839
rect 29917 19799 29975 19805
rect 30282 19796 30288 19848
rect 30340 19836 30346 19848
rect 31941 19839 31999 19845
rect 30340 19808 31754 19836
rect 30340 19796 30346 19808
rect 19705 19771 19763 19777
rect 19705 19737 19717 19771
rect 19751 19768 19763 19771
rect 19751 19740 21220 19768
rect 19751 19737 19763 19740
rect 19705 19731 19763 19737
rect 17218 19700 17224 19712
rect 15580 19672 17224 19700
rect 17218 19660 17224 19672
rect 17276 19660 17282 19712
rect 17402 19660 17408 19712
rect 17460 19660 17466 19712
rect 18141 19703 18199 19709
rect 18141 19669 18153 19703
rect 18187 19700 18199 19703
rect 18322 19700 18328 19712
rect 18187 19672 18328 19700
rect 18187 19669 18199 19672
rect 18141 19663 18199 19669
rect 18322 19660 18328 19672
rect 18380 19660 18386 19712
rect 18506 19660 18512 19712
rect 18564 19660 18570 19712
rect 21192 19700 21220 19740
rect 21266 19728 21272 19780
rect 21324 19728 21330 19780
rect 25961 19771 26019 19777
rect 25961 19737 25973 19771
rect 26007 19768 26019 19771
rect 26007 19740 26464 19768
rect 26007 19737 26019 19740
rect 25961 19731 26019 19737
rect 21450 19700 21456 19712
rect 21192 19672 21456 19700
rect 21450 19660 21456 19672
rect 21508 19660 21514 19712
rect 22738 19660 22744 19712
rect 22796 19660 22802 19712
rect 22830 19660 22836 19712
rect 22888 19700 22894 19712
rect 26436 19709 26464 19740
rect 26786 19728 26792 19780
rect 26844 19728 26850 19780
rect 27614 19728 27620 19780
rect 27672 19728 27678 19780
rect 28445 19771 28503 19777
rect 28445 19737 28457 19771
rect 28491 19768 28503 19771
rect 30926 19768 30932 19780
rect 28491 19740 30932 19768
rect 28491 19737 28503 19740
rect 28445 19731 28503 19737
rect 30926 19728 30932 19740
rect 30984 19728 30990 19780
rect 31726 19768 31754 19808
rect 31941 19805 31953 19839
rect 31987 19836 31999 19839
rect 32030 19836 32036 19848
rect 31987 19808 32036 19836
rect 31987 19805 31999 19808
rect 31941 19799 31999 19805
rect 32030 19796 32036 19808
rect 32088 19836 32094 19848
rect 33781 19839 33839 19845
rect 33781 19836 33793 19839
rect 32088 19808 33793 19836
rect 32088 19796 32094 19808
rect 33781 19805 33793 19808
rect 33827 19805 33839 19839
rect 33781 19799 33839 19805
rect 33873 19839 33931 19845
rect 33873 19805 33885 19839
rect 33919 19836 33931 19839
rect 34054 19836 34060 19848
rect 33919 19808 34060 19836
rect 33919 19805 33931 19808
rect 33873 19799 33931 19805
rect 34054 19796 34060 19808
rect 34112 19796 34118 19848
rect 37366 19796 37372 19848
rect 37424 19836 37430 19848
rect 38197 19839 38255 19845
rect 38197 19836 38209 19839
rect 37424 19808 38209 19836
rect 37424 19796 37430 19808
rect 38197 19805 38209 19808
rect 38243 19836 38255 19839
rect 39114 19836 39120 19848
rect 38243 19808 39120 19836
rect 38243 19805 38255 19808
rect 38197 19799 38255 19805
rect 39114 19796 39120 19808
rect 39172 19796 39178 19848
rect 39209 19839 39267 19845
rect 39209 19805 39221 19839
rect 39255 19836 39267 19839
rect 39255 19808 40356 19836
rect 39255 19805 39267 19808
rect 39209 19799 39267 19805
rect 31726 19740 35020 19768
rect 23109 19703 23167 19709
rect 23109 19700 23121 19703
rect 22888 19672 23121 19700
rect 22888 19660 22894 19672
rect 23109 19669 23121 19672
rect 23155 19669 23167 19703
rect 23109 19663 23167 19669
rect 23201 19703 23259 19709
rect 23201 19669 23213 19703
rect 23247 19700 23259 19703
rect 25593 19703 25651 19709
rect 25593 19700 25605 19703
rect 23247 19672 25605 19700
rect 23247 19669 23259 19672
rect 23201 19663 23259 19669
rect 25593 19669 25605 19672
rect 25639 19669 25651 19703
rect 25593 19663 25651 19669
rect 26421 19703 26479 19709
rect 26421 19669 26433 19703
rect 26467 19669 26479 19703
rect 26421 19663 26479 19669
rect 26881 19703 26939 19709
rect 26881 19669 26893 19703
rect 26927 19700 26939 19703
rect 26970 19700 26976 19712
rect 26927 19672 26976 19700
rect 26927 19669 26939 19672
rect 26881 19663 26939 19669
rect 26970 19660 26976 19672
rect 27028 19660 27034 19712
rect 27246 19660 27252 19712
rect 27304 19660 27310 19712
rect 27709 19703 27767 19709
rect 27709 19669 27721 19703
rect 27755 19700 27767 19703
rect 28902 19700 28908 19712
rect 27755 19672 28908 19700
rect 27755 19669 27767 19672
rect 27709 19663 27767 19669
rect 28902 19660 28908 19672
rect 28960 19660 28966 19712
rect 30650 19660 30656 19712
rect 30708 19700 30714 19712
rect 30745 19703 30803 19709
rect 30745 19700 30757 19703
rect 30708 19672 30757 19700
rect 30708 19660 30714 19672
rect 30745 19669 30757 19672
rect 30791 19669 30803 19703
rect 30745 19663 30803 19669
rect 30834 19660 30840 19712
rect 30892 19660 30898 19712
rect 32033 19703 32091 19709
rect 32033 19669 32045 19703
rect 32079 19700 32091 19703
rect 34054 19700 34060 19712
rect 32079 19672 34060 19700
rect 32079 19669 32091 19672
rect 32033 19663 32091 19669
rect 34054 19660 34060 19672
rect 34112 19660 34118 19712
rect 34992 19700 35020 19740
rect 35066 19728 35072 19780
rect 35124 19768 35130 19780
rect 35253 19771 35311 19777
rect 35253 19768 35265 19771
rect 35124 19740 35265 19768
rect 35124 19728 35130 19740
rect 35253 19737 35265 19740
rect 35299 19737 35311 19771
rect 35253 19731 35311 19737
rect 36449 19771 36507 19777
rect 36449 19737 36461 19771
rect 36495 19768 36507 19771
rect 39942 19768 39948 19780
rect 36495 19740 39948 19768
rect 36495 19737 36507 19740
rect 36449 19731 36507 19737
rect 39942 19728 39948 19740
rect 40000 19728 40006 19780
rect 40328 19768 40356 19808
rect 40405 19771 40463 19777
rect 40405 19768 40417 19771
rect 40328 19740 40417 19768
rect 40405 19737 40417 19740
rect 40451 19737 40463 19771
rect 40405 19731 40463 19737
rect 41601 19771 41659 19777
rect 41601 19737 41613 19771
rect 41647 19768 41659 19771
rect 48406 19768 48412 19780
rect 41647 19740 48412 19768
rect 41647 19737 41659 19740
rect 41601 19731 41659 19737
rect 48406 19728 48412 19740
rect 48464 19728 48470 19780
rect 49145 19771 49203 19777
rect 49145 19737 49157 19771
rect 49191 19768 49203 19771
rect 49326 19768 49332 19780
rect 49191 19740 49332 19768
rect 49191 19737 49203 19740
rect 49145 19731 49203 19737
rect 49326 19728 49332 19740
rect 49384 19728 49390 19780
rect 35894 19700 35900 19712
rect 34992 19672 35900 19700
rect 35894 19660 35900 19672
rect 35952 19660 35958 19712
rect 35986 19660 35992 19712
rect 36044 19700 36050 19712
rect 36081 19703 36139 19709
rect 36081 19700 36093 19703
rect 36044 19672 36093 19700
rect 36044 19660 36050 19672
rect 36081 19669 36093 19672
rect 36127 19669 36139 19703
rect 36081 19663 36139 19669
rect 36538 19660 36544 19712
rect 36596 19660 36602 19712
rect 37829 19703 37887 19709
rect 37829 19669 37841 19703
rect 37875 19700 37887 19703
rect 40954 19700 40960 19712
rect 37875 19672 40960 19700
rect 37875 19669 37887 19672
rect 37829 19663 37887 19669
rect 40954 19660 40960 19672
rect 41012 19660 41018 19712
rect 41138 19660 41144 19712
rect 41196 19700 41202 19712
rect 41233 19703 41291 19709
rect 41233 19700 41245 19703
rect 41196 19672 41245 19700
rect 41196 19660 41202 19672
rect 41233 19669 41245 19672
rect 41279 19669 41291 19703
rect 41233 19663 41291 19669
rect 1104 19610 49864 19632
rect 1104 19558 7950 19610
rect 8002 19558 8014 19610
rect 8066 19558 8078 19610
rect 8130 19558 8142 19610
rect 8194 19558 8206 19610
rect 8258 19558 17950 19610
rect 18002 19558 18014 19610
rect 18066 19558 18078 19610
rect 18130 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 27950 19610
rect 28002 19558 28014 19610
rect 28066 19558 28078 19610
rect 28130 19558 28142 19610
rect 28194 19558 28206 19610
rect 28258 19558 37950 19610
rect 38002 19558 38014 19610
rect 38066 19558 38078 19610
rect 38130 19558 38142 19610
rect 38194 19558 38206 19610
rect 38258 19558 47950 19610
rect 48002 19558 48014 19610
rect 48066 19558 48078 19610
rect 48130 19558 48142 19610
rect 48194 19558 48206 19610
rect 48258 19558 49864 19610
rect 1104 19536 49864 19558
rect 9306 19496 9312 19508
rect 1780 19468 9312 19496
rect 1780 19369 1808 19468
rect 9306 19456 9312 19468
rect 9364 19456 9370 19508
rect 10965 19499 11023 19505
rect 10965 19465 10977 19499
rect 11011 19465 11023 19499
rect 10965 19459 11023 19465
rect 4338 19388 4344 19440
rect 4396 19388 4402 19440
rect 10870 19428 10876 19440
rect 5276 19400 10876 19428
rect 1765 19363 1823 19369
rect 1765 19329 1777 19363
rect 1811 19329 1823 19363
rect 1765 19323 1823 19329
rect 2777 19363 2835 19369
rect 2777 19329 2789 19363
rect 2823 19360 2835 19363
rect 2866 19360 2872 19372
rect 2823 19332 2872 19360
rect 2823 19329 2835 19332
rect 2777 19323 2835 19329
rect 2866 19320 2872 19332
rect 2924 19320 2930 19372
rect 3605 19363 3663 19369
rect 3605 19329 3617 19363
rect 3651 19360 3663 19363
rect 5276 19360 5304 19400
rect 10870 19388 10876 19400
rect 10928 19388 10934 19440
rect 3651 19332 5304 19360
rect 3651 19329 3663 19332
rect 3605 19323 3663 19329
rect 5350 19320 5356 19372
rect 5408 19320 5414 19372
rect 7558 19320 7564 19372
rect 7616 19360 7622 19372
rect 10980 19360 11008 19459
rect 11054 19456 11060 19508
rect 11112 19496 11118 19508
rect 12618 19496 12624 19508
rect 11112 19468 12624 19496
rect 11112 19456 11118 19468
rect 12618 19456 12624 19468
rect 12676 19456 12682 19508
rect 13354 19456 13360 19508
rect 13412 19496 13418 19508
rect 14461 19499 14519 19505
rect 14461 19496 14473 19499
rect 13412 19468 14473 19496
rect 13412 19456 13418 19468
rect 14461 19465 14473 19468
rect 14507 19465 14519 19499
rect 14461 19459 14519 19465
rect 15286 19456 15292 19508
rect 15344 19496 15350 19508
rect 15381 19499 15439 19505
rect 15381 19496 15393 19499
rect 15344 19468 15393 19496
rect 15344 19456 15350 19468
rect 15381 19465 15393 19468
rect 15427 19465 15439 19499
rect 15381 19459 15439 19465
rect 16850 19456 16856 19508
rect 16908 19456 16914 19508
rect 17313 19499 17371 19505
rect 17313 19465 17325 19499
rect 17359 19496 17371 19499
rect 19242 19496 19248 19508
rect 17359 19468 19248 19496
rect 17359 19465 17371 19468
rect 17313 19459 17371 19465
rect 19242 19456 19248 19468
rect 19300 19456 19306 19508
rect 20717 19499 20775 19505
rect 20717 19465 20729 19499
rect 20763 19496 20775 19499
rect 20806 19496 20812 19508
rect 20763 19468 20812 19496
rect 20763 19465 20775 19468
rect 20717 19459 20775 19465
rect 20806 19456 20812 19468
rect 20864 19456 20870 19508
rect 21177 19499 21235 19505
rect 21177 19465 21189 19499
rect 21223 19496 21235 19499
rect 23934 19496 23940 19508
rect 21223 19468 23940 19496
rect 21223 19465 21235 19468
rect 21177 19459 21235 19465
rect 23934 19456 23940 19468
rect 23992 19456 23998 19508
rect 25130 19456 25136 19508
rect 25188 19456 25194 19508
rect 26602 19496 26608 19508
rect 25976 19468 26608 19496
rect 13262 19428 13268 19440
rect 11164 19400 13268 19428
rect 11164 19369 11192 19400
rect 13262 19388 13268 19400
rect 13320 19388 13326 19440
rect 14274 19428 14280 19440
rect 14214 19400 14280 19428
rect 14274 19388 14280 19400
rect 14332 19428 14338 19440
rect 15746 19428 15752 19440
rect 14332 19400 15752 19428
rect 14332 19388 14338 19400
rect 15746 19388 15752 19400
rect 15804 19388 15810 19440
rect 17034 19388 17040 19440
rect 17092 19428 17098 19440
rect 18598 19428 18604 19440
rect 17092 19400 18604 19428
rect 17092 19388 17098 19400
rect 7616 19332 11008 19360
rect 11149 19363 11207 19369
rect 7616 19320 7622 19332
rect 11149 19329 11161 19363
rect 11195 19329 11207 19363
rect 11149 19323 11207 19329
rect 12066 19320 12072 19372
rect 12124 19320 12130 19372
rect 12702 19363 12760 19369
rect 12702 19329 12714 19363
rect 12748 19329 12760 19363
rect 12702 19323 12760 19329
rect 15565 19363 15623 19369
rect 15565 19329 15577 19363
rect 15611 19360 15623 19363
rect 15838 19360 15844 19372
rect 15611 19332 15844 19360
rect 15611 19329 15623 19332
rect 15565 19323 15623 19329
rect 12717 19306 12756 19323
rect 15838 19320 15844 19332
rect 15896 19320 15902 19372
rect 16117 19363 16175 19369
rect 16117 19329 16129 19363
rect 16163 19360 16175 19363
rect 16482 19360 16488 19372
rect 16163 19332 16488 19360
rect 16163 19329 16175 19332
rect 16117 19323 16175 19329
rect 16482 19320 16488 19332
rect 16540 19320 16546 19372
rect 17218 19320 17224 19372
rect 17276 19320 17282 19372
rect 18064 19369 18092 19400
rect 18598 19388 18604 19400
rect 18656 19388 18662 19440
rect 19610 19388 19616 19440
rect 19668 19428 19674 19440
rect 25976 19428 26004 19468
rect 26602 19456 26608 19468
rect 26660 19456 26666 19508
rect 27522 19456 27528 19508
rect 27580 19496 27586 19508
rect 27982 19496 27988 19508
rect 27580 19468 27988 19496
rect 27580 19456 27586 19468
rect 27982 19456 27988 19468
rect 28040 19456 28046 19508
rect 28445 19499 28503 19505
rect 28445 19465 28457 19499
rect 28491 19496 28503 19499
rect 28718 19496 28724 19508
rect 28491 19468 28724 19496
rect 28491 19465 28503 19468
rect 28445 19459 28503 19465
rect 28718 19456 28724 19468
rect 28776 19456 28782 19508
rect 28810 19456 28816 19508
rect 28868 19456 28874 19508
rect 29638 19456 29644 19508
rect 29696 19456 29702 19508
rect 30101 19499 30159 19505
rect 30101 19465 30113 19499
rect 30147 19496 30159 19499
rect 31754 19496 31760 19508
rect 30147 19468 31760 19496
rect 30147 19465 30159 19468
rect 30101 19459 30159 19465
rect 31754 19456 31760 19468
rect 31812 19456 31818 19508
rect 32309 19499 32367 19505
rect 32309 19465 32321 19499
rect 32355 19496 32367 19499
rect 32582 19496 32588 19508
rect 32355 19468 32588 19496
rect 32355 19465 32367 19468
rect 32309 19459 32367 19465
rect 32582 19456 32588 19468
rect 32640 19456 32646 19508
rect 32674 19456 32680 19508
rect 32732 19456 32738 19508
rect 32769 19499 32827 19505
rect 32769 19465 32781 19499
rect 32815 19496 32827 19499
rect 32858 19496 32864 19508
rect 32815 19468 32864 19496
rect 32815 19465 32827 19468
rect 32769 19459 32827 19465
rect 32858 19456 32864 19468
rect 32916 19456 32922 19508
rect 33502 19456 33508 19508
rect 33560 19456 33566 19508
rect 33873 19499 33931 19505
rect 33873 19465 33885 19499
rect 33919 19496 33931 19499
rect 34330 19496 34336 19508
rect 33919 19468 34336 19496
rect 33919 19465 33931 19468
rect 33873 19459 33931 19465
rect 34330 19456 34336 19468
rect 34388 19456 34394 19508
rect 34701 19499 34759 19505
rect 34701 19465 34713 19499
rect 34747 19496 34759 19499
rect 36538 19496 36544 19508
rect 34747 19468 36544 19496
rect 34747 19465 34759 19468
rect 34701 19459 34759 19465
rect 36538 19456 36544 19468
rect 36596 19456 36602 19508
rect 40402 19456 40408 19508
rect 40460 19496 40466 19508
rect 40497 19499 40555 19505
rect 40497 19496 40509 19499
rect 40460 19468 40509 19496
rect 40460 19456 40466 19468
rect 40497 19465 40509 19468
rect 40543 19465 40555 19499
rect 40497 19459 40555 19465
rect 40589 19499 40647 19505
rect 40589 19465 40601 19499
rect 40635 19496 40647 19499
rect 41046 19496 41052 19508
rect 40635 19468 41052 19496
rect 40635 19465 40647 19468
rect 40589 19459 40647 19465
rect 41046 19456 41052 19468
rect 41104 19456 41110 19508
rect 19668 19400 22876 19428
rect 24886 19400 26004 19428
rect 19668 19388 19674 19400
rect 18049 19363 18107 19369
rect 18049 19329 18061 19363
rect 18095 19329 18107 19363
rect 18049 19323 18107 19329
rect 19426 19320 19432 19372
rect 19484 19360 19490 19372
rect 19886 19360 19892 19372
rect 19484 19332 19892 19360
rect 19484 19320 19490 19332
rect 19886 19320 19892 19332
rect 19944 19320 19950 19372
rect 20073 19363 20131 19369
rect 20073 19329 20085 19363
rect 20119 19360 20131 19363
rect 20346 19360 20352 19372
rect 20119 19332 20352 19360
rect 20119 19329 20131 19332
rect 20073 19323 20131 19329
rect 20346 19320 20352 19332
rect 20404 19320 20410 19372
rect 21085 19363 21143 19369
rect 21085 19329 21097 19363
rect 21131 19360 21143 19363
rect 21542 19360 21548 19372
rect 21131 19332 21548 19360
rect 21131 19329 21143 19332
rect 21085 19323 21143 19329
rect 21542 19320 21548 19332
rect 21600 19320 21606 19372
rect 22848 19369 22876 19400
rect 26142 19388 26148 19440
rect 26200 19388 26206 19440
rect 26234 19388 26240 19440
rect 26292 19428 26298 19440
rect 27154 19428 27160 19440
rect 26292 19400 27160 19428
rect 26292 19388 26298 19400
rect 27154 19388 27160 19400
rect 27212 19388 27218 19440
rect 27706 19388 27712 19440
rect 27764 19428 27770 19440
rect 27893 19431 27951 19437
rect 27893 19428 27905 19431
rect 27764 19400 27905 19428
rect 27764 19388 27770 19400
rect 27893 19397 27905 19400
rect 27939 19428 27951 19431
rect 28905 19431 28963 19437
rect 28905 19428 28917 19431
rect 27939 19400 28917 19428
rect 27939 19397 27951 19400
rect 27893 19391 27951 19397
rect 28905 19397 28917 19400
rect 28951 19397 28963 19431
rect 28905 19391 28963 19397
rect 29914 19388 29920 19440
rect 29972 19428 29978 19440
rect 30190 19428 30196 19440
rect 29972 19400 30196 19428
rect 29972 19388 29978 19400
rect 30190 19388 30196 19400
rect 30248 19388 30254 19440
rect 30650 19388 30656 19440
rect 30708 19428 30714 19440
rect 31294 19428 31300 19440
rect 30708 19400 31300 19428
rect 30708 19388 30714 19400
rect 31294 19388 31300 19400
rect 31352 19388 31358 19440
rect 31570 19388 31576 19440
rect 31628 19428 31634 19440
rect 35250 19428 35256 19440
rect 31628 19400 35256 19428
rect 31628 19388 31634 19400
rect 35250 19388 35256 19400
rect 35308 19388 35314 19440
rect 36170 19428 36176 19440
rect 35820 19400 36176 19428
rect 22005 19363 22063 19369
rect 22005 19329 22017 19363
rect 22051 19360 22063 19363
rect 22833 19363 22891 19369
rect 22051 19332 22784 19360
rect 22051 19329 22063 19332
rect 22005 19323 22063 19329
rect 9122 19252 9128 19304
rect 9180 19292 9186 19304
rect 12717 19292 12745 19306
rect 9180 19264 12745 19292
rect 9180 19252 9186 19264
rect 12717 19236 12745 19264
rect 12989 19295 13047 19301
rect 12989 19261 13001 19295
rect 13035 19292 13047 19295
rect 15930 19292 15936 19304
rect 13035 19264 15936 19292
rect 13035 19261 13047 19264
rect 12989 19255 13047 19261
rect 15930 19252 15936 19264
rect 15988 19252 15994 19304
rect 17497 19295 17555 19301
rect 17497 19261 17509 19295
rect 17543 19261 17555 19295
rect 17497 19255 17555 19261
rect 18325 19295 18383 19301
rect 18325 19261 18337 19295
rect 18371 19292 18383 19295
rect 21269 19295 21327 19301
rect 18371 19264 20024 19292
rect 18371 19261 18383 19264
rect 18325 19255 18383 19261
rect 11606 19184 11612 19236
rect 11664 19224 11670 19236
rect 11974 19224 11980 19236
rect 11664 19196 11980 19224
rect 11664 19184 11670 19196
rect 11974 19184 11980 19196
rect 12032 19224 12038 19236
rect 12032 19196 12434 19224
rect 12032 19184 12038 19196
rect 2314 19116 2320 19168
rect 2372 19156 2378 19168
rect 5445 19159 5503 19165
rect 5445 19156 5457 19159
rect 2372 19128 5457 19156
rect 2372 19116 2378 19128
rect 5445 19125 5457 19128
rect 5491 19125 5503 19159
rect 5445 19119 5503 19125
rect 9861 19159 9919 19165
rect 9861 19125 9873 19159
rect 9907 19156 9919 19159
rect 10410 19156 10416 19168
rect 9907 19128 10416 19156
rect 9907 19125 9919 19128
rect 9861 19119 9919 19125
rect 10410 19116 10416 19128
rect 10468 19116 10474 19168
rect 10505 19159 10563 19165
rect 10505 19125 10517 19159
rect 10551 19156 10563 19159
rect 11330 19156 11336 19168
rect 10551 19128 11336 19156
rect 10551 19125 10563 19128
rect 10505 19119 10563 19125
rect 11330 19116 11336 19128
rect 11388 19116 11394 19168
rect 11514 19116 11520 19168
rect 11572 19156 11578 19168
rect 12161 19159 12219 19165
rect 12161 19156 12173 19159
rect 11572 19128 12173 19156
rect 11572 19116 11578 19128
rect 12161 19125 12173 19128
rect 12207 19125 12219 19159
rect 12406 19156 12434 19196
rect 12710 19184 12716 19236
rect 12768 19184 12774 19236
rect 13998 19156 14004 19168
rect 12406 19128 14004 19156
rect 12161 19119 12219 19125
rect 13998 19116 14004 19128
rect 14056 19116 14062 19168
rect 16206 19116 16212 19168
rect 16264 19116 16270 19168
rect 17512 19156 17540 19255
rect 19996 19224 20024 19264
rect 21269 19261 21281 19295
rect 21315 19261 21327 19295
rect 22756 19292 22784 19332
rect 22833 19329 22845 19363
rect 22879 19360 22891 19363
rect 23382 19360 23388 19372
rect 22879 19332 23388 19360
rect 22879 19329 22891 19332
rect 22833 19323 22891 19329
rect 23382 19320 23388 19332
rect 23440 19320 23446 19372
rect 25866 19320 25872 19372
rect 25924 19360 25930 19372
rect 28626 19360 28632 19372
rect 25924 19332 28632 19360
rect 25924 19320 25930 19332
rect 23290 19292 23296 19304
rect 22756 19264 23296 19292
rect 21269 19255 21327 19261
rect 21284 19224 21312 19255
rect 23290 19252 23296 19264
rect 23348 19252 23354 19304
rect 23658 19252 23664 19304
rect 23716 19252 23722 19304
rect 26436 19301 26464 19332
rect 28626 19320 28632 19332
rect 28684 19320 28690 19372
rect 28828 19332 29040 19360
rect 26237 19295 26295 19301
rect 26237 19261 26249 19295
rect 26283 19261 26295 19295
rect 26237 19255 26295 19261
rect 26421 19295 26479 19301
rect 26421 19261 26433 19295
rect 26467 19261 26479 19295
rect 26421 19255 26479 19261
rect 22462 19224 22468 19236
rect 19996 19196 22468 19224
rect 22462 19184 22468 19196
rect 22520 19184 22526 19236
rect 26252 19224 26280 19255
rect 27798 19252 27804 19304
rect 27856 19292 27862 19304
rect 28828 19292 28856 19332
rect 29012 19301 29040 19332
rect 30006 19320 30012 19372
rect 30064 19320 30070 19372
rect 30834 19320 30840 19372
rect 30892 19320 30898 19372
rect 30926 19320 30932 19372
rect 30984 19360 30990 19372
rect 31938 19360 31944 19372
rect 30984 19332 31944 19360
rect 30984 19320 30990 19332
rect 31938 19320 31944 19332
rect 31996 19320 32002 19372
rect 32398 19320 32404 19372
rect 32456 19360 32462 19372
rect 34606 19360 34612 19372
rect 32456 19332 34612 19360
rect 32456 19320 32462 19332
rect 34606 19320 34612 19332
rect 34664 19320 34670 19372
rect 35066 19360 35072 19372
rect 34716 19332 35072 19360
rect 27856 19264 28856 19292
rect 28997 19295 29055 19301
rect 27856 19252 27862 19264
rect 28997 19261 29009 19295
rect 29043 19261 29055 19295
rect 28997 19255 29055 19261
rect 30285 19295 30343 19301
rect 30285 19261 30297 19295
rect 30331 19292 30343 19295
rect 32122 19292 32128 19304
rect 30331 19264 32128 19292
rect 30331 19261 30343 19264
rect 30285 19255 30343 19261
rect 26878 19224 26884 19236
rect 26252 19196 26884 19224
rect 26878 19184 26884 19196
rect 26936 19184 26942 19236
rect 27522 19184 27528 19236
rect 27580 19224 27586 19236
rect 30300 19224 30328 19255
rect 32122 19252 32128 19264
rect 32180 19252 32186 19304
rect 32858 19252 32864 19304
rect 32916 19252 32922 19304
rect 33962 19252 33968 19304
rect 34020 19252 34026 19304
rect 34149 19295 34207 19301
rect 34149 19261 34161 19295
rect 34195 19261 34207 19295
rect 34149 19255 34207 19261
rect 27580 19196 30328 19224
rect 34164 19224 34192 19255
rect 34514 19252 34520 19304
rect 34572 19292 34578 19304
rect 34716 19292 34744 19332
rect 35066 19320 35072 19332
rect 35124 19320 35130 19372
rect 35158 19320 35164 19372
rect 35216 19320 35222 19372
rect 35820 19360 35848 19400
rect 36170 19388 36176 19400
rect 36228 19388 36234 19440
rect 36265 19431 36323 19437
rect 36265 19397 36277 19431
rect 36311 19428 36323 19431
rect 36630 19428 36636 19440
rect 36311 19400 36636 19428
rect 36311 19397 36323 19400
rect 36265 19391 36323 19397
rect 36630 19388 36636 19400
rect 36688 19388 36694 19440
rect 39482 19428 39488 19440
rect 39422 19400 39488 19428
rect 39482 19388 39488 19400
rect 39540 19388 39546 19440
rect 39942 19388 39948 19440
rect 40000 19428 40006 19440
rect 41138 19428 41144 19440
rect 40000 19400 41144 19428
rect 40000 19388 40006 19400
rect 41138 19388 41144 19400
rect 41196 19388 41202 19440
rect 35268 19332 35848 19360
rect 34572 19264 34744 19292
rect 34572 19252 34578 19264
rect 35268 19224 35296 19332
rect 35894 19320 35900 19372
rect 35952 19320 35958 19372
rect 36357 19363 36415 19369
rect 36357 19329 36369 19363
rect 36403 19360 36415 19363
rect 37182 19360 37188 19372
rect 36403 19332 37188 19360
rect 36403 19329 36415 19332
rect 36357 19323 36415 19329
rect 37182 19320 37188 19332
rect 37240 19320 37246 19372
rect 37734 19320 37740 19372
rect 37792 19360 37798 19372
rect 37921 19363 37979 19369
rect 37921 19360 37933 19363
rect 37792 19332 37933 19360
rect 37792 19320 37798 19332
rect 37921 19329 37933 19332
rect 37967 19329 37979 19363
rect 37921 19323 37979 19329
rect 49142 19320 49148 19372
rect 49200 19320 49206 19372
rect 35345 19295 35403 19301
rect 35345 19261 35357 19295
rect 35391 19261 35403 19295
rect 35345 19255 35403 19261
rect 34164 19196 35296 19224
rect 27580 19184 27586 19196
rect 18782 19156 18788 19168
rect 17512 19128 18788 19156
rect 18782 19116 18788 19128
rect 18840 19116 18846 19168
rect 21082 19116 21088 19168
rect 21140 19156 21146 19168
rect 23474 19156 23480 19168
rect 21140 19128 23480 19156
rect 21140 19116 21146 19128
rect 23474 19116 23480 19128
rect 23532 19116 23538 19168
rect 25774 19116 25780 19168
rect 25832 19116 25838 19168
rect 26510 19116 26516 19168
rect 26568 19156 26574 19168
rect 33318 19156 33324 19168
rect 26568 19128 33324 19156
rect 26568 19116 26574 19128
rect 33318 19116 33324 19128
rect 33376 19116 33382 19168
rect 35360 19156 35388 19255
rect 35912 19233 35940 19320
rect 36541 19295 36599 19301
rect 36541 19261 36553 19295
rect 36587 19292 36599 19295
rect 37826 19292 37832 19304
rect 36587 19264 37832 19292
rect 36587 19261 36599 19264
rect 36541 19255 36599 19261
rect 37826 19252 37832 19264
rect 37884 19252 37890 19304
rect 38654 19292 38660 19304
rect 37936 19264 38660 19292
rect 35897 19227 35955 19233
rect 35897 19193 35909 19227
rect 35943 19193 35955 19227
rect 36170 19224 36176 19236
rect 35897 19187 35955 19193
rect 36004 19196 36176 19224
rect 36004 19156 36032 19196
rect 36170 19184 36176 19196
rect 36228 19224 36234 19236
rect 37936 19224 37964 19264
rect 38654 19252 38660 19264
rect 38712 19252 38718 19304
rect 39206 19252 39212 19304
rect 39264 19292 39270 19304
rect 40681 19295 40739 19301
rect 40681 19292 40693 19295
rect 39264 19264 40693 19292
rect 39264 19252 39270 19264
rect 40681 19261 40693 19264
rect 40727 19292 40739 19295
rect 40727 19264 41414 19292
rect 40727 19261 40739 19264
rect 40681 19255 40739 19261
rect 40494 19224 40500 19236
rect 36228 19196 37964 19224
rect 39224 19196 40500 19224
rect 36228 19184 36234 19196
rect 35360 19128 36032 19156
rect 36998 19116 37004 19168
rect 37056 19156 37062 19168
rect 38184 19159 38242 19165
rect 38184 19156 38196 19159
rect 37056 19128 38196 19156
rect 37056 19116 37062 19128
rect 38184 19125 38196 19128
rect 38230 19156 38242 19159
rect 39224 19156 39252 19196
rect 40494 19184 40500 19196
rect 40552 19184 40558 19236
rect 41386 19224 41414 19264
rect 41782 19224 41788 19236
rect 41386 19196 41788 19224
rect 41782 19184 41788 19196
rect 41840 19184 41846 19236
rect 38230 19128 39252 19156
rect 38230 19125 38242 19128
rect 38184 19119 38242 19125
rect 39666 19116 39672 19168
rect 39724 19116 39730 19168
rect 40126 19116 40132 19168
rect 40184 19116 40190 19168
rect 47394 19116 47400 19168
rect 47452 19156 47458 19168
rect 49237 19159 49295 19165
rect 49237 19156 49249 19159
rect 47452 19128 49249 19156
rect 47452 19116 47458 19128
rect 49237 19125 49249 19128
rect 49283 19125 49295 19159
rect 49237 19119 49295 19125
rect 1104 19066 49864 19088
rect 1104 19014 2950 19066
rect 3002 19014 3014 19066
rect 3066 19014 3078 19066
rect 3130 19014 3142 19066
rect 3194 19014 3206 19066
rect 3258 19014 12950 19066
rect 13002 19014 13014 19066
rect 13066 19014 13078 19066
rect 13130 19014 13142 19066
rect 13194 19014 13206 19066
rect 13258 19014 22950 19066
rect 23002 19014 23014 19066
rect 23066 19014 23078 19066
rect 23130 19014 23142 19066
rect 23194 19014 23206 19066
rect 23258 19014 32950 19066
rect 33002 19014 33014 19066
rect 33066 19014 33078 19066
rect 33130 19014 33142 19066
rect 33194 19014 33206 19066
rect 33258 19014 42950 19066
rect 43002 19014 43014 19066
rect 43066 19014 43078 19066
rect 43130 19014 43142 19066
rect 43194 19014 43206 19066
rect 43258 19014 49864 19066
rect 1104 18992 49864 19014
rect 9858 18952 9864 18964
rect 7760 18924 9864 18952
rect 1780 18788 3648 18816
rect 1780 18757 1808 18788
rect 1765 18751 1823 18757
rect 1765 18717 1777 18751
rect 1811 18717 1823 18751
rect 1765 18711 1823 18717
rect 2774 18640 2780 18692
rect 2832 18640 2838 18692
rect 3620 18680 3648 18788
rect 3694 18776 3700 18828
rect 3752 18816 3758 18828
rect 4433 18819 4491 18825
rect 4433 18816 4445 18819
rect 3752 18788 4445 18816
rect 3752 18776 3758 18788
rect 4433 18785 4445 18788
rect 4479 18785 4491 18819
rect 4433 18779 4491 18785
rect 4065 18751 4123 18757
rect 4065 18717 4077 18751
rect 4111 18748 4123 18751
rect 7760 18748 7788 18924
rect 9858 18912 9864 18924
rect 9916 18912 9922 18964
rect 10870 18912 10876 18964
rect 10928 18912 10934 18964
rect 10962 18912 10968 18964
rect 11020 18952 11026 18964
rect 11885 18955 11943 18961
rect 11885 18952 11897 18955
rect 11020 18924 11897 18952
rect 11020 18912 11026 18924
rect 11885 18921 11897 18924
rect 11931 18952 11943 18955
rect 11974 18952 11980 18964
rect 11931 18924 11980 18952
rect 11931 18921 11943 18924
rect 11885 18915 11943 18921
rect 11974 18912 11980 18924
rect 12032 18912 12038 18964
rect 12084 18924 15884 18952
rect 9122 18776 9128 18828
rect 9180 18776 9186 18828
rect 9401 18819 9459 18825
rect 9401 18785 9413 18819
rect 9447 18816 9459 18819
rect 11054 18816 11060 18828
rect 9447 18788 11060 18816
rect 9447 18785 9459 18788
rect 9401 18779 9459 18785
rect 11054 18776 11060 18788
rect 11112 18776 11118 18828
rect 4111 18720 7788 18748
rect 4111 18717 4123 18720
rect 4065 18711 4123 18717
rect 7834 18708 7840 18760
rect 7892 18748 7898 18760
rect 12084 18757 12112 18924
rect 12158 18844 12164 18896
rect 12216 18884 12222 18896
rect 12529 18887 12587 18893
rect 12529 18884 12541 18887
rect 12216 18856 12541 18884
rect 12216 18844 12222 18856
rect 12529 18853 12541 18856
rect 12575 18853 12587 18887
rect 12529 18847 12587 18853
rect 12989 18819 13047 18825
rect 12989 18785 13001 18819
rect 13035 18816 13047 18819
rect 13078 18816 13084 18828
rect 13035 18788 13084 18816
rect 13035 18785 13047 18788
rect 12989 18779 13047 18785
rect 13078 18776 13084 18788
rect 13136 18776 13142 18828
rect 13173 18819 13231 18825
rect 13173 18785 13185 18819
rect 13219 18816 13231 18819
rect 13354 18816 13360 18828
rect 13219 18788 13360 18816
rect 13219 18785 13231 18788
rect 13173 18779 13231 18785
rect 13354 18776 13360 18788
rect 13412 18776 13418 18828
rect 13722 18776 13728 18828
rect 13780 18816 13786 18828
rect 14277 18819 14335 18825
rect 14277 18816 14289 18819
rect 13780 18788 14289 18816
rect 13780 18776 13786 18788
rect 14277 18785 14289 18788
rect 14323 18785 14335 18819
rect 14277 18779 14335 18785
rect 14553 18819 14611 18825
rect 14553 18785 14565 18819
rect 14599 18816 14611 18819
rect 15194 18816 15200 18828
rect 14599 18788 15200 18816
rect 14599 18785 14611 18788
rect 14553 18779 14611 18785
rect 15194 18776 15200 18788
rect 15252 18776 15258 18828
rect 15286 18776 15292 18828
rect 15344 18816 15350 18828
rect 15746 18816 15752 18828
rect 15344 18788 15752 18816
rect 15344 18776 15350 18788
rect 8205 18751 8263 18757
rect 8205 18748 8217 18751
rect 7892 18720 8217 18748
rect 7892 18708 7898 18720
rect 8205 18717 8217 18720
rect 8251 18717 8263 18751
rect 8205 18711 8263 18717
rect 12069 18751 12127 18757
rect 12069 18717 12081 18751
rect 12115 18717 12127 18751
rect 15672 18734 15700 18788
rect 15746 18776 15752 18788
rect 15804 18776 15810 18828
rect 12069 18711 12127 18717
rect 11238 18680 11244 18692
rect 3620 18652 8432 18680
rect 10626 18652 11244 18680
rect 8294 18572 8300 18624
rect 8352 18572 8358 18624
rect 8404 18612 8432 18652
rect 11238 18640 11244 18652
rect 11296 18640 11302 18692
rect 11330 18640 11336 18692
rect 11388 18680 11394 18692
rect 12897 18683 12955 18689
rect 12897 18680 12909 18683
rect 11388 18652 11836 18680
rect 11388 18640 11394 18652
rect 11514 18612 11520 18624
rect 8404 18584 11520 18612
rect 11514 18572 11520 18584
rect 11572 18572 11578 18624
rect 11808 18612 11836 18652
rect 12084 18652 12909 18680
rect 12084 18612 12112 18652
rect 12897 18649 12909 18652
rect 12943 18649 12955 18683
rect 14826 18680 14832 18692
rect 12897 18643 12955 18649
rect 13004 18652 14832 18680
rect 11808 18584 12112 18612
rect 12158 18572 12164 18624
rect 12216 18612 12222 18624
rect 13004 18612 13032 18652
rect 14826 18640 14832 18652
rect 14884 18640 14890 18692
rect 15856 18680 15884 18924
rect 15930 18912 15936 18964
rect 15988 18952 15994 18964
rect 16025 18955 16083 18961
rect 16025 18952 16037 18955
rect 15988 18924 16037 18952
rect 15988 18912 15994 18924
rect 16025 18921 16037 18924
rect 16071 18921 16083 18955
rect 16025 18915 16083 18921
rect 16574 18912 16580 18964
rect 16632 18952 16638 18964
rect 16761 18955 16819 18961
rect 16761 18952 16773 18955
rect 16632 18924 16773 18952
rect 16632 18912 16638 18924
rect 16761 18921 16773 18924
rect 16807 18921 16819 18955
rect 16761 18915 16819 18921
rect 17218 18912 17224 18964
rect 17276 18952 17282 18964
rect 17957 18955 18015 18961
rect 17957 18952 17969 18955
rect 17276 18924 17969 18952
rect 17276 18912 17282 18924
rect 17957 18921 17969 18924
rect 18003 18921 18015 18955
rect 17957 18915 18015 18921
rect 18506 18912 18512 18964
rect 18564 18952 18570 18964
rect 19797 18955 19855 18961
rect 19797 18952 19809 18955
rect 18564 18924 19809 18952
rect 18564 18912 18570 18924
rect 19797 18921 19809 18924
rect 19843 18921 19855 18955
rect 19797 18915 19855 18921
rect 21560 18924 23980 18952
rect 21082 18884 21088 18896
rect 17236 18856 21088 18884
rect 17236 18825 17264 18856
rect 21082 18844 21088 18856
rect 21140 18844 21146 18896
rect 17221 18819 17279 18825
rect 17221 18785 17233 18819
rect 17267 18785 17279 18819
rect 17221 18779 17279 18785
rect 17313 18819 17371 18825
rect 17313 18785 17325 18819
rect 17359 18785 17371 18819
rect 17313 18779 17371 18785
rect 16022 18708 16028 18760
rect 16080 18748 16086 18760
rect 17129 18751 17187 18757
rect 17129 18748 17141 18751
rect 16080 18720 17141 18748
rect 16080 18708 16086 18720
rect 17129 18717 17141 18720
rect 17175 18717 17187 18751
rect 17328 18748 17356 18779
rect 17402 18776 17408 18828
rect 17460 18816 17466 18828
rect 18601 18819 18659 18825
rect 17460 18788 18460 18816
rect 17460 18776 17466 18788
rect 18432 18748 18460 18788
rect 18601 18785 18613 18819
rect 18647 18816 18659 18819
rect 18966 18816 18972 18828
rect 18647 18788 18972 18816
rect 18647 18785 18659 18788
rect 18601 18779 18659 18785
rect 18966 18776 18972 18788
rect 19024 18776 19030 18828
rect 20441 18819 20499 18825
rect 20441 18785 20453 18819
rect 20487 18816 20499 18819
rect 20990 18816 20996 18828
rect 20487 18788 20996 18816
rect 20487 18785 20499 18788
rect 20441 18779 20499 18785
rect 20990 18776 20996 18788
rect 21048 18776 21054 18828
rect 21560 18825 21588 18924
rect 21818 18884 21824 18896
rect 21652 18856 21824 18884
rect 21652 18825 21680 18856
rect 21818 18844 21824 18856
rect 21876 18844 21882 18896
rect 23952 18884 23980 18924
rect 24578 18912 24584 18964
rect 24636 18912 24642 18964
rect 24670 18912 24676 18964
rect 24728 18952 24734 18964
rect 28997 18955 29055 18961
rect 28997 18952 29009 18955
rect 24728 18924 29009 18952
rect 24728 18912 24734 18924
rect 28997 18921 29009 18924
rect 29043 18921 29055 18955
rect 28997 18915 29055 18921
rect 29730 18912 29736 18964
rect 29788 18952 29794 18964
rect 31481 18955 31539 18961
rect 31481 18952 31493 18955
rect 29788 18924 31493 18952
rect 29788 18912 29794 18924
rect 31481 18921 31493 18924
rect 31527 18921 31539 18955
rect 32490 18952 32496 18964
rect 31481 18915 31539 18921
rect 31588 18924 32496 18952
rect 25314 18884 25320 18896
rect 23952 18856 25320 18884
rect 25314 18844 25320 18856
rect 25372 18844 25378 18896
rect 25424 18856 25912 18884
rect 21545 18819 21603 18825
rect 21545 18785 21557 18819
rect 21591 18785 21603 18819
rect 21545 18779 21603 18785
rect 21637 18819 21695 18825
rect 21637 18785 21649 18819
rect 21683 18785 21695 18819
rect 21637 18779 21695 18785
rect 22186 18776 22192 18828
rect 22244 18816 22250 18828
rect 22557 18819 22615 18825
rect 22557 18816 22569 18819
rect 22244 18788 22569 18816
rect 22244 18776 22250 18788
rect 22557 18785 22569 18788
rect 22603 18816 22615 18819
rect 24486 18816 24492 18828
rect 22603 18788 24492 18816
rect 22603 18785 22615 18788
rect 22557 18779 22615 18785
rect 24486 18776 24492 18788
rect 24544 18776 24550 18828
rect 25038 18776 25044 18828
rect 25096 18776 25102 18828
rect 25225 18819 25283 18825
rect 25225 18785 25237 18819
rect 25271 18816 25283 18819
rect 25424 18816 25452 18856
rect 25271 18788 25452 18816
rect 25271 18785 25283 18788
rect 25225 18779 25283 18785
rect 20165 18751 20223 18757
rect 20165 18748 20177 18751
rect 17328 18720 18276 18748
rect 18432 18720 20177 18748
rect 17129 18711 17187 18717
rect 18138 18680 18144 18692
rect 15856 18652 18144 18680
rect 18138 18640 18144 18652
rect 18196 18640 18202 18692
rect 18248 18680 18276 18720
rect 20165 18717 20177 18720
rect 20211 18717 20223 18751
rect 20165 18711 20223 18717
rect 22278 18708 22284 18760
rect 22336 18708 22342 18760
rect 25240 18748 25268 18779
rect 25682 18776 25688 18828
rect 25740 18816 25746 18828
rect 25777 18819 25835 18825
rect 25777 18816 25789 18819
rect 25740 18788 25789 18816
rect 25740 18776 25746 18788
rect 25777 18785 25789 18788
rect 25823 18785 25835 18819
rect 25884 18816 25912 18856
rect 27154 18844 27160 18896
rect 27212 18844 27218 18896
rect 27522 18844 27528 18896
rect 27580 18844 27586 18896
rect 31588 18884 31616 18924
rect 32490 18912 32496 18924
rect 32548 18912 32554 18964
rect 32677 18955 32735 18961
rect 32677 18921 32689 18955
rect 32723 18952 32735 18955
rect 32766 18952 32772 18964
rect 32723 18924 32772 18952
rect 32723 18921 32735 18924
rect 32677 18915 32735 18921
rect 32766 18912 32772 18924
rect 32824 18912 32830 18964
rect 32950 18912 32956 18964
rect 33008 18952 33014 18964
rect 35986 18952 35992 18964
rect 33008 18924 35992 18952
rect 33008 18912 33014 18924
rect 35986 18912 35992 18924
rect 36044 18912 36050 18964
rect 36998 18912 37004 18964
rect 37056 18912 37062 18964
rect 41322 18952 41328 18964
rect 37108 18924 41328 18952
rect 28966 18856 31616 18884
rect 31956 18856 32260 18884
rect 27062 18816 27068 18828
rect 25884 18788 27068 18816
rect 25777 18779 25835 18785
rect 27062 18776 27068 18788
rect 27120 18776 27126 18828
rect 27172 18816 27200 18844
rect 28966 18816 28994 18856
rect 27172 18788 28994 18816
rect 30190 18776 30196 18828
rect 30248 18776 30254 18828
rect 30282 18776 30288 18828
rect 30340 18776 30346 18828
rect 31956 18825 31984 18856
rect 31941 18819 31999 18825
rect 31941 18785 31953 18819
rect 31987 18785 31999 18819
rect 31941 18779 31999 18785
rect 32125 18819 32183 18825
rect 32125 18785 32137 18819
rect 32171 18785 32183 18819
rect 32232 18816 32260 18856
rect 33244 18856 35388 18884
rect 32950 18816 32956 18828
rect 32232 18788 32956 18816
rect 32125 18779 32183 18785
rect 24688 18720 25268 18748
rect 29181 18751 29239 18757
rect 19058 18680 19064 18692
rect 18248 18652 19064 18680
rect 19058 18640 19064 18652
rect 19116 18640 19122 18692
rect 21266 18640 21272 18692
rect 21324 18680 21330 18692
rect 23014 18680 23020 18692
rect 21324 18652 23020 18680
rect 21324 18640 21330 18652
rect 23014 18640 23020 18652
rect 23072 18640 23078 18692
rect 12216 18584 13032 18612
rect 12216 18572 12222 18584
rect 13078 18572 13084 18624
rect 13136 18612 13142 18624
rect 15562 18612 15568 18624
rect 13136 18584 15568 18612
rect 13136 18572 13142 18584
rect 15562 18572 15568 18584
rect 15620 18572 15626 18624
rect 18322 18572 18328 18624
rect 18380 18572 18386 18624
rect 18417 18615 18475 18621
rect 18417 18581 18429 18615
rect 18463 18612 18475 18615
rect 19242 18612 19248 18624
rect 18463 18584 19248 18612
rect 18463 18581 18475 18584
rect 18417 18575 18475 18581
rect 19242 18572 19248 18584
rect 19300 18572 19306 18624
rect 20257 18615 20315 18621
rect 20257 18581 20269 18615
rect 20303 18612 20315 18615
rect 20438 18612 20444 18624
rect 20303 18584 20444 18612
rect 20303 18581 20315 18584
rect 20257 18575 20315 18581
rect 20438 18572 20444 18584
rect 20496 18572 20502 18624
rect 20714 18572 20720 18624
rect 20772 18612 20778 18624
rect 21085 18615 21143 18621
rect 21085 18612 21097 18615
rect 20772 18584 21097 18612
rect 20772 18572 20778 18584
rect 21085 18581 21097 18584
rect 21131 18581 21143 18615
rect 21085 18575 21143 18581
rect 21453 18615 21511 18621
rect 21453 18581 21465 18615
rect 21499 18612 21511 18615
rect 21542 18612 21548 18624
rect 21499 18584 21548 18612
rect 21499 18581 21511 18584
rect 21453 18575 21511 18581
rect 21542 18572 21548 18584
rect 21600 18572 21606 18624
rect 23842 18572 23848 18624
rect 23900 18612 23906 18624
rect 24029 18615 24087 18621
rect 24029 18612 24041 18615
rect 23900 18584 24041 18612
rect 23900 18572 23906 18584
rect 24029 18581 24041 18584
rect 24075 18612 24087 18615
rect 24688 18612 24716 18720
rect 29181 18717 29193 18751
rect 29227 18748 29239 18751
rect 30466 18748 30472 18760
rect 29227 18720 30472 18748
rect 29227 18717 29239 18720
rect 29181 18711 29239 18717
rect 30466 18708 30472 18720
rect 30524 18708 30530 18760
rect 25130 18640 25136 18692
rect 25188 18680 25194 18692
rect 26053 18683 26111 18689
rect 26053 18680 26065 18683
rect 25188 18652 26065 18680
rect 25188 18640 25194 18652
rect 26053 18649 26065 18652
rect 26099 18649 26111 18683
rect 26053 18643 26111 18649
rect 26602 18640 26608 18692
rect 26660 18640 26666 18692
rect 29270 18640 29276 18692
rect 29328 18680 29334 18692
rect 30101 18683 30159 18689
rect 30101 18680 30113 18683
rect 29328 18652 30113 18680
rect 29328 18640 29334 18652
rect 30101 18649 30113 18652
rect 30147 18649 30159 18683
rect 32140 18680 32168 18779
rect 32950 18776 32956 18788
rect 33008 18776 33014 18828
rect 33042 18776 33048 18828
rect 33100 18816 33106 18828
rect 33137 18819 33195 18825
rect 33137 18816 33149 18819
rect 33100 18788 33149 18816
rect 33100 18776 33106 18788
rect 33137 18785 33149 18788
rect 33183 18785 33195 18819
rect 33137 18779 33195 18785
rect 32490 18708 32496 18760
rect 32548 18748 32554 18760
rect 33244 18748 33272 18856
rect 33321 18819 33379 18825
rect 33321 18785 33333 18819
rect 33367 18816 33379 18819
rect 34882 18816 34888 18828
rect 33367 18788 34888 18816
rect 33367 18785 33379 18788
rect 33321 18779 33379 18785
rect 34882 18776 34888 18788
rect 34940 18776 34946 18828
rect 35250 18776 35256 18828
rect 35308 18776 35314 18828
rect 35360 18816 35388 18856
rect 37108 18816 37136 18924
rect 41322 18912 41328 18924
rect 41380 18912 41386 18964
rect 41782 18912 41788 18964
rect 41840 18912 41846 18964
rect 38013 18887 38071 18893
rect 38013 18853 38025 18887
rect 38059 18884 38071 18887
rect 40034 18884 40040 18896
rect 38059 18856 40040 18884
rect 38059 18853 38071 18856
rect 38013 18847 38071 18853
rect 40034 18844 40040 18856
rect 40092 18844 40098 18896
rect 35360 18788 37136 18816
rect 38286 18776 38292 18828
rect 38344 18816 38350 18828
rect 38565 18819 38623 18825
rect 38565 18816 38577 18819
rect 38344 18788 38577 18816
rect 38344 18776 38350 18788
rect 38565 18785 38577 18788
rect 38611 18785 38623 18819
rect 38565 18779 38623 18785
rect 39482 18776 39488 18828
rect 39540 18816 39546 18828
rect 39540 18788 41368 18816
rect 39540 18776 39546 18788
rect 32548 18720 33272 18748
rect 32548 18708 32554 18720
rect 37458 18708 37464 18760
rect 37516 18748 37522 18760
rect 38473 18751 38531 18757
rect 38473 18748 38485 18751
rect 37516 18720 38485 18748
rect 37516 18708 37522 18720
rect 38473 18717 38485 18720
rect 38519 18717 38531 18751
rect 38473 18711 38531 18717
rect 38654 18708 38660 18760
rect 38712 18748 38718 18760
rect 40037 18751 40095 18757
rect 40037 18748 40049 18751
rect 38712 18720 40049 18748
rect 38712 18708 38718 18720
rect 40037 18717 40049 18720
rect 40083 18717 40095 18751
rect 40037 18711 40095 18717
rect 35529 18683 35587 18689
rect 35529 18680 35541 18683
rect 32140 18652 35541 18680
rect 30101 18643 30159 18649
rect 35360 18624 35388 18652
rect 35529 18649 35541 18652
rect 35575 18649 35587 18683
rect 35529 18643 35587 18649
rect 36538 18640 36544 18692
rect 36596 18640 36602 18692
rect 37642 18640 37648 18692
rect 37700 18680 37706 18692
rect 39850 18680 39856 18692
rect 37700 18652 39856 18680
rect 37700 18640 37706 18652
rect 39850 18640 39856 18652
rect 39908 18680 39914 18692
rect 40313 18683 40371 18689
rect 40313 18680 40325 18683
rect 39908 18652 40325 18680
rect 39908 18640 39914 18652
rect 40313 18649 40325 18652
rect 40359 18649 40371 18683
rect 41340 18666 41368 18788
rect 48590 18708 48596 18760
rect 48648 18708 48654 18760
rect 49053 18751 49111 18757
rect 49053 18717 49065 18751
rect 49099 18748 49111 18751
rect 49142 18748 49148 18760
rect 49099 18720 49148 18748
rect 49099 18717 49111 18720
rect 49053 18711 49111 18717
rect 49142 18708 49148 18720
rect 49200 18708 49206 18760
rect 40313 18643 40371 18649
rect 24075 18584 24716 18612
rect 24075 18581 24087 18584
rect 24029 18575 24087 18581
rect 24854 18572 24860 18624
rect 24912 18612 24918 18624
rect 24949 18615 25007 18621
rect 24949 18612 24961 18615
rect 24912 18584 24961 18612
rect 24912 18572 24918 18584
rect 24949 18581 24961 18584
rect 24995 18581 25007 18615
rect 24949 18575 25007 18581
rect 27614 18572 27620 18624
rect 27672 18612 27678 18624
rect 29178 18612 29184 18624
rect 27672 18584 29184 18612
rect 27672 18572 27678 18584
rect 29178 18572 29184 18584
rect 29236 18572 29242 18624
rect 29733 18615 29791 18621
rect 29733 18581 29745 18615
rect 29779 18612 29791 18615
rect 29822 18612 29828 18624
rect 29779 18584 29828 18612
rect 29779 18581 29791 18584
rect 29733 18575 29791 18581
rect 29822 18572 29828 18584
rect 29880 18572 29886 18624
rect 31846 18572 31852 18624
rect 31904 18572 31910 18624
rect 32490 18572 32496 18624
rect 32548 18612 32554 18624
rect 33045 18615 33103 18621
rect 33045 18612 33057 18615
rect 32548 18584 33057 18612
rect 32548 18572 32554 18584
rect 33045 18581 33057 18584
rect 33091 18581 33103 18615
rect 33045 18575 33103 18581
rect 33410 18572 33416 18624
rect 33468 18612 33474 18624
rect 33686 18612 33692 18624
rect 33468 18584 33692 18612
rect 33468 18572 33474 18584
rect 33686 18572 33692 18584
rect 33744 18572 33750 18624
rect 35342 18572 35348 18624
rect 35400 18572 35406 18624
rect 38378 18572 38384 18624
rect 38436 18612 38442 18624
rect 47394 18612 47400 18624
rect 38436 18584 47400 18612
rect 38436 18572 38442 18584
rect 47394 18572 47400 18584
rect 47452 18572 47458 18624
rect 48406 18572 48412 18624
rect 48464 18572 48470 18624
rect 49234 18572 49240 18624
rect 49292 18572 49298 18624
rect 1104 18522 49864 18544
rect 1104 18470 7950 18522
rect 8002 18470 8014 18522
rect 8066 18470 8078 18522
rect 8130 18470 8142 18522
rect 8194 18470 8206 18522
rect 8258 18470 17950 18522
rect 18002 18470 18014 18522
rect 18066 18470 18078 18522
rect 18130 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 27950 18522
rect 28002 18470 28014 18522
rect 28066 18470 28078 18522
rect 28130 18470 28142 18522
rect 28194 18470 28206 18522
rect 28258 18470 37950 18522
rect 38002 18470 38014 18522
rect 38066 18470 38078 18522
rect 38130 18470 38142 18522
rect 38194 18470 38206 18522
rect 38258 18470 47950 18522
rect 48002 18470 48014 18522
rect 48066 18470 48078 18522
rect 48130 18470 48142 18522
rect 48194 18470 48206 18522
rect 48258 18470 49864 18522
rect 1104 18448 49864 18470
rect 5626 18368 5632 18420
rect 5684 18408 5690 18420
rect 7837 18411 7895 18417
rect 7837 18408 7849 18411
rect 5684 18380 7849 18408
rect 5684 18368 5690 18380
rect 7837 18377 7849 18380
rect 7883 18377 7895 18411
rect 7837 18371 7895 18377
rect 9766 18368 9772 18420
rect 9824 18368 9830 18420
rect 10410 18368 10416 18420
rect 10468 18408 10474 18420
rect 10781 18411 10839 18417
rect 10781 18408 10793 18411
rect 10468 18380 10793 18408
rect 10468 18368 10474 18380
rect 10781 18377 10793 18380
rect 10827 18377 10839 18411
rect 11146 18408 11152 18420
rect 10781 18371 10839 18377
rect 10888 18380 11152 18408
rect 10888 18340 10916 18380
rect 11146 18368 11152 18380
rect 11204 18368 11210 18420
rect 11238 18368 11244 18420
rect 11296 18408 11302 18420
rect 11974 18408 11980 18420
rect 11296 18380 11980 18408
rect 11296 18368 11302 18380
rect 11974 18368 11980 18380
rect 12032 18408 12038 18420
rect 12032 18380 12434 18408
rect 12032 18368 12038 18380
rect 12250 18340 12256 18352
rect 2746 18312 10916 18340
rect 10980 18312 12256 18340
rect 1765 18275 1823 18281
rect 1765 18241 1777 18275
rect 1811 18272 1823 18275
rect 2746 18272 2774 18312
rect 1811 18244 2774 18272
rect 1811 18241 1823 18244
rect 1765 18235 1823 18241
rect 3510 18232 3516 18284
rect 3568 18272 3574 18284
rect 4433 18275 4491 18281
rect 4433 18272 4445 18275
rect 3568 18244 4445 18272
rect 3568 18232 3574 18244
rect 4433 18241 4445 18244
rect 4479 18241 4491 18275
rect 4433 18235 4491 18241
rect 7745 18275 7803 18281
rect 7745 18241 7757 18275
rect 7791 18272 7803 18275
rect 9858 18272 9864 18284
rect 7791 18244 9864 18272
rect 7791 18241 7803 18244
rect 7745 18235 7803 18241
rect 9858 18232 9864 18244
rect 9916 18232 9922 18284
rect 9953 18275 10011 18281
rect 9953 18241 9965 18275
rect 9999 18241 10011 18275
rect 9953 18235 10011 18241
rect 2774 18164 2780 18216
rect 2832 18164 2838 18216
rect 4154 18164 4160 18216
rect 4212 18164 4218 18216
rect 9968 18068 9996 18235
rect 10980 18213 11008 18312
rect 12250 18300 12256 18312
rect 12308 18300 12314 18352
rect 12406 18340 12434 18380
rect 12618 18368 12624 18420
rect 12676 18408 12682 18420
rect 14277 18411 14335 18417
rect 14277 18408 14289 18411
rect 12676 18380 14289 18408
rect 12676 18368 12682 18380
rect 14277 18377 14289 18380
rect 14323 18377 14335 18411
rect 14277 18371 14335 18377
rect 14826 18368 14832 18420
rect 14884 18408 14890 18420
rect 15378 18408 15384 18420
rect 14884 18380 15384 18408
rect 14884 18368 14890 18380
rect 15378 18368 15384 18380
rect 15436 18368 15442 18420
rect 15470 18368 15476 18420
rect 15528 18368 15534 18420
rect 16114 18368 16120 18420
rect 16172 18368 16178 18420
rect 16758 18368 16764 18420
rect 16816 18408 16822 18420
rect 16853 18411 16911 18417
rect 16853 18408 16865 18411
rect 16816 18380 16865 18408
rect 16816 18368 16822 18380
rect 16853 18377 16865 18380
rect 16899 18377 16911 18411
rect 16853 18371 16911 18377
rect 17221 18411 17279 18417
rect 17221 18377 17233 18411
rect 17267 18408 17279 18411
rect 17310 18408 17316 18420
rect 17267 18380 17316 18408
rect 17267 18377 17279 18380
rect 17221 18371 17279 18377
rect 17310 18368 17316 18380
rect 17368 18368 17374 18420
rect 18598 18368 18604 18420
rect 18656 18368 18662 18420
rect 18693 18411 18751 18417
rect 18693 18377 18705 18411
rect 18739 18408 18751 18411
rect 24673 18411 24731 18417
rect 24673 18408 24685 18411
rect 18739 18380 24685 18408
rect 18739 18377 18751 18380
rect 18693 18371 18751 18377
rect 24673 18377 24685 18380
rect 24719 18377 24731 18411
rect 24673 18371 24731 18377
rect 25041 18411 25099 18417
rect 25041 18377 25053 18411
rect 25087 18408 25099 18411
rect 25774 18408 25780 18420
rect 25087 18380 25780 18408
rect 25087 18377 25099 18380
rect 25041 18371 25099 18377
rect 25774 18368 25780 18380
rect 25832 18368 25838 18420
rect 26237 18411 26295 18417
rect 26237 18377 26249 18411
rect 26283 18408 26295 18411
rect 27246 18408 27252 18420
rect 26283 18380 27252 18408
rect 26283 18377 26295 18380
rect 26237 18371 26295 18377
rect 27246 18368 27252 18380
rect 27304 18368 27310 18420
rect 27525 18411 27583 18417
rect 27525 18377 27537 18411
rect 27571 18408 27583 18411
rect 27614 18408 27620 18420
rect 27571 18380 27620 18408
rect 27571 18377 27583 18380
rect 27525 18371 27583 18377
rect 27614 18368 27620 18380
rect 27672 18368 27678 18420
rect 28905 18411 28963 18417
rect 28905 18377 28917 18411
rect 28951 18408 28963 18411
rect 29638 18408 29644 18420
rect 28951 18380 29644 18408
rect 28951 18377 28963 18380
rect 28905 18371 28963 18377
rect 29638 18368 29644 18380
rect 29696 18368 29702 18420
rect 30101 18411 30159 18417
rect 30101 18377 30113 18411
rect 30147 18408 30159 18411
rect 31202 18408 31208 18420
rect 30147 18380 31208 18408
rect 30147 18377 30159 18380
rect 30101 18371 30159 18377
rect 31202 18368 31208 18380
rect 31260 18368 31266 18420
rect 32309 18411 32367 18417
rect 32309 18377 32321 18411
rect 32355 18408 32367 18411
rect 36173 18411 36231 18417
rect 36173 18408 36185 18411
rect 32355 18380 36185 18408
rect 32355 18377 32367 18380
rect 32309 18371 32367 18377
rect 36173 18377 36185 18380
rect 36219 18377 36231 18411
rect 36173 18371 36231 18377
rect 36262 18368 36268 18420
rect 36320 18368 36326 18420
rect 37550 18368 37556 18420
rect 37608 18408 37614 18420
rect 37608 18380 39712 18408
rect 37608 18368 37614 18380
rect 12406 18312 12466 18340
rect 13814 18300 13820 18352
rect 13872 18340 13878 18352
rect 18616 18340 18644 18368
rect 18966 18340 18972 18352
rect 13872 18312 17448 18340
rect 18616 18312 18972 18340
rect 13872 18300 13878 18312
rect 15657 18275 15715 18281
rect 15657 18241 15669 18275
rect 15703 18272 15715 18275
rect 16301 18275 16359 18281
rect 15703 18244 16252 18272
rect 15703 18241 15715 18244
rect 15657 18235 15715 18241
rect 10873 18207 10931 18213
rect 10873 18173 10885 18207
rect 10919 18173 10931 18207
rect 10873 18167 10931 18173
rect 10965 18207 11023 18213
rect 10965 18173 10977 18207
rect 11011 18173 11023 18207
rect 10965 18167 11023 18173
rect 10042 18096 10048 18148
rect 10100 18136 10106 18148
rect 10413 18139 10471 18145
rect 10413 18136 10425 18139
rect 10100 18108 10425 18136
rect 10100 18096 10106 18108
rect 10413 18105 10425 18108
rect 10459 18105 10471 18139
rect 10888 18136 10916 18167
rect 11606 18164 11612 18216
rect 11664 18204 11670 18216
rect 11701 18207 11759 18213
rect 11701 18204 11713 18207
rect 11664 18176 11713 18204
rect 11664 18164 11670 18176
rect 11701 18173 11713 18176
rect 11747 18173 11759 18207
rect 11701 18167 11759 18173
rect 11977 18207 12035 18213
rect 11977 18173 11989 18207
rect 12023 18204 12035 18207
rect 13354 18204 13360 18216
rect 12023 18176 13360 18204
rect 12023 18173 12035 18176
rect 11977 18167 12035 18173
rect 13354 18164 13360 18176
rect 13412 18164 13418 18216
rect 13446 18164 13452 18216
rect 13504 18204 13510 18216
rect 14369 18207 14427 18213
rect 13504 18176 13952 18204
rect 13504 18164 13510 18176
rect 11422 18136 11428 18148
rect 10888 18108 11428 18136
rect 10413 18099 10471 18105
rect 11422 18096 11428 18108
rect 11480 18096 11486 18148
rect 13924 18145 13952 18176
rect 14369 18173 14381 18207
rect 14415 18173 14427 18207
rect 14369 18167 14427 18173
rect 14553 18207 14611 18213
rect 14553 18173 14565 18207
rect 14599 18204 14611 18207
rect 15194 18204 15200 18216
rect 14599 18176 15200 18204
rect 14599 18173 14611 18176
rect 14553 18167 14611 18173
rect 13909 18139 13967 18145
rect 13909 18105 13921 18139
rect 13955 18105 13967 18139
rect 14384 18136 14412 18167
rect 15194 18164 15200 18176
rect 15252 18204 15258 18216
rect 16022 18204 16028 18216
rect 15252 18176 16028 18204
rect 15252 18164 15258 18176
rect 16022 18164 16028 18176
rect 16080 18164 16086 18216
rect 16224 18204 16252 18244
rect 16301 18241 16313 18275
rect 16347 18272 16359 18275
rect 16347 18244 16528 18272
rect 16347 18241 16359 18244
rect 16301 18235 16359 18241
rect 16500 18216 16528 18244
rect 16390 18204 16396 18216
rect 16224 18176 16396 18204
rect 16390 18164 16396 18176
rect 16448 18164 16454 18216
rect 16482 18164 16488 18216
rect 16540 18164 16546 18216
rect 17420 18213 17448 18312
rect 18966 18300 18972 18312
rect 19024 18340 19030 18352
rect 19024 18312 19656 18340
rect 19024 18300 19030 18312
rect 18601 18275 18659 18281
rect 18601 18241 18613 18275
rect 18647 18272 18659 18275
rect 19518 18272 19524 18284
rect 18647 18244 19524 18272
rect 18647 18241 18659 18244
rect 18601 18235 18659 18241
rect 19518 18232 19524 18244
rect 19576 18232 19582 18284
rect 19628 18281 19656 18312
rect 22278 18300 22284 18352
rect 22336 18340 22342 18352
rect 22738 18340 22744 18352
rect 22336 18312 22744 18340
rect 22336 18300 22342 18312
rect 22738 18300 22744 18312
rect 22796 18340 22802 18352
rect 24121 18343 24179 18349
rect 24121 18340 24133 18343
rect 22796 18312 24133 18340
rect 22796 18300 22802 18312
rect 24121 18309 24133 18312
rect 24167 18340 24179 18343
rect 25682 18340 25688 18352
rect 24167 18312 25688 18340
rect 24167 18309 24179 18312
rect 24121 18303 24179 18309
rect 25682 18300 25688 18312
rect 25740 18300 25746 18352
rect 26344 18312 28764 18340
rect 19613 18275 19671 18281
rect 19613 18241 19625 18275
rect 19659 18241 19671 18275
rect 19613 18235 19671 18241
rect 20990 18232 20996 18284
rect 21048 18272 21054 18284
rect 21358 18272 21364 18284
rect 21048 18244 21364 18272
rect 21048 18232 21054 18244
rect 21358 18232 21364 18244
rect 21416 18232 21422 18284
rect 22370 18232 22376 18284
rect 22428 18232 22434 18284
rect 23290 18232 23296 18284
rect 23348 18232 23354 18284
rect 25133 18275 25191 18281
rect 25133 18241 25145 18275
rect 25179 18272 25191 18275
rect 26234 18272 26240 18284
rect 25179 18244 26240 18272
rect 25179 18241 25191 18244
rect 25133 18235 25191 18241
rect 26234 18232 26240 18244
rect 26292 18232 26298 18284
rect 26344 18281 26372 18312
rect 26329 18275 26387 18281
rect 26329 18241 26341 18275
rect 26375 18241 26387 18275
rect 26329 18235 26387 18241
rect 26786 18232 26792 18284
rect 26844 18272 26850 18284
rect 27522 18272 27528 18284
rect 26844 18244 27528 18272
rect 26844 18232 26850 18244
rect 27522 18232 27528 18244
rect 27580 18232 27586 18284
rect 27617 18275 27675 18281
rect 27617 18241 27629 18275
rect 27663 18272 27675 18275
rect 28736 18272 28764 18312
rect 28994 18300 29000 18352
rect 29052 18300 29058 18352
rect 30561 18343 30619 18349
rect 30561 18309 30573 18343
rect 30607 18340 30619 18343
rect 30742 18340 30748 18352
rect 30607 18312 30748 18340
rect 30607 18309 30619 18312
rect 30561 18303 30619 18309
rect 30742 18300 30748 18312
rect 30800 18300 30806 18352
rect 31570 18300 31576 18352
rect 31628 18340 31634 18352
rect 35250 18340 35256 18352
rect 31628 18312 33548 18340
rect 35098 18312 35256 18340
rect 31628 18300 31634 18312
rect 30374 18272 30380 18284
rect 27663 18244 28672 18272
rect 28736 18244 30380 18272
rect 27663 18241 27675 18244
rect 27617 18235 27675 18241
rect 17313 18207 17371 18213
rect 17313 18173 17325 18207
rect 17359 18173 17371 18207
rect 17313 18167 17371 18173
rect 17405 18207 17463 18213
rect 17405 18173 17417 18207
rect 17451 18173 17463 18207
rect 17405 18167 17463 18173
rect 18877 18207 18935 18213
rect 18877 18173 18889 18207
rect 18923 18204 18935 18207
rect 19889 18207 19947 18213
rect 19889 18204 19901 18207
rect 18923 18176 19901 18204
rect 18923 18173 18935 18176
rect 18877 18167 18935 18173
rect 19889 18173 19901 18176
rect 19935 18204 19947 18207
rect 20898 18204 20904 18216
rect 19935 18176 20904 18204
rect 19935 18173 19947 18176
rect 19889 18167 19947 18173
rect 16758 18136 16764 18148
rect 14384 18108 16764 18136
rect 13909 18099 13967 18105
rect 16758 18096 16764 18108
rect 16816 18096 16822 18148
rect 17328 18136 17356 18167
rect 20898 18164 20904 18176
rect 20956 18164 20962 18216
rect 21542 18164 21548 18216
rect 21600 18204 21606 18216
rect 21600 18176 22140 18204
rect 21600 18164 21606 18176
rect 18141 18139 18199 18145
rect 18141 18136 18153 18139
rect 17328 18108 18153 18136
rect 18141 18105 18153 18108
rect 18187 18136 18199 18139
rect 18187 18108 18552 18136
rect 18187 18105 18199 18108
rect 18141 18099 18199 18105
rect 11238 18068 11244 18080
rect 9968 18040 11244 18068
rect 11238 18028 11244 18040
rect 11296 18028 11302 18080
rect 12710 18028 12716 18080
rect 12768 18068 12774 18080
rect 13449 18071 13507 18077
rect 13449 18068 13461 18071
rect 12768 18040 13461 18068
rect 12768 18028 12774 18040
rect 13449 18037 13461 18040
rect 13495 18037 13507 18071
rect 13449 18031 13507 18037
rect 18230 18028 18236 18080
rect 18288 18028 18294 18080
rect 18524 18068 18552 18108
rect 21174 18068 21180 18080
rect 18524 18040 21180 18068
rect 21174 18028 21180 18040
rect 21232 18028 21238 18080
rect 21361 18071 21419 18077
rect 21361 18037 21373 18071
rect 21407 18068 21419 18071
rect 21450 18068 21456 18080
rect 21407 18040 21456 18068
rect 21407 18037 21419 18040
rect 21361 18031 21419 18037
rect 21450 18028 21456 18040
rect 21508 18028 21514 18080
rect 22002 18028 22008 18080
rect 22060 18028 22066 18080
rect 22112 18068 22140 18176
rect 22462 18164 22468 18216
rect 22520 18164 22526 18216
rect 22646 18164 22652 18216
rect 22704 18164 22710 18216
rect 25317 18207 25375 18213
rect 25317 18173 25329 18207
rect 25363 18204 25375 18207
rect 25498 18204 25504 18216
rect 25363 18176 25504 18204
rect 25363 18173 25375 18176
rect 25317 18167 25375 18173
rect 25498 18164 25504 18176
rect 25556 18164 25562 18216
rect 25958 18164 25964 18216
rect 26016 18204 26022 18216
rect 26421 18207 26479 18213
rect 26421 18204 26433 18207
rect 26016 18176 26433 18204
rect 26016 18164 26022 18176
rect 26421 18173 26433 18176
rect 26467 18173 26479 18207
rect 26421 18167 26479 18173
rect 26510 18164 26516 18216
rect 26568 18204 26574 18216
rect 27709 18207 27767 18213
rect 27709 18204 27721 18207
rect 26568 18176 27721 18204
rect 26568 18164 26574 18176
rect 27709 18173 27721 18176
rect 27755 18173 27767 18207
rect 27709 18167 27767 18173
rect 23014 18096 23020 18148
rect 23072 18136 23078 18148
rect 23474 18136 23480 18148
rect 23072 18108 23480 18136
rect 23072 18096 23078 18108
rect 23474 18096 23480 18108
rect 23532 18096 23538 18148
rect 23750 18096 23756 18148
rect 23808 18136 23814 18148
rect 25869 18139 25927 18145
rect 25869 18136 25881 18139
rect 23808 18108 25881 18136
rect 23808 18096 23814 18108
rect 25869 18105 25881 18108
rect 25915 18105 25927 18139
rect 28537 18139 28595 18145
rect 28537 18136 28549 18139
rect 25869 18099 25927 18105
rect 25976 18108 28549 18136
rect 23842 18068 23848 18080
rect 22112 18040 23848 18068
rect 23842 18028 23848 18040
rect 23900 18028 23906 18080
rect 23934 18028 23940 18080
rect 23992 18068 23998 18080
rect 25976 18068 26004 18108
rect 28537 18105 28549 18108
rect 28583 18105 28595 18139
rect 28537 18099 28595 18105
rect 23992 18040 26004 18068
rect 23992 18028 23998 18040
rect 26050 18028 26056 18080
rect 26108 18068 26114 18080
rect 27157 18071 27215 18077
rect 27157 18068 27169 18071
rect 26108 18040 27169 18068
rect 26108 18028 26114 18040
rect 27157 18037 27169 18040
rect 27203 18037 27215 18071
rect 27157 18031 27215 18037
rect 27614 18028 27620 18080
rect 27672 18068 27678 18080
rect 27798 18068 27804 18080
rect 27672 18040 27804 18068
rect 27672 18028 27678 18040
rect 27798 18028 27804 18040
rect 27856 18028 27862 18080
rect 28445 18071 28503 18077
rect 28445 18037 28457 18071
rect 28491 18068 28503 18071
rect 28644 18068 28672 18244
rect 30374 18232 30380 18244
rect 30432 18232 30438 18284
rect 30469 18275 30527 18281
rect 30469 18241 30481 18275
rect 30515 18272 30527 18275
rect 31481 18275 31539 18281
rect 31481 18272 31493 18275
rect 30515 18244 31493 18272
rect 30515 18241 30527 18244
rect 30469 18235 30527 18241
rect 31481 18241 31493 18244
rect 31527 18241 31539 18275
rect 31481 18235 31539 18241
rect 32030 18232 32036 18284
rect 32088 18272 32094 18284
rect 32677 18275 32735 18281
rect 32677 18272 32689 18275
rect 32088 18244 32689 18272
rect 32088 18232 32094 18244
rect 32677 18241 32689 18244
rect 32723 18241 32735 18275
rect 32677 18235 32735 18241
rect 28810 18164 28816 18216
rect 28868 18204 28874 18216
rect 29089 18207 29147 18213
rect 29089 18204 29101 18207
rect 28868 18176 29101 18204
rect 28868 18164 28874 18176
rect 29089 18173 29101 18176
rect 29135 18173 29147 18207
rect 29089 18167 29147 18173
rect 30745 18207 30803 18213
rect 30745 18173 30757 18207
rect 30791 18204 30803 18207
rect 32398 18204 32404 18216
rect 30791 18176 32404 18204
rect 30791 18173 30803 18176
rect 30745 18167 30803 18173
rect 32398 18164 32404 18176
rect 32456 18164 32462 18216
rect 32769 18207 32827 18213
rect 32769 18173 32781 18207
rect 32815 18173 32827 18207
rect 32769 18167 32827 18173
rect 32953 18207 33011 18213
rect 32953 18173 32965 18207
rect 32999 18204 33011 18207
rect 33410 18204 33416 18216
rect 32999 18176 33416 18204
rect 32999 18173 33011 18176
rect 32953 18167 33011 18173
rect 28902 18096 28908 18148
rect 28960 18136 28966 18148
rect 32784 18136 32812 18167
rect 33410 18164 33416 18176
rect 33468 18164 33474 18216
rect 28960 18108 32812 18136
rect 33520 18136 33548 18312
rect 35250 18300 35256 18312
rect 35308 18300 35314 18352
rect 35710 18300 35716 18352
rect 35768 18340 35774 18352
rect 38654 18340 38660 18352
rect 35768 18312 38660 18340
rect 35768 18300 35774 18312
rect 37274 18272 37280 18284
rect 35084 18244 37280 18272
rect 33594 18164 33600 18216
rect 33652 18164 33658 18216
rect 33873 18207 33931 18213
rect 33873 18204 33885 18207
rect 33704 18176 33885 18204
rect 33704 18136 33732 18176
rect 33873 18173 33885 18176
rect 33919 18204 33931 18207
rect 35084 18204 35112 18244
rect 37274 18232 37280 18244
rect 37332 18232 37338 18284
rect 38120 18281 38148 18312
rect 38654 18300 38660 18312
rect 38712 18300 38718 18352
rect 39684 18340 39712 18380
rect 39850 18368 39856 18420
rect 39908 18368 39914 18420
rect 40405 18411 40463 18417
rect 40405 18377 40417 18411
rect 40451 18377 40463 18411
rect 40405 18371 40463 18377
rect 40420 18340 40448 18371
rect 40862 18368 40868 18420
rect 40920 18368 40926 18420
rect 41414 18368 41420 18420
rect 41472 18408 41478 18420
rect 49234 18408 49240 18420
rect 41472 18380 49240 18408
rect 41472 18368 41478 18380
rect 49234 18368 49240 18380
rect 49292 18368 49298 18420
rect 39684 18312 40448 18340
rect 40773 18343 40831 18349
rect 40773 18309 40785 18343
rect 40819 18340 40831 18343
rect 48406 18340 48412 18352
rect 40819 18312 48412 18340
rect 40819 18309 40831 18312
rect 40773 18303 40831 18309
rect 48406 18300 48412 18312
rect 48464 18300 48470 18352
rect 38105 18275 38163 18281
rect 38105 18241 38117 18275
rect 38151 18241 38163 18275
rect 38105 18235 38163 18241
rect 39482 18232 39488 18284
rect 39540 18232 39546 18284
rect 49050 18232 49056 18284
rect 49108 18232 49114 18284
rect 33919 18176 35112 18204
rect 33919 18173 33931 18176
rect 33873 18167 33931 18173
rect 35342 18164 35348 18216
rect 35400 18164 35406 18216
rect 36354 18164 36360 18216
rect 36412 18164 36418 18216
rect 37550 18164 37556 18216
rect 37608 18204 37614 18216
rect 38381 18207 38439 18213
rect 38381 18204 38393 18207
rect 37608 18176 38393 18204
rect 37608 18164 37614 18176
rect 38381 18173 38393 18176
rect 38427 18204 38439 18207
rect 39666 18204 39672 18216
rect 38427 18176 39672 18204
rect 38427 18173 38439 18176
rect 38381 18167 38439 18173
rect 39666 18164 39672 18176
rect 39724 18204 39730 18216
rect 40957 18207 41015 18213
rect 40957 18204 40969 18207
rect 39724 18176 40969 18204
rect 39724 18164 39730 18176
rect 40957 18173 40969 18176
rect 41003 18173 41015 18207
rect 40957 18167 41015 18173
rect 36446 18136 36452 18148
rect 33520 18108 33732 18136
rect 35636 18108 36452 18136
rect 28960 18096 28966 18108
rect 30190 18068 30196 18080
rect 28491 18040 30196 18068
rect 28491 18037 28503 18040
rect 28445 18031 28503 18037
rect 30190 18028 30196 18040
rect 30248 18028 30254 18080
rect 30466 18028 30472 18080
rect 30524 18068 30530 18080
rect 35636 18068 35664 18108
rect 36446 18096 36452 18108
rect 36504 18096 36510 18148
rect 30524 18040 35664 18068
rect 35805 18071 35863 18077
rect 30524 18028 30530 18040
rect 35805 18037 35817 18071
rect 35851 18068 35863 18071
rect 38470 18068 38476 18080
rect 35851 18040 38476 18068
rect 35851 18037 35863 18040
rect 35805 18031 35863 18037
rect 38470 18028 38476 18040
rect 38528 18028 38534 18080
rect 45554 18028 45560 18080
rect 45612 18068 45618 18080
rect 49237 18071 49295 18077
rect 49237 18068 49249 18071
rect 45612 18040 49249 18068
rect 45612 18028 45618 18040
rect 49237 18037 49249 18040
rect 49283 18037 49295 18071
rect 49237 18031 49295 18037
rect 1104 17978 49864 18000
rect 1104 17926 2950 17978
rect 3002 17926 3014 17978
rect 3066 17926 3078 17978
rect 3130 17926 3142 17978
rect 3194 17926 3206 17978
rect 3258 17926 12950 17978
rect 13002 17926 13014 17978
rect 13066 17926 13078 17978
rect 13130 17926 13142 17978
rect 13194 17926 13206 17978
rect 13258 17926 22950 17978
rect 23002 17926 23014 17978
rect 23066 17926 23078 17978
rect 23130 17926 23142 17978
rect 23194 17926 23206 17978
rect 23258 17926 32950 17978
rect 33002 17926 33014 17978
rect 33066 17926 33078 17978
rect 33130 17926 33142 17978
rect 33194 17926 33206 17978
rect 33258 17926 42950 17978
rect 43002 17926 43014 17978
rect 43066 17926 43078 17978
rect 43130 17926 43142 17978
rect 43194 17926 43206 17978
rect 43258 17926 49864 17978
rect 1104 17904 49864 17926
rect 12250 17824 12256 17876
rect 12308 17864 12314 17876
rect 12345 17867 12403 17873
rect 12345 17864 12357 17867
rect 12308 17836 12357 17864
rect 12308 17824 12314 17836
rect 12345 17833 12357 17836
rect 12391 17833 12403 17867
rect 12345 17827 12403 17833
rect 12802 17824 12808 17876
rect 12860 17864 12866 17876
rect 12897 17867 12955 17873
rect 12897 17864 12909 17867
rect 12860 17836 12909 17864
rect 12860 17824 12866 17836
rect 12897 17833 12909 17836
rect 12943 17833 12955 17867
rect 12897 17827 12955 17833
rect 15102 17824 15108 17876
rect 15160 17864 15166 17876
rect 15160 17836 15976 17864
rect 15160 17824 15166 17836
rect 12526 17756 12532 17808
rect 12584 17796 12590 17808
rect 13541 17799 13599 17805
rect 13541 17796 13553 17799
rect 12584 17768 13553 17796
rect 12584 17756 12590 17768
rect 13541 17765 13553 17768
rect 13587 17765 13599 17799
rect 15948 17796 15976 17836
rect 16022 17824 16028 17876
rect 16080 17824 16086 17876
rect 16761 17867 16819 17873
rect 16761 17833 16773 17867
rect 16807 17864 16819 17867
rect 18322 17864 18328 17876
rect 16807 17836 18328 17864
rect 16807 17833 16819 17836
rect 16761 17827 16819 17833
rect 18322 17824 18328 17836
rect 18380 17824 18386 17876
rect 21910 17864 21916 17876
rect 19536 17836 21916 17864
rect 19429 17799 19487 17805
rect 19429 17796 19441 17799
rect 15948 17768 19441 17796
rect 13541 17759 13599 17765
rect 19429 17765 19441 17768
rect 19475 17765 19487 17799
rect 19429 17759 19487 17765
rect 1210 17688 1216 17740
rect 1268 17728 1274 17740
rect 2041 17731 2099 17737
rect 2041 17728 2053 17731
rect 1268 17700 2053 17728
rect 1268 17688 1274 17700
rect 2041 17697 2053 17700
rect 2087 17697 2099 17731
rect 11606 17728 11612 17740
rect 2041 17691 2099 17697
rect 10612 17700 11612 17728
rect 10612 17672 10640 17700
rect 11606 17688 11612 17700
rect 11664 17688 11670 17740
rect 13814 17688 13820 17740
rect 13872 17728 13878 17740
rect 13998 17728 14004 17740
rect 13872 17700 14004 17728
rect 13872 17688 13878 17700
rect 13998 17688 14004 17700
rect 14056 17728 14062 17740
rect 14277 17731 14335 17737
rect 14277 17728 14289 17731
rect 14056 17700 14289 17728
rect 14056 17688 14062 17700
rect 14277 17697 14289 17700
rect 14323 17728 14335 17731
rect 14323 17700 16068 17728
rect 14323 17697 14335 17700
rect 14277 17691 14335 17697
rect 1765 17663 1823 17669
rect 1765 17629 1777 17663
rect 1811 17660 1823 17663
rect 10502 17660 10508 17672
rect 1811 17632 10508 17660
rect 1811 17629 1823 17632
rect 1765 17623 1823 17629
rect 10502 17620 10508 17632
rect 10560 17620 10566 17672
rect 10594 17620 10600 17672
rect 10652 17620 10658 17672
rect 11974 17620 11980 17672
rect 12032 17620 12038 17672
rect 13081 17663 13139 17669
rect 13081 17629 13093 17663
rect 13127 17629 13139 17663
rect 13081 17623 13139 17629
rect 10873 17595 10931 17601
rect 10873 17561 10885 17595
rect 10919 17561 10931 17595
rect 10873 17555 10931 17561
rect 10888 17524 10916 17555
rect 12158 17524 12164 17536
rect 10888 17496 12164 17524
rect 12158 17484 12164 17496
rect 12216 17524 12222 17536
rect 12710 17524 12716 17536
rect 12216 17496 12716 17524
rect 12216 17484 12222 17496
rect 12710 17484 12716 17496
rect 12768 17484 12774 17536
rect 13096 17524 13124 17623
rect 13630 17620 13636 17672
rect 13688 17660 13694 17672
rect 13725 17663 13783 17669
rect 13725 17660 13737 17663
rect 13688 17632 13737 17660
rect 13688 17620 13694 17632
rect 13725 17629 13737 17632
rect 13771 17629 13783 17663
rect 16040 17660 16068 17700
rect 17126 17688 17132 17740
rect 17184 17728 17190 17740
rect 18693 17731 18751 17737
rect 18693 17728 18705 17731
rect 17184 17700 18705 17728
rect 17184 17688 17190 17700
rect 18693 17697 18705 17700
rect 18739 17728 18751 17731
rect 18966 17728 18972 17740
rect 18739 17700 18972 17728
rect 18739 17697 18751 17700
rect 18693 17691 18751 17697
rect 18966 17688 18972 17700
rect 19024 17688 19030 17740
rect 16040 17632 18736 17660
rect 13725 17623 13783 17629
rect 18708 17604 18736 17632
rect 14550 17552 14556 17604
rect 14608 17552 14614 17604
rect 15286 17552 15292 17604
rect 15344 17552 15350 17604
rect 17313 17595 17371 17601
rect 17313 17561 17325 17595
rect 17359 17592 17371 17595
rect 17359 17564 17724 17592
rect 17359 17561 17371 17564
rect 17313 17555 17371 17561
rect 16666 17524 16672 17536
rect 13096 17496 16672 17524
rect 16666 17484 16672 17496
rect 16724 17484 16730 17536
rect 17218 17484 17224 17536
rect 17276 17524 17282 17536
rect 17405 17527 17463 17533
rect 17405 17524 17417 17527
rect 17276 17496 17417 17524
rect 17276 17484 17282 17496
rect 17405 17493 17417 17496
rect 17451 17493 17463 17527
rect 17696 17524 17724 17564
rect 17770 17552 17776 17604
rect 17828 17592 17834 17604
rect 17957 17595 18015 17601
rect 17957 17592 17969 17595
rect 17828 17564 17969 17592
rect 17828 17552 17834 17564
rect 17957 17561 17969 17564
rect 18003 17561 18015 17595
rect 17957 17555 18015 17561
rect 18690 17552 18696 17604
rect 18748 17552 18754 17604
rect 19536 17524 19564 17836
rect 21910 17824 21916 17836
rect 21968 17824 21974 17876
rect 22830 17824 22836 17876
rect 22888 17864 22894 17876
rect 23293 17867 23351 17873
rect 23293 17864 23305 17867
rect 22888 17836 23305 17864
rect 22888 17824 22894 17836
rect 23293 17833 23305 17836
rect 23339 17833 23351 17867
rect 23293 17827 23351 17833
rect 23842 17824 23848 17876
rect 23900 17864 23906 17876
rect 25225 17867 25283 17873
rect 25225 17864 25237 17867
rect 23900 17836 25237 17864
rect 23900 17824 23906 17836
rect 25225 17833 25237 17836
rect 25271 17833 25283 17867
rect 30098 17864 30104 17876
rect 25225 17827 25283 17833
rect 25792 17836 30104 17864
rect 21634 17756 21640 17808
rect 21692 17796 21698 17808
rect 24581 17799 24639 17805
rect 24581 17796 24593 17799
rect 21692 17768 24593 17796
rect 21692 17756 21698 17768
rect 24581 17765 24593 17768
rect 24627 17765 24639 17799
rect 24581 17759 24639 17765
rect 20257 17731 20315 17737
rect 20257 17697 20269 17731
rect 20303 17728 20315 17731
rect 20530 17728 20536 17740
rect 20303 17700 20536 17728
rect 20303 17697 20315 17700
rect 20257 17691 20315 17697
rect 20530 17688 20536 17700
rect 20588 17688 20594 17740
rect 23658 17688 23664 17740
rect 23716 17728 23722 17740
rect 23845 17731 23903 17737
rect 23845 17728 23857 17731
rect 23716 17700 23857 17728
rect 23716 17688 23722 17700
rect 23845 17697 23857 17700
rect 23891 17697 23903 17731
rect 25792 17728 25820 17836
rect 30098 17824 30104 17836
rect 30156 17824 30162 17876
rect 30374 17824 30380 17876
rect 30432 17864 30438 17876
rect 32766 17864 32772 17876
rect 30432 17836 32772 17864
rect 30432 17824 30438 17836
rect 32766 17824 32772 17836
rect 32824 17824 32830 17876
rect 34606 17864 34612 17876
rect 32876 17836 34612 17864
rect 28350 17756 28356 17808
rect 28408 17796 28414 17808
rect 32674 17796 32680 17808
rect 28408 17768 32680 17796
rect 28408 17756 28414 17768
rect 32674 17756 32680 17768
rect 32732 17756 32738 17808
rect 23845 17691 23903 17697
rect 24780 17700 25820 17728
rect 25869 17731 25927 17737
rect 19613 17663 19671 17669
rect 19613 17629 19625 17663
rect 19659 17629 19671 17663
rect 19613 17623 19671 17629
rect 17696 17496 19564 17524
rect 19628 17524 19656 17623
rect 22646 17620 22652 17672
rect 22704 17620 22710 17672
rect 24780 17669 24808 17700
rect 25869 17697 25881 17731
rect 25915 17728 25927 17731
rect 26326 17728 26332 17740
rect 25915 17700 26332 17728
rect 25915 17697 25927 17700
rect 25869 17691 25927 17697
rect 26326 17688 26332 17700
rect 26384 17688 26390 17740
rect 28534 17728 28540 17740
rect 27080 17700 28540 17728
rect 24765 17663 24823 17669
rect 24765 17629 24777 17663
rect 24811 17629 24823 17663
rect 24765 17623 24823 17629
rect 25406 17620 25412 17672
rect 25464 17660 25470 17672
rect 27080 17669 27108 17700
rect 28534 17688 28540 17700
rect 28592 17728 28598 17740
rect 30926 17728 30932 17740
rect 28592 17700 30932 17728
rect 28592 17688 28598 17700
rect 30926 17688 30932 17700
rect 30984 17688 30990 17740
rect 31662 17688 31668 17740
rect 31720 17728 31726 17740
rect 32125 17731 32183 17737
rect 32125 17728 32137 17731
rect 31720 17700 32137 17728
rect 31720 17688 31726 17700
rect 32125 17697 32137 17700
rect 32171 17697 32183 17731
rect 32876 17728 32904 17836
rect 34606 17824 34612 17836
rect 34664 17824 34670 17876
rect 36814 17864 36820 17876
rect 35636 17836 36820 17864
rect 34882 17796 34888 17808
rect 32125 17691 32183 17697
rect 32600 17700 32904 17728
rect 32968 17768 34888 17796
rect 27065 17663 27123 17669
rect 27065 17660 27077 17663
rect 25464 17632 27077 17660
rect 25464 17620 25470 17632
rect 27065 17629 27077 17632
rect 27111 17629 27123 17663
rect 27065 17623 27123 17629
rect 30193 17663 30251 17669
rect 30193 17629 30205 17663
rect 30239 17660 30251 17663
rect 30834 17660 30840 17672
rect 30239 17632 30840 17660
rect 30239 17629 30251 17632
rect 30193 17623 30251 17629
rect 30834 17620 30840 17632
rect 30892 17660 30898 17672
rect 32600 17660 32628 17700
rect 30892 17632 32628 17660
rect 30892 17620 30898 17632
rect 20254 17552 20260 17604
rect 20312 17592 20318 17604
rect 20533 17595 20591 17601
rect 20533 17592 20545 17595
rect 20312 17564 20545 17592
rect 20312 17552 20318 17564
rect 20533 17561 20545 17564
rect 20579 17592 20591 17595
rect 20622 17592 20628 17604
rect 20579 17564 20628 17592
rect 20579 17561 20591 17564
rect 20533 17555 20591 17561
rect 20622 17552 20628 17564
rect 20680 17552 20686 17604
rect 20990 17552 20996 17604
rect 21048 17552 21054 17604
rect 22186 17592 22192 17604
rect 21836 17564 22192 17592
rect 21836 17524 21864 17564
rect 22186 17552 22192 17564
rect 22244 17552 22250 17604
rect 23106 17552 23112 17604
rect 23164 17592 23170 17604
rect 25682 17592 25688 17604
rect 23164 17564 25688 17592
rect 23164 17552 23170 17564
rect 25682 17552 25688 17564
rect 25740 17552 25746 17604
rect 26786 17552 26792 17604
rect 26844 17592 26850 17604
rect 27341 17595 27399 17601
rect 27341 17592 27353 17595
rect 26844 17564 27353 17592
rect 26844 17552 26850 17564
rect 27341 17561 27353 17564
rect 27387 17561 27399 17595
rect 27341 17555 27399 17561
rect 27798 17552 27804 17604
rect 27856 17552 27862 17604
rect 28626 17552 28632 17604
rect 28684 17592 28690 17604
rect 28684 17564 31754 17592
rect 28684 17552 28690 17564
rect 19628 17496 21864 17524
rect 17405 17487 17463 17493
rect 21910 17484 21916 17536
rect 21968 17524 21974 17536
rect 22005 17527 22063 17533
rect 22005 17524 22017 17527
rect 21968 17496 22017 17524
rect 21968 17484 21974 17496
rect 22005 17493 22017 17496
rect 22051 17493 22063 17527
rect 22005 17487 22063 17493
rect 22462 17484 22468 17536
rect 22520 17484 22526 17536
rect 23658 17484 23664 17536
rect 23716 17484 23722 17536
rect 23750 17484 23756 17536
rect 23808 17484 23814 17536
rect 25590 17484 25596 17536
rect 25648 17484 25654 17536
rect 25866 17484 25872 17536
rect 25924 17524 25930 17536
rect 28810 17524 28816 17536
rect 25924 17496 28816 17524
rect 25924 17484 25930 17496
rect 28810 17484 28816 17496
rect 28868 17484 28874 17536
rect 28902 17484 28908 17536
rect 28960 17524 28966 17536
rect 30374 17524 30380 17536
rect 28960 17496 30380 17524
rect 28960 17484 28966 17496
rect 30374 17484 30380 17496
rect 30432 17484 30438 17536
rect 31478 17484 31484 17536
rect 31536 17524 31542 17536
rect 31573 17527 31631 17533
rect 31573 17524 31585 17527
rect 31536 17496 31585 17524
rect 31536 17484 31542 17496
rect 31573 17493 31585 17496
rect 31619 17493 31631 17527
rect 31726 17524 31754 17564
rect 31938 17552 31944 17604
rect 31996 17552 32002 17604
rect 32033 17595 32091 17601
rect 32033 17561 32045 17595
rect 32079 17592 32091 17595
rect 32214 17592 32220 17604
rect 32079 17564 32220 17592
rect 32079 17561 32091 17564
rect 32033 17555 32091 17561
rect 32214 17552 32220 17564
rect 32272 17552 32278 17604
rect 32968 17592 32996 17768
rect 34882 17756 34888 17768
rect 34940 17756 34946 17808
rect 33226 17688 33232 17740
rect 33284 17688 33290 17740
rect 33413 17731 33471 17737
rect 33413 17697 33425 17731
rect 33459 17728 33471 17731
rect 35636 17728 35664 17836
rect 36814 17824 36820 17836
rect 36872 17824 36878 17876
rect 37182 17824 37188 17876
rect 37240 17864 37246 17876
rect 40497 17867 40555 17873
rect 40497 17864 40509 17867
rect 37240 17836 40509 17864
rect 37240 17824 37246 17836
rect 40497 17833 40509 17836
rect 40543 17833 40555 17867
rect 40497 17827 40555 17833
rect 37274 17756 37280 17808
rect 37332 17796 37338 17808
rect 37553 17799 37611 17805
rect 37553 17796 37565 17799
rect 37332 17768 37565 17796
rect 37332 17756 37338 17768
rect 37553 17765 37565 17768
rect 37599 17765 37611 17799
rect 37553 17759 37611 17765
rect 38013 17799 38071 17805
rect 38013 17765 38025 17799
rect 38059 17796 38071 17799
rect 40862 17796 40868 17808
rect 38059 17768 40868 17796
rect 38059 17765 38071 17768
rect 38013 17759 38071 17765
rect 40862 17756 40868 17768
rect 40920 17756 40926 17808
rect 33459 17700 35664 17728
rect 33459 17697 33471 17700
rect 33413 17691 33471 17697
rect 35710 17688 35716 17740
rect 35768 17728 35774 17740
rect 35805 17731 35863 17737
rect 35805 17728 35817 17731
rect 35768 17700 35817 17728
rect 35768 17688 35774 17700
rect 35805 17697 35817 17700
rect 35851 17697 35863 17731
rect 35805 17691 35863 17697
rect 36081 17731 36139 17737
rect 36081 17697 36093 17731
rect 36127 17728 36139 17731
rect 36170 17728 36176 17740
rect 36127 17700 36176 17728
rect 36127 17697 36139 17700
rect 36081 17691 36139 17697
rect 36170 17688 36176 17700
rect 36228 17688 36234 17740
rect 38470 17688 38476 17740
rect 38528 17688 38534 17740
rect 38565 17731 38623 17737
rect 38565 17697 38577 17731
rect 38611 17697 38623 17731
rect 38565 17691 38623 17697
rect 35066 17620 35072 17672
rect 35124 17620 35130 17672
rect 37366 17620 37372 17672
rect 37424 17660 37430 17672
rect 38580 17660 38608 17691
rect 40126 17688 40132 17740
rect 40184 17728 40190 17740
rect 40957 17731 41015 17737
rect 40957 17728 40969 17731
rect 40184 17700 40969 17728
rect 40184 17688 40190 17700
rect 40957 17697 40969 17700
rect 41003 17697 41015 17731
rect 40957 17691 41015 17697
rect 41049 17731 41107 17737
rect 41049 17697 41061 17731
rect 41095 17697 41107 17731
rect 41049 17691 41107 17697
rect 37424 17632 38608 17660
rect 37424 17620 37430 17632
rect 40678 17620 40684 17672
rect 40736 17660 40742 17672
rect 41064 17660 41092 17691
rect 40736 17632 41092 17660
rect 40736 17620 40742 17632
rect 49050 17620 49056 17672
rect 49108 17620 49114 17672
rect 35986 17592 35992 17604
rect 32692 17564 32996 17592
rect 33060 17564 35992 17592
rect 32692 17524 32720 17564
rect 31726 17496 32720 17524
rect 32769 17527 32827 17533
rect 31573 17487 31631 17493
rect 32769 17493 32781 17527
rect 32815 17524 32827 17527
rect 33060 17524 33088 17564
rect 35986 17552 35992 17564
rect 36044 17552 36050 17604
rect 36538 17552 36544 17604
rect 36596 17552 36602 17604
rect 38381 17595 38439 17601
rect 38381 17592 38393 17595
rect 37384 17564 38393 17592
rect 32815 17496 33088 17524
rect 33137 17527 33195 17533
rect 32815 17493 32827 17496
rect 32769 17487 32827 17493
rect 33137 17493 33149 17527
rect 33183 17524 33195 17527
rect 34238 17524 34244 17536
rect 33183 17496 34244 17524
rect 33183 17493 33195 17496
rect 33137 17487 33195 17493
rect 34238 17484 34244 17496
rect 34296 17484 34302 17536
rect 34514 17484 34520 17536
rect 34572 17524 34578 17536
rect 37384 17524 37412 17564
rect 38381 17561 38393 17564
rect 38427 17561 38439 17595
rect 38381 17555 38439 17561
rect 40865 17595 40923 17601
rect 40865 17561 40877 17595
rect 40911 17592 40923 17595
rect 48406 17592 48412 17604
rect 40911 17564 48412 17592
rect 40911 17561 40923 17564
rect 40865 17555 40923 17561
rect 48406 17552 48412 17564
rect 48464 17552 48470 17604
rect 34572 17496 37412 17524
rect 34572 17484 34578 17496
rect 47394 17484 47400 17536
rect 47452 17524 47458 17536
rect 49237 17527 49295 17533
rect 49237 17524 49249 17527
rect 47452 17496 49249 17524
rect 47452 17484 47458 17496
rect 49237 17493 49249 17496
rect 49283 17493 49295 17527
rect 49237 17487 49295 17493
rect 1104 17434 49864 17456
rect 1104 17382 7950 17434
rect 8002 17382 8014 17434
rect 8066 17382 8078 17434
rect 8130 17382 8142 17434
rect 8194 17382 8206 17434
rect 8258 17382 17950 17434
rect 18002 17382 18014 17434
rect 18066 17382 18078 17434
rect 18130 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 27950 17434
rect 28002 17382 28014 17434
rect 28066 17382 28078 17434
rect 28130 17382 28142 17434
rect 28194 17382 28206 17434
rect 28258 17382 37950 17434
rect 38002 17382 38014 17434
rect 38066 17382 38078 17434
rect 38130 17382 38142 17434
rect 38194 17382 38206 17434
rect 38258 17382 47950 17434
rect 48002 17382 48014 17434
rect 48066 17382 48078 17434
rect 48130 17382 48142 17434
rect 48194 17382 48206 17434
rect 48258 17382 49864 17434
rect 1104 17360 49864 17382
rect 10413 17323 10471 17329
rect 10413 17289 10425 17323
rect 10459 17320 10471 17323
rect 12618 17320 12624 17332
rect 10459 17292 12624 17320
rect 10459 17289 10471 17292
rect 10413 17283 10471 17289
rect 12618 17280 12624 17292
rect 12676 17280 12682 17332
rect 12713 17323 12771 17329
rect 12713 17289 12725 17323
rect 12759 17320 12771 17323
rect 13354 17320 13360 17332
rect 12759 17292 13360 17320
rect 12759 17289 12771 17292
rect 12713 17283 12771 17289
rect 13354 17280 13360 17292
rect 13412 17280 13418 17332
rect 15562 17280 15568 17332
rect 15620 17280 15626 17332
rect 18782 17280 18788 17332
rect 18840 17320 18846 17332
rect 18840 17292 20852 17320
rect 18840 17280 18846 17292
rect 5350 17212 5356 17264
rect 5408 17252 5414 17264
rect 13173 17255 13231 17261
rect 13173 17252 13185 17255
rect 5408 17224 13185 17252
rect 5408 17212 5414 17224
rect 13173 17221 13185 17224
rect 13219 17221 13231 17255
rect 13173 17215 13231 17221
rect 14182 17212 14188 17264
rect 14240 17212 14246 17264
rect 14458 17212 14464 17264
rect 14516 17252 14522 17264
rect 16945 17255 17003 17261
rect 14516 17224 16712 17252
rect 14516 17212 14522 17224
rect 1765 17187 1823 17193
rect 1765 17153 1777 17187
rect 1811 17184 1823 17187
rect 8294 17184 8300 17196
rect 1811 17156 8300 17184
rect 1811 17153 1823 17156
rect 1765 17147 1823 17153
rect 8294 17144 8300 17156
rect 8352 17144 8358 17196
rect 10686 17144 10692 17196
rect 10744 17184 10750 17196
rect 10781 17187 10839 17193
rect 10781 17184 10793 17187
rect 10744 17156 10793 17184
rect 10744 17144 10750 17156
rect 10781 17153 10793 17156
rect 10827 17153 10839 17187
rect 10781 17147 10839 17153
rect 11514 17144 11520 17196
rect 11572 17184 11578 17196
rect 11793 17187 11851 17193
rect 11572 17156 11744 17184
rect 11572 17144 11578 17156
rect 1302 17076 1308 17128
rect 1360 17116 1366 17128
rect 2041 17119 2099 17125
rect 2041 17116 2053 17119
rect 1360 17088 2053 17116
rect 1360 17076 1366 17088
rect 2041 17085 2053 17088
rect 2087 17085 2099 17119
rect 2041 17079 2099 17085
rect 10226 17076 10232 17128
rect 10284 17116 10290 17128
rect 10410 17116 10416 17128
rect 10284 17088 10416 17116
rect 10284 17076 10290 17088
rect 10410 17076 10416 17088
rect 10468 17116 10474 17128
rect 10873 17119 10931 17125
rect 10873 17116 10885 17119
rect 10468 17088 10885 17116
rect 10468 17076 10474 17088
rect 10873 17085 10885 17088
rect 10919 17085 10931 17119
rect 10873 17079 10931 17085
rect 10962 17076 10968 17128
rect 11020 17076 11026 17128
rect 11716 17116 11744 17156
rect 11793 17153 11805 17187
rect 11839 17184 11851 17187
rect 12066 17184 12072 17196
rect 11839 17156 12072 17184
rect 11839 17153 11851 17156
rect 11793 17147 11851 17153
rect 12066 17144 12072 17156
rect 12124 17144 12130 17196
rect 12434 17144 12440 17196
rect 12492 17184 12498 17196
rect 13081 17187 13139 17193
rect 13081 17184 13093 17187
rect 12492 17156 13093 17184
rect 12492 17144 12498 17156
rect 13081 17153 13093 17156
rect 13127 17153 13139 17187
rect 13081 17147 13139 17153
rect 15381 17187 15439 17193
rect 15381 17153 15393 17187
rect 15427 17184 15439 17187
rect 15654 17184 15660 17196
rect 15427 17156 15660 17184
rect 15427 17153 15439 17156
rect 15381 17147 15439 17153
rect 15654 17144 15660 17156
rect 15712 17144 15718 17196
rect 15746 17144 15752 17196
rect 15804 17184 15810 17196
rect 15933 17187 15991 17193
rect 15933 17184 15945 17187
rect 15804 17156 15945 17184
rect 15804 17144 15810 17156
rect 15933 17153 15945 17156
rect 15979 17153 15991 17187
rect 15933 17147 15991 17153
rect 16025 17187 16083 17193
rect 16025 17153 16037 17187
rect 16071 17184 16083 17187
rect 16574 17184 16580 17196
rect 16071 17156 16580 17184
rect 16071 17153 16083 17156
rect 16025 17147 16083 17153
rect 11977 17119 12035 17125
rect 11977 17116 11989 17119
rect 11716 17088 11989 17116
rect 11977 17085 11989 17088
rect 12023 17085 12035 17119
rect 11977 17079 12035 17085
rect 12250 17076 12256 17128
rect 12308 17116 12314 17128
rect 13265 17119 13323 17125
rect 13265 17116 13277 17119
rect 12308 17088 13277 17116
rect 12308 17076 12314 17088
rect 13265 17085 13277 17088
rect 13311 17116 13323 17119
rect 15010 17116 15016 17128
rect 13311 17088 15016 17116
rect 13311 17085 13323 17088
rect 13265 17079 13323 17085
rect 15010 17076 15016 17088
rect 15068 17076 15074 17128
rect 15105 17119 15163 17125
rect 15105 17085 15117 17119
rect 15151 17116 15163 17119
rect 16040 17116 16068 17147
rect 16574 17144 16580 17156
rect 16632 17144 16638 17196
rect 16684 17184 16712 17224
rect 16945 17221 16957 17255
rect 16991 17252 17003 17255
rect 19150 17252 19156 17264
rect 16991 17224 19156 17252
rect 16991 17221 17003 17224
rect 16945 17215 17003 17221
rect 19150 17212 19156 17224
rect 19208 17212 19214 17264
rect 19610 17252 19616 17264
rect 19260 17224 19616 17252
rect 16684 17156 17172 17184
rect 15151 17088 16068 17116
rect 16117 17119 16175 17125
rect 15151 17085 15163 17088
rect 15105 17079 15163 17085
rect 16117 17085 16129 17119
rect 16163 17085 16175 17119
rect 16117 17079 16175 17085
rect 6822 17008 6828 17060
rect 6880 17048 6886 17060
rect 14369 17051 14427 17057
rect 14369 17048 14381 17051
rect 6880 17020 14381 17048
rect 6880 17008 6886 17020
rect 14369 17017 14381 17020
rect 14415 17017 14427 17051
rect 14369 17011 14427 17017
rect 15286 17008 15292 17060
rect 15344 17048 15350 17060
rect 15344 17020 15608 17048
rect 15344 17008 15350 17020
rect 9858 16940 9864 16992
rect 9916 16980 9922 16992
rect 15197 16983 15255 16989
rect 15197 16980 15209 16983
rect 9916 16952 15209 16980
rect 9916 16940 9922 16952
rect 15197 16949 15209 16952
rect 15243 16980 15255 16983
rect 15470 16980 15476 16992
rect 15243 16952 15476 16980
rect 15243 16949 15255 16952
rect 15197 16943 15255 16949
rect 15470 16940 15476 16952
rect 15528 16940 15534 16992
rect 15580 16980 15608 17020
rect 15930 17008 15936 17060
rect 15988 17048 15994 17060
rect 16132 17048 16160 17079
rect 15988 17020 16160 17048
rect 15988 17008 15994 17020
rect 17037 16983 17095 16989
rect 17037 16980 17049 16983
rect 15580 16952 17049 16980
rect 17037 16949 17049 16952
rect 17083 16949 17095 16983
rect 17144 16980 17172 17156
rect 17770 17144 17776 17196
rect 17828 17184 17834 17196
rect 19260 17193 19288 17224
rect 19610 17212 19616 17224
rect 19668 17212 19674 17264
rect 19978 17212 19984 17264
rect 20036 17212 20042 17264
rect 20824 17252 20852 17292
rect 20898 17280 20904 17332
rect 20956 17320 20962 17332
rect 20993 17323 21051 17329
rect 20993 17320 21005 17323
rect 20956 17292 21005 17320
rect 20956 17280 20962 17292
rect 20993 17289 21005 17292
rect 21039 17289 21051 17323
rect 20993 17283 21051 17289
rect 22646 17280 22652 17332
rect 22704 17320 22710 17332
rect 24949 17323 25007 17329
rect 24949 17320 24961 17323
rect 22704 17292 24961 17320
rect 22704 17280 22710 17292
rect 24949 17289 24961 17292
rect 24995 17289 25007 17323
rect 24949 17283 25007 17289
rect 25409 17323 25467 17329
rect 25409 17289 25421 17323
rect 25455 17320 25467 17323
rect 27341 17323 27399 17329
rect 27341 17320 27353 17323
rect 25455 17292 27353 17320
rect 25455 17289 25467 17292
rect 25409 17283 25467 17289
rect 27341 17289 27353 17292
rect 27387 17289 27399 17323
rect 27341 17283 27399 17289
rect 27430 17280 27436 17332
rect 27488 17320 27494 17332
rect 28902 17320 28908 17332
rect 27488 17292 28908 17320
rect 27488 17280 27494 17292
rect 28902 17280 28908 17292
rect 28960 17280 28966 17332
rect 29086 17280 29092 17332
rect 29144 17280 29150 17332
rect 29181 17323 29239 17329
rect 29181 17289 29193 17323
rect 29227 17320 29239 17323
rect 29454 17320 29460 17332
rect 29227 17292 29460 17320
rect 29227 17289 29239 17292
rect 29181 17283 29239 17289
rect 29454 17280 29460 17292
rect 29512 17280 29518 17332
rect 30193 17323 30251 17329
rect 30193 17289 30205 17323
rect 30239 17320 30251 17323
rect 32030 17320 32036 17332
rect 30239 17292 32036 17320
rect 30239 17289 30251 17292
rect 30193 17283 30251 17289
rect 32030 17280 32036 17292
rect 32088 17280 32094 17332
rect 33594 17320 33600 17332
rect 32324 17292 33600 17320
rect 23106 17252 23112 17264
rect 20824 17224 23112 17252
rect 23106 17212 23112 17224
rect 23164 17212 23170 17264
rect 23474 17212 23480 17264
rect 23532 17212 23538 17264
rect 24302 17212 24308 17264
rect 24360 17252 24366 17264
rect 24360 17224 25636 17252
rect 24360 17212 24366 17224
rect 17865 17187 17923 17193
rect 17865 17184 17877 17187
rect 17828 17156 17877 17184
rect 17828 17144 17834 17156
rect 17865 17153 17877 17156
rect 17911 17153 17923 17187
rect 17865 17147 17923 17153
rect 19245 17187 19303 17193
rect 19245 17153 19257 17187
rect 19291 17153 19303 17187
rect 19245 17147 19303 17153
rect 22738 17144 22744 17196
rect 22796 17144 22802 17196
rect 25314 17144 25320 17196
rect 25372 17144 25378 17196
rect 18690 17076 18696 17128
rect 18748 17076 18754 17128
rect 19521 17119 19579 17125
rect 19521 17085 19533 17119
rect 19567 17116 19579 17119
rect 20070 17116 20076 17128
rect 19567 17088 20076 17116
rect 19567 17085 19579 17088
rect 19521 17079 19579 17085
rect 20070 17076 20076 17088
rect 20128 17076 20134 17128
rect 24486 17076 24492 17128
rect 24544 17076 24550 17128
rect 25222 17076 25228 17128
rect 25280 17116 25286 17128
rect 25501 17119 25559 17125
rect 25501 17116 25513 17119
rect 25280 17088 25513 17116
rect 25280 17076 25286 17088
rect 25501 17085 25513 17088
rect 25547 17085 25559 17119
rect 25608 17116 25636 17224
rect 26142 17212 26148 17264
rect 26200 17252 26206 17264
rect 30285 17255 30343 17261
rect 30285 17252 30297 17255
rect 26200 17224 30297 17252
rect 26200 17212 26206 17224
rect 30285 17221 30297 17224
rect 30331 17221 30343 17255
rect 30285 17215 30343 17221
rect 30926 17212 30932 17264
rect 30984 17252 30990 17264
rect 32324 17252 32352 17292
rect 33594 17280 33600 17292
rect 33652 17280 33658 17332
rect 35066 17280 35072 17332
rect 35124 17320 35130 17332
rect 36357 17323 36415 17329
rect 36357 17320 36369 17323
rect 35124 17292 36369 17320
rect 35124 17280 35130 17292
rect 36357 17289 36369 17292
rect 36403 17289 36415 17323
rect 36357 17283 36415 17289
rect 36446 17280 36452 17332
rect 36504 17320 36510 17332
rect 37461 17323 37519 17329
rect 37461 17320 37473 17323
rect 36504 17292 37473 17320
rect 36504 17280 36510 17292
rect 37461 17289 37473 17292
rect 37507 17289 37519 17323
rect 37461 17283 37519 17289
rect 48406 17280 48412 17332
rect 48464 17280 48470 17332
rect 34422 17252 34428 17264
rect 30984 17224 32352 17252
rect 33810 17224 34428 17252
rect 30984 17212 30990 17224
rect 32324 17196 32352 17224
rect 34422 17212 34428 17224
rect 34480 17212 34486 17264
rect 34606 17212 34612 17264
rect 34664 17212 34670 17264
rect 37829 17255 37887 17261
rect 37829 17221 37841 17255
rect 37875 17252 37887 17255
rect 38378 17252 38384 17264
rect 37875 17224 38384 17252
rect 37875 17221 37887 17224
rect 37829 17215 37887 17221
rect 38378 17212 38384 17224
rect 38436 17212 38442 17264
rect 39206 17212 39212 17264
rect 39264 17212 39270 17264
rect 39666 17212 39672 17264
rect 39724 17212 39730 17264
rect 48222 17212 48228 17264
rect 48280 17252 48286 17264
rect 49145 17255 49203 17261
rect 49145 17252 49157 17255
rect 48280 17224 49157 17252
rect 48280 17212 48286 17224
rect 49145 17221 49157 17224
rect 49191 17221 49203 17255
rect 49145 17215 49203 17221
rect 26970 17144 26976 17196
rect 27028 17184 27034 17196
rect 27430 17184 27436 17196
rect 27028 17156 27436 17184
rect 27028 17144 27034 17156
rect 27430 17144 27436 17156
rect 27488 17144 27494 17196
rect 27706 17144 27712 17196
rect 27764 17144 27770 17196
rect 28537 17187 28595 17193
rect 28537 17184 28549 17187
rect 27816 17156 28549 17184
rect 27724 17116 27752 17144
rect 27816 17128 27844 17156
rect 28537 17153 28549 17156
rect 28583 17184 28595 17187
rect 28626 17184 28632 17196
rect 28583 17156 28632 17184
rect 28583 17153 28595 17156
rect 28537 17147 28595 17153
rect 28626 17144 28632 17156
rect 28684 17144 28690 17196
rect 29546 17144 29552 17196
rect 29604 17184 29610 17196
rect 31294 17184 31300 17196
rect 29604 17156 31300 17184
rect 29604 17144 29610 17156
rect 31294 17144 31300 17156
rect 31352 17144 31358 17196
rect 31389 17187 31447 17193
rect 31389 17153 31401 17187
rect 31435 17184 31447 17187
rect 31435 17156 31754 17184
rect 31435 17153 31447 17156
rect 31389 17147 31447 17153
rect 25608 17088 27752 17116
rect 25501 17079 25559 17085
rect 27798 17076 27804 17128
rect 27856 17076 27862 17128
rect 27982 17076 27988 17128
rect 28040 17076 28046 17128
rect 29273 17119 29331 17125
rect 29273 17085 29285 17119
rect 29319 17085 29331 17119
rect 29273 17079 29331 17085
rect 25774 17048 25780 17060
rect 24044 17020 25780 17048
rect 22002 16980 22008 16992
rect 17144 16952 22008 16980
rect 17037 16943 17095 16949
rect 22002 16940 22008 16952
rect 22060 16940 22066 16992
rect 22738 16940 22744 16992
rect 22796 16980 22802 16992
rect 23004 16983 23062 16989
rect 23004 16980 23016 16983
rect 22796 16952 23016 16980
rect 22796 16940 22802 16952
rect 23004 16949 23016 16952
rect 23050 16980 23062 16983
rect 23382 16980 23388 16992
rect 23050 16952 23388 16980
rect 23050 16949 23062 16952
rect 23004 16943 23062 16949
rect 23382 16940 23388 16952
rect 23440 16940 23446 16992
rect 23566 16940 23572 16992
rect 23624 16980 23630 16992
rect 24044 16980 24072 17020
rect 25774 17008 25780 17020
rect 25832 17008 25838 17060
rect 29086 17008 29092 17060
rect 29144 17048 29150 17060
rect 29288 17048 29316 17079
rect 29914 17076 29920 17128
rect 29972 17116 29978 17128
rect 30377 17119 30435 17125
rect 30377 17116 30389 17119
rect 29972 17088 30389 17116
rect 29972 17076 29978 17088
rect 30377 17085 30389 17088
rect 30423 17085 30435 17119
rect 30377 17079 30435 17085
rect 30558 17076 30564 17128
rect 30616 17116 30622 17128
rect 31481 17119 31539 17125
rect 31481 17116 31493 17119
rect 30616 17088 31493 17116
rect 30616 17076 30622 17088
rect 31481 17085 31493 17088
rect 31527 17085 31539 17119
rect 31481 17079 31539 17085
rect 31573 17119 31631 17125
rect 31573 17085 31585 17119
rect 31619 17085 31631 17119
rect 31573 17079 31631 17085
rect 29144 17020 29316 17048
rect 29144 17008 29150 17020
rect 30466 17008 30472 17060
rect 30524 17048 30530 17060
rect 31588 17048 31616 17079
rect 30524 17020 31616 17048
rect 30524 17008 30530 17020
rect 23624 16952 24072 16980
rect 23624 16940 23630 16952
rect 25590 16940 25596 16992
rect 25648 16980 25654 16992
rect 28350 16980 28356 16992
rect 25648 16952 28356 16980
rect 25648 16940 25654 16952
rect 28350 16940 28356 16952
rect 28408 16940 28414 16992
rect 28718 16940 28724 16992
rect 28776 16940 28782 16992
rect 29825 16983 29883 16989
rect 29825 16949 29837 16983
rect 29871 16980 29883 16983
rect 30926 16980 30932 16992
rect 29871 16952 30932 16980
rect 29871 16949 29883 16952
rect 29825 16943 29883 16949
rect 30926 16940 30932 16952
rect 30984 16940 30990 16992
rect 31018 16940 31024 16992
rect 31076 16940 31082 16992
rect 31726 16980 31754 17156
rect 32306 17144 32312 17196
rect 32364 17144 32370 17196
rect 37921 17187 37979 17193
rect 37921 17153 37933 17187
rect 37967 17184 37979 17187
rect 38838 17184 38844 17196
rect 37967 17156 38844 17184
rect 37967 17153 37979 17156
rect 37921 17147 37979 17153
rect 38838 17144 38844 17156
rect 38896 17144 38902 17196
rect 48590 17144 48596 17196
rect 48648 17144 48654 17196
rect 32214 17076 32220 17128
rect 32272 17116 32278 17128
rect 32585 17119 32643 17125
rect 32585 17116 32597 17119
rect 32272 17088 32597 17116
rect 32272 17076 32278 17088
rect 32585 17085 32597 17088
rect 32631 17085 32643 17119
rect 32585 17079 32643 17085
rect 32674 17076 32680 17128
rect 32732 17116 32738 17128
rect 34790 17116 34796 17128
rect 32732 17088 34796 17116
rect 32732 17076 32738 17088
rect 34790 17076 34796 17088
rect 34848 17076 34854 17128
rect 34882 17076 34888 17128
rect 34940 17116 34946 17128
rect 35345 17119 35403 17125
rect 35345 17116 35357 17119
rect 34940 17088 35357 17116
rect 34940 17076 34946 17088
rect 35345 17085 35357 17088
rect 35391 17085 35403 17119
rect 35345 17079 35403 17085
rect 36170 17076 36176 17128
rect 36228 17116 36234 17128
rect 36449 17119 36507 17125
rect 36449 17116 36461 17119
rect 36228 17088 36461 17116
rect 36228 17076 36234 17088
rect 36449 17085 36461 17088
rect 36495 17085 36507 17119
rect 36449 17079 36507 17085
rect 36633 17119 36691 17125
rect 36633 17085 36645 17119
rect 36679 17116 36691 17119
rect 37550 17116 37556 17128
rect 36679 17088 37556 17116
rect 36679 17085 36691 17088
rect 36633 17079 36691 17085
rect 37550 17076 37556 17088
rect 37608 17076 37614 17128
rect 37642 17076 37648 17128
rect 37700 17116 37706 17128
rect 38013 17119 38071 17125
rect 38013 17116 38025 17119
rect 37700 17088 38025 17116
rect 37700 17076 37706 17088
rect 38013 17085 38025 17088
rect 38059 17085 38071 17119
rect 38013 17079 38071 17085
rect 38933 17119 38991 17125
rect 38933 17085 38945 17119
rect 38979 17085 38991 17119
rect 38933 17079 38991 17085
rect 35989 17051 36047 17057
rect 35989 17017 36001 17051
rect 36035 17048 36047 17051
rect 36078 17048 36084 17060
rect 36035 17020 36084 17048
rect 36035 17017 36047 17020
rect 35989 17011 36047 17017
rect 36078 17008 36084 17020
rect 36136 17008 36142 17060
rect 37734 17008 37740 17060
rect 37792 17048 37798 17060
rect 38948 17048 38976 17079
rect 47394 17048 47400 17060
rect 37792 17020 38976 17048
rect 40236 17020 47400 17048
rect 37792 17008 37798 17020
rect 33870 16980 33876 16992
rect 31726 16952 33876 16980
rect 33870 16940 33876 16952
rect 33928 16940 33934 16992
rect 34054 16940 34060 16992
rect 34112 16940 34118 16992
rect 37550 16940 37556 16992
rect 37608 16980 37614 16992
rect 40236 16980 40264 17020
rect 47394 17008 47400 17020
rect 47452 17008 47458 17060
rect 37608 16952 40264 16980
rect 37608 16940 37614 16952
rect 40678 16940 40684 16992
rect 40736 16940 40742 16992
rect 49234 16940 49240 16992
rect 49292 16940 49298 16992
rect 1104 16890 49864 16912
rect 1104 16838 2950 16890
rect 3002 16838 3014 16890
rect 3066 16838 3078 16890
rect 3130 16838 3142 16890
rect 3194 16838 3206 16890
rect 3258 16838 12950 16890
rect 13002 16838 13014 16890
rect 13066 16838 13078 16890
rect 13130 16838 13142 16890
rect 13194 16838 13206 16890
rect 13258 16838 22950 16890
rect 23002 16838 23014 16890
rect 23066 16838 23078 16890
rect 23130 16838 23142 16890
rect 23194 16838 23206 16890
rect 23258 16838 32950 16890
rect 33002 16838 33014 16890
rect 33066 16838 33078 16890
rect 33130 16838 33142 16890
rect 33194 16838 33206 16890
rect 33258 16838 42950 16890
rect 43002 16838 43014 16890
rect 43066 16838 43078 16890
rect 43130 16838 43142 16890
rect 43194 16838 43206 16890
rect 43258 16838 49864 16890
rect 1104 16816 49864 16838
rect 10502 16736 10508 16788
rect 10560 16736 10566 16788
rect 11882 16736 11888 16788
rect 11940 16776 11946 16788
rect 16022 16776 16028 16788
rect 11940 16748 16028 16776
rect 11940 16736 11946 16748
rect 16022 16736 16028 16748
rect 16080 16736 16086 16788
rect 16114 16736 16120 16788
rect 16172 16776 16178 16788
rect 17218 16776 17224 16788
rect 16172 16748 17224 16776
rect 16172 16736 16178 16748
rect 17218 16736 17224 16748
rect 17276 16736 17282 16788
rect 17392 16779 17450 16785
rect 17392 16745 17404 16779
rect 17438 16776 17450 16779
rect 18506 16776 18512 16788
rect 17438 16748 18512 16776
rect 17438 16745 17450 16748
rect 17392 16739 17450 16745
rect 18506 16736 18512 16748
rect 18564 16776 18570 16788
rect 21910 16776 21916 16788
rect 18564 16748 21916 16776
rect 18564 16736 18570 16748
rect 21910 16736 21916 16748
rect 21968 16736 21974 16788
rect 22002 16736 22008 16788
rect 22060 16776 22066 16788
rect 22462 16776 22468 16788
rect 22060 16748 22468 16776
rect 22060 16736 22066 16748
rect 22462 16736 22468 16748
rect 22520 16736 22526 16788
rect 23658 16736 23664 16788
rect 23716 16776 23722 16788
rect 24765 16779 24823 16785
rect 24765 16776 24777 16779
rect 23716 16748 24777 16776
rect 23716 16736 23722 16748
rect 24765 16745 24777 16748
rect 24811 16745 24823 16779
rect 27338 16776 27344 16788
rect 24765 16739 24823 16745
rect 25332 16748 27344 16776
rect 10962 16668 10968 16720
rect 11020 16708 11026 16720
rect 12250 16708 12256 16720
rect 11020 16680 12256 16708
rect 11020 16668 11026 16680
rect 12250 16668 12256 16680
rect 12308 16668 12314 16720
rect 12526 16668 12532 16720
rect 12584 16708 12590 16720
rect 15657 16711 15715 16717
rect 12584 16680 14872 16708
rect 12584 16668 12590 16680
rect 4430 16600 4436 16652
rect 4488 16640 4494 16652
rect 5442 16640 5448 16652
rect 4488 16612 5448 16640
rect 4488 16600 4494 16612
rect 5442 16600 5448 16612
rect 5500 16640 5506 16652
rect 8205 16643 8263 16649
rect 8205 16640 8217 16643
rect 5500 16612 8217 16640
rect 5500 16600 5506 16612
rect 8205 16609 8217 16612
rect 8251 16609 8263 16643
rect 8205 16603 8263 16609
rect 8389 16643 8447 16649
rect 8389 16609 8401 16643
rect 8435 16640 8447 16643
rect 8570 16640 8576 16652
rect 8435 16612 8576 16640
rect 8435 16609 8447 16612
rect 8389 16603 8447 16609
rect 8570 16600 8576 16612
rect 8628 16600 8634 16652
rect 10870 16600 10876 16652
rect 10928 16640 10934 16652
rect 13464 16649 13492 16680
rect 14844 16652 14872 16680
rect 15657 16677 15669 16711
rect 15703 16677 15715 16711
rect 16942 16708 16948 16720
rect 15657 16671 15715 16677
rect 16132 16680 16948 16708
rect 11609 16643 11667 16649
rect 11609 16640 11621 16643
rect 10928 16612 11621 16640
rect 10928 16600 10934 16612
rect 11609 16609 11621 16612
rect 11655 16609 11667 16643
rect 11609 16603 11667 16609
rect 13449 16643 13507 16649
rect 13449 16609 13461 16643
rect 13495 16609 13507 16643
rect 13449 16603 13507 16609
rect 13633 16643 13691 16649
rect 13633 16609 13645 16643
rect 13679 16640 13691 16643
rect 13906 16640 13912 16652
rect 13679 16612 13912 16640
rect 13679 16609 13691 16612
rect 13633 16603 13691 16609
rect 13906 16600 13912 16612
rect 13964 16600 13970 16652
rect 14826 16600 14832 16652
rect 14884 16640 14890 16652
rect 14921 16643 14979 16649
rect 14921 16640 14933 16643
rect 14884 16612 14933 16640
rect 14884 16600 14890 16612
rect 14921 16609 14933 16612
rect 14967 16609 14979 16643
rect 14921 16603 14979 16609
rect 15102 16600 15108 16652
rect 15160 16600 15166 16652
rect 15672 16584 15700 16671
rect 15838 16600 15844 16652
rect 15896 16640 15902 16652
rect 16132 16649 16160 16680
rect 16942 16668 16948 16680
rect 17000 16668 17006 16720
rect 23934 16708 23940 16720
rect 23768 16680 23940 16708
rect 16117 16643 16175 16649
rect 16117 16640 16129 16643
rect 15896 16612 16129 16640
rect 15896 16600 15902 16612
rect 16117 16609 16129 16612
rect 16163 16609 16175 16643
rect 16117 16603 16175 16609
rect 16298 16600 16304 16652
rect 16356 16600 16362 16652
rect 17126 16600 17132 16652
rect 17184 16600 17190 16652
rect 18690 16600 18696 16652
rect 18748 16600 18754 16652
rect 19610 16600 19616 16652
rect 19668 16600 19674 16652
rect 20530 16600 20536 16652
rect 20588 16640 20594 16652
rect 20993 16643 21051 16649
rect 20993 16640 21005 16643
rect 20588 16612 21005 16640
rect 20588 16600 20594 16612
rect 20993 16609 21005 16612
rect 21039 16609 21051 16643
rect 20993 16603 21051 16609
rect 21269 16643 21327 16649
rect 21269 16609 21281 16643
rect 21315 16640 21327 16643
rect 22462 16640 22468 16652
rect 21315 16612 22468 16640
rect 21315 16609 21327 16612
rect 21269 16603 21327 16609
rect 22462 16600 22468 16612
rect 22520 16640 22526 16652
rect 23566 16640 23572 16652
rect 22520 16612 23572 16640
rect 22520 16600 22526 16612
rect 23566 16600 23572 16612
rect 23624 16600 23630 16652
rect 23768 16649 23796 16680
rect 23934 16668 23940 16680
rect 23992 16668 23998 16720
rect 23753 16643 23811 16649
rect 23753 16609 23765 16643
rect 23799 16609 23811 16643
rect 23753 16603 23811 16609
rect 23845 16643 23903 16649
rect 23845 16609 23857 16643
rect 23891 16640 23903 16643
rect 25332 16640 25360 16748
rect 27338 16736 27344 16748
rect 27396 16736 27402 16788
rect 27614 16736 27620 16788
rect 27672 16776 27678 16788
rect 27982 16776 27988 16788
rect 27672 16748 27988 16776
rect 27672 16736 27678 16748
rect 27982 16736 27988 16748
rect 28040 16736 28046 16788
rect 29270 16736 29276 16788
rect 29328 16776 29334 16788
rect 29328 16748 30972 16776
rect 29328 16736 29334 16748
rect 30650 16708 30656 16720
rect 26896 16680 30656 16708
rect 23891 16612 25360 16640
rect 23891 16609 23903 16612
rect 23845 16603 23903 16609
rect 25406 16600 25412 16652
rect 25464 16640 25470 16652
rect 25593 16643 25651 16649
rect 25593 16640 25605 16643
rect 25464 16612 25605 16640
rect 25464 16600 25470 16612
rect 25593 16609 25605 16612
rect 25639 16609 25651 16643
rect 25593 16603 25651 16609
rect 25866 16600 25872 16652
rect 25924 16600 25930 16652
rect 26234 16600 26240 16652
rect 26292 16640 26298 16652
rect 26896 16640 26924 16680
rect 30650 16668 30656 16680
rect 30708 16668 30714 16720
rect 30944 16708 30972 16748
rect 31018 16736 31024 16788
rect 31076 16776 31082 16788
rect 33962 16776 33968 16788
rect 31076 16748 33968 16776
rect 31076 16736 31082 16748
rect 33962 16736 33968 16748
rect 34020 16736 34026 16788
rect 34790 16736 34796 16788
rect 34848 16776 34854 16788
rect 49234 16776 49240 16788
rect 34848 16748 49240 16776
rect 34848 16736 34854 16748
rect 49234 16736 49240 16748
rect 49292 16736 49298 16788
rect 30944 16680 32444 16708
rect 26292 16612 26924 16640
rect 26292 16600 26298 16612
rect 30006 16600 30012 16652
rect 30064 16640 30070 16652
rect 30285 16643 30343 16649
rect 30285 16640 30297 16643
rect 30064 16612 30297 16640
rect 30064 16600 30070 16612
rect 30285 16609 30297 16612
rect 30331 16609 30343 16643
rect 30285 16603 30343 16609
rect 31386 16600 31392 16652
rect 31444 16600 31450 16652
rect 31570 16600 31576 16652
rect 31628 16600 31634 16652
rect 32306 16600 32312 16652
rect 32364 16600 32370 16652
rect 32416 16640 32444 16680
rect 35618 16668 35624 16720
rect 35676 16708 35682 16720
rect 35676 16680 36768 16708
rect 35676 16668 35682 16680
rect 32585 16643 32643 16649
rect 32585 16640 32597 16643
rect 32416 16612 32597 16640
rect 32585 16609 32597 16612
rect 32631 16640 32643 16643
rect 33318 16640 33324 16652
rect 32631 16612 33324 16640
rect 32631 16609 32643 16612
rect 32585 16603 32643 16609
rect 33318 16600 33324 16612
rect 33376 16640 33382 16652
rect 34054 16640 34060 16652
rect 33376 16612 34060 16640
rect 33376 16600 33382 16612
rect 34054 16600 34060 16612
rect 34112 16600 34118 16652
rect 35710 16600 35716 16652
rect 35768 16600 35774 16652
rect 36740 16649 36768 16680
rect 36725 16643 36783 16649
rect 36725 16609 36737 16643
rect 36771 16609 36783 16643
rect 36725 16603 36783 16609
rect 36814 16600 36820 16652
rect 36872 16600 36878 16652
rect 37182 16600 37188 16652
rect 37240 16640 37246 16652
rect 38013 16643 38071 16649
rect 38013 16640 38025 16643
rect 37240 16612 38025 16640
rect 37240 16600 37246 16612
rect 38013 16609 38025 16612
rect 38059 16640 38071 16643
rect 40678 16640 40684 16652
rect 38059 16612 40684 16640
rect 38059 16609 38071 16612
rect 38013 16603 38071 16609
rect 40678 16600 40684 16612
rect 40736 16600 40742 16652
rect 1765 16575 1823 16581
rect 1765 16541 1777 16575
rect 1811 16572 1823 16575
rect 6822 16572 6828 16584
rect 1811 16544 6828 16572
rect 1811 16541 1823 16544
rect 1765 16535 1823 16541
rect 6822 16532 6828 16544
rect 6880 16532 6886 16584
rect 7558 16532 7564 16584
rect 7616 16572 7622 16584
rect 8113 16575 8171 16581
rect 8113 16572 8125 16575
rect 7616 16544 8125 16572
rect 7616 16532 7622 16544
rect 8113 16541 8125 16544
rect 8159 16541 8171 16575
rect 8113 16535 8171 16541
rect 11054 16532 11060 16584
rect 11112 16572 11118 16584
rect 12434 16572 12440 16584
rect 11112 16544 12440 16572
rect 11112 16532 11118 16544
rect 12434 16532 12440 16544
rect 12492 16532 12498 16584
rect 12529 16575 12587 16581
rect 12529 16541 12541 16575
rect 12575 16572 12587 16575
rect 12575 16544 15424 16572
rect 12575 16541 12587 16544
rect 12529 16535 12587 16541
rect 1302 16464 1308 16516
rect 1360 16504 1366 16516
rect 2501 16507 2559 16513
rect 2501 16504 2513 16507
rect 1360 16476 2513 16504
rect 1360 16464 1366 16476
rect 2501 16473 2513 16476
rect 2547 16473 2559 16507
rect 9582 16504 9588 16516
rect 2501 16467 2559 16473
rect 7760 16476 9588 16504
rect 7760 16445 7788 16476
rect 9582 16464 9588 16476
rect 9640 16464 9646 16516
rect 10413 16507 10471 16513
rect 10413 16473 10425 16507
rect 10459 16504 10471 16507
rect 11330 16504 11336 16516
rect 10459 16476 11336 16504
rect 10459 16473 10471 16476
rect 10413 16467 10471 16473
rect 11330 16464 11336 16476
rect 11388 16464 11394 16516
rect 11425 16507 11483 16513
rect 11425 16473 11437 16507
rect 11471 16504 11483 16507
rect 12618 16504 12624 16516
rect 11471 16476 12624 16504
rect 11471 16473 11483 16476
rect 11425 16467 11483 16473
rect 12618 16464 12624 16476
rect 12676 16464 12682 16516
rect 13357 16507 13415 16513
rect 13357 16473 13369 16507
rect 13403 16504 13415 16507
rect 13538 16504 13544 16516
rect 13403 16476 13544 16504
rect 13403 16473 13415 16476
rect 13357 16467 13415 16473
rect 13538 16464 13544 16476
rect 13596 16504 13602 16516
rect 15396 16504 15424 16544
rect 15654 16532 15660 16584
rect 15712 16532 15718 16584
rect 16022 16532 16028 16584
rect 16080 16532 16086 16584
rect 16132 16544 16436 16572
rect 16132 16504 16160 16544
rect 13596 16476 14872 16504
rect 15396 16476 16160 16504
rect 13596 16464 13602 16476
rect 7745 16439 7803 16445
rect 7745 16405 7757 16439
rect 7791 16405 7803 16439
rect 7745 16399 7803 16405
rect 11054 16396 11060 16448
rect 11112 16396 11118 16448
rect 11514 16396 11520 16448
rect 11572 16396 11578 16448
rect 12066 16396 12072 16448
rect 12124 16436 12130 16448
rect 12345 16439 12403 16445
rect 12345 16436 12357 16439
rect 12124 16408 12357 16436
rect 12124 16396 12130 16408
rect 12345 16405 12357 16408
rect 12391 16405 12403 16439
rect 12345 16399 12403 16405
rect 12989 16439 13047 16445
rect 12989 16405 13001 16439
rect 13035 16436 13047 16439
rect 13262 16436 13268 16448
rect 13035 16408 13268 16436
rect 13035 16405 13047 16408
rect 12989 16399 13047 16405
rect 13262 16396 13268 16408
rect 13320 16396 13326 16448
rect 14458 16396 14464 16448
rect 14516 16396 14522 16448
rect 14844 16445 14872 16476
rect 14829 16439 14887 16445
rect 14829 16405 14841 16439
rect 14875 16436 14887 16439
rect 16114 16436 16120 16448
rect 14875 16408 16120 16436
rect 14875 16405 14887 16408
rect 14829 16399 14887 16405
rect 16114 16396 16120 16408
rect 16172 16396 16178 16448
rect 16408 16436 16436 16544
rect 17678 16464 17684 16516
rect 17736 16504 17742 16516
rect 17736 16476 17894 16504
rect 17736 16464 17742 16476
rect 18708 16448 18736 16600
rect 20254 16532 20260 16584
rect 20312 16532 20318 16584
rect 25498 16572 25504 16584
rect 23308 16544 25504 16572
rect 20714 16504 20720 16516
rect 18800 16476 20720 16504
rect 18800 16448 18828 16476
rect 20714 16464 20720 16476
rect 20772 16464 20778 16516
rect 20990 16464 20996 16516
rect 21048 16504 21054 16516
rect 23308 16504 23336 16544
rect 25498 16532 25504 16544
rect 25556 16532 25562 16584
rect 30760 16544 32352 16572
rect 21048 16476 21758 16504
rect 22756 16476 23336 16504
rect 23661 16507 23719 16513
rect 21048 16464 21054 16476
rect 18322 16436 18328 16448
rect 16408 16408 18328 16436
rect 18322 16396 18328 16408
rect 18380 16396 18386 16448
rect 18690 16396 18696 16448
rect 18748 16396 18754 16448
rect 18782 16396 18788 16448
rect 18840 16396 18846 16448
rect 18874 16396 18880 16448
rect 18932 16396 18938 16448
rect 19794 16396 19800 16448
rect 19852 16436 19858 16448
rect 20073 16439 20131 16445
rect 20073 16436 20085 16439
rect 19852 16408 20085 16436
rect 19852 16396 19858 16408
rect 20073 16405 20085 16408
rect 20119 16405 20131 16439
rect 20073 16399 20131 16405
rect 20162 16396 20168 16448
rect 20220 16436 20226 16448
rect 22756 16445 22784 16476
rect 23661 16473 23673 16507
rect 23707 16504 23719 16507
rect 25130 16504 25136 16516
rect 23707 16476 25136 16504
rect 23707 16473 23719 16476
rect 23661 16467 23719 16473
rect 25130 16464 25136 16476
rect 25188 16464 25194 16516
rect 26602 16464 26608 16516
rect 26660 16464 26666 16516
rect 29178 16464 29184 16516
rect 29236 16504 29242 16516
rect 30101 16507 30159 16513
rect 30101 16504 30113 16507
rect 29236 16476 30113 16504
rect 29236 16464 29242 16476
rect 30101 16473 30113 16476
rect 30147 16473 30159 16507
rect 30101 16467 30159 16473
rect 30190 16464 30196 16516
rect 30248 16464 30254 16516
rect 22741 16439 22799 16445
rect 22741 16436 22753 16439
rect 20220 16408 22753 16436
rect 20220 16396 20226 16408
rect 22741 16405 22753 16408
rect 22787 16405 22799 16439
rect 22741 16399 22799 16405
rect 22830 16396 22836 16448
rect 22888 16436 22894 16448
rect 23293 16439 23351 16445
rect 23293 16436 23305 16439
rect 22888 16408 23305 16436
rect 22888 16396 22894 16408
rect 23293 16405 23305 16408
rect 23339 16405 23351 16439
rect 23293 16399 23351 16405
rect 23382 16396 23388 16448
rect 23440 16436 23446 16448
rect 25958 16436 25964 16448
rect 23440 16408 25964 16436
rect 23440 16396 23446 16408
rect 25958 16396 25964 16408
rect 26016 16396 26022 16448
rect 29733 16439 29791 16445
rect 29733 16405 29745 16439
rect 29779 16436 29791 16439
rect 30760 16436 30788 16544
rect 31846 16504 31852 16516
rect 30944 16476 31852 16504
rect 30944 16445 30972 16476
rect 31846 16464 31852 16476
rect 31904 16464 31910 16516
rect 29779 16408 30788 16436
rect 30929 16439 30987 16445
rect 29779 16405 29791 16408
rect 29733 16399 29791 16405
rect 30929 16405 30941 16439
rect 30975 16405 30987 16439
rect 30929 16399 30987 16405
rect 31294 16396 31300 16448
rect 31352 16396 31358 16448
rect 32324 16436 32352 16544
rect 34606 16532 34612 16584
rect 34664 16572 34670 16584
rect 34885 16575 34943 16581
rect 34885 16572 34897 16575
rect 34664 16544 34897 16572
rect 34664 16532 34670 16544
rect 34885 16541 34897 16544
rect 34931 16541 34943 16575
rect 34885 16535 34943 16541
rect 35986 16532 35992 16584
rect 36044 16572 36050 16584
rect 36633 16575 36691 16581
rect 36633 16572 36645 16575
rect 36044 16544 36645 16572
rect 36044 16532 36050 16544
rect 36633 16541 36645 16544
rect 36679 16541 36691 16575
rect 36633 16535 36691 16541
rect 37734 16532 37740 16584
rect 37792 16532 37798 16584
rect 49053 16575 49111 16581
rect 49053 16541 49065 16575
rect 49099 16572 49111 16575
rect 49142 16572 49148 16584
rect 49099 16544 49148 16572
rect 49099 16541 49111 16544
rect 49053 16535 49111 16541
rect 49142 16532 49148 16544
rect 49200 16532 49206 16584
rect 34422 16504 34428 16516
rect 33810 16476 34428 16504
rect 34422 16464 34428 16476
rect 34480 16464 34486 16516
rect 39574 16504 39580 16516
rect 39238 16476 39580 16504
rect 39574 16464 39580 16476
rect 39632 16464 39638 16516
rect 33594 16436 33600 16448
rect 32324 16408 33600 16436
rect 33594 16396 33600 16408
rect 33652 16396 33658 16448
rect 34054 16396 34060 16448
rect 34112 16396 34118 16448
rect 36262 16396 36268 16448
rect 36320 16396 36326 16448
rect 37826 16396 37832 16448
rect 37884 16436 37890 16448
rect 39485 16439 39543 16445
rect 39485 16436 39497 16439
rect 37884 16408 39497 16436
rect 37884 16396 37890 16408
rect 39485 16405 39497 16408
rect 39531 16405 39543 16439
rect 39485 16399 39543 16405
rect 49234 16396 49240 16448
rect 49292 16396 49298 16448
rect 1104 16346 49864 16368
rect 1104 16294 7950 16346
rect 8002 16294 8014 16346
rect 8066 16294 8078 16346
rect 8130 16294 8142 16346
rect 8194 16294 8206 16346
rect 8258 16294 17950 16346
rect 18002 16294 18014 16346
rect 18066 16294 18078 16346
rect 18130 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 27950 16346
rect 28002 16294 28014 16346
rect 28066 16294 28078 16346
rect 28130 16294 28142 16346
rect 28194 16294 28206 16346
rect 28258 16294 37950 16346
rect 38002 16294 38014 16346
rect 38066 16294 38078 16346
rect 38130 16294 38142 16346
rect 38194 16294 38206 16346
rect 38258 16294 47950 16346
rect 48002 16294 48014 16346
rect 48066 16294 48078 16346
rect 48130 16294 48142 16346
rect 48194 16294 48206 16346
rect 48258 16294 49864 16346
rect 1104 16272 49864 16294
rect 6362 16192 6368 16244
rect 6420 16232 6426 16244
rect 8297 16235 8355 16241
rect 8297 16232 8309 16235
rect 6420 16204 8309 16232
rect 6420 16192 6426 16204
rect 8297 16201 8309 16204
rect 8343 16201 8355 16235
rect 8297 16195 8355 16201
rect 1762 16056 1768 16108
rect 1820 16056 1826 16108
rect 8312 16096 8340 16195
rect 9306 16192 9312 16244
rect 9364 16192 9370 16244
rect 11057 16235 11115 16241
rect 11057 16201 11069 16235
rect 11103 16232 11115 16235
rect 11146 16232 11152 16244
rect 11103 16204 11152 16232
rect 11103 16201 11115 16204
rect 11057 16195 11115 16201
rect 11146 16192 11152 16204
rect 11204 16192 11210 16244
rect 11514 16192 11520 16244
rect 11572 16232 11578 16244
rect 11793 16235 11851 16241
rect 11793 16232 11805 16235
rect 11572 16204 11805 16232
rect 11572 16192 11578 16204
rect 11793 16201 11805 16204
rect 11839 16201 11851 16235
rect 11793 16195 11851 16201
rect 12989 16235 13047 16241
rect 12989 16201 13001 16235
rect 13035 16232 13047 16235
rect 13354 16232 13360 16244
rect 13035 16204 13360 16232
rect 13035 16201 13047 16204
rect 12989 16195 13047 16201
rect 13354 16192 13360 16204
rect 13412 16192 13418 16244
rect 15378 16192 15384 16244
rect 15436 16232 15442 16244
rect 15933 16235 15991 16241
rect 15933 16232 15945 16235
rect 15436 16204 15945 16232
rect 15436 16192 15442 16204
rect 15933 16201 15945 16204
rect 15979 16201 15991 16235
rect 15933 16195 15991 16201
rect 16025 16235 16083 16241
rect 16025 16201 16037 16235
rect 16071 16232 16083 16235
rect 16071 16204 16436 16232
rect 16071 16201 16083 16204
rect 16025 16195 16083 16201
rect 9217 16167 9275 16173
rect 9217 16133 9229 16167
rect 9263 16164 9275 16167
rect 12342 16164 12348 16176
rect 9263 16136 12348 16164
rect 9263 16133 9275 16136
rect 9217 16127 9275 16133
rect 12342 16124 12348 16136
rect 12400 16124 12406 16176
rect 12710 16124 12716 16176
rect 12768 16164 12774 16176
rect 13081 16167 13139 16173
rect 13081 16164 13093 16167
rect 12768 16136 13093 16164
rect 12768 16124 12774 16136
rect 13081 16133 13093 16136
rect 13127 16133 13139 16167
rect 13081 16127 13139 16133
rect 14366 16124 14372 16176
rect 14424 16164 14430 16176
rect 14737 16167 14795 16173
rect 14737 16164 14749 16167
rect 14424 16136 14749 16164
rect 14424 16124 14430 16136
rect 14737 16133 14749 16136
rect 14783 16164 14795 16167
rect 15286 16164 15292 16176
rect 14783 16136 15292 16164
rect 14783 16133 14795 16136
rect 14737 16127 14795 16133
rect 15286 16124 15292 16136
rect 15344 16124 15350 16176
rect 16408 16164 16436 16204
rect 16482 16192 16488 16244
rect 16540 16232 16546 16244
rect 19794 16232 19800 16244
rect 16540 16204 19800 16232
rect 16540 16192 16546 16204
rect 19794 16192 19800 16204
rect 19852 16192 19858 16244
rect 20254 16192 20260 16244
rect 20312 16232 20318 16244
rect 23017 16235 23075 16241
rect 23017 16232 23029 16235
rect 20312 16204 23029 16232
rect 20312 16192 20318 16204
rect 23017 16201 23029 16204
rect 23063 16201 23075 16235
rect 25406 16232 25412 16244
rect 23017 16195 23075 16201
rect 24136 16204 25412 16232
rect 16850 16164 16856 16176
rect 16408 16136 16856 16164
rect 16850 16124 16856 16136
rect 16908 16124 16914 16176
rect 17773 16167 17831 16173
rect 17773 16133 17785 16167
rect 17819 16164 17831 16167
rect 17862 16164 17868 16176
rect 17819 16136 17868 16164
rect 17819 16133 17831 16136
rect 17773 16127 17831 16133
rect 17862 16124 17868 16136
rect 17920 16124 17926 16176
rect 18782 16164 18788 16176
rect 17972 16136 18788 16164
rect 10965 16099 11023 16105
rect 8312 16068 10916 16096
rect 1302 15988 1308 16040
rect 1360 16028 1366 16040
rect 2041 16031 2099 16037
rect 2041 16028 2053 16031
rect 1360 16000 2053 16028
rect 1360 15988 1366 16000
rect 2041 15997 2053 16000
rect 2087 15997 2099 16031
rect 2041 15991 2099 15997
rect 4154 15988 4160 16040
rect 4212 16028 4218 16040
rect 8389 16031 8447 16037
rect 8389 16028 8401 16031
rect 4212 16000 8401 16028
rect 4212 15988 4218 16000
rect 8389 15997 8401 16000
rect 8435 15997 8447 16031
rect 8389 15991 8447 15997
rect 8570 15988 8576 16040
rect 8628 15988 8634 16040
rect 10888 16028 10916 16068
rect 10965 16065 10977 16099
rect 11011 16096 11023 16099
rect 11698 16096 11704 16108
rect 11011 16068 11704 16096
rect 11011 16065 11023 16068
rect 10965 16059 11023 16065
rect 11698 16056 11704 16068
rect 11756 16056 11762 16108
rect 12161 16099 12219 16105
rect 12161 16065 12173 16099
rect 12207 16096 12219 16099
rect 13722 16096 13728 16108
rect 12207 16068 13728 16096
rect 12207 16065 12219 16068
rect 12161 16059 12219 16065
rect 13722 16056 13728 16068
rect 13780 16056 13786 16108
rect 13998 16056 14004 16108
rect 14056 16096 14062 16108
rect 16298 16096 16304 16108
rect 14056 16068 16304 16096
rect 14056 16056 14062 16068
rect 12066 16028 12072 16040
rect 10888 16000 12072 16028
rect 12066 15988 12072 16000
rect 12124 15988 12130 16040
rect 12250 15988 12256 16040
rect 12308 15988 12314 16040
rect 12434 15988 12440 16040
rect 12492 15988 12498 16040
rect 12802 15988 12808 16040
rect 12860 16028 12866 16040
rect 13173 16031 13231 16037
rect 13173 16028 13185 16031
rect 12860 16000 13185 16028
rect 12860 15988 12866 16000
rect 13173 15997 13185 16000
rect 13219 15997 13231 16031
rect 13173 15991 13231 15997
rect 13909 16031 13967 16037
rect 13909 15997 13921 16031
rect 13955 16028 13967 16031
rect 14090 16028 14096 16040
rect 13955 16000 14096 16028
rect 13955 15997 13967 16000
rect 13909 15991 13967 15997
rect 14090 15988 14096 16000
rect 14148 16028 14154 16040
rect 14826 16028 14832 16040
rect 14148 16000 14832 16028
rect 14148 15988 14154 16000
rect 14826 15988 14832 16000
rect 14884 15988 14890 16040
rect 14936 16037 14964 16068
rect 16298 16056 16304 16068
rect 16356 16056 16362 16108
rect 14921 16031 14979 16037
rect 14921 15997 14933 16031
rect 14967 15997 14979 16031
rect 14921 15991 14979 15997
rect 15102 15988 15108 16040
rect 15160 16028 15166 16040
rect 16114 16028 16120 16040
rect 15160 16000 16120 16028
rect 15160 15988 15166 16000
rect 16114 15988 16120 16000
rect 16172 15988 16178 16040
rect 17865 16031 17923 16037
rect 17865 15997 17877 16031
rect 17911 16028 17923 16031
rect 17972 16028 18000 16136
rect 18782 16124 18788 16136
rect 18840 16124 18846 16176
rect 18874 16124 18880 16176
rect 18932 16164 18938 16176
rect 19429 16167 19487 16173
rect 19429 16164 19441 16167
rect 18932 16136 19441 16164
rect 18932 16124 18938 16136
rect 19429 16133 19441 16136
rect 19475 16133 19487 16167
rect 19429 16127 19487 16133
rect 19886 16124 19892 16176
rect 19944 16124 19950 16176
rect 18892 16096 18920 16124
rect 18064 16068 18920 16096
rect 18064 16037 18092 16068
rect 23382 16056 23388 16108
rect 23440 16056 23446 16108
rect 24136 16105 24164 16204
rect 25406 16192 25412 16204
rect 25464 16192 25470 16244
rect 25869 16235 25927 16241
rect 25869 16201 25881 16235
rect 25915 16232 25927 16235
rect 25958 16232 25964 16244
rect 25915 16204 25964 16232
rect 25915 16201 25927 16204
rect 25869 16195 25927 16201
rect 25958 16192 25964 16204
rect 26016 16192 26022 16244
rect 26326 16192 26332 16244
rect 26384 16232 26390 16244
rect 27154 16232 27160 16244
rect 26384 16204 27160 16232
rect 26384 16192 26390 16204
rect 27154 16192 27160 16204
rect 27212 16232 27218 16244
rect 27617 16235 27675 16241
rect 27617 16232 27629 16235
rect 27212 16204 27629 16232
rect 27212 16192 27218 16204
rect 27617 16201 27629 16204
rect 27663 16201 27675 16235
rect 27617 16195 27675 16201
rect 30285 16235 30343 16241
rect 30285 16201 30297 16235
rect 30331 16232 30343 16235
rect 30466 16232 30472 16244
rect 30331 16204 30472 16232
rect 30331 16201 30343 16204
rect 30285 16195 30343 16201
rect 30466 16192 30472 16204
rect 30524 16192 30530 16244
rect 30926 16192 30932 16244
rect 30984 16232 30990 16244
rect 31021 16235 31079 16241
rect 31021 16232 31033 16235
rect 30984 16204 31033 16232
rect 30984 16192 30990 16204
rect 31021 16201 31033 16204
rect 31067 16201 31079 16235
rect 31021 16195 31079 16201
rect 31110 16192 31116 16244
rect 31168 16192 31174 16244
rect 31754 16192 31760 16244
rect 31812 16232 31818 16244
rect 32398 16232 32404 16244
rect 31812 16204 32404 16232
rect 31812 16192 31818 16204
rect 32398 16192 32404 16204
rect 32456 16192 32462 16244
rect 32766 16192 32772 16244
rect 32824 16192 32830 16244
rect 33962 16192 33968 16244
rect 34020 16192 34026 16244
rect 37550 16232 37556 16244
rect 35728 16204 37556 16232
rect 24397 16167 24455 16173
rect 24397 16133 24409 16167
rect 24443 16164 24455 16167
rect 24486 16164 24492 16176
rect 24443 16136 24492 16164
rect 24443 16133 24455 16136
rect 24397 16127 24455 16133
rect 24486 16124 24492 16136
rect 24544 16124 24550 16176
rect 25774 16164 25780 16176
rect 25622 16136 25780 16164
rect 25774 16124 25780 16136
rect 25832 16164 25838 16176
rect 26602 16164 26608 16176
rect 25832 16136 26608 16164
rect 25832 16124 25838 16136
rect 26602 16124 26608 16136
rect 26660 16124 26666 16176
rect 28810 16124 28816 16176
rect 28868 16124 28874 16176
rect 30650 16164 30656 16176
rect 30038 16136 30656 16164
rect 30650 16124 30656 16136
rect 30708 16124 30714 16176
rect 35728 16164 35756 16204
rect 37550 16192 37556 16204
rect 37608 16192 37614 16244
rect 38838 16192 38844 16244
rect 38896 16232 38902 16244
rect 40497 16235 40555 16241
rect 40497 16232 40509 16235
rect 38896 16204 40509 16232
rect 38896 16192 38902 16204
rect 40497 16201 40509 16204
rect 40543 16201 40555 16235
rect 40497 16195 40555 16201
rect 40954 16192 40960 16244
rect 41012 16192 41018 16244
rect 30760 16136 35756 16164
rect 24121 16099 24179 16105
rect 24121 16065 24133 16099
rect 24167 16065 24179 16099
rect 24121 16059 24179 16065
rect 26142 16056 26148 16108
rect 26200 16096 26206 16108
rect 27525 16099 27583 16105
rect 27525 16096 27537 16099
rect 26200 16068 27537 16096
rect 26200 16056 26206 16068
rect 27525 16065 27537 16068
rect 27571 16096 27583 16099
rect 28353 16099 28411 16105
rect 28353 16096 28365 16099
rect 27571 16068 28365 16096
rect 27571 16065 27583 16068
rect 27525 16059 27583 16065
rect 28353 16065 28365 16068
rect 28399 16065 28411 16099
rect 28353 16059 28411 16065
rect 17911 16000 18000 16028
rect 18049 16031 18107 16037
rect 17911 15997 17923 16000
rect 17865 15991 17923 15997
rect 18049 15997 18061 16031
rect 18095 15997 18107 16031
rect 18049 15991 18107 15997
rect 18690 15988 18696 16040
rect 18748 16028 18754 16040
rect 19153 16031 19211 16037
rect 19153 16028 19165 16031
rect 18748 16000 19165 16028
rect 18748 15988 18754 16000
rect 19153 15997 19165 16000
rect 19199 16028 19211 16031
rect 20714 16028 20720 16040
rect 19199 16000 20720 16028
rect 19199 15997 19211 16000
rect 19153 15991 19211 15997
rect 20714 15988 20720 16000
rect 20772 15988 20778 16040
rect 23474 15988 23480 16040
rect 23532 15988 23538 16040
rect 23661 16031 23719 16037
rect 23661 15997 23673 16031
rect 23707 16028 23719 16031
rect 25038 16028 25044 16040
rect 23707 16000 25044 16028
rect 23707 15997 23719 16000
rect 23661 15991 23719 15997
rect 25038 15988 25044 16000
rect 25096 15988 25102 16040
rect 27709 16031 27767 16037
rect 27709 15997 27721 16031
rect 27755 15997 27767 16031
rect 28368 16028 28396 16059
rect 28534 16056 28540 16108
rect 28592 16056 28598 16108
rect 30760 16028 30788 16136
rect 37826 16124 37832 16176
rect 37884 16164 37890 16176
rect 38473 16167 38531 16173
rect 38473 16164 38485 16167
rect 37884 16136 38485 16164
rect 37884 16124 37890 16136
rect 38473 16133 38485 16136
rect 38519 16133 38531 16167
rect 38473 16127 38531 16133
rect 32677 16099 32735 16105
rect 32677 16065 32689 16099
rect 32723 16096 32735 16099
rect 32723 16068 33272 16096
rect 32723 16065 32735 16068
rect 32677 16059 32735 16065
rect 28368 16000 30788 16028
rect 27709 15991 27767 15997
rect 9490 15920 9496 15972
rect 9548 15960 9554 15972
rect 11882 15960 11888 15972
rect 9548 15932 11888 15960
rect 9548 15920 9554 15932
rect 11882 15920 11888 15932
rect 11940 15920 11946 15972
rect 14458 15920 14464 15972
rect 14516 15960 14522 15972
rect 15378 15960 15384 15972
rect 14516 15932 15384 15960
rect 14516 15920 14522 15932
rect 15378 15920 15384 15932
rect 15436 15920 15442 15972
rect 15565 15963 15623 15969
rect 15565 15929 15577 15963
rect 15611 15960 15623 15963
rect 17586 15960 17592 15972
rect 15611 15932 17592 15960
rect 15611 15929 15623 15932
rect 15565 15923 15623 15929
rect 17586 15920 17592 15932
rect 17644 15920 17650 15972
rect 25424 15932 26464 15960
rect 7929 15895 7987 15901
rect 7929 15861 7941 15895
rect 7975 15892 7987 15895
rect 9214 15892 9220 15904
rect 7975 15864 9220 15892
rect 7975 15861 7987 15864
rect 7929 15855 7987 15861
rect 9214 15852 9220 15864
rect 9272 15852 9278 15904
rect 12621 15895 12679 15901
rect 12621 15861 12633 15895
rect 12667 15892 12679 15895
rect 12710 15892 12716 15904
rect 12667 15864 12716 15892
rect 12667 15861 12679 15864
rect 12621 15855 12679 15861
rect 12710 15852 12716 15864
rect 12768 15852 12774 15904
rect 14366 15852 14372 15904
rect 14424 15852 14430 15904
rect 14734 15852 14740 15904
rect 14792 15892 14798 15904
rect 17405 15895 17463 15901
rect 17405 15892 17417 15895
rect 14792 15864 17417 15892
rect 14792 15852 14798 15864
rect 17405 15861 17417 15864
rect 17451 15861 17463 15895
rect 17405 15855 17463 15861
rect 17678 15852 17684 15904
rect 17736 15892 17742 15904
rect 19886 15892 19892 15904
rect 17736 15864 19892 15892
rect 17736 15852 17742 15864
rect 19886 15852 19892 15864
rect 19944 15852 19950 15904
rect 20898 15852 20904 15904
rect 20956 15852 20962 15904
rect 23842 15852 23848 15904
rect 23900 15892 23906 15904
rect 25424 15892 25452 15932
rect 23900 15864 25452 15892
rect 26436 15892 26464 15932
rect 26786 15920 26792 15972
rect 26844 15960 26850 15972
rect 27724 15960 27752 15991
rect 31202 15988 31208 16040
rect 31260 15988 31266 16040
rect 31938 15988 31944 16040
rect 31996 16028 32002 16040
rect 32858 16028 32864 16040
rect 31996 16000 32864 16028
rect 31996 15988 32002 16000
rect 32858 15988 32864 16000
rect 32916 15988 32922 16040
rect 33244 16028 33272 16068
rect 33318 16056 33324 16108
rect 33376 16096 33382 16108
rect 33873 16099 33931 16105
rect 33873 16096 33885 16099
rect 33376 16068 33885 16096
rect 33376 16056 33382 16068
rect 33873 16065 33885 16068
rect 33919 16065 33931 16099
rect 33873 16059 33931 16065
rect 36446 16056 36452 16108
rect 36504 16056 36510 16108
rect 39574 16056 39580 16108
rect 39632 16056 39638 16108
rect 40865 16099 40923 16105
rect 40865 16065 40877 16099
rect 40911 16096 40923 16099
rect 48958 16096 48964 16108
rect 40911 16068 48964 16096
rect 40911 16065 40923 16068
rect 40865 16059 40923 16065
rect 48958 16056 48964 16068
rect 49016 16056 49022 16108
rect 49050 16056 49056 16108
rect 49108 16056 49114 16108
rect 33778 16028 33784 16040
rect 33244 16000 33784 16028
rect 33778 15988 33784 16000
rect 33836 15988 33842 16040
rect 34057 16031 34115 16037
rect 34057 15997 34069 16031
rect 34103 15997 34115 16031
rect 34057 15991 34115 15997
rect 26844 15932 27752 15960
rect 26844 15920 26850 15932
rect 29914 15920 29920 15972
rect 29972 15960 29978 15972
rect 30190 15960 30196 15972
rect 29972 15932 30196 15960
rect 29972 15920 29978 15932
rect 30190 15920 30196 15932
rect 30248 15920 30254 15972
rect 32214 15920 32220 15972
rect 32272 15960 32278 15972
rect 34072 15960 34100 15991
rect 34882 15988 34888 16040
rect 34940 16028 34946 16040
rect 35069 16031 35127 16037
rect 35069 16028 35081 16031
rect 34940 16000 35081 16028
rect 34940 15988 34946 16000
rect 35069 15997 35081 16000
rect 35115 15997 35127 16031
rect 35069 15991 35127 15997
rect 35345 16031 35403 16037
rect 35345 15997 35357 16031
rect 35391 16028 35403 16031
rect 37366 16028 37372 16040
rect 35391 16000 37372 16028
rect 35391 15997 35403 16000
rect 35345 15991 35403 15997
rect 37366 15988 37372 16000
rect 37424 15988 37430 16040
rect 37734 15988 37740 16040
rect 37792 16028 37798 16040
rect 38197 16031 38255 16037
rect 38197 16028 38209 16031
rect 37792 16000 38209 16028
rect 37792 15988 37798 16000
rect 38197 15997 38209 16000
rect 38243 15997 38255 16031
rect 41049 16031 41107 16037
rect 41049 16028 41061 16031
rect 38197 15991 38255 15997
rect 38304 16000 41061 16028
rect 32272 15932 34100 15960
rect 36817 15963 36875 15969
rect 32272 15920 32278 15932
rect 36817 15929 36829 15963
rect 36863 15960 36875 15963
rect 36906 15960 36912 15972
rect 36863 15932 36912 15960
rect 36863 15929 36875 15932
rect 36817 15923 36875 15929
rect 27157 15895 27215 15901
rect 27157 15892 27169 15895
rect 26436 15864 27169 15892
rect 23900 15852 23906 15864
rect 27157 15861 27169 15864
rect 27203 15861 27215 15895
rect 27157 15855 27215 15861
rect 30653 15895 30711 15901
rect 30653 15861 30665 15895
rect 30699 15892 30711 15895
rect 32122 15892 32128 15904
rect 30699 15864 32128 15892
rect 30699 15861 30711 15864
rect 30653 15855 30711 15861
rect 32122 15852 32128 15864
rect 32180 15852 32186 15904
rect 32306 15852 32312 15904
rect 32364 15852 32370 15904
rect 33505 15895 33563 15901
rect 33505 15861 33517 15895
rect 33551 15892 33563 15895
rect 35802 15892 35808 15904
rect 33551 15864 35808 15892
rect 33551 15861 33563 15864
rect 33505 15855 33563 15861
rect 35802 15852 35808 15864
rect 35860 15852 35866 15904
rect 35894 15852 35900 15904
rect 35952 15892 35958 15904
rect 36832 15892 36860 15923
rect 36906 15920 36912 15932
rect 36964 15920 36970 15972
rect 38010 15920 38016 15972
rect 38068 15960 38074 15972
rect 38304 15960 38332 16000
rect 41049 15997 41061 16000
rect 41095 16028 41107 16031
rect 41782 16028 41788 16040
rect 41095 16000 41788 16028
rect 41095 15997 41107 16000
rect 41049 15991 41107 15997
rect 41782 15988 41788 16000
rect 41840 15988 41846 16040
rect 38068 15932 38332 15960
rect 38068 15920 38074 15932
rect 35952 15864 36860 15892
rect 35952 15852 35958 15864
rect 38654 15852 38660 15904
rect 38712 15892 38718 15904
rect 39942 15892 39948 15904
rect 38712 15864 39948 15892
rect 38712 15852 38718 15864
rect 39942 15852 39948 15864
rect 40000 15852 40006 15904
rect 48682 15852 48688 15904
rect 48740 15892 48746 15904
rect 49237 15895 49295 15901
rect 49237 15892 49249 15895
rect 48740 15864 49249 15892
rect 48740 15852 48746 15864
rect 49237 15861 49249 15864
rect 49283 15861 49295 15895
rect 49237 15855 49295 15861
rect 1104 15802 49864 15824
rect 1104 15750 2950 15802
rect 3002 15750 3014 15802
rect 3066 15750 3078 15802
rect 3130 15750 3142 15802
rect 3194 15750 3206 15802
rect 3258 15750 12950 15802
rect 13002 15750 13014 15802
rect 13066 15750 13078 15802
rect 13130 15750 13142 15802
rect 13194 15750 13206 15802
rect 13258 15750 22950 15802
rect 23002 15750 23014 15802
rect 23066 15750 23078 15802
rect 23130 15750 23142 15802
rect 23194 15750 23206 15802
rect 23258 15750 32950 15802
rect 33002 15750 33014 15802
rect 33066 15750 33078 15802
rect 33130 15750 33142 15802
rect 33194 15750 33206 15802
rect 33258 15750 42950 15802
rect 43002 15750 43014 15802
rect 43066 15750 43078 15802
rect 43130 15750 43142 15802
rect 43194 15750 43206 15802
rect 43258 15750 49864 15802
rect 1104 15728 49864 15750
rect 1762 15648 1768 15700
rect 1820 15688 1826 15700
rect 1820 15660 10916 15688
rect 1820 15648 1826 15660
rect 1302 15512 1308 15564
rect 1360 15552 1366 15564
rect 2041 15555 2099 15561
rect 2041 15552 2053 15555
rect 1360 15524 2053 15552
rect 1360 15512 1366 15524
rect 2041 15521 2053 15524
rect 2087 15521 2099 15555
rect 2041 15515 2099 15521
rect 10594 15512 10600 15564
rect 10652 15552 10658 15564
rect 10781 15555 10839 15561
rect 10781 15552 10793 15555
rect 10652 15524 10793 15552
rect 10652 15512 10658 15524
rect 10781 15521 10793 15524
rect 10827 15521 10839 15555
rect 10888 15552 10916 15660
rect 11054 15648 11060 15700
rect 11112 15688 11118 15700
rect 11112 15660 12112 15688
rect 11112 15648 11118 15660
rect 12084 15620 12112 15660
rect 12250 15648 12256 15700
rect 12308 15688 12314 15700
rect 13173 15691 13231 15697
rect 13173 15688 13185 15691
rect 12308 15660 13185 15688
rect 12308 15648 12314 15660
rect 13173 15657 13185 15660
rect 13219 15657 13231 15691
rect 13173 15651 13231 15657
rect 13262 15648 13268 15700
rect 13320 15688 13326 15700
rect 13320 15660 13676 15688
rect 13320 15648 13326 15660
rect 13446 15620 13452 15632
rect 12084 15592 13452 15620
rect 13446 15580 13452 15592
rect 13504 15580 13510 15632
rect 13648 15620 13676 15660
rect 15562 15648 15568 15700
rect 15620 15648 15626 15700
rect 16758 15648 16764 15700
rect 16816 15648 16822 15700
rect 16942 15648 16948 15700
rect 17000 15688 17006 15700
rect 18049 15691 18107 15697
rect 17000 15660 17448 15688
rect 17000 15648 17006 15660
rect 13648 15592 13768 15620
rect 11054 15552 11060 15564
rect 10888 15524 11060 15552
rect 10781 15515 10839 15521
rect 11054 15512 11060 15524
rect 11112 15512 11118 15564
rect 13354 15512 13360 15564
rect 13412 15552 13418 15564
rect 13740 15561 13768 15592
rect 14550 15580 14556 15632
rect 14608 15620 14614 15632
rect 17420 15620 17448 15660
rect 18049 15657 18061 15691
rect 18095 15688 18107 15691
rect 18414 15688 18420 15700
rect 18095 15660 18420 15688
rect 18095 15657 18107 15660
rect 18049 15651 18107 15657
rect 18414 15648 18420 15660
rect 18472 15648 18478 15700
rect 19150 15648 19156 15700
rect 19208 15688 19214 15700
rect 19889 15691 19947 15697
rect 19889 15688 19901 15691
rect 19208 15660 19901 15688
rect 19208 15648 19214 15660
rect 19889 15657 19901 15660
rect 19935 15657 19947 15691
rect 19889 15651 19947 15657
rect 20438 15648 20444 15700
rect 20496 15688 20502 15700
rect 21177 15691 21235 15697
rect 21177 15688 21189 15691
rect 20496 15660 21189 15688
rect 20496 15648 20502 15660
rect 21177 15657 21189 15660
rect 21223 15657 21235 15691
rect 21177 15651 21235 15657
rect 23474 15648 23480 15700
rect 23532 15688 23538 15700
rect 25869 15691 25927 15697
rect 25869 15688 25881 15691
rect 23532 15660 25881 15688
rect 23532 15648 23538 15660
rect 25869 15657 25881 15660
rect 25915 15657 25927 15691
rect 26510 15688 26516 15700
rect 25869 15651 25927 15657
rect 25976 15660 26516 15688
rect 21634 15620 21640 15632
rect 14608 15592 17356 15620
rect 17420 15592 21640 15620
rect 14608 15580 14614 15592
rect 13633 15555 13691 15561
rect 13633 15552 13645 15555
rect 13412 15524 13645 15552
rect 13412 15512 13418 15524
rect 13633 15521 13645 15524
rect 13679 15521 13691 15555
rect 13633 15515 13691 15521
rect 13725 15555 13783 15561
rect 13725 15521 13737 15555
rect 13771 15552 13783 15555
rect 15010 15552 15016 15564
rect 13771 15524 15016 15552
rect 13771 15521 13783 15524
rect 13725 15515 13783 15521
rect 15010 15512 15016 15524
rect 15068 15512 15074 15564
rect 16114 15512 16120 15564
rect 16172 15552 16178 15564
rect 16298 15552 16304 15564
rect 16172 15524 16304 15552
rect 16172 15512 16178 15524
rect 16298 15512 16304 15524
rect 16356 15512 16362 15564
rect 17328 15561 17356 15592
rect 21634 15580 21640 15592
rect 21692 15580 21698 15632
rect 17313 15555 17371 15561
rect 17313 15521 17325 15555
rect 17359 15521 17371 15555
rect 17313 15515 17371 15521
rect 18322 15512 18328 15564
rect 18380 15552 18386 15564
rect 19058 15552 19064 15564
rect 18380 15524 19064 15552
rect 18380 15512 18386 15524
rect 19058 15512 19064 15524
rect 19116 15512 19122 15564
rect 20533 15555 20591 15561
rect 20533 15521 20545 15555
rect 20579 15552 20591 15555
rect 21358 15552 21364 15564
rect 20579 15524 21364 15552
rect 20579 15521 20591 15524
rect 20533 15515 20591 15521
rect 21358 15512 21364 15524
rect 21416 15512 21422 15564
rect 21450 15512 21456 15564
rect 21508 15552 21514 15564
rect 21729 15555 21787 15561
rect 21729 15552 21741 15555
rect 21508 15524 21741 15552
rect 21508 15512 21514 15524
rect 21729 15521 21741 15524
rect 21775 15521 21787 15555
rect 21729 15515 21787 15521
rect 23658 15512 23664 15564
rect 23716 15512 23722 15564
rect 24854 15512 24860 15564
rect 24912 15552 24918 15564
rect 25317 15555 25375 15561
rect 25317 15552 25329 15555
rect 24912 15524 25329 15552
rect 24912 15512 24918 15524
rect 25317 15521 25329 15524
rect 25363 15552 25375 15555
rect 25976 15552 26004 15660
rect 26510 15648 26516 15660
rect 26568 15648 26574 15700
rect 29181 15691 29239 15697
rect 29181 15657 29193 15691
rect 29227 15688 29239 15691
rect 31294 15688 31300 15700
rect 29227 15660 31300 15688
rect 29227 15657 29239 15660
rect 29181 15651 29239 15657
rect 31294 15648 31300 15660
rect 31352 15648 31358 15700
rect 32214 15648 32220 15700
rect 32272 15648 32278 15700
rect 34054 15648 34060 15700
rect 34112 15688 34118 15700
rect 35148 15691 35206 15697
rect 35148 15688 35160 15691
rect 34112 15660 35160 15688
rect 34112 15648 34118 15660
rect 35148 15657 35160 15660
rect 35194 15688 35206 15691
rect 36354 15688 36360 15700
rect 35194 15660 36360 15688
rect 35194 15657 35206 15660
rect 35148 15651 35206 15657
rect 36354 15648 36360 15660
rect 36412 15648 36418 15700
rect 36633 15691 36691 15697
rect 36633 15657 36645 15691
rect 36679 15688 36691 15691
rect 37366 15688 37372 15700
rect 36679 15660 37372 15688
rect 36679 15657 36691 15660
rect 36633 15651 36691 15657
rect 37366 15648 37372 15660
rect 37424 15648 37430 15700
rect 37642 15648 37648 15700
rect 37700 15688 37706 15700
rect 39485 15691 39543 15697
rect 39485 15688 39497 15691
rect 37700 15660 39497 15688
rect 37700 15648 37706 15660
rect 39485 15657 39497 15660
rect 39531 15657 39543 15691
rect 39485 15651 39543 15657
rect 41782 15648 41788 15700
rect 41840 15648 41846 15700
rect 48958 15648 48964 15700
rect 49016 15688 49022 15700
rect 49145 15691 49203 15697
rect 49145 15688 49157 15691
rect 49016 15660 49157 15688
rect 49016 15648 49022 15660
rect 49145 15657 49157 15660
rect 49191 15657 49203 15691
rect 49145 15651 49203 15657
rect 29730 15620 29736 15632
rect 25363 15524 26004 15552
rect 26344 15592 29736 15620
rect 25363 15521 25375 15524
rect 25317 15515 25375 15521
rect 1765 15487 1823 15493
rect 1765 15453 1777 15487
rect 1811 15484 1823 15487
rect 10410 15484 10416 15496
rect 1811 15456 10416 15484
rect 1811 15453 1823 15456
rect 1765 15447 1823 15453
rect 10410 15444 10416 15456
rect 10468 15444 10474 15496
rect 12342 15444 12348 15496
rect 12400 15484 12406 15496
rect 13541 15487 13599 15493
rect 12400 15456 13492 15484
rect 12400 15444 12406 15456
rect 6549 15419 6607 15425
rect 6549 15385 6561 15419
rect 6595 15416 6607 15419
rect 10962 15416 10968 15428
rect 6595 15388 10968 15416
rect 6595 15385 6607 15388
rect 6549 15379 6607 15385
rect 10962 15376 10968 15388
rect 11020 15376 11026 15428
rect 11057 15419 11115 15425
rect 11057 15385 11069 15419
rect 11103 15385 11115 15419
rect 11057 15379 11115 15385
rect 6638 15308 6644 15360
rect 6696 15308 6702 15360
rect 11072 15348 11100 15379
rect 12066 15376 12072 15428
rect 12124 15376 12130 15428
rect 13262 15416 13268 15428
rect 12360 15388 13268 15416
rect 12360 15348 12388 15388
rect 13262 15376 13268 15388
rect 13320 15376 13326 15428
rect 13464 15416 13492 15456
rect 13541 15453 13553 15487
rect 13587 15484 13599 15487
rect 14366 15484 14372 15496
rect 13587 15456 14372 15484
rect 13587 15453 13599 15456
rect 13541 15447 13599 15453
rect 14366 15444 14372 15456
rect 14424 15444 14430 15496
rect 15286 15444 15292 15496
rect 15344 15484 15350 15496
rect 15933 15487 15991 15493
rect 15933 15484 15945 15487
rect 15344 15456 15945 15484
rect 15344 15444 15350 15456
rect 15933 15453 15945 15456
rect 15979 15453 15991 15487
rect 15933 15447 15991 15453
rect 17221 15487 17279 15493
rect 17221 15453 17233 15487
rect 17267 15484 17279 15487
rect 18414 15484 18420 15496
rect 17267 15456 18420 15484
rect 17267 15453 17279 15456
rect 17221 15447 17279 15453
rect 18414 15444 18420 15456
rect 18472 15444 18478 15496
rect 18601 15487 18659 15493
rect 18601 15453 18613 15487
rect 18647 15484 18659 15487
rect 22830 15484 22836 15496
rect 18647 15456 22836 15484
rect 18647 15453 18659 15456
rect 18601 15447 18659 15453
rect 22830 15444 22836 15456
rect 22888 15444 22894 15496
rect 23569 15487 23627 15493
rect 23569 15453 23581 15487
rect 23615 15484 23627 15487
rect 24670 15484 24676 15496
rect 23615 15456 24676 15484
rect 23615 15453 23627 15456
rect 23569 15447 23627 15453
rect 24670 15444 24676 15456
rect 24728 15444 24734 15496
rect 25133 15487 25191 15493
rect 25133 15453 25145 15487
rect 25179 15484 25191 15487
rect 26050 15484 26056 15496
rect 25179 15456 26056 15484
rect 25179 15453 25191 15456
rect 25133 15447 25191 15453
rect 26050 15444 26056 15456
rect 26108 15444 26114 15496
rect 26234 15444 26240 15496
rect 26292 15444 26298 15496
rect 16114 15416 16120 15428
rect 13464 15388 16120 15416
rect 16114 15376 16120 15388
rect 16172 15416 16178 15428
rect 20349 15419 20407 15425
rect 16172 15388 17264 15416
rect 16172 15376 16178 15388
rect 11072 15320 12388 15348
rect 12434 15308 12440 15360
rect 12492 15348 12498 15360
rect 12529 15351 12587 15357
rect 12529 15348 12541 15351
rect 12492 15320 12541 15348
rect 12492 15308 12498 15320
rect 12529 15317 12541 15320
rect 12575 15348 12587 15351
rect 13538 15348 13544 15360
rect 12575 15320 13544 15348
rect 12575 15317 12587 15320
rect 12529 15311 12587 15317
rect 13538 15308 13544 15320
rect 13596 15308 13602 15360
rect 14826 15308 14832 15360
rect 14884 15348 14890 15360
rect 15105 15351 15163 15357
rect 15105 15348 15117 15351
rect 14884 15320 15117 15348
rect 14884 15308 14890 15320
rect 15105 15317 15117 15320
rect 15151 15348 15163 15351
rect 16025 15351 16083 15357
rect 16025 15348 16037 15351
rect 15151 15320 16037 15348
rect 15151 15317 15163 15320
rect 15105 15311 15163 15317
rect 16025 15317 16037 15320
rect 16071 15348 16083 15351
rect 16942 15348 16948 15360
rect 16071 15320 16948 15348
rect 16071 15317 16083 15320
rect 16025 15311 16083 15317
rect 16942 15308 16948 15320
rect 17000 15308 17006 15360
rect 17034 15308 17040 15360
rect 17092 15348 17098 15360
rect 17129 15351 17187 15357
rect 17129 15348 17141 15351
rect 17092 15320 17141 15348
rect 17092 15308 17098 15320
rect 17129 15317 17141 15320
rect 17175 15317 17187 15351
rect 17236 15348 17264 15388
rect 20349 15385 20361 15419
rect 20395 15416 20407 15419
rect 23477 15419 23535 15425
rect 20395 15388 22094 15416
rect 20395 15385 20407 15388
rect 20349 15379 20407 15385
rect 18417 15351 18475 15357
rect 18417 15348 18429 15351
rect 17236 15320 18429 15348
rect 17129 15311 17187 15317
rect 18417 15317 18429 15320
rect 18463 15317 18475 15351
rect 18417 15311 18475 15317
rect 19978 15308 19984 15360
rect 20036 15348 20042 15360
rect 20257 15351 20315 15357
rect 20257 15348 20269 15351
rect 20036 15320 20269 15348
rect 20036 15308 20042 15320
rect 20257 15317 20269 15320
rect 20303 15317 20315 15351
rect 20257 15311 20315 15317
rect 21542 15308 21548 15360
rect 21600 15308 21606 15360
rect 21637 15351 21695 15357
rect 21637 15317 21649 15351
rect 21683 15348 21695 15351
rect 21726 15348 21732 15360
rect 21683 15320 21732 15348
rect 21683 15317 21695 15320
rect 21637 15311 21695 15317
rect 21726 15308 21732 15320
rect 21784 15308 21790 15360
rect 22066 15348 22094 15388
rect 23477 15385 23489 15419
rect 23523 15385 23535 15419
rect 23477 15379 23535 15385
rect 25041 15419 25099 15425
rect 25041 15385 25053 15419
rect 25087 15416 25099 15419
rect 25406 15416 25412 15428
rect 25087 15388 25412 15416
rect 25087 15385 25099 15388
rect 25041 15379 25099 15385
rect 23109 15351 23167 15357
rect 23109 15348 23121 15351
rect 22066 15320 23121 15348
rect 23109 15317 23121 15320
rect 23155 15317 23167 15351
rect 23492 15348 23520 15379
rect 25406 15376 25412 15388
rect 25464 15376 25470 15428
rect 26142 15376 26148 15428
rect 26200 15416 26206 15428
rect 26344 15425 26372 15592
rect 29730 15580 29736 15592
rect 29788 15580 29794 15632
rect 32677 15623 32735 15629
rect 32677 15589 32689 15623
rect 32723 15620 32735 15623
rect 34790 15620 34796 15632
rect 32723 15592 34796 15620
rect 32723 15589 32735 15592
rect 32677 15583 32735 15589
rect 34790 15580 34796 15592
rect 34848 15580 34854 15632
rect 26418 15512 26424 15564
rect 26476 15512 26482 15564
rect 26510 15512 26516 15564
rect 26568 15552 26574 15564
rect 27985 15555 28043 15561
rect 27985 15552 27997 15555
rect 26568 15524 27997 15552
rect 26568 15512 26574 15524
rect 27985 15521 27997 15524
rect 28031 15521 28043 15555
rect 27985 15515 28043 15521
rect 28534 15512 28540 15564
rect 28592 15552 28598 15564
rect 30469 15555 30527 15561
rect 30469 15552 30481 15555
rect 28592 15524 30481 15552
rect 28592 15512 28598 15524
rect 30469 15521 30481 15524
rect 30515 15521 30527 15555
rect 30469 15515 30527 15521
rect 32398 15512 32404 15564
rect 32456 15552 32462 15564
rect 33137 15555 33195 15561
rect 33137 15552 33149 15555
rect 32456 15524 33149 15552
rect 32456 15512 32462 15524
rect 33137 15521 33149 15524
rect 33183 15521 33195 15555
rect 33137 15515 33195 15521
rect 33321 15555 33379 15561
rect 33321 15521 33333 15555
rect 33367 15552 33379 15555
rect 33502 15552 33508 15564
rect 33367 15524 33508 15552
rect 33367 15521 33379 15524
rect 33321 15515 33379 15521
rect 33502 15512 33508 15524
rect 33560 15512 33566 15564
rect 35158 15512 35164 15564
rect 35216 15552 35222 15564
rect 37277 15555 37335 15561
rect 37277 15552 37289 15555
rect 35216 15524 37289 15552
rect 35216 15512 35222 15524
rect 37277 15521 37289 15524
rect 37323 15521 37335 15555
rect 40037 15555 40095 15561
rect 40037 15552 40049 15555
rect 37277 15515 37335 15521
rect 37752 15524 40049 15552
rect 37752 15496 37780 15524
rect 40037 15521 40049 15524
rect 40083 15521 40095 15555
rect 40037 15515 40095 15521
rect 27801 15487 27859 15493
rect 27801 15453 27813 15487
rect 27847 15484 27859 15487
rect 28350 15484 28356 15496
rect 27847 15456 28356 15484
rect 27847 15453 27859 15456
rect 27801 15447 27859 15453
rect 28350 15444 28356 15456
rect 28408 15444 28414 15496
rect 30006 15444 30012 15496
rect 30064 15444 30070 15496
rect 34054 15444 34060 15496
rect 34112 15444 34118 15496
rect 34882 15444 34888 15496
rect 34940 15444 34946 15496
rect 37090 15444 37096 15496
rect 37148 15484 37154 15496
rect 37734 15484 37740 15496
rect 37148 15456 37740 15484
rect 37148 15444 37154 15456
rect 37734 15444 37740 15456
rect 37792 15444 37798 15496
rect 49326 15444 49332 15496
rect 49384 15444 49390 15496
rect 26329 15419 26387 15425
rect 26329 15416 26341 15419
rect 26200 15388 26341 15416
rect 26200 15376 26206 15388
rect 26329 15385 26341 15388
rect 26375 15385 26387 15419
rect 26329 15379 26387 15385
rect 27893 15419 27951 15425
rect 27893 15385 27905 15419
rect 27939 15416 27951 15419
rect 28442 15416 28448 15428
rect 27939 15388 28448 15416
rect 27939 15385 27951 15388
rect 27893 15379 27951 15385
rect 28442 15376 28448 15388
rect 28500 15376 28506 15428
rect 30282 15376 30288 15428
rect 30340 15416 30346 15428
rect 30466 15416 30472 15428
rect 30340 15388 30472 15416
rect 30340 15376 30346 15388
rect 30466 15376 30472 15388
rect 30524 15416 30530 15428
rect 30745 15419 30803 15425
rect 30745 15416 30757 15419
rect 30524 15388 30757 15416
rect 30524 15376 30530 15388
rect 30745 15385 30757 15388
rect 30791 15385 30803 15419
rect 34422 15416 34428 15428
rect 31970 15388 34428 15416
rect 30745 15379 30803 15385
rect 34422 15376 34428 15388
rect 34480 15376 34486 15428
rect 36446 15416 36452 15428
rect 36386 15388 36452 15416
rect 36446 15376 36452 15388
rect 36504 15376 36510 15428
rect 37550 15376 37556 15428
rect 37608 15416 37614 15428
rect 38010 15416 38016 15428
rect 37608 15388 38016 15416
rect 37608 15376 37614 15388
rect 38010 15376 38016 15388
rect 38068 15376 38074 15428
rect 39238 15388 39344 15416
rect 24673 15351 24731 15357
rect 24673 15348 24685 15351
rect 23492 15320 24685 15348
rect 23109 15311 23167 15317
rect 24673 15317 24685 15320
rect 24719 15317 24731 15351
rect 24673 15311 24731 15317
rect 26602 15308 26608 15360
rect 26660 15348 26666 15360
rect 27433 15351 27491 15357
rect 27433 15348 27445 15351
rect 26660 15320 27445 15348
rect 26660 15308 26666 15320
rect 27433 15317 27445 15320
rect 27479 15317 27491 15351
rect 27433 15311 27491 15317
rect 29638 15308 29644 15360
rect 29696 15348 29702 15360
rect 30374 15348 30380 15360
rect 29696 15320 30380 15348
rect 29696 15308 29702 15320
rect 30374 15308 30380 15320
rect 30432 15308 30438 15360
rect 31110 15308 31116 15360
rect 31168 15348 31174 15360
rect 31754 15348 31760 15360
rect 31168 15320 31760 15348
rect 31168 15308 31174 15320
rect 31754 15308 31760 15320
rect 31812 15308 31818 15360
rect 32030 15308 32036 15360
rect 32088 15348 32094 15360
rect 32398 15348 32404 15360
rect 32088 15320 32404 15348
rect 32088 15308 32094 15320
rect 32398 15308 32404 15320
rect 32456 15348 32462 15360
rect 33045 15351 33103 15357
rect 33045 15348 33057 15351
rect 32456 15320 33057 15348
rect 32456 15308 32462 15320
rect 33045 15317 33057 15320
rect 33091 15317 33103 15351
rect 33045 15311 33103 15317
rect 33686 15308 33692 15360
rect 33744 15348 33750 15360
rect 34514 15348 34520 15360
rect 33744 15320 34520 15348
rect 33744 15308 33750 15320
rect 34514 15308 34520 15320
rect 34572 15308 34578 15360
rect 35250 15308 35256 15360
rect 35308 15348 35314 15360
rect 35894 15348 35900 15360
rect 35308 15320 35900 15348
rect 35308 15308 35314 15320
rect 35894 15308 35900 15320
rect 35952 15308 35958 15360
rect 39316 15348 39344 15388
rect 39942 15376 39948 15428
rect 40000 15416 40006 15428
rect 40313 15419 40371 15425
rect 40313 15416 40325 15419
rect 40000 15388 40325 15416
rect 40000 15376 40006 15388
rect 40313 15385 40325 15388
rect 40359 15385 40371 15419
rect 40313 15379 40371 15385
rect 40420 15388 40802 15416
rect 39574 15348 39580 15360
rect 39316 15320 39580 15348
rect 39574 15308 39580 15320
rect 39632 15348 39638 15360
rect 40420 15348 40448 15388
rect 39632 15320 40448 15348
rect 39632 15308 39638 15320
rect 1104 15258 49864 15280
rect 1104 15206 7950 15258
rect 8002 15206 8014 15258
rect 8066 15206 8078 15258
rect 8130 15206 8142 15258
rect 8194 15206 8206 15258
rect 8258 15206 17950 15258
rect 18002 15206 18014 15258
rect 18066 15206 18078 15258
rect 18130 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 27950 15258
rect 28002 15206 28014 15258
rect 28066 15206 28078 15258
rect 28130 15206 28142 15258
rect 28194 15206 28206 15258
rect 28258 15206 37950 15258
rect 38002 15206 38014 15258
rect 38066 15206 38078 15258
rect 38130 15206 38142 15258
rect 38194 15206 38206 15258
rect 38258 15206 47950 15258
rect 48002 15206 48014 15258
rect 48066 15206 48078 15258
rect 48130 15206 48142 15258
rect 48194 15206 48206 15258
rect 48258 15206 49864 15258
rect 1104 15184 49864 15206
rect 9214 15104 9220 15156
rect 9272 15144 9278 15156
rect 9769 15147 9827 15153
rect 9769 15144 9781 15147
rect 9272 15116 9781 15144
rect 9272 15104 9278 15116
rect 9769 15113 9781 15116
rect 9815 15113 9827 15147
rect 9769 15107 9827 15113
rect 11054 15104 11060 15156
rect 11112 15104 11118 15156
rect 11422 15104 11428 15156
rect 11480 15144 11486 15156
rect 11885 15147 11943 15153
rect 11885 15144 11897 15147
rect 11480 15116 11897 15144
rect 11480 15104 11486 15116
rect 11885 15113 11897 15116
rect 11931 15113 11943 15147
rect 11885 15107 11943 15113
rect 12250 15104 12256 15156
rect 12308 15104 12314 15156
rect 12406 15116 13124 15144
rect 9582 15036 9588 15088
rect 9640 15076 9646 15088
rect 9861 15079 9919 15085
rect 9861 15076 9873 15079
rect 9640 15048 9873 15076
rect 9640 15036 9646 15048
rect 9861 15045 9873 15048
rect 9907 15045 9919 15079
rect 9861 15039 9919 15045
rect 10965 15079 11023 15085
rect 10965 15045 10977 15079
rect 11011 15076 11023 15079
rect 12406 15076 12434 15116
rect 11011 15048 12434 15076
rect 11011 15045 11023 15048
rect 10965 15039 11023 15045
rect 1765 15011 1823 15017
rect 1765 14977 1777 15011
rect 1811 15008 1823 15011
rect 6638 15008 6644 15020
rect 1811 14980 6644 15008
rect 1811 14977 1823 14980
rect 1765 14971 1823 14977
rect 6638 14968 6644 14980
rect 6696 14968 6702 15020
rect 11054 14968 11060 15020
rect 11112 15008 11118 15020
rect 11790 15008 11796 15020
rect 11112 14980 11796 15008
rect 11112 14968 11118 14980
rect 11790 14968 11796 14980
rect 11848 14968 11854 15020
rect 12158 14968 12164 15020
rect 12216 15008 12222 15020
rect 12216 14980 12480 15008
rect 12216 14968 12222 14980
rect 1302 14900 1308 14952
rect 1360 14940 1366 14952
rect 2041 14943 2099 14949
rect 2041 14940 2053 14943
rect 1360 14912 2053 14940
rect 1360 14900 1366 14912
rect 2041 14909 2053 14912
rect 2087 14909 2099 14943
rect 2041 14903 2099 14909
rect 10045 14943 10103 14949
rect 10045 14909 10057 14943
rect 10091 14940 10103 14943
rect 10778 14940 10784 14952
rect 10091 14912 10784 14940
rect 10091 14909 10103 14912
rect 10045 14903 10103 14909
rect 10778 14900 10784 14912
rect 10836 14900 10842 14952
rect 12452 14949 12480 14980
rect 12345 14943 12403 14949
rect 12345 14909 12357 14943
rect 12391 14909 12403 14943
rect 12345 14903 12403 14909
rect 12437 14943 12495 14949
rect 12437 14909 12449 14943
rect 12483 14909 12495 14943
rect 13096 14940 13124 15116
rect 13722 15104 13728 15156
rect 13780 15144 13786 15156
rect 15565 15147 15623 15153
rect 15565 15144 15577 15147
rect 13780 15116 15577 15144
rect 13780 15104 13786 15116
rect 15565 15113 15577 15116
rect 15611 15113 15623 15147
rect 15565 15107 15623 15113
rect 15654 15104 15660 15156
rect 15712 15144 15718 15156
rect 16025 15147 16083 15153
rect 16025 15144 16037 15147
rect 15712 15116 16037 15144
rect 15712 15104 15718 15116
rect 16025 15113 16037 15116
rect 16071 15113 16083 15147
rect 16025 15107 16083 15113
rect 18874 15104 18880 15156
rect 18932 15144 18938 15156
rect 18932 15116 19472 15144
rect 18932 15104 18938 15116
rect 13814 15076 13820 15088
rect 13280 15048 13820 15076
rect 13170 14968 13176 15020
rect 13228 14968 13234 15020
rect 13280 15017 13308 15048
rect 13814 15036 13820 15048
rect 13872 15036 13878 15088
rect 14182 15036 14188 15088
rect 14240 15036 14246 15088
rect 15933 15079 15991 15085
rect 15933 15045 15945 15079
rect 15979 15076 15991 15079
rect 18046 15076 18052 15088
rect 15979 15048 18052 15076
rect 15979 15045 15991 15048
rect 15933 15039 15991 15045
rect 18046 15036 18052 15048
rect 18104 15036 18110 15088
rect 18690 15036 18696 15088
rect 18748 15036 18754 15088
rect 19444 15076 19472 15116
rect 19518 15104 19524 15156
rect 19576 15104 19582 15156
rect 20346 15144 20352 15156
rect 19628 15116 20352 15144
rect 19628 15076 19656 15116
rect 20346 15104 20352 15116
rect 20404 15104 20410 15156
rect 20438 15104 20444 15156
rect 20496 15144 20502 15156
rect 21726 15144 21732 15156
rect 20496 15116 21732 15144
rect 20496 15104 20502 15116
rect 21726 15104 21732 15116
rect 21784 15104 21790 15156
rect 22554 15104 22560 15156
rect 22612 15144 22618 15156
rect 22925 15147 22983 15153
rect 22925 15144 22937 15147
rect 22612 15116 22937 15144
rect 22612 15104 22618 15116
rect 22925 15113 22937 15116
rect 22971 15113 22983 15147
rect 22925 15107 22983 15113
rect 23750 15104 23756 15156
rect 23808 15144 23814 15156
rect 24121 15147 24179 15153
rect 24121 15144 24133 15147
rect 23808 15116 24133 15144
rect 23808 15104 23814 15116
rect 24121 15113 24133 15116
rect 24167 15113 24179 15147
rect 24121 15107 24179 15113
rect 25130 15104 25136 15156
rect 25188 15104 25194 15156
rect 26421 15147 26479 15153
rect 25240 15116 25820 15144
rect 19444 15048 19656 15076
rect 19889 15079 19947 15085
rect 19889 15045 19901 15079
rect 19935 15076 19947 15079
rect 20806 15076 20812 15088
rect 19935 15048 20812 15076
rect 19935 15045 19947 15048
rect 19889 15039 19947 15045
rect 20806 15036 20812 15048
rect 20864 15036 20870 15088
rect 21082 15036 21088 15088
rect 21140 15036 21146 15088
rect 21174 15036 21180 15088
rect 21232 15076 21238 15088
rect 21232 15048 24624 15076
rect 21232 15036 21238 15048
rect 13265 15011 13323 15017
rect 13265 14977 13277 15011
rect 13311 14977 13323 15011
rect 17221 15011 17279 15017
rect 13265 14971 13323 14977
rect 14936 14980 17172 15008
rect 14936 14940 14964 14980
rect 13096 14912 14964 14940
rect 12437 14903 12495 14909
rect 2314 14832 2320 14884
rect 2372 14872 2378 14884
rect 12250 14872 12256 14884
rect 2372 14844 12256 14872
rect 2372 14832 2378 14844
rect 12250 14832 12256 14844
rect 12308 14832 12314 14884
rect 12360 14872 12388 14903
rect 15010 14900 15016 14952
rect 15068 14940 15074 14952
rect 16117 14943 16175 14949
rect 16117 14940 16129 14943
rect 15068 14912 16129 14940
rect 15068 14900 15074 14912
rect 16117 14909 16129 14912
rect 16163 14909 16175 14943
rect 16117 14903 16175 14909
rect 13170 14872 13176 14884
rect 12360 14844 13176 14872
rect 13170 14832 13176 14844
rect 13228 14832 13234 14884
rect 16132 14872 16160 14903
rect 16942 14872 16948 14884
rect 16132 14844 16948 14872
rect 16942 14832 16948 14844
rect 17000 14832 17006 14884
rect 17144 14872 17172 14980
rect 17221 14977 17233 15011
rect 17267 15008 17279 15011
rect 18141 15011 18199 15017
rect 18141 15008 18153 15011
rect 17267 14980 18153 15008
rect 17267 14977 17279 14980
rect 17221 14971 17279 14977
rect 18141 14977 18153 14980
rect 18187 15008 18199 15011
rect 18230 15008 18236 15020
rect 18187 14980 18236 15008
rect 18187 14977 18199 14980
rect 18141 14971 18199 14977
rect 18230 14968 18236 14980
rect 18288 14968 18294 15020
rect 18322 14968 18328 15020
rect 18380 15008 18386 15020
rect 18380 14980 18552 15008
rect 18380 14968 18386 14980
rect 17310 14900 17316 14952
rect 17368 14900 17374 14952
rect 17402 14900 17408 14952
rect 17460 14940 17466 14952
rect 18414 14940 18420 14952
rect 17460 14912 18420 14940
rect 17460 14900 17466 14912
rect 18414 14900 18420 14912
rect 18472 14900 18478 14952
rect 18524 14940 18552 14980
rect 18782 14968 18788 15020
rect 18840 14968 18846 15020
rect 19981 15011 20039 15017
rect 19981 14977 19993 15011
rect 20027 15008 20039 15011
rect 20898 15008 20904 15020
rect 20027 14980 20904 15008
rect 20027 14977 20039 14980
rect 19981 14971 20039 14977
rect 20898 14968 20904 14980
rect 20956 14968 20962 15020
rect 22094 14968 22100 15020
rect 22152 15008 22158 15020
rect 23293 15011 23351 15017
rect 23293 15008 23305 15011
rect 22152 14980 23305 15008
rect 22152 14968 22158 14980
rect 23293 14977 23305 14980
rect 23339 14977 23351 15011
rect 23293 14971 23351 14977
rect 24394 14968 24400 15020
rect 24452 15008 24458 15020
rect 24596 15017 24624 15048
rect 24854 15036 24860 15088
rect 24912 15076 24918 15088
rect 25240 15076 25268 15116
rect 24912 15048 25268 15076
rect 25593 15079 25651 15085
rect 24912 15036 24918 15048
rect 25593 15045 25605 15079
rect 25639 15076 25651 15079
rect 25682 15076 25688 15088
rect 25639 15048 25688 15076
rect 25639 15045 25651 15048
rect 25593 15039 25651 15045
rect 25682 15036 25688 15048
rect 25740 15036 25746 15088
rect 25792 15076 25820 15116
rect 26421 15113 26433 15147
rect 26467 15144 26479 15147
rect 26694 15144 26700 15156
rect 26467 15116 26700 15144
rect 26467 15113 26479 15116
rect 26421 15107 26479 15113
rect 26694 15104 26700 15116
rect 26752 15144 26758 15156
rect 27617 15147 27675 15153
rect 27617 15144 27629 15147
rect 26752 15116 27629 15144
rect 26752 15104 26758 15116
rect 27617 15113 27629 15116
rect 27663 15113 27675 15147
rect 30101 15147 30159 15153
rect 27617 15107 27675 15113
rect 27724 15116 29776 15144
rect 27724 15076 27752 15116
rect 28813 15079 28871 15085
rect 28813 15076 28825 15079
rect 25792 15048 27752 15076
rect 28276 15048 28825 15076
rect 24489 15011 24547 15017
rect 24489 15008 24501 15011
rect 24452 14980 24501 15008
rect 24452 14968 24458 14980
rect 24489 14977 24501 14980
rect 24535 14977 24547 15011
rect 24489 14971 24547 14977
rect 24581 15011 24639 15017
rect 24581 14977 24593 15011
rect 24627 15008 24639 15011
rect 24627 14980 25452 15008
rect 24627 14977 24639 14980
rect 24581 14971 24639 14977
rect 18877 14943 18935 14949
rect 18877 14940 18889 14943
rect 18524 14912 18889 14940
rect 18877 14909 18889 14912
rect 18923 14909 18935 14943
rect 18877 14903 18935 14909
rect 20070 14900 20076 14952
rect 20128 14900 20134 14952
rect 20346 14900 20352 14952
rect 20404 14940 20410 14952
rect 20404 14912 20944 14940
rect 20404 14900 20410 14912
rect 17218 14872 17224 14884
rect 17144 14844 17224 14872
rect 17218 14832 17224 14844
rect 17276 14832 17282 14884
rect 17494 14832 17500 14884
rect 17552 14872 17558 14884
rect 20717 14875 20775 14881
rect 20717 14872 20729 14875
rect 17552 14844 20729 14872
rect 17552 14832 17558 14844
rect 20717 14841 20729 14844
rect 20763 14841 20775 14875
rect 20916 14872 20944 14912
rect 20990 14900 20996 14952
rect 21048 14940 21054 14952
rect 21177 14943 21235 14949
rect 21177 14940 21189 14943
rect 21048 14912 21189 14940
rect 21048 14900 21054 14912
rect 21177 14909 21189 14912
rect 21223 14909 21235 14943
rect 21177 14903 21235 14909
rect 21269 14943 21327 14949
rect 21269 14909 21281 14943
rect 21315 14909 21327 14943
rect 21269 14903 21327 14909
rect 21284 14872 21312 14903
rect 22646 14900 22652 14952
rect 22704 14940 22710 14952
rect 23385 14943 23443 14949
rect 23385 14940 23397 14943
rect 22704 14912 23397 14940
rect 22704 14900 22710 14912
rect 23385 14909 23397 14912
rect 23431 14909 23443 14943
rect 23385 14903 23443 14909
rect 23477 14943 23535 14949
rect 23477 14909 23489 14943
rect 23523 14909 23535 14943
rect 23477 14903 23535 14909
rect 20916 14844 21312 14872
rect 20717 14835 20775 14841
rect 22738 14832 22744 14884
rect 22796 14872 22802 14884
rect 23492 14872 23520 14903
rect 24118 14900 24124 14952
rect 24176 14940 24182 14952
rect 24673 14943 24731 14949
rect 24673 14940 24685 14943
rect 24176 14912 24685 14940
rect 24176 14900 24182 14912
rect 24673 14909 24685 14912
rect 24719 14909 24731 14943
rect 25424 14940 25452 14980
rect 25498 14968 25504 15020
rect 25556 14968 25562 15020
rect 27522 15008 27528 15020
rect 25608 14980 27528 15008
rect 25608 14940 25636 14980
rect 27522 14968 27528 14980
rect 27580 14968 27586 15020
rect 28276 15008 28304 15048
rect 28813 15045 28825 15048
rect 28859 15076 28871 15079
rect 29748 15076 29776 15116
rect 30101 15113 30113 15147
rect 30147 15144 30159 15147
rect 31110 15144 31116 15156
rect 30147 15116 31116 15144
rect 30147 15113 30159 15116
rect 30101 15107 30159 15113
rect 31110 15104 31116 15116
rect 31168 15104 31174 15156
rect 31389 15147 31447 15153
rect 31389 15113 31401 15147
rect 31435 15144 31447 15147
rect 32030 15144 32036 15156
rect 31435 15116 32036 15144
rect 31435 15113 31447 15116
rect 31389 15107 31447 15113
rect 32030 15104 32036 15116
rect 32088 15104 32094 15156
rect 32306 15104 32312 15156
rect 32364 15144 32370 15156
rect 32677 15147 32735 15153
rect 32677 15144 32689 15147
rect 32364 15116 32689 15144
rect 32364 15104 32370 15116
rect 32677 15113 32689 15116
rect 32723 15113 32735 15147
rect 32677 15107 32735 15113
rect 33505 15147 33563 15153
rect 33505 15113 33517 15147
rect 33551 15144 33563 15147
rect 33686 15144 33692 15156
rect 33551 15116 33692 15144
rect 33551 15113 33563 15116
rect 33505 15107 33563 15113
rect 33686 15104 33692 15116
rect 33744 15104 33750 15156
rect 33873 15147 33931 15153
rect 33873 15113 33885 15147
rect 33919 15144 33931 15147
rect 34054 15144 34060 15156
rect 33919 15116 34060 15144
rect 33919 15113 33931 15116
rect 33873 15107 33931 15113
rect 34054 15104 34060 15116
rect 34112 15104 34118 15156
rect 35069 15147 35127 15153
rect 35069 15113 35081 15147
rect 35115 15144 35127 15147
rect 35158 15144 35164 15156
rect 35115 15116 35164 15144
rect 35115 15113 35127 15116
rect 35069 15107 35127 15113
rect 35158 15104 35164 15116
rect 35216 15104 35222 15156
rect 39669 15147 39727 15153
rect 39669 15144 39681 15147
rect 35728 15116 39681 15144
rect 30742 15076 30748 15088
rect 28859 15048 29592 15076
rect 29748 15048 30748 15076
rect 28859 15045 28871 15048
rect 28813 15039 28871 15045
rect 27632 14980 28304 15008
rect 25424 14912 25636 14940
rect 25777 14943 25835 14949
rect 24673 14903 24731 14909
rect 25777 14909 25789 14943
rect 25823 14940 25835 14943
rect 25866 14940 25872 14952
rect 25823 14912 25872 14940
rect 25823 14909 25835 14912
rect 25777 14903 25835 14909
rect 25866 14900 25872 14912
rect 25924 14900 25930 14952
rect 26142 14900 26148 14952
rect 26200 14940 26206 14952
rect 27632 14940 27660 14980
rect 28350 14968 28356 15020
rect 28408 15008 28414 15020
rect 28721 15011 28779 15017
rect 28721 15008 28733 15011
rect 28408 14980 28733 15008
rect 28408 14968 28414 14980
rect 28721 14977 28733 14980
rect 28767 14977 28779 15011
rect 28721 14971 28779 14977
rect 29564 14952 29592 15048
rect 30742 15036 30748 15048
rect 30800 15036 30806 15088
rect 31481 15079 31539 15085
rect 31481 15045 31493 15079
rect 31527 15076 31539 15079
rect 31527 15048 32536 15076
rect 31527 15045 31539 15048
rect 31481 15039 31539 15045
rect 29730 14968 29736 15020
rect 29788 14968 29794 15020
rect 31754 14968 31760 15020
rect 31812 15008 31818 15020
rect 31864 15008 31984 15012
rect 31812 14984 31984 15008
rect 31812 14980 31892 14984
rect 31812 14968 31818 14980
rect 26200 14912 27660 14940
rect 27709 14943 27767 14949
rect 26200 14900 26206 14912
rect 27709 14909 27721 14943
rect 27755 14909 27767 14943
rect 27709 14903 27767 14909
rect 28905 14943 28963 14949
rect 28905 14909 28917 14943
rect 28951 14940 28963 14943
rect 29270 14940 29276 14952
rect 28951 14912 29276 14940
rect 28951 14909 28963 14912
rect 28905 14903 28963 14909
rect 22796 14844 23520 14872
rect 22796 14832 22802 14844
rect 24762 14832 24768 14884
rect 24820 14872 24826 14884
rect 27724 14872 27752 14903
rect 29270 14900 29276 14912
rect 29328 14900 29334 14952
rect 29546 14900 29552 14952
rect 29604 14900 29610 14952
rect 24820 14844 27752 14872
rect 28353 14875 28411 14881
rect 24820 14832 24826 14844
rect 28353 14841 28365 14875
rect 28399 14872 28411 14875
rect 29454 14872 29460 14884
rect 28399 14844 29460 14872
rect 28399 14841 28411 14844
rect 28353 14835 28411 14841
rect 29454 14832 29460 14844
rect 29512 14832 29518 14884
rect 29748 14881 29776 14968
rect 30193 14943 30251 14949
rect 30193 14909 30205 14943
rect 30239 14909 30251 14943
rect 30193 14903 30251 14909
rect 30285 14943 30343 14949
rect 30285 14909 30297 14943
rect 30331 14940 30343 14943
rect 30374 14940 30380 14952
rect 30331 14912 30380 14940
rect 30331 14909 30343 14912
rect 30285 14903 30343 14909
rect 29733 14875 29791 14881
rect 29733 14841 29745 14875
rect 29779 14841 29791 14875
rect 30208 14872 30236 14903
rect 30374 14900 30380 14912
rect 30432 14900 30438 14952
rect 31110 14900 31116 14952
rect 31168 14940 31174 14952
rect 31573 14943 31631 14949
rect 31573 14940 31585 14943
rect 31168 14912 31585 14940
rect 31168 14900 31174 14912
rect 31573 14909 31585 14912
rect 31619 14909 31631 14943
rect 31956 14940 31984 14984
rect 32508 15008 32536 15048
rect 32582 15036 32588 15088
rect 32640 15076 32646 15088
rect 32769 15079 32827 15085
rect 32769 15076 32781 15079
rect 32640 15048 32781 15076
rect 32640 15036 32646 15048
rect 32769 15045 32781 15048
rect 32815 15045 32827 15079
rect 35728 15076 35756 15116
rect 39669 15113 39681 15116
rect 39715 15113 39727 15147
rect 39669 15107 39727 15113
rect 40034 15104 40040 15156
rect 40092 15144 40098 15156
rect 40129 15147 40187 15153
rect 40129 15144 40141 15147
rect 40092 15116 40141 15144
rect 40092 15104 40098 15116
rect 40129 15113 40141 15116
rect 40175 15113 40187 15147
rect 40129 15107 40187 15113
rect 32769 15039 32827 15045
rect 32876 15048 35756 15076
rect 36357 15079 36415 15085
rect 32876 15008 32904 15048
rect 36357 15045 36369 15079
rect 36403 15076 36415 15079
rect 36722 15076 36728 15088
rect 36403 15048 36728 15076
rect 36403 15045 36415 15048
rect 36357 15039 36415 15045
rect 36722 15036 36728 15048
rect 36780 15036 36786 15088
rect 37642 15036 37648 15088
rect 37700 15076 37706 15088
rect 37737 15079 37795 15085
rect 37737 15076 37749 15079
rect 37700 15048 37749 15076
rect 37700 15036 37706 15048
rect 37737 15045 37749 15048
rect 37783 15045 37795 15079
rect 37737 15039 37795 15045
rect 37826 15036 37832 15088
rect 37884 15076 37890 15088
rect 37884 15048 38226 15076
rect 37884 15036 37890 15048
rect 32508 14980 32904 15008
rect 33410 14968 33416 15020
rect 33468 15008 33474 15020
rect 36265 15011 36323 15017
rect 36265 15008 36277 15011
rect 33468 14980 36277 15008
rect 33468 14968 33474 14980
rect 36265 14977 36277 14980
rect 36311 14977 36323 15011
rect 37182 15008 37188 15020
rect 36265 14971 36323 14977
rect 36372 14980 37188 15008
rect 32674 14940 32680 14952
rect 31956 14912 32680 14940
rect 31573 14903 31631 14909
rect 32674 14900 32680 14912
rect 32732 14900 32738 14952
rect 32766 14900 32772 14952
rect 32824 14940 32830 14952
rect 32861 14943 32919 14949
rect 32861 14940 32873 14943
rect 32824 14912 32873 14940
rect 32824 14900 32830 14912
rect 32861 14909 32873 14912
rect 32907 14909 32919 14943
rect 32861 14903 32919 14909
rect 33965 14943 34023 14949
rect 33965 14909 33977 14943
rect 34011 14909 34023 14943
rect 33965 14903 34023 14909
rect 29733 14835 29791 14841
rect 30024 14844 30236 14872
rect 9401 14807 9459 14813
rect 9401 14773 9413 14807
rect 9447 14804 9459 14807
rect 10870 14804 10876 14816
rect 9447 14776 10876 14804
rect 9447 14773 9459 14776
rect 9401 14767 9459 14773
rect 10870 14764 10876 14776
rect 10928 14764 10934 14816
rect 13528 14807 13586 14813
rect 13528 14773 13540 14807
rect 13574 14804 13586 14807
rect 13722 14804 13728 14816
rect 13574 14776 13728 14804
rect 13574 14773 13586 14776
rect 13528 14767 13586 14773
rect 13722 14764 13728 14776
rect 13780 14764 13786 14816
rect 15930 14764 15936 14816
rect 15988 14804 15994 14816
rect 16853 14807 16911 14813
rect 16853 14804 16865 14807
rect 15988 14776 16865 14804
rect 15988 14764 15994 14776
rect 16853 14773 16865 14776
rect 16899 14773 16911 14807
rect 16853 14767 16911 14773
rect 18046 14764 18052 14816
rect 18104 14804 18110 14816
rect 18325 14807 18383 14813
rect 18325 14804 18337 14807
rect 18104 14776 18337 14804
rect 18104 14764 18110 14776
rect 18325 14773 18337 14776
rect 18371 14773 18383 14807
rect 18325 14767 18383 14773
rect 18414 14764 18420 14816
rect 18472 14804 18478 14816
rect 19242 14804 19248 14816
rect 18472 14776 19248 14804
rect 18472 14764 18478 14776
rect 19242 14764 19248 14776
rect 19300 14764 19306 14816
rect 20622 14764 20628 14816
rect 20680 14804 20686 14816
rect 24854 14804 24860 14816
rect 20680 14776 24860 14804
rect 20680 14764 20686 14776
rect 24854 14764 24860 14776
rect 24912 14764 24918 14816
rect 24946 14764 24952 14816
rect 25004 14804 25010 14816
rect 25130 14804 25136 14816
rect 25004 14776 25136 14804
rect 25004 14764 25010 14776
rect 25130 14764 25136 14776
rect 25188 14804 25194 14816
rect 25406 14804 25412 14816
rect 25188 14776 25412 14804
rect 25188 14764 25194 14776
rect 25406 14764 25412 14776
rect 25464 14764 25470 14816
rect 26326 14764 26332 14816
rect 26384 14804 26390 14816
rect 27157 14807 27215 14813
rect 27157 14804 27169 14807
rect 26384 14776 27169 14804
rect 26384 14764 26390 14776
rect 27157 14773 27169 14776
rect 27203 14773 27215 14807
rect 27157 14767 27215 14773
rect 27430 14764 27436 14816
rect 27488 14804 27494 14816
rect 30024 14804 30052 14844
rect 32214 14832 32220 14884
rect 32272 14872 32278 14884
rect 33980 14872 34008 14903
rect 34146 14900 34152 14952
rect 34204 14900 34210 14952
rect 34974 14900 34980 14952
rect 35032 14940 35038 14952
rect 35161 14943 35219 14949
rect 35161 14940 35173 14943
rect 35032 14912 35173 14940
rect 35032 14900 35038 14912
rect 35161 14909 35173 14912
rect 35207 14909 35219 14943
rect 35161 14903 35219 14909
rect 35345 14943 35403 14949
rect 35345 14909 35357 14943
rect 35391 14940 35403 14943
rect 36372 14940 36400 14980
rect 37182 14968 37188 14980
rect 37240 14968 37246 15020
rect 40037 15011 40095 15017
rect 40037 14977 40049 15011
rect 40083 15008 40095 15011
rect 40083 14980 40724 15008
rect 40083 14977 40095 14980
rect 40037 14971 40095 14977
rect 35391 14912 36400 14940
rect 35391 14909 35403 14912
rect 35345 14903 35403 14909
rect 36446 14900 36452 14952
rect 36504 14900 36510 14952
rect 37090 14900 37096 14952
rect 37148 14940 37154 14952
rect 37461 14943 37519 14949
rect 37461 14940 37473 14943
rect 37148 14912 37473 14940
rect 37148 14900 37154 14912
rect 37461 14909 37473 14912
rect 37507 14909 37519 14943
rect 37461 14903 37519 14909
rect 38286 14900 38292 14952
rect 38344 14940 38350 14952
rect 39209 14943 39267 14949
rect 39209 14940 39221 14943
rect 38344 14912 39221 14940
rect 38344 14900 38350 14912
rect 39209 14909 39221 14912
rect 39255 14909 39267 14943
rect 39209 14903 39267 14909
rect 39298 14900 39304 14952
rect 39356 14940 39362 14952
rect 40221 14943 40279 14949
rect 40221 14940 40233 14943
rect 39356 14912 40233 14940
rect 39356 14900 39362 14912
rect 40221 14909 40233 14912
rect 40267 14909 40279 14943
rect 40696 14940 40724 14980
rect 40862 14968 40868 15020
rect 40920 15008 40926 15020
rect 41049 15011 41107 15017
rect 41049 15008 41061 15011
rect 40920 14980 41061 15008
rect 40920 14968 40926 14980
rect 41049 14977 41061 14980
rect 41095 14977 41107 15011
rect 41049 14971 41107 14977
rect 49050 14968 49056 15020
rect 49108 14968 49114 15020
rect 48406 14940 48412 14952
rect 40696 14912 48412 14940
rect 40221 14903 40279 14909
rect 48406 14900 48412 14912
rect 48464 14900 48470 14952
rect 32272 14844 34008 14872
rect 34701 14875 34759 14881
rect 32272 14832 32278 14844
rect 34701 14841 34713 14875
rect 34747 14872 34759 14875
rect 36630 14872 36636 14884
rect 34747 14844 36636 14872
rect 34747 14841 34759 14844
rect 34701 14835 34759 14841
rect 36630 14832 36636 14844
rect 36688 14832 36694 14884
rect 48314 14832 48320 14884
rect 48372 14872 48378 14884
rect 49237 14875 49295 14881
rect 49237 14872 49249 14875
rect 48372 14844 49249 14872
rect 48372 14832 48378 14844
rect 49237 14841 49249 14844
rect 49283 14841 49295 14875
rect 49237 14835 49295 14841
rect 27488 14776 30052 14804
rect 27488 14764 27494 14776
rect 30098 14764 30104 14816
rect 30156 14804 30162 14816
rect 31021 14807 31079 14813
rect 31021 14804 31033 14807
rect 30156 14776 31033 14804
rect 30156 14764 30162 14776
rect 31021 14773 31033 14776
rect 31067 14773 31079 14807
rect 31021 14767 31079 14773
rect 31294 14764 31300 14816
rect 31352 14804 31358 14816
rect 31662 14804 31668 14816
rect 31352 14776 31668 14804
rect 31352 14764 31358 14776
rect 31662 14764 31668 14776
rect 31720 14764 31726 14816
rect 32309 14807 32367 14813
rect 32309 14773 32321 14807
rect 32355 14804 32367 14807
rect 35710 14804 35716 14816
rect 32355 14776 35716 14804
rect 32355 14773 32367 14776
rect 32309 14767 32367 14773
rect 35710 14764 35716 14776
rect 35768 14764 35774 14816
rect 35897 14807 35955 14813
rect 35897 14773 35909 14807
rect 35943 14804 35955 14807
rect 37274 14804 37280 14816
rect 35943 14776 37280 14804
rect 35943 14773 35955 14776
rect 35897 14767 35955 14773
rect 37274 14764 37280 14776
rect 37332 14764 37338 14816
rect 38470 14764 38476 14816
rect 38528 14804 38534 14816
rect 39298 14804 39304 14816
rect 38528 14776 39304 14804
rect 38528 14764 38534 14776
rect 39298 14764 39304 14776
rect 39356 14764 39362 14816
rect 40865 14807 40923 14813
rect 40865 14773 40877 14807
rect 40911 14804 40923 14807
rect 45830 14804 45836 14816
rect 40911 14776 45836 14804
rect 40911 14773 40923 14776
rect 40865 14767 40923 14773
rect 45830 14764 45836 14776
rect 45888 14764 45894 14816
rect 1104 14714 49864 14736
rect 1104 14662 2950 14714
rect 3002 14662 3014 14714
rect 3066 14662 3078 14714
rect 3130 14662 3142 14714
rect 3194 14662 3206 14714
rect 3258 14662 12950 14714
rect 13002 14662 13014 14714
rect 13066 14662 13078 14714
rect 13130 14662 13142 14714
rect 13194 14662 13206 14714
rect 13258 14662 22950 14714
rect 23002 14662 23014 14714
rect 23066 14662 23078 14714
rect 23130 14662 23142 14714
rect 23194 14662 23206 14714
rect 23258 14662 32950 14714
rect 33002 14662 33014 14714
rect 33066 14662 33078 14714
rect 33130 14662 33142 14714
rect 33194 14662 33206 14714
rect 33258 14662 42950 14714
rect 43002 14662 43014 14714
rect 43066 14662 43078 14714
rect 43130 14662 43142 14714
rect 43194 14662 43206 14714
rect 43258 14662 49864 14714
rect 1104 14640 49864 14662
rect 10410 14560 10416 14612
rect 10468 14560 10474 14612
rect 11238 14560 11244 14612
rect 11296 14600 11302 14612
rect 11793 14603 11851 14609
rect 11793 14600 11805 14603
rect 11296 14572 11805 14600
rect 11296 14560 11302 14572
rect 11793 14569 11805 14572
rect 11839 14569 11851 14603
rect 11793 14563 11851 14569
rect 12250 14560 12256 14612
rect 12308 14600 12314 14612
rect 14277 14603 14335 14609
rect 14277 14600 14289 14603
rect 12308 14572 14289 14600
rect 12308 14560 12314 14572
rect 14277 14569 14289 14572
rect 14323 14569 14335 14603
rect 16850 14600 16856 14612
rect 14277 14563 14335 14569
rect 14660 14572 16856 14600
rect 3602 14492 3608 14544
rect 3660 14532 3666 14544
rect 12526 14532 12532 14544
rect 3660 14504 12532 14532
rect 3660 14492 3666 14504
rect 12526 14492 12532 14504
rect 12584 14492 12590 14544
rect 12618 14492 12624 14544
rect 12676 14532 12682 14544
rect 12989 14535 13047 14541
rect 12989 14532 13001 14535
rect 12676 14504 13001 14532
rect 12676 14492 12682 14504
rect 12989 14501 13001 14504
rect 13035 14501 13047 14535
rect 14660 14532 14688 14572
rect 16850 14560 16856 14572
rect 16908 14560 16914 14612
rect 17218 14560 17224 14612
rect 17276 14600 17282 14612
rect 20530 14600 20536 14612
rect 17276 14572 20536 14600
rect 17276 14560 17282 14572
rect 20530 14560 20536 14572
rect 20588 14600 20594 14612
rect 24029 14603 24087 14609
rect 20588 14572 23980 14600
rect 20588 14560 20594 14572
rect 18141 14535 18199 14541
rect 18141 14532 18153 14535
rect 12989 14495 13047 14501
rect 13280 14504 14688 14532
rect 14752 14504 18153 14532
rect 1302 14424 1308 14476
rect 1360 14464 1366 14476
rect 2041 14467 2099 14473
rect 2041 14464 2053 14467
rect 1360 14436 2053 14464
rect 1360 14424 1366 14436
rect 2041 14433 2053 14436
rect 2087 14433 2099 14467
rect 2041 14427 2099 14433
rect 11698 14424 11704 14476
rect 11756 14464 11762 14476
rect 12345 14467 12403 14473
rect 11756 14436 12204 14464
rect 11756 14424 11762 14436
rect 1765 14399 1823 14405
rect 1765 14365 1777 14399
rect 1811 14396 1823 14399
rect 9769 14399 9827 14405
rect 9769 14396 9781 14399
rect 1811 14368 9781 14396
rect 1811 14365 1823 14368
rect 1765 14359 1823 14365
rect 9769 14365 9781 14368
rect 9815 14365 9827 14399
rect 12176 14396 12204 14436
rect 12345 14433 12357 14467
rect 12391 14464 12403 14467
rect 13170 14464 13176 14476
rect 12391 14436 13176 14464
rect 12391 14433 12403 14436
rect 12345 14427 12403 14433
rect 13170 14424 13176 14436
rect 13228 14424 13234 14476
rect 13280 14396 13308 14504
rect 13538 14424 13544 14476
rect 13596 14424 13602 14476
rect 14752 14473 14780 14504
rect 18141 14501 18153 14504
rect 18187 14501 18199 14535
rect 19426 14532 19432 14544
rect 18141 14495 18199 14501
rect 18248 14504 19432 14532
rect 14737 14467 14795 14473
rect 14737 14433 14749 14467
rect 14783 14433 14795 14467
rect 14737 14427 14795 14433
rect 14918 14424 14924 14476
rect 14976 14424 14982 14476
rect 15749 14467 15807 14473
rect 15749 14433 15761 14467
rect 15795 14464 15807 14467
rect 16206 14464 16212 14476
rect 15795 14436 16212 14464
rect 15795 14433 15807 14436
rect 15749 14427 15807 14433
rect 16206 14424 16212 14436
rect 16264 14424 16270 14476
rect 16942 14424 16948 14476
rect 17000 14424 17006 14476
rect 18248 14464 18276 14504
rect 19426 14492 19432 14504
rect 19484 14532 19490 14544
rect 20438 14532 20444 14544
rect 19484 14504 20444 14532
rect 19484 14492 19490 14504
rect 20438 14492 20444 14504
rect 20496 14492 20502 14544
rect 22462 14492 22468 14544
rect 22520 14532 22526 14544
rect 22833 14535 22891 14541
rect 22833 14532 22845 14535
rect 22520 14504 22845 14532
rect 22520 14492 22526 14504
rect 22833 14501 22845 14504
rect 22879 14501 22891 14535
rect 23952 14532 23980 14572
rect 24029 14569 24041 14603
rect 24075 14600 24087 14603
rect 25498 14600 25504 14612
rect 24075 14572 25504 14600
rect 24075 14569 24087 14572
rect 24029 14563 24087 14569
rect 25498 14560 25504 14572
rect 25556 14560 25562 14612
rect 26050 14560 26056 14612
rect 26108 14600 26114 14612
rect 27249 14603 27307 14609
rect 27249 14600 27261 14603
rect 26108 14572 27261 14600
rect 26108 14560 26114 14572
rect 27249 14569 27261 14572
rect 27295 14600 27307 14603
rect 27798 14600 27804 14612
rect 27295 14572 27804 14600
rect 27295 14569 27307 14572
rect 27249 14563 27307 14569
rect 27798 14560 27804 14572
rect 27856 14600 27862 14612
rect 28258 14600 28264 14612
rect 27856 14572 28264 14600
rect 27856 14560 27862 14572
rect 28258 14560 28264 14572
rect 28316 14600 28322 14612
rect 28442 14600 28448 14612
rect 28316 14572 28448 14600
rect 28316 14560 28322 14572
rect 28442 14560 28448 14572
rect 28500 14560 28506 14612
rect 29733 14603 29791 14609
rect 29733 14569 29745 14603
rect 29779 14600 29791 14603
rect 33318 14600 33324 14612
rect 29779 14572 33324 14600
rect 29779 14569 29791 14572
rect 29733 14563 29791 14569
rect 33318 14560 33324 14572
rect 33376 14560 33382 14612
rect 33410 14560 33416 14612
rect 33468 14560 33474 14612
rect 35342 14600 35348 14612
rect 34808 14572 35348 14600
rect 24946 14532 24952 14544
rect 23952 14504 24952 14532
rect 22833 14495 22891 14501
rect 24946 14492 24952 14504
rect 25004 14492 25010 14544
rect 26878 14492 26884 14544
rect 26936 14532 26942 14544
rect 26936 14504 30236 14532
rect 26936 14492 26942 14504
rect 17420 14436 18276 14464
rect 18693 14467 18751 14473
rect 12176 14368 13308 14396
rect 13357 14399 13415 14405
rect 9769 14359 9827 14365
rect 13357 14365 13369 14399
rect 13403 14396 13415 14399
rect 13403 14368 15240 14396
rect 13403 14365 13415 14368
rect 13357 14359 13415 14365
rect 9585 14331 9643 14337
rect 9585 14297 9597 14331
rect 9631 14328 9643 14331
rect 10134 14328 10140 14340
rect 9631 14300 10140 14328
rect 9631 14297 9643 14300
rect 9585 14291 9643 14297
rect 10134 14288 10140 14300
rect 10192 14288 10198 14340
rect 10318 14288 10324 14340
rect 10376 14288 10382 14340
rect 11146 14288 11152 14340
rect 11204 14288 11210 14340
rect 12161 14331 12219 14337
rect 12161 14297 12173 14331
rect 12207 14328 12219 14331
rect 12618 14328 12624 14340
rect 12207 14300 12624 14328
rect 12207 14297 12219 14300
rect 12161 14291 12219 14297
rect 12618 14288 12624 14300
rect 12676 14288 12682 14340
rect 14645 14331 14703 14337
rect 14645 14297 14657 14331
rect 14691 14328 14703 14331
rect 15212 14328 15240 14368
rect 15470 14356 15476 14408
rect 15528 14356 15534 14408
rect 16117 14399 16175 14405
rect 16117 14365 16129 14399
rect 16163 14396 16175 14399
rect 16761 14399 16819 14405
rect 16761 14396 16773 14399
rect 16163 14368 16773 14396
rect 16163 14365 16175 14368
rect 16117 14359 16175 14365
rect 16761 14365 16773 14368
rect 16807 14365 16819 14399
rect 17420 14396 17448 14436
rect 18693 14433 18705 14467
rect 18739 14433 18751 14467
rect 18693 14427 18751 14433
rect 16761 14359 16819 14365
rect 16868 14368 17448 14396
rect 14691 14300 15148 14328
rect 15212 14300 16436 14328
rect 14691 14297 14703 14300
rect 14645 14291 14703 14297
rect 11238 14220 11244 14272
rect 11296 14220 11302 14272
rect 12253 14263 12311 14269
rect 12253 14229 12265 14263
rect 12299 14260 12311 14263
rect 12526 14260 12532 14272
rect 12299 14232 12532 14260
rect 12299 14229 12311 14232
rect 12253 14223 12311 14229
rect 12526 14220 12532 14232
rect 12584 14220 12590 14272
rect 13449 14263 13507 14269
rect 13449 14229 13461 14263
rect 13495 14260 13507 14263
rect 13722 14260 13728 14272
rect 13495 14232 13728 14260
rect 13495 14229 13507 14232
rect 13449 14223 13507 14229
rect 13722 14220 13728 14232
rect 13780 14220 13786 14272
rect 15120 14269 15148 14300
rect 15105 14263 15163 14269
rect 15105 14229 15117 14263
rect 15151 14229 15163 14263
rect 15105 14223 15163 14229
rect 15565 14263 15623 14269
rect 15565 14229 15577 14263
rect 15611 14260 15623 14263
rect 15654 14260 15660 14272
rect 15611 14232 15660 14260
rect 15611 14229 15623 14232
rect 15565 14223 15623 14229
rect 15654 14220 15660 14232
rect 15712 14220 15718 14272
rect 16408 14269 16436 14300
rect 16393 14263 16451 14269
rect 16393 14229 16405 14263
rect 16439 14229 16451 14263
rect 16393 14223 16451 14229
rect 16758 14220 16764 14272
rect 16816 14260 16822 14272
rect 16868 14269 16896 14368
rect 17954 14356 17960 14408
rect 18012 14396 18018 14408
rect 18708 14396 18736 14427
rect 19242 14424 19248 14476
rect 19300 14464 19306 14476
rect 20073 14467 20131 14473
rect 20073 14464 20085 14467
rect 19300 14436 20085 14464
rect 19300 14424 19306 14436
rect 20073 14433 20085 14436
rect 20119 14433 20131 14467
rect 20073 14427 20131 14433
rect 20714 14424 20720 14476
rect 20772 14464 20778 14476
rect 21085 14467 21143 14473
rect 21085 14464 21097 14467
rect 20772 14436 21097 14464
rect 20772 14424 20778 14436
rect 21085 14433 21097 14436
rect 21131 14433 21143 14467
rect 21085 14427 21143 14433
rect 21358 14424 21364 14476
rect 21416 14424 21422 14476
rect 21450 14424 21456 14476
rect 21508 14464 21514 14476
rect 24394 14464 24400 14476
rect 21508 14436 24400 14464
rect 21508 14424 21514 14436
rect 24394 14424 24400 14436
rect 24452 14424 24458 14476
rect 25406 14424 25412 14476
rect 25464 14464 25470 14476
rect 26789 14467 26847 14473
rect 26789 14464 26801 14467
rect 25464 14436 26801 14464
rect 25464 14424 25470 14436
rect 26789 14433 26801 14436
rect 26835 14433 26847 14467
rect 26789 14427 26847 14433
rect 28258 14424 28264 14476
rect 28316 14424 28322 14476
rect 28445 14467 28503 14473
rect 28445 14433 28457 14467
rect 28491 14464 28503 14467
rect 28810 14464 28816 14476
rect 28491 14436 28816 14464
rect 28491 14433 28503 14436
rect 28445 14427 28503 14433
rect 28810 14424 28816 14436
rect 28868 14424 28874 14476
rect 18012 14368 18736 14396
rect 18012 14356 18018 14368
rect 19886 14356 19892 14408
rect 19944 14396 19950 14408
rect 19981 14399 20039 14405
rect 19981 14396 19993 14399
rect 19944 14368 19993 14396
rect 19944 14356 19950 14368
rect 19981 14365 19993 14368
rect 20027 14396 20039 14399
rect 20622 14396 20628 14408
rect 20027 14368 20628 14396
rect 20027 14365 20039 14368
rect 19981 14359 20039 14365
rect 20622 14356 20628 14368
rect 20680 14396 20686 14408
rect 20809 14399 20867 14405
rect 20809 14396 20821 14399
rect 20680 14368 20821 14396
rect 20680 14356 20686 14368
rect 20809 14365 20821 14368
rect 20855 14365 20867 14399
rect 20809 14359 20867 14365
rect 24946 14356 24952 14408
rect 25004 14356 25010 14408
rect 25041 14399 25099 14405
rect 25041 14365 25053 14399
rect 25087 14365 25099 14399
rect 25041 14359 25099 14365
rect 18598 14328 18604 14340
rect 17604 14300 18604 14328
rect 16853 14263 16911 14269
rect 16853 14260 16865 14263
rect 16816 14232 16865 14260
rect 16816 14220 16822 14232
rect 16853 14229 16865 14232
rect 16899 14229 16911 14263
rect 16853 14223 16911 14229
rect 17402 14220 17408 14272
rect 17460 14260 17466 14272
rect 17604 14269 17632 14300
rect 18598 14288 18604 14300
rect 18656 14288 18662 14340
rect 19334 14288 19340 14340
rect 19392 14328 19398 14340
rect 19794 14328 19800 14340
rect 19392 14300 19800 14328
rect 19392 14288 19398 14300
rect 19794 14288 19800 14300
rect 19852 14328 19858 14340
rect 21450 14328 21456 14340
rect 19852 14300 21456 14328
rect 19852 14288 19858 14300
rect 21450 14288 21456 14300
rect 21508 14288 21514 14340
rect 22738 14328 22744 14340
rect 22586 14300 22744 14328
rect 22738 14288 22744 14300
rect 22796 14328 22802 14340
rect 23566 14328 23572 14340
rect 22796 14300 23572 14328
rect 22796 14288 22802 14300
rect 23566 14288 23572 14300
rect 23624 14288 23630 14340
rect 24854 14288 24860 14340
rect 24912 14328 24918 14340
rect 25056 14328 25084 14359
rect 27706 14356 27712 14408
rect 27764 14396 27770 14408
rect 28169 14399 28227 14405
rect 28169 14396 28181 14399
rect 27764 14368 28181 14396
rect 27764 14356 27770 14368
rect 28169 14365 28181 14368
rect 28215 14365 28227 14399
rect 28169 14359 28227 14365
rect 30006 14356 30012 14408
rect 30064 14396 30070 14408
rect 30101 14399 30159 14405
rect 30101 14396 30113 14399
rect 30064 14368 30113 14396
rect 30064 14356 30070 14368
rect 30101 14365 30113 14368
rect 30147 14365 30159 14399
rect 30208 14396 30236 14504
rect 30374 14492 30380 14544
rect 30432 14532 30438 14544
rect 31662 14532 31668 14544
rect 30432 14504 31668 14532
rect 30432 14492 30438 14504
rect 31662 14492 31668 14504
rect 31720 14492 31726 14544
rect 34054 14532 34060 14544
rect 32140 14504 34060 14532
rect 30282 14424 30288 14476
rect 30340 14424 30346 14476
rect 31294 14424 31300 14476
rect 31352 14464 31358 14476
rect 31573 14467 31631 14473
rect 31573 14464 31585 14467
rect 31352 14436 31585 14464
rect 31352 14424 31358 14436
rect 31573 14433 31585 14436
rect 31619 14433 31631 14467
rect 31573 14427 31631 14433
rect 30208 14368 30328 14396
rect 30101 14359 30159 14365
rect 24912 14300 25084 14328
rect 24912 14288 24918 14300
rect 17589 14263 17647 14269
rect 17589 14260 17601 14263
rect 17460 14232 17601 14260
rect 17460 14220 17466 14232
rect 17589 14229 17601 14232
rect 17635 14229 17647 14263
rect 17589 14223 17647 14229
rect 18509 14263 18567 14269
rect 18509 14229 18521 14263
rect 18555 14260 18567 14263
rect 18690 14260 18696 14272
rect 18555 14232 18696 14260
rect 18555 14229 18567 14232
rect 18509 14223 18567 14229
rect 18690 14220 18696 14232
rect 18748 14220 18754 14272
rect 19518 14220 19524 14272
rect 19576 14220 19582 14272
rect 19702 14220 19708 14272
rect 19760 14260 19766 14272
rect 19889 14263 19947 14269
rect 19889 14260 19901 14263
rect 19760 14232 19901 14260
rect 19760 14220 19766 14232
rect 19889 14229 19901 14232
rect 19935 14229 19947 14263
rect 25056 14260 25084 14300
rect 25317 14331 25375 14337
rect 25317 14297 25329 14331
rect 25363 14328 25375 14331
rect 25590 14328 25596 14340
rect 25363 14300 25596 14328
rect 25363 14297 25375 14300
rect 25317 14291 25375 14297
rect 25590 14288 25596 14300
rect 25648 14288 25654 14340
rect 25774 14288 25780 14340
rect 25832 14288 25838 14340
rect 30193 14331 30251 14337
rect 30193 14328 30205 14331
rect 27816 14300 30205 14328
rect 26694 14260 26700 14272
rect 25056 14232 26700 14260
rect 19889 14223 19947 14229
rect 26694 14220 26700 14232
rect 26752 14220 26758 14272
rect 27816 14269 27844 14300
rect 30193 14297 30205 14300
rect 30239 14297 30251 14331
rect 30300 14328 30328 14368
rect 30926 14356 30932 14408
rect 30984 14396 30990 14408
rect 31110 14396 31116 14408
rect 30984 14368 31116 14396
rect 30984 14356 30990 14368
rect 31110 14356 31116 14368
rect 31168 14396 31174 14408
rect 32140 14396 32168 14504
rect 34054 14492 34060 14504
rect 34112 14492 34118 14544
rect 32306 14424 32312 14476
rect 32364 14464 32370 14476
rect 32677 14467 32735 14473
rect 32677 14464 32689 14467
rect 32364 14436 32689 14464
rect 32364 14424 32370 14436
rect 32677 14433 32689 14436
rect 32723 14433 32735 14467
rect 32677 14427 32735 14433
rect 32858 14424 32864 14476
rect 32916 14424 32922 14476
rect 33410 14424 33416 14476
rect 33468 14464 33474 14476
rect 33594 14464 33600 14476
rect 33468 14436 33600 14464
rect 33468 14424 33474 14436
rect 33594 14424 33600 14436
rect 33652 14424 33658 14476
rect 33965 14467 34023 14473
rect 33965 14433 33977 14467
rect 34011 14464 34023 14467
rect 34808 14464 34836 14572
rect 35342 14560 35348 14572
rect 35400 14560 35406 14612
rect 35802 14560 35808 14612
rect 35860 14600 35866 14612
rect 36633 14603 36691 14609
rect 35860 14572 36584 14600
rect 35860 14560 35866 14572
rect 36556 14532 36584 14572
rect 36633 14569 36645 14603
rect 36679 14600 36691 14603
rect 36814 14600 36820 14612
rect 36679 14572 36820 14600
rect 36679 14569 36691 14572
rect 36633 14563 36691 14569
rect 36814 14560 36820 14572
rect 36872 14560 36878 14612
rect 37200 14572 39528 14600
rect 37200 14532 37228 14572
rect 36556 14504 37228 14532
rect 38841 14535 38899 14541
rect 38841 14501 38853 14535
rect 38887 14532 38899 14535
rect 39298 14532 39304 14544
rect 38887 14504 39304 14532
rect 38887 14501 38899 14504
rect 38841 14495 38899 14501
rect 39298 14492 39304 14504
rect 39356 14492 39362 14544
rect 34011 14436 34836 14464
rect 34011 14433 34023 14436
rect 33965 14427 34023 14433
rect 34882 14424 34888 14476
rect 34940 14464 34946 14476
rect 37090 14464 37096 14476
rect 34940 14436 37096 14464
rect 34940 14424 34946 14436
rect 37090 14424 37096 14436
rect 37148 14424 37154 14476
rect 37369 14467 37427 14473
rect 37369 14433 37381 14467
rect 37415 14464 37427 14467
rect 38102 14464 38108 14476
rect 37415 14436 38108 14464
rect 37415 14433 37427 14436
rect 37369 14427 37427 14433
rect 38102 14424 38108 14436
rect 38160 14424 38166 14476
rect 31168 14368 32168 14396
rect 31168 14356 31174 14368
rect 32214 14356 32220 14408
rect 32272 14396 32278 14408
rect 39500 14405 39528 14572
rect 33873 14399 33931 14405
rect 33873 14396 33885 14399
rect 32272 14368 33885 14396
rect 32272 14356 32278 14368
rect 33873 14365 33885 14368
rect 33919 14365 33931 14399
rect 33873 14359 33931 14365
rect 39485 14399 39543 14405
rect 39485 14365 39497 14399
rect 39531 14365 39543 14399
rect 39485 14359 39543 14365
rect 49050 14356 49056 14408
rect 49108 14356 49114 14408
rect 31389 14331 31447 14337
rect 30300 14300 31156 14328
rect 30193 14291 30251 14297
rect 27801 14263 27859 14269
rect 27801 14229 27813 14263
rect 27847 14229 27859 14263
rect 27801 14223 27859 14229
rect 31018 14220 31024 14272
rect 31076 14220 31082 14272
rect 31128 14260 31156 14300
rect 31389 14297 31401 14331
rect 31435 14328 31447 14331
rect 31435 14300 31616 14328
rect 31435 14297 31447 14300
rect 31389 14291 31447 14297
rect 31481 14263 31539 14269
rect 31481 14260 31493 14263
rect 31128 14232 31493 14260
rect 31481 14229 31493 14232
rect 31527 14229 31539 14263
rect 31588 14260 31616 14300
rect 31662 14288 31668 14340
rect 31720 14328 31726 14340
rect 32585 14331 32643 14337
rect 32585 14328 32597 14331
rect 31720 14300 32597 14328
rect 31720 14288 31726 14300
rect 32585 14297 32597 14300
rect 32631 14297 32643 14331
rect 32585 14291 32643 14297
rect 33778 14288 33784 14340
rect 33836 14288 33842 14340
rect 34514 14288 34520 14340
rect 34572 14328 34578 14340
rect 35161 14331 35219 14337
rect 35161 14328 35173 14331
rect 34572 14300 35173 14328
rect 34572 14288 34578 14300
rect 35161 14297 35173 14300
rect 35207 14328 35219 14331
rect 35250 14328 35256 14340
rect 35207 14300 35256 14328
rect 35207 14297 35219 14300
rect 35161 14291 35219 14297
rect 35250 14288 35256 14300
rect 35308 14288 35314 14340
rect 36538 14328 36544 14340
rect 36386 14300 36544 14328
rect 36538 14288 36544 14300
rect 36596 14288 36602 14340
rect 37826 14328 37832 14340
rect 37476 14300 37832 14328
rect 32030 14260 32036 14272
rect 31588 14232 32036 14260
rect 31481 14223 31539 14229
rect 32030 14220 32036 14232
rect 32088 14220 32094 14272
rect 32217 14263 32275 14269
rect 32217 14229 32229 14263
rect 32263 14260 32275 14263
rect 32490 14260 32496 14272
rect 32263 14232 32496 14260
rect 32263 14229 32275 14232
rect 32217 14223 32275 14229
rect 32490 14220 32496 14232
rect 32548 14220 32554 14272
rect 32674 14220 32680 14272
rect 32732 14260 32738 14272
rect 34238 14260 34244 14272
rect 32732 14232 34244 14260
rect 32732 14220 32738 14232
rect 34238 14220 34244 14232
rect 34296 14220 34302 14272
rect 36556 14260 36584 14288
rect 37476 14260 37504 14300
rect 37826 14288 37832 14300
rect 37884 14288 37890 14340
rect 36556 14232 37504 14260
rect 39301 14263 39359 14269
rect 39301 14229 39313 14263
rect 39347 14260 39359 14263
rect 45002 14260 45008 14272
rect 39347 14232 45008 14260
rect 39347 14229 39359 14232
rect 39301 14223 39359 14229
rect 45002 14220 45008 14232
rect 45060 14220 45066 14272
rect 49234 14220 49240 14272
rect 49292 14220 49298 14272
rect 1104 14170 49864 14192
rect 1104 14118 7950 14170
rect 8002 14118 8014 14170
rect 8066 14118 8078 14170
rect 8130 14118 8142 14170
rect 8194 14118 8206 14170
rect 8258 14118 17950 14170
rect 18002 14118 18014 14170
rect 18066 14118 18078 14170
rect 18130 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 27950 14170
rect 28002 14118 28014 14170
rect 28066 14118 28078 14170
rect 28130 14118 28142 14170
rect 28194 14118 28206 14170
rect 28258 14118 37950 14170
rect 38002 14118 38014 14170
rect 38066 14118 38078 14170
rect 38130 14118 38142 14170
rect 38194 14118 38206 14170
rect 38258 14118 47950 14170
rect 48002 14118 48014 14170
rect 48066 14118 48078 14170
rect 48130 14118 48142 14170
rect 48194 14118 48206 14170
rect 48258 14118 49864 14170
rect 1104 14096 49864 14118
rect 3602 14016 3608 14068
rect 3660 14016 3666 14068
rect 11701 14059 11759 14065
rect 11701 14025 11713 14059
rect 11747 14056 11759 14059
rect 11974 14056 11980 14068
rect 11747 14028 11980 14056
rect 11747 14025 11759 14028
rect 11701 14019 11759 14025
rect 11974 14016 11980 14028
rect 12032 14016 12038 14068
rect 14550 14016 14556 14068
rect 14608 14056 14614 14068
rect 14645 14059 14703 14065
rect 14645 14056 14657 14059
rect 14608 14028 14657 14056
rect 14608 14016 14614 14028
rect 14645 14025 14657 14028
rect 14691 14025 14703 14059
rect 14645 14019 14703 14025
rect 15286 14016 15292 14068
rect 15344 14056 15350 14068
rect 15565 14059 15623 14065
rect 15565 14056 15577 14059
rect 15344 14028 15577 14056
rect 15344 14016 15350 14028
rect 15565 14025 15577 14028
rect 15611 14025 15623 14059
rect 15565 14019 15623 14025
rect 15930 14016 15936 14068
rect 15988 14016 15994 14068
rect 16758 14016 16764 14068
rect 16816 14056 16822 14068
rect 17129 14059 17187 14065
rect 17129 14056 17141 14059
rect 16816 14028 17141 14056
rect 16816 14016 16822 14028
rect 17129 14025 17141 14028
rect 17175 14025 17187 14059
rect 17129 14019 17187 14025
rect 17494 14016 17500 14068
rect 17552 14016 17558 14068
rect 17586 14016 17592 14068
rect 17644 14016 17650 14068
rect 17862 14016 17868 14068
rect 17920 14056 17926 14068
rect 18325 14059 18383 14065
rect 18325 14056 18337 14059
rect 17920 14028 18337 14056
rect 17920 14016 17926 14028
rect 18325 14025 18337 14028
rect 18371 14025 18383 14059
rect 18325 14019 18383 14025
rect 18693 14059 18751 14065
rect 18693 14025 18705 14059
rect 18739 14056 18751 14059
rect 19610 14056 19616 14068
rect 18739 14028 19616 14056
rect 18739 14025 18751 14028
rect 18693 14019 18751 14025
rect 19610 14016 19616 14028
rect 19668 14016 19674 14068
rect 21358 14016 21364 14068
rect 21416 14056 21422 14068
rect 21453 14059 21511 14065
rect 21453 14056 21465 14059
rect 21416 14028 21465 14056
rect 21416 14016 21422 14028
rect 21453 14025 21465 14028
rect 21499 14025 21511 14059
rect 21453 14019 21511 14025
rect 21634 14016 21640 14068
rect 21692 14056 21698 14068
rect 26050 14056 26056 14068
rect 21692 14028 26056 14056
rect 21692 14016 21698 14028
rect 26050 14016 26056 14028
rect 26108 14016 26114 14068
rect 26418 14016 26424 14068
rect 26476 14056 26482 14068
rect 26605 14059 26663 14065
rect 26605 14056 26617 14059
rect 26476 14028 26617 14056
rect 26476 14016 26482 14028
rect 26605 14025 26617 14028
rect 26651 14025 26663 14059
rect 26605 14019 26663 14025
rect 27614 14016 27620 14068
rect 27672 14056 27678 14068
rect 31113 14059 31171 14065
rect 31113 14056 31125 14059
rect 27672 14028 31125 14056
rect 27672 14016 27678 14028
rect 31113 14025 31125 14028
rect 31159 14025 31171 14059
rect 31113 14019 31171 14025
rect 31294 14016 31300 14068
rect 31352 14056 31358 14068
rect 31662 14056 31668 14068
rect 31352 14028 31668 14056
rect 31352 14016 31358 14028
rect 31662 14016 31668 14028
rect 31720 14016 31726 14068
rect 31772 14028 33916 14056
rect 11238 13988 11244 14000
rect 2746 13960 11244 13988
rect 1765 13923 1823 13929
rect 1765 13889 1777 13923
rect 1811 13920 1823 13923
rect 2746 13920 2774 13960
rect 11238 13948 11244 13960
rect 11296 13948 11302 14000
rect 14182 13948 14188 14000
rect 14240 13948 14246 14000
rect 16025 13991 16083 13997
rect 16025 13957 16037 13991
rect 16071 13988 16083 13991
rect 19518 13988 19524 14000
rect 16071 13960 19524 13988
rect 16071 13957 16083 13960
rect 16025 13951 16083 13957
rect 19518 13948 19524 13960
rect 19576 13948 19582 14000
rect 19981 13991 20039 13997
rect 19981 13957 19993 13991
rect 20027 13988 20039 13991
rect 20070 13988 20076 14000
rect 20027 13960 20076 13988
rect 20027 13957 20039 13960
rect 19981 13951 20039 13957
rect 20070 13948 20076 13960
rect 20128 13948 20134 14000
rect 22738 13988 22744 14000
rect 21206 13960 22744 13988
rect 22738 13948 22744 13960
rect 22796 13948 22802 14000
rect 23566 13988 23572 14000
rect 23506 13960 23572 13988
rect 23566 13948 23572 13960
rect 23624 13988 23630 14000
rect 24670 13988 24676 14000
rect 23624 13960 24676 13988
rect 23624 13948 23630 13960
rect 24670 13948 24676 13960
rect 24728 13948 24734 14000
rect 25133 13991 25191 13997
rect 25133 13957 25145 13991
rect 25179 13988 25191 13991
rect 25222 13988 25228 14000
rect 25179 13960 25228 13988
rect 25179 13957 25191 13960
rect 25133 13951 25191 13957
rect 25222 13948 25228 13960
rect 25280 13988 25286 14000
rect 25406 13988 25412 14000
rect 25280 13960 25412 13988
rect 25280 13948 25286 13960
rect 25406 13948 25412 13960
rect 25464 13948 25470 14000
rect 25774 13948 25780 14000
rect 25832 13948 25838 14000
rect 26694 13948 26700 14000
rect 26752 13988 26758 14000
rect 26752 13960 29408 13988
rect 26752 13948 26758 13960
rect 1811 13892 2774 13920
rect 1811 13889 1823 13892
rect 1765 13883 1823 13889
rect 3510 13880 3516 13932
rect 3568 13880 3574 13932
rect 11149 13923 11207 13929
rect 11149 13889 11161 13923
rect 11195 13920 11207 13923
rect 12069 13923 12127 13929
rect 12069 13920 12081 13923
rect 11195 13892 12081 13920
rect 11195 13889 11207 13892
rect 11149 13883 11207 13889
rect 12069 13889 12081 13892
rect 12115 13889 12127 13923
rect 12069 13883 12127 13889
rect 18785 13923 18843 13929
rect 18785 13889 18797 13923
rect 18831 13920 18843 13923
rect 19334 13920 19340 13932
rect 18831 13892 19340 13920
rect 18831 13889 18843 13892
rect 18785 13883 18843 13889
rect 19334 13880 19340 13892
rect 19392 13880 19398 13932
rect 24854 13880 24860 13932
rect 24912 13880 24918 13932
rect 27154 13880 27160 13932
rect 27212 13880 27218 13932
rect 29380 13929 29408 13960
rect 30650 13948 30656 14000
rect 30708 13948 30714 14000
rect 31772 13929 31800 14028
rect 32030 13948 32036 14000
rect 32088 13988 32094 14000
rect 32674 13988 32680 14000
rect 32088 13960 32680 13988
rect 32088 13948 32094 13960
rect 32674 13948 32680 13960
rect 32732 13948 32738 14000
rect 33888 13988 33916 14028
rect 34054 14016 34060 14068
rect 34112 14016 34118 14068
rect 34790 14016 34796 14068
rect 34848 14056 34854 14068
rect 34885 14059 34943 14065
rect 34885 14056 34897 14059
rect 34848 14028 34897 14056
rect 34848 14016 34854 14028
rect 34885 14025 34897 14028
rect 34931 14025 34943 14059
rect 34885 14019 34943 14025
rect 35713 14059 35771 14065
rect 35713 14025 35725 14059
rect 35759 14056 35771 14059
rect 37829 14059 37887 14065
rect 37829 14056 37841 14059
rect 35759 14028 37841 14056
rect 35759 14025 35771 14028
rect 35713 14019 35771 14025
rect 37829 14025 37841 14028
rect 37875 14025 37887 14059
rect 41506 14056 41512 14068
rect 37829 14019 37887 14025
rect 41386 14028 41512 14056
rect 36081 13991 36139 13997
rect 36081 13988 36093 13991
rect 33888 13960 36093 13988
rect 36081 13957 36093 13960
rect 36127 13957 36139 13991
rect 36081 13951 36139 13957
rect 36262 13948 36268 14000
rect 36320 13988 36326 14000
rect 37921 13991 37979 13997
rect 37921 13988 37933 13991
rect 36320 13960 37933 13988
rect 36320 13948 36326 13960
rect 37921 13957 37933 13960
rect 37967 13957 37979 13991
rect 37921 13951 37979 13957
rect 29365 13923 29423 13929
rect 29365 13889 29377 13923
rect 29411 13889 29423 13923
rect 29365 13883 29423 13889
rect 31757 13923 31815 13929
rect 31757 13889 31769 13923
rect 31803 13889 31815 13923
rect 31757 13883 31815 13889
rect 33686 13880 33692 13932
rect 33744 13920 33750 13932
rect 34422 13920 34428 13932
rect 33744 13892 34428 13920
rect 33744 13880 33750 13892
rect 34422 13880 34428 13892
rect 34480 13880 34486 13932
rect 37366 13920 37372 13932
rect 34532 13892 37372 13920
rect 1302 13812 1308 13864
rect 1360 13852 1366 13864
rect 2041 13855 2099 13861
rect 2041 13852 2053 13855
rect 1360 13824 2053 13852
rect 1360 13812 1366 13824
rect 2041 13821 2053 13824
rect 2087 13821 2099 13855
rect 2041 13815 2099 13821
rect 11790 13812 11796 13864
rect 11848 13852 11854 13864
rect 12161 13855 12219 13861
rect 12161 13852 12173 13855
rect 11848 13824 12173 13852
rect 11848 13812 11854 13824
rect 12161 13821 12173 13824
rect 12207 13821 12219 13855
rect 12161 13815 12219 13821
rect 12345 13855 12403 13861
rect 12345 13821 12357 13855
rect 12391 13821 12403 13855
rect 12345 13815 12403 13821
rect 12360 13784 12388 13815
rect 12802 13812 12808 13864
rect 12860 13852 12866 13864
rect 12897 13855 12955 13861
rect 12897 13852 12909 13855
rect 12860 13824 12909 13852
rect 12860 13812 12866 13824
rect 12897 13821 12909 13824
rect 12943 13821 12955 13855
rect 12897 13815 12955 13821
rect 13170 13812 13176 13864
rect 13228 13852 13234 13864
rect 13630 13852 13636 13864
rect 13228 13824 13636 13852
rect 13228 13812 13234 13824
rect 13630 13812 13636 13824
rect 13688 13812 13694 13864
rect 16117 13855 16175 13861
rect 16117 13821 16129 13855
rect 16163 13821 16175 13855
rect 16117 13815 16175 13821
rect 12434 13784 12440 13796
rect 12360 13756 12440 13784
rect 12434 13744 12440 13756
rect 12492 13744 12498 13796
rect 16132 13784 16160 13815
rect 16574 13812 16580 13864
rect 16632 13852 16638 13864
rect 17310 13852 17316 13864
rect 16632 13824 17316 13852
rect 16632 13812 16638 13824
rect 17310 13812 17316 13824
rect 17368 13812 17374 13864
rect 17773 13855 17831 13861
rect 17773 13821 17785 13855
rect 17819 13821 17831 13855
rect 17773 13815 17831 13821
rect 18877 13855 18935 13861
rect 18877 13821 18889 13855
rect 18923 13821 18935 13855
rect 18877 13815 18935 13821
rect 16040 13756 16160 13784
rect 12894 13676 12900 13728
rect 12952 13716 12958 13728
rect 15930 13716 15936 13728
rect 12952 13688 15936 13716
rect 12952 13676 12958 13688
rect 15930 13676 15936 13688
rect 15988 13716 15994 13728
rect 16040 13716 16068 13756
rect 17678 13744 17684 13796
rect 17736 13784 17742 13796
rect 17788 13784 17816 13815
rect 17736 13756 17816 13784
rect 17736 13744 17742 13756
rect 18506 13744 18512 13796
rect 18564 13784 18570 13796
rect 18892 13784 18920 13815
rect 18966 13812 18972 13864
rect 19024 13852 19030 13864
rect 19705 13855 19763 13861
rect 19705 13852 19717 13855
rect 19024 13824 19717 13852
rect 19024 13812 19030 13824
rect 19705 13821 19717 13824
rect 19751 13821 19763 13855
rect 19705 13815 19763 13821
rect 19812 13824 21036 13852
rect 18564 13756 18920 13784
rect 18564 13744 18570 13756
rect 15988 13688 16068 13716
rect 15988 13676 15994 13688
rect 16482 13676 16488 13728
rect 16540 13716 16546 13728
rect 19812 13716 19840 13824
rect 16540 13688 19840 13716
rect 21008 13716 21036 13824
rect 22002 13812 22008 13864
rect 22060 13812 22066 13864
rect 22278 13812 22284 13864
rect 22336 13812 22342 13864
rect 23658 13812 23664 13864
rect 23716 13852 23722 13864
rect 24397 13855 24455 13861
rect 24397 13852 24409 13855
rect 23716 13824 24409 13852
rect 23716 13812 23722 13824
rect 24397 13821 24409 13824
rect 24443 13821 24455 13855
rect 24397 13815 24455 13821
rect 25498 13812 25504 13864
rect 25556 13852 25562 13864
rect 27614 13852 27620 13864
rect 25556 13824 27620 13852
rect 25556 13812 25562 13824
rect 27614 13812 27620 13824
rect 27672 13812 27678 13864
rect 28902 13812 28908 13864
rect 28960 13812 28966 13864
rect 30834 13812 30840 13864
rect 30892 13852 30898 13864
rect 32214 13852 32220 13864
rect 30892 13824 32220 13852
rect 30892 13812 30898 13824
rect 32214 13812 32220 13824
rect 32272 13812 32278 13864
rect 32309 13855 32367 13861
rect 32309 13821 32321 13855
rect 32355 13821 32367 13855
rect 32309 13815 32367 13821
rect 23750 13744 23756 13796
rect 23808 13744 23814 13796
rect 31754 13744 31760 13796
rect 31812 13784 31818 13796
rect 32324 13784 32352 13815
rect 32582 13812 32588 13864
rect 32640 13812 32646 13864
rect 32674 13812 32680 13864
rect 32732 13852 32738 13864
rect 33594 13852 33600 13864
rect 32732 13824 33600 13852
rect 32732 13812 32738 13824
rect 33594 13812 33600 13824
rect 33652 13812 33658 13864
rect 34532 13793 34560 13892
rect 37366 13880 37372 13892
rect 37424 13880 37430 13932
rect 41386 13920 41414 14028
rect 41506 14016 41512 14028
rect 41564 14016 41570 14068
rect 45649 14059 45707 14065
rect 45649 14025 45661 14059
rect 45695 14056 45707 14059
rect 47026 14056 47032 14068
rect 45695 14028 47032 14056
rect 45695 14025 45707 14028
rect 45649 14019 45707 14025
rect 47026 14016 47032 14028
rect 47084 14016 47090 14068
rect 48406 14016 48412 14068
rect 48464 14016 48470 14068
rect 48498 14016 48504 14068
rect 48556 14056 48562 14068
rect 49237 14059 49295 14065
rect 49237 14056 49249 14059
rect 48556 14028 49249 14056
rect 48556 14016 48562 14028
rect 49237 14025 49249 14028
rect 49283 14025 49295 14059
rect 49237 14019 49295 14025
rect 45002 13948 45008 14000
rect 45060 13948 45066 14000
rect 46842 13948 46848 14000
rect 46900 13988 46906 14000
rect 48682 13988 48688 14000
rect 46900 13960 48688 13988
rect 46900 13948 46906 13960
rect 48682 13948 48688 13960
rect 48740 13948 48746 14000
rect 49142 13948 49148 14000
rect 49200 13948 49206 14000
rect 37476 13892 41414 13920
rect 34698 13812 34704 13864
rect 34756 13852 34762 13864
rect 34977 13855 35035 13861
rect 34977 13852 34989 13855
rect 34756 13824 34989 13852
rect 34756 13812 34762 13824
rect 34977 13821 34989 13824
rect 35023 13821 35035 13855
rect 34977 13815 35035 13821
rect 35069 13855 35127 13861
rect 35069 13821 35081 13855
rect 35115 13821 35127 13855
rect 35069 13815 35127 13821
rect 31812 13756 32352 13784
rect 34517 13787 34575 13793
rect 31812 13744 31818 13756
rect 34517 13753 34529 13787
rect 34563 13753 34575 13787
rect 34517 13747 34575 13753
rect 35084 13728 35112 13815
rect 35986 13812 35992 13864
rect 36044 13852 36050 13864
rect 36173 13855 36231 13861
rect 36173 13852 36185 13855
rect 36044 13824 36185 13852
rect 36044 13812 36050 13824
rect 36173 13821 36185 13824
rect 36219 13821 36231 13855
rect 36173 13815 36231 13821
rect 36357 13855 36415 13861
rect 36357 13821 36369 13855
rect 36403 13852 36415 13855
rect 36630 13852 36636 13864
rect 36403 13824 36636 13852
rect 36403 13821 36415 13824
rect 36357 13815 36415 13821
rect 36630 13812 36636 13824
rect 36688 13852 36694 13864
rect 36814 13852 36820 13864
rect 36688 13824 36820 13852
rect 36688 13812 36694 13824
rect 36814 13812 36820 13824
rect 36872 13812 36878 13864
rect 37476 13793 37504 13892
rect 45830 13880 45836 13932
rect 45888 13880 45894 13932
rect 48222 13880 48228 13932
rect 48280 13920 48286 13932
rect 48593 13923 48651 13929
rect 48593 13920 48605 13923
rect 48280 13892 48605 13920
rect 48280 13880 48286 13892
rect 48593 13889 48605 13892
rect 48639 13889 48651 13923
rect 48593 13883 48651 13889
rect 38013 13855 38071 13861
rect 38013 13821 38025 13855
rect 38059 13821 38071 13855
rect 38013 13815 38071 13821
rect 45189 13855 45247 13861
rect 45189 13821 45201 13855
rect 45235 13852 45247 13855
rect 46290 13852 46296 13864
rect 45235 13824 46296 13852
rect 45235 13821 45247 13824
rect 45189 13815 45247 13821
rect 37461 13787 37519 13793
rect 37461 13753 37473 13787
rect 37507 13753 37519 13787
rect 37461 13747 37519 13753
rect 37826 13744 37832 13796
rect 37884 13784 37890 13796
rect 38028 13784 38056 13815
rect 46290 13812 46296 13824
rect 46348 13812 46354 13864
rect 37884 13756 38056 13784
rect 37884 13744 37890 13756
rect 22830 13716 22836 13728
rect 21008 13688 22836 13716
rect 16540 13676 16546 13688
rect 22830 13676 22836 13688
rect 22888 13676 22894 13728
rect 23934 13676 23940 13728
rect 23992 13716 23998 13728
rect 26234 13716 26240 13728
rect 23992 13688 26240 13716
rect 23992 13676 23998 13688
rect 26234 13676 26240 13688
rect 26292 13676 26298 13728
rect 29628 13719 29686 13725
rect 29628 13685 29640 13719
rect 29674 13716 29686 13719
rect 30926 13716 30932 13728
rect 29674 13688 30932 13716
rect 29674 13685 29686 13688
rect 29628 13679 29686 13685
rect 30926 13676 30932 13688
rect 30984 13676 30990 13728
rect 31110 13676 31116 13728
rect 31168 13716 31174 13728
rect 34790 13716 34796 13728
rect 31168 13688 34796 13716
rect 31168 13676 31174 13688
rect 34790 13676 34796 13688
rect 34848 13676 34854 13728
rect 35066 13676 35072 13728
rect 35124 13676 35130 13728
rect 35526 13676 35532 13728
rect 35584 13716 35590 13728
rect 37550 13716 37556 13728
rect 35584 13688 37556 13716
rect 35584 13676 35590 13688
rect 37550 13676 37556 13688
rect 37608 13676 37614 13728
rect 38838 13676 38844 13728
rect 38896 13676 38902 13728
rect 1104 13626 49864 13648
rect 1104 13574 2950 13626
rect 3002 13574 3014 13626
rect 3066 13574 3078 13626
rect 3130 13574 3142 13626
rect 3194 13574 3206 13626
rect 3258 13574 12950 13626
rect 13002 13574 13014 13626
rect 13066 13574 13078 13626
rect 13130 13574 13142 13626
rect 13194 13574 13206 13626
rect 13258 13574 22950 13626
rect 23002 13574 23014 13626
rect 23066 13574 23078 13626
rect 23130 13574 23142 13626
rect 23194 13574 23206 13626
rect 23258 13574 32950 13626
rect 33002 13574 33014 13626
rect 33066 13574 33078 13626
rect 33130 13574 33142 13626
rect 33194 13574 33206 13626
rect 33258 13574 42950 13626
rect 43002 13574 43014 13626
rect 43066 13574 43078 13626
rect 43130 13574 43142 13626
rect 43194 13574 43206 13626
rect 43258 13574 49864 13626
rect 1104 13552 49864 13574
rect 2746 13484 12434 13512
rect 2746 13376 2774 13484
rect 12406 13444 12434 13484
rect 12618 13472 12624 13524
rect 12676 13512 12682 13524
rect 13265 13515 13323 13521
rect 13265 13512 13277 13515
rect 12676 13484 13277 13512
rect 12676 13472 12682 13484
rect 13265 13481 13277 13484
rect 13311 13481 13323 13515
rect 17678 13512 17684 13524
rect 13265 13475 13323 13481
rect 15856 13484 17684 13512
rect 14553 13447 14611 13453
rect 14553 13444 14565 13447
rect 12406 13416 14565 13444
rect 14553 13413 14565 13416
rect 14599 13413 14611 13447
rect 14553 13407 14611 13413
rect 12802 13376 12808 13388
rect 1780 13348 2774 13376
rect 10796 13348 12808 13376
rect 1780 13317 1808 13348
rect 1765 13311 1823 13317
rect 1765 13277 1777 13311
rect 1811 13277 1823 13311
rect 1765 13271 1823 13277
rect 2774 13268 2780 13320
rect 2832 13268 2838 13320
rect 10502 13268 10508 13320
rect 10560 13308 10566 13320
rect 10796 13317 10824 13348
rect 12802 13336 12808 13348
rect 12860 13336 12866 13388
rect 15102 13376 15108 13388
rect 14384 13348 15108 13376
rect 10781 13311 10839 13317
rect 10781 13308 10793 13311
rect 10560 13280 10793 13308
rect 10560 13268 10566 13280
rect 10781 13277 10793 13280
rect 10827 13277 10839 13311
rect 10781 13271 10839 13277
rect 12158 13268 12164 13320
rect 12216 13268 12222 13320
rect 12894 13268 12900 13320
rect 12952 13308 12958 13320
rect 14384 13317 14412 13348
rect 15102 13336 15108 13348
rect 15160 13336 15166 13388
rect 15378 13336 15384 13388
rect 15436 13376 15442 13388
rect 15856 13385 15884 13484
rect 17678 13472 17684 13484
rect 17736 13512 17742 13524
rect 18141 13515 18199 13521
rect 18141 13512 18153 13515
rect 17736 13484 18153 13512
rect 17736 13472 17742 13484
rect 18141 13481 18153 13484
rect 18187 13481 18199 13515
rect 18141 13475 18199 13481
rect 20898 13472 20904 13524
rect 20956 13472 20962 13524
rect 22097 13515 22155 13521
rect 22097 13481 22109 13515
rect 22143 13512 22155 13515
rect 22186 13512 22192 13524
rect 22143 13484 22192 13512
rect 22143 13481 22155 13484
rect 22097 13475 22155 13481
rect 22186 13472 22192 13484
rect 22244 13472 22250 13524
rect 22830 13472 22836 13524
rect 22888 13512 22894 13524
rect 23293 13515 23351 13521
rect 23293 13512 23305 13515
rect 22888 13484 23305 13512
rect 22888 13472 22894 13484
rect 23293 13481 23305 13484
rect 23339 13481 23351 13515
rect 23293 13475 23351 13481
rect 24857 13515 24915 13521
rect 24857 13481 24869 13515
rect 24903 13512 24915 13515
rect 25314 13512 25320 13524
rect 24903 13484 25320 13512
rect 24903 13481 24915 13484
rect 24857 13475 24915 13481
rect 25314 13472 25320 13484
rect 25372 13472 25378 13524
rect 27798 13472 27804 13524
rect 27856 13512 27862 13524
rect 29733 13515 29791 13521
rect 27856 13484 28764 13512
rect 27856 13472 27862 13484
rect 26602 13444 26608 13456
rect 22572 13416 26608 13444
rect 15657 13379 15715 13385
rect 15657 13376 15669 13379
rect 15436 13348 15669 13376
rect 15436 13336 15442 13348
rect 15657 13345 15669 13348
rect 15703 13345 15715 13379
rect 15657 13339 15715 13345
rect 15841 13379 15899 13385
rect 15841 13345 15853 13379
rect 15887 13345 15899 13379
rect 15841 13339 15899 13345
rect 16393 13379 16451 13385
rect 16393 13345 16405 13379
rect 16439 13376 16451 13379
rect 18966 13376 18972 13388
rect 16439 13348 18972 13376
rect 16439 13345 16451 13348
rect 16393 13339 16451 13345
rect 14369 13311 14427 13317
rect 12952 13280 14228 13308
rect 12952 13268 12958 13280
rect 8570 13200 8576 13252
rect 8628 13240 8634 13252
rect 11054 13240 11060 13252
rect 8628 13212 11060 13240
rect 8628 13200 8634 13212
rect 11054 13200 11060 13212
rect 11112 13200 11118 13252
rect 14200 13240 14228 13280
rect 14369 13277 14381 13311
rect 14415 13277 14427 13311
rect 14369 13271 14427 13277
rect 14550 13268 14556 13320
rect 14608 13308 14614 13320
rect 16408 13308 16436 13339
rect 18966 13336 18972 13348
rect 19024 13336 19030 13388
rect 21450 13336 21456 13388
rect 21508 13376 21514 13388
rect 22462 13376 22468 13388
rect 21508 13348 22468 13376
rect 21508 13336 21514 13348
rect 22462 13336 22468 13348
rect 22520 13336 22526 13388
rect 22572 13385 22600 13416
rect 26602 13404 26608 13416
rect 26660 13404 26666 13456
rect 22557 13379 22615 13385
rect 22557 13345 22569 13379
rect 22603 13345 22615 13379
rect 22557 13339 22615 13345
rect 22741 13379 22799 13385
rect 22741 13345 22753 13379
rect 22787 13376 22799 13379
rect 23566 13376 23572 13388
rect 22787 13348 23572 13376
rect 22787 13345 22799 13348
rect 22741 13339 22799 13345
rect 23566 13336 23572 13348
rect 23624 13336 23630 13388
rect 23753 13379 23811 13385
rect 23753 13345 23765 13379
rect 23799 13376 23811 13379
rect 23842 13376 23848 13388
rect 23799 13348 23848 13376
rect 23799 13345 23811 13348
rect 23753 13339 23811 13345
rect 23842 13336 23848 13348
rect 23900 13336 23906 13388
rect 23937 13379 23995 13385
rect 23937 13345 23949 13379
rect 23983 13376 23995 13379
rect 24854 13376 24860 13388
rect 23983 13348 24860 13376
rect 23983 13345 23995 13348
rect 23937 13339 23995 13345
rect 24854 13336 24860 13348
rect 24912 13336 24918 13388
rect 25498 13336 25504 13388
rect 25556 13336 25562 13388
rect 26694 13336 26700 13388
rect 26752 13376 26758 13388
rect 26789 13379 26847 13385
rect 26789 13376 26801 13379
rect 26752 13348 26801 13376
rect 26752 13336 26758 13348
rect 26789 13345 26801 13348
rect 26835 13345 26847 13379
rect 26789 13339 26847 13345
rect 27065 13379 27123 13385
rect 27065 13345 27077 13379
rect 27111 13376 27123 13379
rect 28626 13376 28632 13388
rect 27111 13348 28632 13376
rect 27111 13345 27123 13348
rect 27065 13339 27123 13345
rect 28626 13336 28632 13348
rect 28684 13336 28690 13388
rect 28736 13376 28764 13484
rect 29733 13481 29745 13515
rect 29779 13512 29791 13515
rect 32030 13512 32036 13524
rect 29779 13484 32036 13512
rect 29779 13481 29791 13484
rect 29733 13475 29791 13481
rect 32030 13472 32036 13484
rect 32088 13472 32094 13524
rect 33321 13515 33379 13521
rect 33321 13481 33333 13515
rect 33367 13512 33379 13515
rect 33870 13512 33876 13524
rect 33367 13484 33876 13512
rect 33367 13481 33379 13484
rect 33321 13475 33379 13481
rect 33870 13472 33876 13484
rect 33928 13472 33934 13524
rect 34885 13515 34943 13521
rect 34885 13481 34897 13515
rect 34931 13512 34943 13515
rect 38378 13512 38384 13524
rect 34931 13484 38384 13512
rect 34931 13481 34943 13484
rect 34885 13475 34943 13481
rect 38378 13472 38384 13484
rect 38436 13472 38442 13524
rect 28994 13404 29000 13456
rect 29052 13444 29058 13456
rect 30098 13444 30104 13456
rect 29052 13416 30104 13444
rect 29052 13404 29058 13416
rect 30098 13404 30104 13416
rect 30156 13404 30162 13456
rect 33686 13444 33692 13456
rect 32876 13416 33692 13444
rect 28813 13379 28871 13385
rect 28813 13376 28825 13379
rect 28736 13348 28825 13376
rect 28813 13345 28825 13348
rect 28859 13345 28871 13379
rect 28813 13339 28871 13345
rect 29822 13336 29828 13388
rect 29880 13376 29886 13388
rect 30193 13379 30251 13385
rect 30193 13376 30205 13379
rect 29880 13348 30205 13376
rect 29880 13336 29886 13348
rect 30193 13345 30205 13348
rect 30239 13345 30251 13379
rect 30193 13339 30251 13345
rect 30282 13336 30288 13388
rect 30340 13336 30346 13388
rect 31021 13379 31079 13385
rect 31021 13345 31033 13379
rect 31067 13376 31079 13379
rect 31754 13376 31760 13388
rect 31067 13348 31760 13376
rect 31067 13345 31079 13348
rect 31021 13339 31079 13345
rect 31754 13336 31760 13348
rect 31812 13336 31818 13388
rect 31846 13336 31852 13388
rect 31904 13376 31910 13388
rect 32769 13379 32827 13385
rect 32769 13376 32781 13379
rect 31904 13348 32781 13376
rect 31904 13336 31910 13348
rect 32769 13345 32781 13348
rect 32815 13345 32827 13379
rect 32769 13339 32827 13345
rect 14608 13280 16436 13308
rect 18877 13311 18935 13317
rect 14608 13268 14614 13280
rect 14200 13212 15516 13240
rect 10778 13132 10784 13184
rect 10836 13172 10842 13184
rect 12434 13172 12440 13184
rect 10836 13144 12440 13172
rect 10836 13132 10842 13144
rect 12434 13132 12440 13144
rect 12492 13172 12498 13184
rect 12529 13175 12587 13181
rect 12529 13172 12541 13175
rect 12492 13144 12541 13172
rect 12492 13132 12498 13144
rect 12529 13141 12541 13144
rect 12575 13172 12587 13175
rect 14918 13172 14924 13184
rect 12575 13144 14924 13172
rect 12575 13141 12587 13144
rect 12529 13135 12587 13141
rect 14918 13132 14924 13144
rect 14976 13132 14982 13184
rect 15194 13132 15200 13184
rect 15252 13132 15258 13184
rect 15488 13172 15516 13212
rect 15562 13200 15568 13252
rect 15620 13200 15626 13252
rect 15654 13200 15660 13252
rect 15712 13240 15718 13252
rect 15838 13240 15844 13252
rect 15712 13212 15844 13240
rect 15712 13200 15718 13212
rect 15838 13200 15844 13212
rect 15896 13200 15902 13252
rect 16298 13200 16304 13252
rect 16356 13240 16362 13252
rect 16669 13243 16727 13249
rect 16669 13240 16681 13243
rect 16356 13212 16681 13240
rect 16356 13200 16362 13212
rect 16669 13209 16681 13212
rect 16715 13209 16727 13243
rect 16669 13203 16727 13209
rect 17402 13172 17408 13184
rect 15488 13144 17408 13172
rect 17402 13132 17408 13144
rect 17460 13132 17466 13184
rect 17586 13132 17592 13184
rect 17644 13172 17650 13184
rect 17788 13172 17816 13294
rect 18877 13277 18889 13311
rect 18923 13308 18935 13311
rect 20070 13308 20076 13320
rect 18923 13280 20076 13308
rect 18923 13277 18935 13280
rect 18877 13271 18935 13277
rect 20070 13268 20076 13280
rect 20128 13268 20134 13320
rect 21266 13268 21272 13320
rect 21324 13308 21330 13320
rect 21634 13308 21640 13320
rect 21324 13280 21640 13308
rect 21324 13268 21330 13280
rect 21634 13268 21640 13280
rect 21692 13268 21698 13320
rect 23198 13268 23204 13320
rect 23256 13308 23262 13320
rect 23256 13280 24348 13308
rect 23256 13268 23262 13280
rect 21361 13243 21419 13249
rect 21361 13209 21373 13243
rect 21407 13209 21419 13243
rect 21361 13203 21419 13209
rect 22465 13243 22523 13249
rect 22465 13209 22477 13243
rect 22511 13240 22523 13243
rect 24210 13240 24216 13252
rect 22511 13212 24216 13240
rect 22511 13209 22523 13212
rect 22465 13203 22523 13209
rect 17644 13144 17816 13172
rect 17644 13132 17650 13144
rect 17954 13132 17960 13184
rect 18012 13172 18018 13184
rect 18598 13172 18604 13184
rect 18012 13144 18604 13172
rect 18012 13132 18018 13144
rect 18598 13132 18604 13144
rect 18656 13172 18662 13184
rect 20349 13175 20407 13181
rect 20349 13172 20361 13175
rect 18656 13144 20361 13172
rect 18656 13132 18662 13144
rect 20349 13141 20361 13144
rect 20395 13172 20407 13175
rect 21376 13172 21404 13203
rect 24210 13200 24216 13212
rect 24268 13200 24274 13252
rect 24320 13240 24348 13280
rect 24946 13268 24952 13320
rect 25004 13308 25010 13320
rect 25225 13311 25283 13317
rect 25225 13308 25237 13311
rect 25004 13280 25237 13308
rect 25004 13268 25010 13280
rect 25225 13277 25237 13280
rect 25271 13277 25283 13311
rect 25225 13271 25283 13277
rect 25590 13268 25596 13320
rect 25648 13308 25654 13320
rect 26237 13311 26295 13317
rect 26237 13308 26249 13311
rect 25648 13280 26249 13308
rect 25648 13268 25654 13280
rect 26237 13277 26249 13280
rect 26283 13277 26295 13311
rect 26237 13271 26295 13277
rect 28442 13268 28448 13320
rect 28500 13308 28506 13320
rect 28500 13280 29684 13308
rect 28500 13268 28506 13280
rect 29546 13240 29552 13252
rect 24320 13212 25452 13240
rect 28290 13212 29552 13240
rect 22370 13172 22376 13184
rect 20395 13144 22376 13172
rect 20395 13141 20407 13144
rect 20349 13135 20407 13141
rect 22370 13132 22376 13144
rect 22428 13132 22434 13184
rect 23474 13132 23480 13184
rect 23532 13172 23538 13184
rect 23661 13175 23719 13181
rect 23661 13172 23673 13175
rect 23532 13144 23673 13172
rect 23532 13132 23538 13144
rect 23661 13141 23673 13144
rect 23707 13141 23719 13175
rect 23661 13135 23719 13141
rect 25314 13132 25320 13184
rect 25372 13132 25378 13184
rect 25424 13172 25452 13212
rect 29546 13200 29552 13212
rect 29604 13200 29610 13252
rect 27798 13172 27804 13184
rect 25424 13144 27804 13172
rect 27798 13132 27804 13144
rect 27856 13132 27862 13184
rect 29656 13172 29684 13280
rect 29730 13268 29736 13320
rect 29788 13308 29794 13320
rect 30101 13311 30159 13317
rect 30101 13308 30113 13311
rect 29788 13280 30113 13308
rect 29788 13268 29794 13280
rect 30101 13277 30113 13280
rect 30147 13277 30159 13311
rect 32876 13308 32904 13416
rect 33686 13404 33692 13416
rect 33744 13404 33750 13456
rect 38838 13444 38844 13456
rect 37660 13416 38844 13444
rect 33778 13336 33784 13388
rect 33836 13336 33842 13388
rect 33870 13336 33876 13388
rect 33928 13336 33934 13388
rect 34054 13336 34060 13388
rect 34112 13376 34118 13388
rect 35158 13376 35164 13388
rect 34112 13348 35164 13376
rect 34112 13336 34118 13348
rect 35158 13336 35164 13348
rect 35216 13336 35222 13388
rect 35526 13336 35532 13388
rect 35584 13336 35590 13388
rect 37660 13376 37688 13416
rect 38838 13404 38844 13416
rect 38896 13404 38902 13456
rect 35728 13348 37688 13376
rect 32430 13280 32904 13308
rect 30101 13271 30159 13277
rect 33594 13268 33600 13320
rect 33652 13308 33658 13320
rect 33689 13311 33747 13317
rect 33689 13308 33701 13311
rect 33652 13280 33701 13308
rect 33652 13268 33658 13280
rect 33689 13277 33701 13280
rect 33735 13277 33747 13311
rect 33796 13308 33824 13336
rect 34146 13308 34152 13320
rect 33796 13280 34152 13308
rect 33689 13271 33747 13277
rect 34146 13268 34152 13280
rect 34204 13268 34210 13320
rect 35253 13311 35311 13317
rect 35253 13277 35265 13311
rect 35299 13308 35311 13311
rect 35728 13308 35756 13348
rect 37826 13336 37832 13388
rect 37884 13376 37890 13388
rect 38105 13379 38163 13385
rect 38105 13376 38117 13379
rect 37884 13348 38117 13376
rect 37884 13336 37890 13348
rect 38105 13345 38117 13348
rect 38151 13345 38163 13379
rect 38105 13339 38163 13345
rect 35299 13280 35756 13308
rect 35299 13277 35311 13280
rect 35253 13271 35311 13277
rect 35802 13268 35808 13320
rect 35860 13308 35866 13320
rect 36357 13311 36415 13317
rect 36357 13308 36369 13311
rect 35860 13280 36369 13308
rect 35860 13268 35866 13280
rect 36357 13277 36369 13280
rect 36403 13277 36415 13311
rect 36357 13271 36415 13277
rect 41506 13268 41512 13320
rect 41564 13268 41570 13320
rect 46290 13268 46296 13320
rect 46348 13308 46354 13320
rect 47949 13311 48007 13317
rect 47949 13308 47961 13311
rect 46348 13280 47961 13308
rect 46348 13268 46354 13280
rect 47949 13277 47961 13280
rect 47995 13277 48007 13311
rect 47949 13271 48007 13277
rect 49142 13268 49148 13320
rect 49200 13268 49206 13320
rect 30190 13200 30196 13252
rect 30248 13240 30254 13252
rect 30650 13240 30656 13252
rect 30248 13212 30656 13240
rect 30248 13200 30254 13212
rect 30650 13200 30656 13212
rect 30708 13200 30714 13252
rect 31297 13243 31355 13249
rect 31297 13209 31309 13243
rect 31343 13209 31355 13243
rect 33870 13240 33876 13252
rect 31297 13203 31355 13209
rect 33244 13212 33876 13240
rect 31110 13172 31116 13184
rect 29656 13144 31116 13172
rect 31110 13132 31116 13144
rect 31168 13132 31174 13184
rect 31312 13172 31340 13203
rect 33244 13172 33272 13212
rect 33870 13200 33876 13212
rect 33928 13240 33934 13252
rect 33928 13212 34652 13240
rect 33928 13200 33934 13212
rect 31312 13144 33272 13172
rect 34624 13172 34652 13212
rect 34698 13200 34704 13252
rect 34756 13240 34762 13252
rect 35345 13243 35403 13249
rect 35345 13240 35357 13243
rect 34756 13212 35357 13240
rect 34756 13200 34762 13212
rect 35345 13209 35357 13212
rect 35391 13209 35403 13243
rect 35345 13203 35403 13209
rect 36630 13200 36636 13252
rect 36688 13200 36694 13252
rect 36740 13212 37122 13240
rect 36354 13172 36360 13184
rect 34624 13144 36360 13172
rect 36354 13132 36360 13144
rect 36412 13132 36418 13184
rect 36538 13132 36544 13184
rect 36596 13172 36602 13184
rect 36740 13172 36768 13212
rect 36596 13144 36768 13172
rect 41325 13175 41383 13181
rect 36596 13132 36602 13144
rect 41325 13141 41337 13175
rect 41371 13172 41383 13175
rect 46106 13172 46112 13184
rect 41371 13144 46112 13172
rect 41371 13141 41383 13144
rect 41325 13135 41383 13141
rect 46106 13132 46112 13144
rect 46164 13132 46170 13184
rect 1104 13082 49864 13104
rect 1104 13030 7950 13082
rect 8002 13030 8014 13082
rect 8066 13030 8078 13082
rect 8130 13030 8142 13082
rect 8194 13030 8206 13082
rect 8258 13030 17950 13082
rect 18002 13030 18014 13082
rect 18066 13030 18078 13082
rect 18130 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 27950 13082
rect 28002 13030 28014 13082
rect 28066 13030 28078 13082
rect 28130 13030 28142 13082
rect 28194 13030 28206 13082
rect 28258 13030 37950 13082
rect 38002 13030 38014 13082
rect 38066 13030 38078 13082
rect 38130 13030 38142 13082
rect 38194 13030 38206 13082
rect 38258 13030 47950 13082
rect 48002 13030 48014 13082
rect 48066 13030 48078 13082
rect 48130 13030 48142 13082
rect 48194 13030 48206 13082
rect 48258 13030 49864 13082
rect 1104 13008 49864 13030
rect 2869 12971 2927 12977
rect 2869 12937 2881 12971
rect 2915 12968 2927 12971
rect 5442 12968 5448 12980
rect 2915 12940 5448 12968
rect 2915 12937 2927 12940
rect 2869 12931 2927 12937
rect 5442 12928 5448 12940
rect 5500 12928 5506 12980
rect 10870 12928 10876 12980
rect 10928 12968 10934 12980
rect 12161 12971 12219 12977
rect 12161 12968 12173 12971
rect 10928 12940 12173 12968
rect 10928 12928 10934 12940
rect 12161 12937 12173 12940
rect 12207 12937 12219 12971
rect 12161 12931 12219 12937
rect 12250 12928 12256 12980
rect 12308 12928 12314 12980
rect 14182 12928 14188 12980
rect 14240 12968 14246 12980
rect 15933 12971 15991 12977
rect 14240 12940 14412 12968
rect 14240 12928 14246 12940
rect 934 12860 940 12912
rect 992 12900 998 12912
rect 1673 12903 1731 12909
rect 1673 12900 1685 12903
rect 992 12872 1685 12900
rect 992 12860 998 12872
rect 1673 12869 1685 12872
rect 1719 12869 1731 12903
rect 1673 12863 1731 12869
rect 1857 12903 1915 12909
rect 1857 12869 1869 12903
rect 1903 12900 1915 12903
rect 10226 12900 10232 12912
rect 1903 12872 10232 12900
rect 1903 12869 1915 12872
rect 1857 12863 1915 12869
rect 10226 12860 10232 12872
rect 10284 12860 10290 12912
rect 12069 12903 12127 12909
rect 12069 12869 12081 12903
rect 12115 12900 12127 12903
rect 12268 12900 12296 12928
rect 12115 12872 12296 12900
rect 12115 12869 12127 12872
rect 12069 12863 12127 12869
rect 1302 12792 1308 12844
rect 1360 12832 1366 12844
rect 3053 12835 3111 12841
rect 3053 12832 3065 12835
rect 1360 12804 3065 12832
rect 1360 12792 1366 12804
rect 3053 12801 3065 12804
rect 3099 12801 3111 12835
rect 14384 12832 14412 12940
rect 15933 12937 15945 12971
rect 15979 12968 15991 12971
rect 16114 12968 16120 12980
rect 15979 12940 16120 12968
rect 15979 12937 15991 12940
rect 15933 12931 15991 12937
rect 16114 12928 16120 12940
rect 16172 12928 16178 12980
rect 18877 12971 18935 12977
rect 18877 12968 18889 12971
rect 16224 12940 18889 12968
rect 14642 12860 14648 12912
rect 14700 12900 14706 12912
rect 16224 12900 16252 12940
rect 18877 12937 18889 12940
rect 18923 12937 18935 12971
rect 18877 12931 18935 12937
rect 19705 12971 19763 12977
rect 19705 12937 19717 12971
rect 19751 12968 19763 12971
rect 19978 12968 19984 12980
rect 19751 12940 19984 12968
rect 19751 12937 19763 12940
rect 19705 12931 19763 12937
rect 19978 12928 19984 12940
rect 20036 12928 20042 12980
rect 20070 12928 20076 12980
rect 20128 12928 20134 12980
rect 23109 12971 23167 12977
rect 23109 12937 23121 12971
rect 23155 12968 23167 12971
rect 23934 12968 23940 12980
rect 23155 12940 23940 12968
rect 23155 12937 23167 12940
rect 23109 12931 23167 12937
rect 18693 12903 18751 12909
rect 14700 12872 16252 12900
rect 16776 12872 18184 12900
rect 14700 12860 14706 12872
rect 15378 12832 15384 12844
rect 14384 12818 15384 12832
rect 14398 12804 15384 12818
rect 3053 12795 3111 12801
rect 15378 12792 15384 12804
rect 15436 12792 15442 12844
rect 15838 12792 15844 12844
rect 15896 12832 15902 12844
rect 16025 12835 16083 12841
rect 16025 12832 16037 12835
rect 15896 12804 16037 12832
rect 15896 12792 15902 12804
rect 16025 12801 16037 12804
rect 16071 12801 16083 12835
rect 16482 12832 16488 12844
rect 16025 12795 16083 12801
rect 16132 12804 16488 12832
rect 12158 12724 12164 12776
rect 12216 12764 12222 12776
rect 12253 12767 12311 12773
rect 12253 12764 12265 12767
rect 12216 12736 12265 12764
rect 12216 12724 12222 12736
rect 12253 12733 12265 12736
rect 12299 12733 12311 12767
rect 12253 12727 12311 12733
rect 12434 12724 12440 12776
rect 12492 12764 12498 12776
rect 12802 12764 12808 12776
rect 12492 12736 12808 12764
rect 12492 12724 12498 12736
rect 12802 12724 12808 12736
rect 12860 12764 12866 12776
rect 12989 12767 13047 12773
rect 12989 12764 13001 12767
rect 12860 12736 13001 12764
rect 12860 12724 12866 12736
rect 12989 12733 13001 12736
rect 13035 12764 13047 12767
rect 13265 12767 13323 12773
rect 13035 12736 13124 12764
rect 13035 12733 13047 12736
rect 12989 12727 13047 12733
rect 11701 12631 11759 12637
rect 11701 12597 11713 12631
rect 11747 12628 11759 12631
rect 12618 12628 12624 12640
rect 11747 12600 12624 12628
rect 11747 12597 11759 12600
rect 11701 12591 11759 12597
rect 12618 12588 12624 12600
rect 12676 12588 12682 12640
rect 13096 12628 13124 12736
rect 13265 12733 13277 12767
rect 13311 12764 13323 12767
rect 13354 12764 13360 12776
rect 13311 12736 13360 12764
rect 13311 12733 13323 12736
rect 13265 12727 13323 12733
rect 13354 12724 13360 12736
rect 13412 12724 13418 12776
rect 13630 12724 13636 12776
rect 13688 12764 13694 12776
rect 16132 12773 16160 12804
rect 16482 12792 16488 12804
rect 16540 12792 16546 12844
rect 14737 12767 14795 12773
rect 14737 12764 14749 12767
rect 13688 12736 14749 12764
rect 13688 12724 13694 12736
rect 14737 12733 14749 12736
rect 14783 12733 14795 12767
rect 14737 12727 14795 12733
rect 16117 12767 16175 12773
rect 16117 12733 16129 12767
rect 16163 12733 16175 12767
rect 16117 12727 16175 12733
rect 16206 12724 16212 12776
rect 16264 12764 16270 12776
rect 16776 12764 16804 12872
rect 17770 12792 17776 12844
rect 17828 12832 17834 12844
rect 17865 12835 17923 12841
rect 17865 12832 17877 12835
rect 17828 12804 17877 12832
rect 17828 12792 17834 12804
rect 17865 12801 17877 12804
rect 17911 12801 17923 12835
rect 18156 12832 18184 12872
rect 18693 12869 18705 12903
rect 18739 12900 18751 12903
rect 18966 12900 18972 12912
rect 18739 12872 18972 12900
rect 18739 12869 18751 12872
rect 18693 12863 18751 12869
rect 18966 12860 18972 12872
rect 19024 12860 19030 12912
rect 23124 12900 23152 12931
rect 23934 12928 23940 12940
rect 23992 12928 23998 12980
rect 25038 12928 25044 12980
rect 25096 12968 25102 12980
rect 25777 12971 25835 12977
rect 25777 12968 25789 12971
rect 25096 12940 25789 12968
rect 25096 12928 25102 12940
rect 25777 12937 25789 12940
rect 25823 12937 25835 12971
rect 25777 12931 25835 12937
rect 27614 12928 27620 12980
rect 27672 12968 27678 12980
rect 30653 12971 30711 12977
rect 30653 12968 30665 12971
rect 27672 12940 30665 12968
rect 27672 12928 27678 12940
rect 30653 12937 30665 12940
rect 30699 12937 30711 12971
rect 30653 12931 30711 12937
rect 31938 12928 31944 12980
rect 31996 12968 32002 12980
rect 31996 12940 32536 12968
rect 31996 12928 32002 12940
rect 29546 12900 29552 12912
rect 21008 12872 23152 12900
rect 29486 12872 29552 12900
rect 18156 12804 18920 12832
rect 17865 12795 17923 12801
rect 16264 12736 16804 12764
rect 16264 12724 16270 12736
rect 16850 12724 16856 12776
rect 16908 12764 16914 12776
rect 16908 12736 18736 12764
rect 16908 12724 16914 12736
rect 14274 12628 14280 12640
rect 13096 12600 14280 12628
rect 14274 12588 14280 12600
rect 14332 12588 14338 12640
rect 15565 12631 15623 12637
rect 15565 12597 15577 12631
rect 15611 12628 15623 12631
rect 16114 12628 16120 12640
rect 15611 12600 16120 12628
rect 15611 12597 15623 12600
rect 15565 12591 15623 12597
rect 16114 12588 16120 12600
rect 16172 12588 16178 12640
rect 17405 12631 17463 12637
rect 17405 12597 17417 12631
rect 17451 12628 17463 12631
rect 18230 12628 18236 12640
rect 17451 12600 18236 12628
rect 17451 12597 17463 12600
rect 17405 12591 17463 12597
rect 18230 12588 18236 12600
rect 18288 12588 18294 12640
rect 18708 12628 18736 12736
rect 18892 12696 18920 12804
rect 19242 12792 19248 12844
rect 19300 12792 19306 12844
rect 19337 12835 19395 12841
rect 19337 12801 19349 12835
rect 19383 12832 19395 12835
rect 20714 12832 20720 12844
rect 19383 12804 20720 12832
rect 19383 12801 19395 12804
rect 19337 12795 19395 12801
rect 20714 12792 20720 12804
rect 20772 12792 20778 12844
rect 19518 12724 19524 12776
rect 19576 12724 19582 12776
rect 20162 12724 20168 12776
rect 20220 12724 20226 12776
rect 20254 12724 20260 12776
rect 20312 12724 20318 12776
rect 20717 12699 20775 12705
rect 20717 12696 20729 12699
rect 18892 12668 20729 12696
rect 20717 12665 20729 12668
rect 20763 12665 20775 12699
rect 20717 12659 20775 12665
rect 21008 12628 21036 12872
rect 29546 12860 29552 12872
rect 29604 12900 29610 12912
rect 30190 12900 30196 12912
rect 29604 12872 30196 12900
rect 29604 12860 29610 12872
rect 30190 12860 30196 12872
rect 30248 12860 30254 12912
rect 31846 12900 31852 12912
rect 30300 12872 31852 12900
rect 21085 12835 21143 12841
rect 21085 12801 21097 12835
rect 21131 12832 21143 12835
rect 21910 12832 21916 12844
rect 21131 12804 21916 12832
rect 21131 12801 21143 12804
rect 21085 12795 21143 12801
rect 21910 12792 21916 12804
rect 21968 12792 21974 12844
rect 22830 12792 22836 12844
rect 22888 12832 22894 12844
rect 23017 12835 23075 12841
rect 23017 12832 23029 12835
rect 22888 12804 23029 12832
rect 22888 12792 22894 12804
rect 23017 12801 23029 12804
rect 23063 12801 23075 12835
rect 23017 12795 23075 12801
rect 25406 12792 25412 12844
rect 25464 12832 25470 12844
rect 25774 12832 25780 12844
rect 25464 12804 25780 12832
rect 25464 12792 25470 12804
rect 25774 12792 25780 12804
rect 25832 12792 25838 12844
rect 26694 12792 26700 12844
rect 26752 12832 26758 12844
rect 27982 12832 27988 12844
rect 26752 12804 27988 12832
rect 26752 12792 26758 12804
rect 27982 12792 27988 12804
rect 28040 12792 28046 12844
rect 30098 12792 30104 12844
rect 30156 12832 30162 12844
rect 30300 12832 30328 12872
rect 31846 12860 31852 12872
rect 31904 12860 31910 12912
rect 32508 12900 32536 12940
rect 32766 12928 32772 12980
rect 32824 12968 32830 12980
rect 34057 12971 34115 12977
rect 34057 12968 34069 12971
rect 32824 12940 34069 12968
rect 32824 12928 32830 12940
rect 34057 12937 34069 12940
rect 34103 12937 34115 12971
rect 34057 12931 34115 12937
rect 35710 12928 35716 12980
rect 35768 12968 35774 12980
rect 36357 12971 36415 12977
rect 36357 12968 36369 12971
rect 35768 12940 36369 12968
rect 35768 12928 35774 12940
rect 36357 12937 36369 12940
rect 36403 12937 36415 12971
rect 36357 12931 36415 12937
rect 32585 12903 32643 12909
rect 32585 12900 32597 12903
rect 31956 12872 32260 12900
rect 32508 12872 32597 12900
rect 30156 12804 30328 12832
rect 30561 12835 30619 12841
rect 30156 12792 30162 12804
rect 30561 12801 30573 12835
rect 30607 12801 30619 12835
rect 30561 12795 30619 12801
rect 21177 12767 21235 12773
rect 21177 12733 21189 12767
rect 21223 12733 21235 12767
rect 21177 12727 21235 12733
rect 21192 12696 21220 12727
rect 21266 12724 21272 12776
rect 21324 12724 21330 12776
rect 22554 12724 22560 12776
rect 22612 12764 22618 12776
rect 23198 12764 23204 12776
rect 22612 12736 23204 12764
rect 22612 12724 22618 12736
rect 23198 12724 23204 12736
rect 23256 12724 23262 12776
rect 23934 12724 23940 12776
rect 23992 12764 23998 12776
rect 24029 12767 24087 12773
rect 24029 12764 24041 12767
rect 23992 12736 24041 12764
rect 23992 12724 23998 12736
rect 24029 12733 24041 12736
rect 24075 12733 24087 12767
rect 24029 12727 24087 12733
rect 24302 12724 24308 12776
rect 24360 12764 24366 12776
rect 26418 12764 26424 12776
rect 24360 12736 26424 12764
rect 24360 12724 24366 12736
rect 26418 12724 26424 12736
rect 26476 12724 26482 12776
rect 27798 12724 27804 12776
rect 27856 12764 27862 12776
rect 28261 12767 28319 12773
rect 28261 12764 28273 12767
rect 27856 12736 28273 12764
rect 27856 12724 27862 12736
rect 28261 12733 28273 12736
rect 28307 12764 28319 12767
rect 28994 12764 29000 12776
rect 28307 12736 29000 12764
rect 28307 12733 28319 12736
rect 28261 12727 28319 12733
rect 28994 12724 29000 12736
rect 29052 12724 29058 12776
rect 30576 12764 30604 12795
rect 30650 12792 30656 12844
rect 30708 12832 30714 12844
rect 31110 12832 31116 12844
rect 30708 12804 31116 12832
rect 30708 12792 30714 12804
rect 31110 12792 31116 12804
rect 31168 12792 31174 12844
rect 31570 12792 31576 12844
rect 31628 12832 31634 12844
rect 31754 12832 31760 12844
rect 31628 12804 31760 12832
rect 31628 12792 31634 12804
rect 31754 12792 31760 12804
rect 31812 12832 31818 12844
rect 31956 12832 31984 12872
rect 31812 12804 31984 12832
rect 32232 12832 32260 12872
rect 32585 12869 32597 12872
rect 32631 12869 32643 12903
rect 32585 12863 32643 12869
rect 34517 12903 34575 12909
rect 34517 12869 34529 12903
rect 34563 12900 34575 12903
rect 34606 12900 34612 12912
rect 34563 12872 34612 12900
rect 34563 12869 34575 12872
rect 34517 12863 34575 12869
rect 34606 12860 34612 12872
rect 34664 12860 34670 12912
rect 34882 12860 34888 12912
rect 34940 12900 34946 12912
rect 38657 12903 38715 12909
rect 38657 12900 38669 12903
rect 34940 12872 38669 12900
rect 34940 12860 34946 12872
rect 38657 12869 38669 12872
rect 38703 12900 38715 12903
rect 39942 12900 39948 12912
rect 38703 12872 39948 12900
rect 38703 12869 38715 12872
rect 38657 12863 38715 12869
rect 39942 12860 39948 12872
rect 40000 12860 40006 12912
rect 32309 12835 32367 12841
rect 32309 12832 32321 12835
rect 32232 12804 32321 12832
rect 31812 12792 31818 12804
rect 29288 12736 30604 12764
rect 30837 12767 30895 12773
rect 21192 12668 24164 12696
rect 18708 12600 21036 12628
rect 22186 12588 22192 12640
rect 22244 12588 22250 12640
rect 22646 12588 22652 12640
rect 22704 12588 22710 12640
rect 24136 12628 24164 12668
rect 26326 12628 26332 12640
rect 24136 12600 26332 12628
rect 26326 12588 26332 12600
rect 26384 12588 26390 12640
rect 27525 12631 27583 12637
rect 27525 12597 27537 12631
rect 27571 12628 27583 12631
rect 29288 12628 29316 12736
rect 30837 12733 30849 12767
rect 30883 12764 30895 12767
rect 31202 12764 31208 12776
rect 30883 12736 31208 12764
rect 30883 12733 30895 12736
rect 30837 12727 30895 12733
rect 30193 12699 30251 12705
rect 30193 12665 30205 12699
rect 30239 12696 30251 12699
rect 30374 12696 30380 12708
rect 30239 12668 30380 12696
rect 30239 12665 30251 12668
rect 30193 12659 30251 12665
rect 30374 12656 30380 12668
rect 30432 12656 30438 12708
rect 27571 12600 29316 12628
rect 29733 12631 29791 12637
rect 27571 12597 27583 12600
rect 27525 12591 27583 12597
rect 29733 12597 29745 12631
rect 29779 12628 29791 12631
rect 30006 12628 30012 12640
rect 29779 12600 30012 12628
rect 29779 12597 29791 12600
rect 29733 12591 29791 12597
rect 30006 12588 30012 12600
rect 30064 12628 30070 12640
rect 30852 12628 30880 12727
rect 31202 12724 31208 12736
rect 31260 12724 31266 12776
rect 32232 12696 32260 12804
rect 32309 12801 32321 12804
rect 32355 12801 32367 12835
rect 32309 12795 32367 12801
rect 33686 12792 33692 12844
rect 33744 12792 33750 12844
rect 36262 12792 36268 12844
rect 36320 12792 36326 12844
rect 39485 12835 39543 12841
rect 39485 12801 39497 12835
rect 39531 12832 39543 12835
rect 40037 12835 40095 12841
rect 40037 12832 40049 12835
rect 39531 12804 40049 12832
rect 39531 12801 39543 12804
rect 39485 12795 39543 12801
rect 40037 12801 40049 12804
rect 40083 12801 40095 12835
rect 40037 12795 40095 12801
rect 34882 12724 34888 12776
rect 34940 12764 34946 12776
rect 35253 12767 35311 12773
rect 35253 12764 35265 12767
rect 34940 12736 35265 12764
rect 34940 12724 34946 12736
rect 35253 12733 35265 12736
rect 35299 12733 35311 12767
rect 35253 12727 35311 12733
rect 36354 12724 36360 12776
rect 36412 12764 36418 12776
rect 36449 12767 36507 12773
rect 36449 12764 36461 12767
rect 36412 12736 36461 12764
rect 36412 12724 36418 12736
rect 36449 12733 36461 12736
rect 36495 12733 36507 12767
rect 36449 12727 36507 12733
rect 34900 12696 34928 12724
rect 32232 12668 32352 12696
rect 30064 12600 30880 12628
rect 31573 12631 31631 12637
rect 30064 12588 30070 12600
rect 31573 12597 31585 12631
rect 31619 12628 31631 12631
rect 32122 12628 32128 12640
rect 31619 12600 32128 12628
rect 31619 12597 31631 12600
rect 31573 12591 31631 12597
rect 32122 12588 32128 12600
rect 32180 12588 32186 12640
rect 32324 12628 32352 12668
rect 33612 12668 34928 12696
rect 35897 12699 35955 12705
rect 33612 12628 33640 12668
rect 35897 12665 35909 12699
rect 35943 12696 35955 12699
rect 39298 12696 39304 12708
rect 35943 12668 39304 12696
rect 35943 12665 35955 12668
rect 35897 12659 35955 12665
rect 39298 12656 39304 12668
rect 39356 12656 39362 12708
rect 32324 12600 33640 12628
rect 34790 12588 34796 12640
rect 34848 12628 34854 12640
rect 39500 12628 39528 12795
rect 46106 12792 46112 12844
rect 46164 12792 46170 12844
rect 47026 12792 47032 12844
rect 47084 12832 47090 12844
rect 47949 12835 48007 12841
rect 47949 12832 47961 12835
rect 47084 12804 47961 12832
rect 47084 12792 47090 12804
rect 47949 12801 47961 12804
rect 47995 12801 48007 12835
rect 47949 12795 48007 12801
rect 49142 12792 49148 12844
rect 49200 12792 49206 12844
rect 34848 12600 39528 12628
rect 40129 12631 40187 12637
rect 34848 12588 34854 12600
rect 40129 12597 40141 12631
rect 40175 12628 40187 12631
rect 42702 12628 42708 12640
rect 40175 12600 42708 12628
rect 40175 12597 40187 12600
rect 40129 12591 40187 12597
rect 42702 12588 42708 12600
rect 42760 12588 42766 12640
rect 45925 12631 45983 12637
rect 45925 12597 45937 12631
rect 45971 12628 45983 12631
rect 47946 12628 47952 12640
rect 45971 12600 47952 12628
rect 45971 12597 45983 12600
rect 45925 12591 45983 12597
rect 47946 12588 47952 12600
rect 48004 12588 48010 12640
rect 1104 12538 49864 12560
rect 1104 12486 2950 12538
rect 3002 12486 3014 12538
rect 3066 12486 3078 12538
rect 3130 12486 3142 12538
rect 3194 12486 3206 12538
rect 3258 12486 12950 12538
rect 13002 12486 13014 12538
rect 13066 12486 13078 12538
rect 13130 12486 13142 12538
rect 13194 12486 13206 12538
rect 13258 12486 22950 12538
rect 23002 12486 23014 12538
rect 23066 12486 23078 12538
rect 23130 12486 23142 12538
rect 23194 12486 23206 12538
rect 23258 12486 32950 12538
rect 33002 12486 33014 12538
rect 33066 12486 33078 12538
rect 33130 12486 33142 12538
rect 33194 12486 33206 12538
rect 33258 12486 42950 12538
rect 43002 12486 43014 12538
rect 43066 12486 43078 12538
rect 43130 12486 43142 12538
rect 43194 12486 43206 12538
rect 43258 12486 49864 12538
rect 1104 12464 49864 12486
rect 12989 12427 13047 12433
rect 12989 12393 13001 12427
rect 13035 12424 13047 12427
rect 16022 12424 16028 12436
rect 13035 12396 16028 12424
rect 13035 12393 13047 12396
rect 12989 12387 13047 12393
rect 16022 12384 16028 12396
rect 16080 12384 16086 12436
rect 16390 12384 16396 12436
rect 16448 12424 16454 12436
rect 20622 12424 20628 12436
rect 16448 12396 20628 12424
rect 16448 12384 16454 12396
rect 20622 12384 20628 12396
rect 20680 12384 20686 12436
rect 20806 12384 20812 12436
rect 20864 12384 20870 12436
rect 22094 12384 22100 12436
rect 22152 12384 22158 12436
rect 23198 12384 23204 12436
rect 23256 12424 23262 12436
rect 25866 12424 25872 12436
rect 23256 12396 25872 12424
rect 23256 12384 23262 12396
rect 25866 12384 25872 12396
rect 25924 12384 25930 12436
rect 26326 12384 26332 12436
rect 26384 12424 26390 12436
rect 26786 12424 26792 12436
rect 26384 12396 26792 12424
rect 26384 12384 26390 12396
rect 26786 12384 26792 12396
rect 26844 12384 26850 12436
rect 28810 12384 28816 12436
rect 28868 12424 28874 12436
rect 29546 12424 29552 12436
rect 28868 12396 29552 12424
rect 28868 12384 28874 12396
rect 29546 12384 29552 12396
rect 29604 12384 29610 12436
rect 31481 12427 31539 12433
rect 31481 12393 31493 12427
rect 31527 12424 31539 12427
rect 31754 12424 31760 12436
rect 31527 12396 31760 12424
rect 31527 12393 31539 12396
rect 31481 12387 31539 12393
rect 31754 12384 31760 12396
rect 31812 12424 31818 12436
rect 32858 12424 32864 12436
rect 31812 12396 32864 12424
rect 31812 12384 31818 12396
rect 32858 12384 32864 12396
rect 32916 12384 32922 12436
rect 33870 12384 33876 12436
rect 33928 12384 33934 12436
rect 39390 12424 39396 12436
rect 34808 12396 39396 12424
rect 15562 12316 15568 12368
rect 15620 12356 15626 12368
rect 19429 12359 19487 12365
rect 19429 12356 19441 12359
rect 15620 12328 19441 12356
rect 15620 12316 15626 12328
rect 19429 12325 19441 12328
rect 19475 12325 19487 12359
rect 19429 12319 19487 12325
rect 19536 12328 23244 12356
rect 1857 12291 1915 12297
rect 1857 12257 1869 12291
rect 1903 12288 1915 12291
rect 5350 12288 5356 12300
rect 1903 12260 5356 12288
rect 1903 12257 1915 12260
rect 1857 12251 1915 12257
rect 5350 12248 5356 12260
rect 5408 12248 5414 12300
rect 10502 12248 10508 12300
rect 10560 12248 10566 12300
rect 10778 12248 10784 12300
rect 10836 12248 10842 12300
rect 12710 12248 12716 12300
rect 12768 12288 12774 12300
rect 13449 12291 13507 12297
rect 13449 12288 13461 12291
rect 12768 12260 13461 12288
rect 12768 12248 12774 12260
rect 13449 12257 13461 12260
rect 13495 12257 13507 12291
rect 13449 12251 13507 12257
rect 13630 12248 13636 12300
rect 13688 12248 13694 12300
rect 14274 12248 14280 12300
rect 14332 12288 14338 12300
rect 14550 12288 14556 12300
rect 14332 12260 14556 12288
rect 14332 12248 14338 12260
rect 14550 12248 14556 12260
rect 14608 12248 14614 12300
rect 16850 12248 16856 12300
rect 16908 12288 16914 12300
rect 16908 12260 17080 12288
rect 16908 12248 16914 12260
rect 934 12180 940 12232
rect 992 12220 998 12232
rect 1581 12223 1639 12229
rect 1581 12220 1593 12223
rect 992 12192 1593 12220
rect 992 12180 998 12192
rect 1581 12189 1593 12192
rect 1627 12189 1639 12223
rect 1581 12183 1639 12189
rect 12250 12180 12256 12232
rect 12308 12180 12314 12232
rect 13354 12180 13360 12232
rect 13412 12220 13418 12232
rect 17052 12229 17080 12260
rect 17218 12248 17224 12300
rect 17276 12248 17282 12300
rect 18690 12248 18696 12300
rect 18748 12288 18754 12300
rect 19536 12288 19564 12328
rect 18748 12260 19564 12288
rect 18748 12248 18754 12260
rect 19978 12248 19984 12300
rect 20036 12248 20042 12300
rect 21450 12248 21456 12300
rect 21508 12248 21514 12300
rect 22554 12248 22560 12300
rect 22612 12288 22618 12300
rect 22649 12291 22707 12297
rect 22649 12288 22661 12291
rect 22612 12260 22661 12288
rect 22612 12248 22618 12260
rect 22649 12257 22661 12260
rect 22695 12257 22707 12291
rect 23216 12288 23244 12328
rect 23290 12316 23296 12368
rect 23348 12356 23354 12368
rect 23348 12328 23980 12356
rect 23348 12316 23354 12328
rect 23750 12288 23756 12300
rect 23216 12260 23756 12288
rect 22649 12251 22707 12257
rect 23750 12248 23756 12260
rect 23808 12248 23814 12300
rect 23845 12291 23903 12297
rect 23845 12257 23857 12291
rect 23891 12257 23903 12291
rect 23952 12288 23980 12328
rect 23952 12260 26096 12288
rect 23845 12251 23903 12257
rect 17037 12223 17095 12229
rect 13412 12192 13584 12220
rect 13412 12180 13418 12192
rect 12268 12152 12296 12180
rect 13446 12152 13452 12164
rect 12006 12124 13452 12152
rect 13446 12112 13452 12124
rect 13504 12112 13510 12164
rect 13556 12152 13584 12192
rect 17037 12189 17049 12223
rect 17083 12189 17095 12223
rect 17037 12183 17095 12189
rect 17770 12180 17776 12232
rect 17828 12220 17834 12232
rect 17865 12223 17923 12229
rect 17865 12220 17877 12223
rect 17828 12192 17877 12220
rect 17828 12180 17834 12192
rect 17865 12189 17877 12192
rect 17911 12189 17923 12223
rect 17865 12183 17923 12189
rect 18230 12180 18236 12232
rect 18288 12220 18294 12232
rect 19797 12223 19855 12229
rect 19797 12220 19809 12223
rect 18288 12192 19809 12220
rect 18288 12180 18294 12192
rect 19797 12189 19809 12192
rect 19843 12189 19855 12223
rect 19797 12183 19855 12189
rect 21177 12223 21235 12229
rect 21177 12189 21189 12223
rect 21223 12220 21235 12223
rect 22186 12220 22192 12232
rect 21223 12192 22192 12220
rect 21223 12189 21235 12192
rect 21177 12183 21235 12189
rect 22186 12180 22192 12192
rect 22244 12180 22250 12232
rect 23658 12180 23664 12232
rect 23716 12180 23722 12232
rect 23860 12220 23888 12251
rect 24302 12220 24308 12232
rect 23860 12192 24308 12220
rect 24302 12180 24308 12192
rect 24360 12180 24366 12232
rect 24578 12180 24584 12232
rect 24636 12180 24642 12232
rect 26068 12220 26096 12260
rect 27522 12248 27528 12300
rect 27580 12248 27586 12300
rect 30006 12248 30012 12300
rect 30064 12248 30070 12300
rect 30742 12248 30748 12300
rect 30800 12288 30806 12300
rect 31202 12288 31208 12300
rect 30800 12260 31208 12288
rect 30800 12248 30806 12260
rect 31202 12248 31208 12260
rect 31260 12288 31266 12300
rect 34808 12288 34836 12396
rect 39390 12384 39396 12396
rect 39448 12384 39454 12436
rect 41233 12359 41291 12365
rect 41233 12325 41245 12359
rect 41279 12356 41291 12359
rect 41279 12328 45554 12356
rect 41279 12325 41291 12328
rect 41233 12319 41291 12325
rect 31260 12260 34836 12288
rect 31260 12248 31266 12260
rect 34882 12248 34888 12300
rect 34940 12288 34946 12300
rect 35802 12288 35808 12300
rect 34940 12260 35808 12288
rect 34940 12248 34946 12260
rect 35802 12248 35808 12260
rect 35860 12288 35866 12300
rect 37461 12291 37519 12297
rect 37461 12288 37473 12291
rect 35860 12260 37473 12288
rect 35860 12248 35866 12260
rect 37461 12257 37473 12260
rect 37507 12257 37519 12291
rect 37461 12251 37519 12257
rect 37737 12291 37795 12297
rect 37737 12257 37749 12291
rect 37783 12288 37795 12291
rect 37826 12288 37832 12300
rect 37783 12260 37832 12288
rect 37783 12257 37795 12260
rect 37737 12251 37795 12257
rect 37826 12248 37832 12260
rect 37884 12248 37890 12300
rect 38286 12248 38292 12300
rect 38344 12288 38350 12300
rect 38344 12260 41460 12288
rect 38344 12248 38350 12260
rect 29733 12223 29791 12229
rect 26068 12192 28304 12220
rect 14458 12152 14464 12164
rect 13556 12124 14464 12152
rect 14458 12112 14464 12124
rect 14516 12112 14522 12164
rect 14553 12155 14611 12161
rect 14553 12121 14565 12155
rect 14599 12152 14611 12155
rect 14642 12152 14648 12164
rect 14599 12124 14648 12152
rect 14599 12121 14611 12124
rect 14553 12115 14611 12121
rect 14642 12112 14648 12124
rect 14700 12112 14706 12164
rect 16390 12152 16396 12164
rect 15778 12124 16396 12152
rect 12158 12044 12164 12096
rect 12216 12084 12222 12096
rect 12253 12087 12311 12093
rect 12253 12084 12265 12087
rect 12216 12056 12265 12084
rect 12216 12044 12222 12056
rect 12253 12053 12265 12056
rect 12299 12053 12311 12087
rect 12253 12047 12311 12053
rect 13357 12087 13415 12093
rect 13357 12053 13369 12087
rect 13403 12084 13415 12087
rect 15286 12084 15292 12096
rect 13403 12056 15292 12084
rect 13403 12053 13415 12056
rect 13357 12047 13415 12053
rect 15286 12044 15292 12056
rect 15344 12044 15350 12096
rect 15378 12044 15384 12096
rect 15436 12084 15442 12096
rect 15856 12084 15884 12124
rect 16390 12112 16396 12124
rect 16448 12112 16454 12164
rect 16850 12112 16856 12164
rect 16908 12152 16914 12164
rect 18601 12155 18659 12161
rect 18601 12152 18613 12155
rect 16908 12124 18613 12152
rect 16908 12112 16914 12124
rect 18601 12121 18613 12124
rect 18647 12121 18659 12155
rect 18601 12115 18659 12121
rect 22465 12155 22523 12161
rect 22465 12121 22477 12155
rect 22511 12152 22523 12155
rect 24857 12155 24915 12161
rect 22511 12124 23888 12152
rect 22511 12121 22523 12124
rect 22465 12115 22523 12121
rect 15436 12056 15884 12084
rect 15436 12044 15442 12056
rect 15930 12044 15936 12096
rect 15988 12084 15994 12096
rect 16025 12087 16083 12093
rect 16025 12084 16037 12087
rect 15988 12056 16037 12084
rect 15988 12044 15994 12056
rect 16025 12053 16037 12056
rect 16071 12053 16083 12087
rect 16025 12047 16083 12053
rect 16206 12044 16212 12096
rect 16264 12084 16270 12096
rect 16669 12087 16727 12093
rect 16669 12084 16681 12087
rect 16264 12056 16681 12084
rect 16264 12044 16270 12056
rect 16669 12053 16681 12056
rect 16715 12053 16727 12087
rect 16669 12047 16727 12053
rect 17129 12087 17187 12093
rect 17129 12053 17141 12087
rect 17175 12084 17187 12087
rect 17218 12084 17224 12096
rect 17175 12056 17224 12084
rect 17175 12053 17187 12056
rect 17129 12047 17187 12053
rect 17218 12044 17224 12056
rect 17276 12044 17282 12096
rect 19889 12087 19947 12093
rect 19889 12053 19901 12087
rect 19935 12084 19947 12087
rect 21174 12084 21180 12096
rect 19935 12056 21180 12084
rect 19935 12053 19947 12056
rect 19889 12047 19947 12053
rect 21174 12044 21180 12056
rect 21232 12044 21238 12096
rect 21269 12087 21327 12093
rect 21269 12053 21281 12087
rect 21315 12084 21327 12087
rect 22557 12087 22615 12093
rect 22557 12084 22569 12087
rect 21315 12056 22569 12084
rect 21315 12053 21327 12056
rect 21269 12047 21327 12053
rect 22557 12053 22569 12056
rect 22603 12084 22615 12087
rect 23198 12084 23204 12096
rect 22603 12056 23204 12084
rect 22603 12053 22615 12056
rect 22557 12047 22615 12053
rect 23198 12044 23204 12056
rect 23256 12044 23262 12096
rect 23293 12087 23351 12093
rect 23293 12053 23305 12087
rect 23339 12084 23351 12087
rect 23382 12084 23388 12096
rect 23339 12056 23388 12084
rect 23339 12053 23351 12056
rect 23293 12047 23351 12053
rect 23382 12044 23388 12056
rect 23440 12044 23446 12096
rect 23750 12044 23756 12096
rect 23808 12044 23814 12096
rect 23860 12084 23888 12124
rect 24857 12121 24869 12155
rect 24903 12152 24915 12155
rect 24946 12152 24952 12164
rect 24903 12124 24952 12152
rect 24903 12121 24915 12124
rect 24857 12115 24915 12121
rect 24946 12112 24952 12124
rect 25004 12112 25010 12164
rect 25406 12112 25412 12164
rect 25464 12112 25470 12164
rect 26234 12112 26240 12164
rect 26292 12152 26298 12164
rect 27062 12152 27068 12164
rect 26292 12124 27068 12152
rect 26292 12112 26298 12124
rect 27062 12112 27068 12124
rect 27120 12152 27126 12164
rect 28276 12161 28304 12192
rect 29733 12189 29745 12223
rect 29779 12189 29791 12223
rect 29733 12183 29791 12189
rect 27433 12155 27491 12161
rect 27433 12152 27445 12155
rect 27120 12124 27445 12152
rect 27120 12112 27126 12124
rect 27433 12121 27445 12124
rect 27479 12121 27491 12155
rect 27433 12115 27491 12121
rect 28261 12155 28319 12161
rect 28261 12121 28273 12155
rect 28307 12152 28319 12155
rect 28902 12152 28908 12164
rect 28307 12124 28908 12152
rect 28307 12121 28319 12124
rect 28261 12115 28319 12121
rect 28902 12112 28908 12124
rect 28960 12112 28966 12164
rect 28997 12155 29055 12161
rect 28997 12121 29009 12155
rect 29043 12152 29055 12155
rect 29748 12152 29776 12183
rect 31110 12180 31116 12232
rect 31168 12180 31174 12232
rect 31570 12180 31576 12232
rect 31628 12220 31634 12232
rect 32125 12223 32183 12229
rect 32125 12220 32137 12223
rect 31628 12192 32137 12220
rect 31628 12180 31634 12192
rect 32125 12189 32137 12192
rect 32171 12189 32183 12223
rect 32125 12183 32183 12189
rect 39298 12180 39304 12232
rect 39356 12220 39362 12232
rect 39356 12192 39620 12220
rect 39356 12180 39362 12192
rect 29043 12124 29776 12152
rect 32401 12155 32459 12161
rect 29043 12121 29055 12124
rect 28997 12115 29055 12121
rect 32401 12121 32413 12155
rect 32447 12152 32459 12155
rect 32490 12152 32496 12164
rect 32447 12124 32496 12152
rect 32447 12121 32459 12124
rect 32401 12115 32459 12121
rect 25590 12084 25596 12096
rect 23860 12056 25596 12084
rect 25590 12044 25596 12056
rect 25648 12044 25654 12096
rect 26973 12087 27031 12093
rect 26973 12053 26985 12087
rect 27019 12084 27031 12087
rect 27246 12084 27252 12096
rect 27019 12056 27252 12084
rect 27019 12053 27031 12056
rect 26973 12047 27031 12053
rect 27246 12044 27252 12056
rect 27304 12044 27310 12096
rect 27338 12044 27344 12096
rect 27396 12044 27402 12096
rect 27982 12044 27988 12096
rect 28040 12084 28046 12096
rect 28442 12084 28448 12096
rect 28040 12056 28448 12084
rect 28040 12044 28046 12056
rect 28442 12044 28448 12056
rect 28500 12084 28506 12096
rect 29012 12084 29040 12115
rect 32490 12112 32496 12124
rect 32548 12112 32554 12164
rect 33686 12152 33692 12164
rect 33626 12124 33692 12152
rect 33686 12112 33692 12124
rect 33744 12112 33750 12164
rect 35161 12155 35219 12161
rect 35161 12121 35173 12155
rect 35207 12121 35219 12155
rect 36538 12152 36544 12164
rect 36386 12124 36544 12152
rect 35161 12115 35219 12121
rect 28500 12056 29040 12084
rect 28500 12044 28506 12056
rect 31386 12044 31392 12096
rect 31444 12084 31450 12096
rect 34514 12084 34520 12096
rect 31444 12056 34520 12084
rect 31444 12044 31450 12056
rect 34514 12044 34520 12056
rect 34572 12044 34578 12096
rect 35176 12084 35204 12115
rect 36538 12112 36544 12124
rect 36596 12152 36602 12164
rect 39485 12155 39543 12161
rect 36596 12124 38226 12152
rect 36596 12112 36602 12124
rect 39485 12121 39497 12155
rect 39531 12121 39543 12155
rect 39592 12152 39620 12192
rect 39942 12180 39948 12232
rect 40000 12180 40006 12232
rect 41432 12229 41460 12260
rect 40405 12223 40463 12229
rect 40405 12220 40417 12223
rect 40052 12192 40417 12220
rect 40052 12152 40080 12192
rect 40405 12189 40417 12192
rect 40451 12189 40463 12223
rect 40405 12183 40463 12189
rect 41417 12223 41475 12229
rect 41417 12189 41429 12223
rect 41463 12189 41475 12223
rect 45526 12220 45554 12328
rect 49142 12248 49148 12300
rect 49200 12248 49206 12300
rect 46109 12223 46167 12229
rect 46109 12220 46121 12223
rect 45526 12192 46121 12220
rect 41417 12183 41475 12189
rect 46109 12189 46121 12192
rect 46155 12189 46167 12223
rect 46109 12183 46167 12189
rect 47946 12180 47952 12232
rect 48004 12180 48010 12232
rect 39592 12124 40080 12152
rect 40129 12155 40187 12161
rect 39485 12115 39543 12121
rect 40129 12121 40141 12155
rect 40175 12152 40187 12155
rect 47026 12152 47032 12164
rect 40175 12124 47032 12152
rect 40175 12121 40187 12124
rect 40129 12115 40187 12121
rect 35434 12084 35440 12096
rect 35176 12056 35440 12084
rect 35434 12044 35440 12056
rect 35492 12084 35498 12096
rect 35802 12084 35808 12096
rect 35492 12056 35808 12084
rect 35492 12044 35498 12056
rect 35802 12044 35808 12056
rect 35860 12044 35866 12096
rect 36446 12044 36452 12096
rect 36504 12084 36510 12096
rect 36633 12087 36691 12093
rect 36633 12084 36645 12087
rect 36504 12056 36645 12084
rect 36504 12044 36510 12056
rect 36633 12053 36645 12056
rect 36679 12084 36691 12087
rect 36722 12084 36728 12096
rect 36679 12056 36728 12084
rect 36679 12053 36691 12056
rect 36633 12047 36691 12053
rect 36722 12044 36728 12056
rect 36780 12044 36786 12096
rect 37642 12044 37648 12096
rect 37700 12084 37706 12096
rect 39500 12084 39528 12115
rect 47026 12112 47032 12124
rect 47084 12112 47090 12164
rect 37700 12056 39528 12084
rect 37700 12044 37706 12056
rect 40218 12044 40224 12096
rect 40276 12044 40282 12096
rect 45922 12044 45928 12096
rect 45980 12044 45986 12096
rect 1104 11994 49864 12016
rect 1104 11942 7950 11994
rect 8002 11942 8014 11994
rect 8066 11942 8078 11994
rect 8130 11942 8142 11994
rect 8194 11942 8206 11994
rect 8258 11942 17950 11994
rect 18002 11942 18014 11994
rect 18066 11942 18078 11994
rect 18130 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 27950 11994
rect 28002 11942 28014 11994
rect 28066 11942 28078 11994
rect 28130 11942 28142 11994
rect 28194 11942 28206 11994
rect 28258 11942 37950 11994
rect 38002 11942 38014 11994
rect 38066 11942 38078 11994
rect 38130 11942 38142 11994
rect 38194 11942 38206 11994
rect 38258 11942 47950 11994
rect 48002 11942 48014 11994
rect 48066 11942 48078 11994
rect 48130 11942 48142 11994
rect 48194 11942 48206 11994
rect 48258 11942 49864 11994
rect 1104 11920 49864 11942
rect 1854 11840 1860 11892
rect 1912 11880 1918 11892
rect 1912 11852 14504 11880
rect 1912 11840 1918 11852
rect 12342 11812 12348 11824
rect 12084 11784 12348 11812
rect 1026 11704 1032 11756
rect 1084 11744 1090 11756
rect 12084 11753 12112 11784
rect 12342 11772 12348 11784
rect 12400 11772 12406 11824
rect 14476 11812 14504 11852
rect 14550 11840 14556 11892
rect 14608 11880 14614 11892
rect 18601 11883 18659 11889
rect 18601 11880 18613 11883
rect 14608 11852 18613 11880
rect 14608 11840 14614 11852
rect 18601 11849 18613 11852
rect 18647 11849 18659 11883
rect 18601 11843 18659 11849
rect 19794 11840 19800 11892
rect 19852 11880 19858 11892
rect 19889 11883 19947 11889
rect 19889 11880 19901 11883
rect 19852 11852 19901 11880
rect 19852 11840 19858 11852
rect 19889 11849 19901 11852
rect 19935 11849 19947 11883
rect 26326 11880 26332 11892
rect 19889 11843 19947 11849
rect 24228 11852 26332 11880
rect 16574 11812 16580 11824
rect 14476 11784 16580 11812
rect 16574 11772 16580 11784
rect 16632 11772 16638 11824
rect 17586 11812 17592 11824
rect 16868 11784 17592 11812
rect 1581 11747 1639 11753
rect 1581 11744 1593 11747
rect 1084 11716 1593 11744
rect 1084 11704 1090 11716
rect 1581 11713 1593 11716
rect 1627 11713 1639 11747
rect 1581 11707 1639 11713
rect 2501 11747 2559 11753
rect 2501 11713 2513 11747
rect 2547 11713 2559 11747
rect 2501 11707 2559 11713
rect 12069 11747 12127 11753
rect 12069 11713 12081 11747
rect 12115 11713 12127 11747
rect 12069 11707 12127 11713
rect 934 11636 940 11688
rect 992 11676 998 11688
rect 2516 11676 2544 11707
rect 13446 11704 13452 11756
rect 13504 11704 13510 11756
rect 13814 11704 13820 11756
rect 13872 11744 13878 11756
rect 14093 11747 14151 11753
rect 14093 11744 14105 11747
rect 13872 11716 14105 11744
rect 13872 11704 13878 11716
rect 14093 11713 14105 11716
rect 14139 11744 14151 11747
rect 14139 11716 15424 11744
rect 14139 11713 14151 11716
rect 14093 11707 14151 11713
rect 992 11648 2544 11676
rect 12345 11679 12403 11685
rect 992 11636 998 11648
rect 12345 11645 12357 11679
rect 12391 11676 12403 11679
rect 12710 11676 12716 11688
rect 12391 11648 12716 11676
rect 12391 11645 12403 11648
rect 12345 11639 12403 11645
rect 12710 11636 12716 11648
rect 12768 11636 12774 11688
rect 1765 11611 1823 11617
rect 1765 11577 1777 11611
rect 1811 11608 1823 11611
rect 13464 11608 13492 11704
rect 15286 11608 15292 11620
rect 1811 11580 6914 11608
rect 13464 11580 15292 11608
rect 1811 11577 1823 11580
rect 1765 11571 1823 11577
rect 2317 11543 2375 11549
rect 2317 11509 2329 11543
rect 2363 11540 2375 11543
rect 4154 11540 4160 11552
rect 2363 11512 4160 11540
rect 2363 11509 2375 11512
rect 2317 11503 2375 11509
rect 4154 11500 4160 11512
rect 4212 11500 4218 11552
rect 6886 11540 6914 11580
rect 15286 11568 15292 11580
rect 15344 11568 15350 11620
rect 15396 11608 15424 11716
rect 15470 11704 15476 11756
rect 15528 11704 15534 11756
rect 15565 11747 15623 11753
rect 15565 11713 15577 11747
rect 15611 11744 15623 11747
rect 15838 11744 15844 11756
rect 15611 11716 15844 11744
rect 15611 11713 15623 11716
rect 15565 11707 15623 11713
rect 15838 11704 15844 11716
rect 15896 11704 15902 11756
rect 16390 11704 16396 11756
rect 16448 11744 16454 11756
rect 16868 11744 16896 11784
rect 17586 11772 17592 11784
rect 17644 11772 17650 11824
rect 22278 11812 22284 11824
rect 20088 11784 22284 11812
rect 16448 11716 16896 11744
rect 16448 11704 16454 11716
rect 15749 11679 15807 11685
rect 15749 11645 15761 11679
rect 15795 11676 15807 11679
rect 15795 11648 15884 11676
rect 15795 11645 15807 11648
rect 15749 11639 15807 11645
rect 15856 11608 15884 11648
rect 16850 11636 16856 11688
rect 16908 11636 16914 11688
rect 17129 11679 17187 11685
rect 17129 11645 17141 11679
rect 17175 11676 17187 11679
rect 19794 11676 19800 11688
rect 17175 11648 19800 11676
rect 17175 11645 17187 11648
rect 17129 11639 17187 11645
rect 19794 11636 19800 11648
rect 19852 11636 19858 11688
rect 20088 11685 20116 11784
rect 22278 11772 22284 11784
rect 22336 11772 22342 11824
rect 22462 11772 22468 11824
rect 22520 11812 22526 11824
rect 22557 11815 22615 11821
rect 22557 11812 22569 11815
rect 22520 11784 22569 11812
rect 22520 11772 22526 11784
rect 22557 11781 22569 11784
rect 22603 11812 22615 11815
rect 23290 11812 23296 11824
rect 22603 11784 23296 11812
rect 22603 11781 22615 11784
rect 22557 11775 22615 11781
rect 23290 11772 23296 11784
rect 23348 11772 23354 11824
rect 23382 11772 23388 11824
rect 23440 11812 23446 11824
rect 24228 11821 24256 11852
rect 26326 11840 26332 11852
rect 26384 11840 26390 11892
rect 27157 11883 27215 11889
rect 27157 11849 27169 11883
rect 27203 11880 27215 11883
rect 27614 11880 27620 11892
rect 27203 11852 27620 11880
rect 27203 11849 27215 11852
rect 27157 11843 27215 11849
rect 27614 11840 27620 11852
rect 27672 11840 27678 11892
rect 28902 11840 28908 11892
rect 28960 11880 28966 11892
rect 37645 11883 37703 11889
rect 28960 11852 33824 11880
rect 28960 11840 28966 11852
rect 24213 11815 24271 11821
rect 24213 11812 24225 11815
rect 23440 11784 24225 11812
rect 23440 11772 23446 11784
rect 24213 11781 24225 11784
rect 24259 11781 24271 11815
rect 24213 11775 24271 11781
rect 26786 11772 26792 11824
rect 26844 11812 26850 11824
rect 27525 11815 27583 11821
rect 27525 11812 27537 11815
rect 26844 11784 27537 11812
rect 26844 11772 26850 11784
rect 27525 11781 27537 11784
rect 27571 11781 27583 11815
rect 27525 11775 27583 11781
rect 28810 11772 28816 11824
rect 28868 11812 28874 11824
rect 31754 11812 31760 11824
rect 28868 11784 29210 11812
rect 30208 11784 31760 11812
rect 28868 11772 28874 11784
rect 20162 11704 20168 11756
rect 20220 11744 20226 11756
rect 21085 11747 21143 11753
rect 21085 11744 21097 11747
rect 20220 11716 21097 11744
rect 20220 11704 20226 11716
rect 21085 11713 21097 11716
rect 21131 11713 21143 11747
rect 21085 11707 21143 11713
rect 21177 11747 21235 11753
rect 21177 11713 21189 11747
rect 21223 11744 21235 11747
rect 23842 11744 23848 11756
rect 21223 11716 23848 11744
rect 21223 11713 21235 11716
rect 21177 11707 21235 11713
rect 23842 11704 23848 11716
rect 23900 11704 23906 11756
rect 25314 11704 25320 11756
rect 25372 11704 25378 11756
rect 26605 11747 26663 11753
rect 26605 11713 26617 11747
rect 26651 11744 26663 11747
rect 27338 11744 27344 11756
rect 26651 11716 27344 11744
rect 26651 11713 26663 11716
rect 26605 11707 26663 11713
rect 27338 11704 27344 11716
rect 27396 11704 27402 11756
rect 28442 11704 28448 11756
rect 28500 11704 28506 11756
rect 19981 11679 20039 11685
rect 19981 11645 19993 11679
rect 20027 11645 20039 11679
rect 19981 11639 20039 11645
rect 20073 11679 20131 11685
rect 20073 11645 20085 11679
rect 20119 11645 20131 11679
rect 20073 11639 20131 11645
rect 21361 11679 21419 11685
rect 21361 11645 21373 11679
rect 21407 11645 21419 11679
rect 21361 11639 21419 11645
rect 15396 11580 15884 11608
rect 14090 11540 14096 11552
rect 6886 11512 14096 11540
rect 14090 11500 14096 11512
rect 14148 11500 14154 11552
rect 14826 11500 14832 11552
rect 14884 11540 14890 11552
rect 15105 11543 15163 11549
rect 15105 11540 15117 11543
rect 14884 11512 15117 11540
rect 14884 11500 14890 11512
rect 15105 11509 15117 11512
rect 15151 11509 15163 11543
rect 15856 11540 15884 11580
rect 18138 11568 18144 11620
rect 18196 11608 18202 11620
rect 19886 11608 19892 11620
rect 18196 11580 19892 11608
rect 18196 11568 18202 11580
rect 19886 11568 19892 11580
rect 19944 11568 19950 11620
rect 19996 11608 20024 11639
rect 21376 11608 21404 11639
rect 21450 11636 21456 11688
rect 21508 11676 21514 11688
rect 22002 11676 22008 11688
rect 21508 11648 22008 11676
rect 21508 11636 21514 11648
rect 22002 11636 22008 11648
rect 22060 11676 22066 11688
rect 23385 11679 23443 11685
rect 23385 11676 23397 11679
rect 22060 11648 23397 11676
rect 22060 11636 22066 11648
rect 23385 11645 23397 11648
rect 23431 11676 23443 11679
rect 23658 11676 23664 11688
rect 23431 11648 23664 11676
rect 23431 11645 23443 11648
rect 23385 11639 23443 11645
rect 23658 11636 23664 11648
rect 23716 11676 23722 11688
rect 23934 11676 23940 11688
rect 23716 11648 23940 11676
rect 23716 11636 23722 11648
rect 23934 11636 23940 11648
rect 23992 11636 23998 11688
rect 24854 11636 24860 11688
rect 24912 11676 24918 11688
rect 25685 11679 25743 11685
rect 25685 11676 25697 11679
rect 24912 11648 25697 11676
rect 24912 11636 24918 11648
rect 25685 11645 25697 11648
rect 25731 11645 25743 11679
rect 25685 11639 25743 11645
rect 27430 11636 27436 11688
rect 27488 11676 27494 11688
rect 27617 11679 27675 11685
rect 27617 11676 27629 11679
rect 27488 11648 27629 11676
rect 27488 11636 27494 11648
rect 27617 11645 27629 11648
rect 27663 11645 27675 11679
rect 27617 11639 27675 11645
rect 27798 11636 27804 11688
rect 27856 11636 27862 11688
rect 28721 11679 28779 11685
rect 28721 11645 28733 11679
rect 28767 11676 28779 11679
rect 30208 11676 30236 11784
rect 31754 11772 31760 11784
rect 31812 11772 31818 11824
rect 32122 11772 32128 11824
rect 32180 11812 32186 11824
rect 33796 11821 33824 11852
rect 37645 11849 37657 11883
rect 37691 11880 37703 11883
rect 38105 11883 38163 11889
rect 38105 11880 38117 11883
rect 37691 11852 38117 11880
rect 37691 11849 37703 11852
rect 37645 11843 37703 11849
rect 38105 11849 38117 11852
rect 38151 11849 38163 11883
rect 38105 11843 38163 11849
rect 32677 11815 32735 11821
rect 32677 11812 32689 11815
rect 32180 11784 32689 11812
rect 32180 11772 32186 11784
rect 32677 11781 32689 11784
rect 32723 11781 32735 11815
rect 32677 11775 32735 11781
rect 33781 11815 33839 11821
rect 33781 11781 33793 11815
rect 33827 11812 33839 11815
rect 34606 11812 34612 11824
rect 33827 11784 34612 11812
rect 33827 11781 33839 11784
rect 33781 11775 33839 11781
rect 34606 11772 34612 11784
rect 34664 11772 34670 11824
rect 37274 11772 37280 11824
rect 37332 11812 37338 11824
rect 37737 11815 37795 11821
rect 37737 11812 37749 11815
rect 37332 11784 37749 11812
rect 37332 11772 37338 11784
rect 37737 11781 37749 11784
rect 37783 11781 37795 11815
rect 37737 11775 37795 11781
rect 37844 11784 38608 11812
rect 30466 11704 30472 11756
rect 30524 11744 30530 11756
rect 31113 11747 31171 11753
rect 31113 11744 31125 11747
rect 30524 11716 31125 11744
rect 30524 11704 30530 11716
rect 31113 11713 31125 11716
rect 31159 11713 31171 11747
rect 31113 11707 31171 11713
rect 31202 11704 31208 11756
rect 31260 11704 31266 11756
rect 34882 11704 34888 11756
rect 34940 11744 34946 11756
rect 35161 11747 35219 11753
rect 35161 11744 35173 11747
rect 34940 11716 35173 11744
rect 34940 11704 34946 11716
rect 35161 11713 35173 11716
rect 35207 11713 35219 11747
rect 35161 11707 35219 11713
rect 36538 11704 36544 11756
rect 36596 11704 36602 11756
rect 36722 11704 36728 11756
rect 36780 11744 36786 11756
rect 37844 11744 37872 11784
rect 36780 11716 37872 11744
rect 36780 11704 36786 11716
rect 38378 11704 38384 11756
rect 38436 11744 38442 11756
rect 38473 11747 38531 11753
rect 38473 11744 38485 11747
rect 38436 11716 38485 11744
rect 38436 11704 38442 11716
rect 38473 11713 38485 11716
rect 38519 11713 38531 11747
rect 38580 11744 38608 11784
rect 39390 11772 39396 11824
rect 39448 11772 39454 11824
rect 40218 11772 40224 11824
rect 40276 11812 40282 11824
rect 45097 11815 45155 11821
rect 45097 11812 45109 11815
rect 40276 11784 45109 11812
rect 40276 11772 40282 11784
rect 45097 11781 45109 11784
rect 45143 11781 45155 11815
rect 45097 11775 45155 11781
rect 49142 11772 49148 11824
rect 49200 11772 49206 11824
rect 38580 11716 38700 11744
rect 38473 11707 38531 11713
rect 28767 11648 30236 11676
rect 28767 11645 28779 11648
rect 28721 11639 28779 11645
rect 31386 11636 31392 11688
rect 31444 11636 31450 11688
rect 31938 11636 31944 11688
rect 31996 11676 32002 11688
rect 32769 11679 32827 11685
rect 32769 11676 32781 11679
rect 31996 11648 32781 11676
rect 31996 11636 32002 11648
rect 32769 11645 32781 11648
rect 32815 11645 32827 11679
rect 32769 11639 32827 11645
rect 32861 11679 32919 11685
rect 32861 11645 32873 11679
rect 32907 11645 32919 11679
rect 32861 11639 32919 11645
rect 22278 11608 22284 11620
rect 19996 11580 21220 11608
rect 21376 11580 22284 11608
rect 18322 11540 18328 11552
rect 15856 11512 18328 11540
rect 15105 11503 15163 11509
rect 18322 11500 18328 11512
rect 18380 11500 18386 11552
rect 19521 11543 19579 11549
rect 19521 11509 19533 11543
rect 19567 11540 19579 11543
rect 20070 11540 20076 11552
rect 19567 11512 20076 11540
rect 19567 11509 19579 11512
rect 19521 11503 19579 11509
rect 20070 11500 20076 11512
rect 20128 11500 20134 11552
rect 20622 11500 20628 11552
rect 20680 11540 20686 11552
rect 20717 11543 20775 11549
rect 20717 11540 20729 11543
rect 20680 11512 20729 11540
rect 20680 11500 20686 11512
rect 20717 11509 20729 11512
rect 20763 11509 20775 11543
rect 21192 11540 21220 11580
rect 22278 11568 22284 11580
rect 22336 11568 22342 11620
rect 28350 11608 28356 11620
rect 25240 11580 28356 11608
rect 21542 11540 21548 11552
rect 21192 11512 21548 11540
rect 20717 11503 20775 11509
rect 21542 11500 21548 11512
rect 21600 11540 21606 11552
rect 22094 11540 22100 11552
rect 21600 11512 22100 11540
rect 21600 11500 21606 11512
rect 22094 11500 22100 11512
rect 22152 11540 22158 11552
rect 22830 11540 22836 11552
rect 22152 11512 22836 11540
rect 22152 11500 22158 11512
rect 22830 11500 22836 11512
rect 22888 11500 22894 11552
rect 23290 11500 23296 11552
rect 23348 11540 23354 11552
rect 25240 11540 25268 11580
rect 28350 11568 28356 11580
rect 28408 11568 28414 11620
rect 32214 11568 32220 11620
rect 32272 11608 32278 11620
rect 32309 11611 32367 11617
rect 32309 11608 32321 11611
rect 32272 11580 32321 11608
rect 32272 11568 32278 11580
rect 32309 11577 32321 11580
rect 32355 11577 32367 11611
rect 32309 11571 32367 11577
rect 32582 11568 32588 11620
rect 32640 11608 32646 11620
rect 32876 11608 32904 11639
rect 33502 11636 33508 11688
rect 33560 11676 33566 11688
rect 34517 11679 34575 11685
rect 34517 11676 34529 11679
rect 33560 11648 34529 11676
rect 33560 11636 33566 11648
rect 34517 11645 34529 11648
rect 34563 11676 34575 11679
rect 34790 11676 34796 11688
rect 34563 11648 34796 11676
rect 34563 11645 34575 11648
rect 34517 11639 34575 11645
rect 34790 11636 34796 11648
rect 34848 11636 34854 11688
rect 35437 11679 35495 11685
rect 35437 11645 35449 11679
rect 35483 11676 35495 11679
rect 36740 11676 36768 11704
rect 38672 11685 38700 11716
rect 45922 11704 45928 11756
rect 45980 11744 45986 11756
rect 47949 11747 48007 11753
rect 47949 11744 47961 11747
rect 45980 11716 47961 11744
rect 45980 11704 45986 11716
rect 47949 11713 47961 11716
rect 47995 11713 48007 11747
rect 47949 11707 48007 11713
rect 37829 11679 37887 11685
rect 37829 11676 37841 11679
rect 35483 11648 36768 11676
rect 36924 11648 37841 11676
rect 35483 11645 35495 11648
rect 35437 11639 35495 11645
rect 32640 11580 32904 11608
rect 32640 11568 32646 11580
rect 32950 11568 32956 11620
rect 33008 11608 33014 11620
rect 33962 11608 33968 11620
rect 33008 11580 33968 11608
rect 33008 11568 33014 11580
rect 33962 11568 33968 11580
rect 34020 11568 34026 11620
rect 23348 11512 25268 11540
rect 23348 11500 23354 11512
rect 27338 11500 27344 11552
rect 27396 11540 27402 11552
rect 29730 11540 29736 11552
rect 27396 11512 29736 11540
rect 27396 11500 27402 11512
rect 29730 11500 29736 11512
rect 29788 11540 29794 11552
rect 30193 11543 30251 11549
rect 30193 11540 30205 11543
rect 29788 11512 30205 11540
rect 29788 11500 29794 11512
rect 30193 11509 30205 11512
rect 30239 11509 30251 11543
rect 30193 11503 30251 11509
rect 30745 11543 30803 11549
rect 30745 11509 30757 11543
rect 30791 11540 30803 11543
rect 35986 11540 35992 11552
rect 30791 11512 35992 11540
rect 30791 11509 30803 11512
rect 30745 11503 30803 11509
rect 35986 11500 35992 11512
rect 36044 11500 36050 11552
rect 36078 11500 36084 11552
rect 36136 11540 36142 11552
rect 36924 11549 36952 11648
rect 37829 11645 37841 11648
rect 37875 11645 37887 11679
rect 37829 11639 37887 11645
rect 38565 11679 38623 11685
rect 38565 11645 38577 11679
rect 38611 11645 38623 11679
rect 38565 11639 38623 11645
rect 38657 11679 38715 11685
rect 38657 11645 38669 11679
rect 38703 11645 38715 11679
rect 38657 11639 38715 11645
rect 36998 11568 37004 11620
rect 37056 11608 37062 11620
rect 38580 11608 38608 11639
rect 37056 11580 38608 11608
rect 39577 11611 39635 11617
rect 37056 11568 37062 11580
rect 39577 11577 39589 11611
rect 39623 11608 39635 11611
rect 44174 11608 44180 11620
rect 39623 11580 44180 11608
rect 39623 11577 39635 11580
rect 39577 11571 39635 11577
rect 44174 11568 44180 11580
rect 44232 11568 44238 11620
rect 45281 11611 45339 11617
rect 45281 11577 45293 11611
rect 45327 11608 45339 11611
rect 46658 11608 46664 11620
rect 45327 11580 46664 11608
rect 45327 11577 45339 11580
rect 45281 11571 45339 11577
rect 46658 11568 46664 11580
rect 46716 11568 46722 11620
rect 36909 11543 36967 11549
rect 36909 11540 36921 11543
rect 36136 11512 36921 11540
rect 36136 11500 36142 11512
rect 36909 11509 36921 11512
rect 36955 11509 36967 11543
rect 36909 11503 36967 11509
rect 37277 11543 37335 11549
rect 37277 11509 37289 11543
rect 37323 11540 37335 11543
rect 38286 11540 38292 11552
rect 37323 11512 38292 11540
rect 37323 11509 37335 11512
rect 37277 11503 37335 11509
rect 38286 11500 38292 11512
rect 38344 11500 38350 11552
rect 1104 11450 49864 11472
rect 1104 11398 2950 11450
rect 3002 11398 3014 11450
rect 3066 11398 3078 11450
rect 3130 11398 3142 11450
rect 3194 11398 3206 11450
rect 3258 11398 12950 11450
rect 13002 11398 13014 11450
rect 13066 11398 13078 11450
rect 13130 11398 13142 11450
rect 13194 11398 13206 11450
rect 13258 11398 22950 11450
rect 23002 11398 23014 11450
rect 23066 11398 23078 11450
rect 23130 11398 23142 11450
rect 23194 11398 23206 11450
rect 23258 11398 32950 11450
rect 33002 11398 33014 11450
rect 33066 11398 33078 11450
rect 33130 11398 33142 11450
rect 33194 11398 33206 11450
rect 33258 11398 42950 11450
rect 43002 11398 43014 11450
rect 43066 11398 43078 11450
rect 43130 11398 43142 11450
rect 43194 11398 43206 11450
rect 43258 11398 49864 11450
rect 1104 11376 49864 11398
rect 6886 11308 13216 11336
rect 1765 11271 1823 11277
rect 1765 11237 1777 11271
rect 1811 11268 1823 11271
rect 6886 11268 6914 11308
rect 1811 11240 6914 11268
rect 1811 11237 1823 11240
rect 1765 11231 1823 11237
rect 12710 11228 12716 11280
rect 12768 11228 12774 11280
rect 13188 11268 13216 11308
rect 13722 11296 13728 11348
rect 13780 11336 13786 11348
rect 14369 11339 14427 11345
rect 14369 11336 14381 11339
rect 13780 11308 14381 11336
rect 13780 11296 13786 11308
rect 14369 11305 14381 11308
rect 14415 11305 14427 11339
rect 14369 11299 14427 11305
rect 16666 11296 16672 11348
rect 16724 11336 16730 11348
rect 16761 11339 16819 11345
rect 16761 11336 16773 11339
rect 16724 11308 16773 11336
rect 16724 11296 16730 11308
rect 16761 11305 16773 11308
rect 16807 11305 16819 11339
rect 19610 11336 19616 11348
rect 16761 11299 16819 11305
rect 17420 11308 19616 11336
rect 13906 11268 13912 11280
rect 13188 11240 13912 11268
rect 13906 11228 13912 11240
rect 13964 11228 13970 11280
rect 15565 11271 15623 11277
rect 15565 11237 15577 11271
rect 15611 11268 15623 11271
rect 16482 11268 16488 11280
rect 15611 11240 16488 11268
rect 15611 11237 15623 11240
rect 15565 11231 15623 11237
rect 16482 11228 16488 11240
rect 16540 11228 16546 11280
rect 10965 11203 11023 11209
rect 10965 11169 10977 11203
rect 11011 11200 11023 11203
rect 13814 11200 13820 11212
rect 11011 11172 13820 11200
rect 11011 11169 11023 11172
rect 10965 11163 11023 11169
rect 13814 11160 13820 11172
rect 13872 11160 13878 11212
rect 14826 11160 14832 11212
rect 14884 11160 14890 11212
rect 15013 11203 15071 11209
rect 15013 11169 15025 11203
rect 15059 11200 15071 11203
rect 15102 11200 15108 11212
rect 15059 11172 15108 11200
rect 15059 11169 15071 11172
rect 15013 11163 15071 11169
rect 15102 11160 15108 11172
rect 15160 11160 15166 11212
rect 15194 11160 15200 11212
rect 15252 11200 15258 11212
rect 17420 11209 17448 11308
rect 19610 11296 19616 11308
rect 19668 11296 19674 11348
rect 19981 11339 20039 11345
rect 19981 11305 19993 11339
rect 20027 11336 20039 11339
rect 20162 11336 20168 11348
rect 20027 11308 20168 11336
rect 20027 11305 20039 11308
rect 19981 11299 20039 11305
rect 20162 11296 20168 11308
rect 20220 11296 20226 11348
rect 21266 11336 21272 11348
rect 20272 11308 21272 11336
rect 17957 11271 18015 11277
rect 17957 11237 17969 11271
rect 18003 11268 18015 11271
rect 18414 11268 18420 11280
rect 18003 11240 18420 11268
rect 18003 11237 18015 11240
rect 17957 11231 18015 11237
rect 18414 11228 18420 11240
rect 18472 11228 18478 11280
rect 19794 11228 19800 11280
rect 19852 11268 19858 11280
rect 20272 11268 20300 11308
rect 21266 11296 21272 11308
rect 21324 11336 21330 11348
rect 22189 11339 22247 11345
rect 22189 11336 22201 11339
rect 21324 11308 22201 11336
rect 21324 11296 21330 11308
rect 22189 11305 22201 11308
rect 22235 11305 22247 11339
rect 22189 11299 22247 11305
rect 22741 11339 22799 11345
rect 22741 11305 22753 11339
rect 22787 11336 22799 11339
rect 23474 11336 23480 11348
rect 22787 11308 23480 11336
rect 22787 11305 22799 11308
rect 22741 11299 22799 11305
rect 23474 11296 23480 11308
rect 23532 11296 23538 11348
rect 26329 11339 26387 11345
rect 26329 11305 26341 11339
rect 26375 11336 26387 11339
rect 26510 11336 26516 11348
rect 26375 11308 26516 11336
rect 26375 11305 26387 11308
rect 26329 11299 26387 11305
rect 26510 11296 26516 11308
rect 26568 11296 26574 11348
rect 27144 11339 27202 11345
rect 27144 11305 27156 11339
rect 27190 11336 27202 11339
rect 27522 11336 27528 11348
rect 27190 11308 27528 11336
rect 27190 11305 27202 11308
rect 27144 11299 27202 11305
rect 27522 11296 27528 11308
rect 27580 11336 27586 11348
rect 29086 11336 29092 11348
rect 27580 11308 29092 11336
rect 27580 11296 27586 11308
rect 29086 11296 29092 11308
rect 29144 11336 29150 11348
rect 29270 11336 29276 11348
rect 29144 11308 29276 11336
rect 29144 11296 29150 11308
rect 29270 11296 29276 11308
rect 29328 11296 29334 11348
rect 29733 11339 29791 11345
rect 29733 11305 29745 11339
rect 29779 11336 29791 11339
rect 32766 11336 32772 11348
rect 29779 11308 32772 11336
rect 29779 11305 29791 11308
rect 29733 11299 29791 11305
rect 32766 11296 32772 11308
rect 32824 11296 32830 11348
rect 32876 11308 33916 11336
rect 19852 11240 20300 11268
rect 28644 11240 30328 11268
rect 19852 11228 19858 11240
rect 28644 11212 28672 11240
rect 16025 11203 16083 11209
rect 16025 11200 16037 11203
rect 15252 11172 16037 11200
rect 15252 11160 15258 11172
rect 16025 11169 16037 11172
rect 16071 11169 16083 11203
rect 16025 11163 16083 11169
rect 16209 11203 16267 11209
rect 16209 11169 16221 11203
rect 16255 11200 16267 11203
rect 17405 11203 17463 11209
rect 16255 11172 17264 11200
rect 16255 11169 16267 11172
rect 16209 11163 16267 11169
rect 1578 11092 1584 11144
rect 1636 11092 1642 11144
rect 14734 11092 14740 11144
rect 14792 11092 14798 11144
rect 15933 11135 15991 11141
rect 15933 11101 15945 11135
rect 15979 11132 15991 11135
rect 16758 11132 16764 11144
rect 15979 11104 16764 11132
rect 15979 11101 15991 11104
rect 15933 11095 15991 11101
rect 16758 11092 16764 11104
rect 16816 11092 16822 11144
rect 16942 11092 16948 11144
rect 17000 11132 17006 11144
rect 17129 11135 17187 11141
rect 17129 11132 17141 11135
rect 17000 11104 17141 11132
rect 17000 11092 17006 11104
rect 17129 11101 17141 11104
rect 17175 11101 17187 11135
rect 17236 11132 17264 11172
rect 17405 11169 17417 11203
rect 17451 11169 17463 11203
rect 17405 11163 17463 11169
rect 18506 11160 18512 11212
rect 18564 11200 18570 11212
rect 18601 11203 18659 11209
rect 18601 11200 18613 11203
rect 18564 11172 18613 11200
rect 18564 11160 18570 11172
rect 18601 11169 18613 11172
rect 18647 11200 18659 11203
rect 18874 11200 18880 11212
rect 18647 11172 18880 11200
rect 18647 11169 18659 11172
rect 18601 11163 18659 11169
rect 18874 11160 18880 11172
rect 18932 11160 18938 11212
rect 20441 11203 20499 11209
rect 20441 11169 20453 11203
rect 20487 11200 20499 11203
rect 21450 11200 21456 11212
rect 20487 11172 21456 11200
rect 20487 11169 20499 11172
rect 20441 11163 20499 11169
rect 21450 11160 21456 11172
rect 21508 11160 21514 11212
rect 23201 11203 23259 11209
rect 23201 11169 23213 11203
rect 23247 11200 23259 11203
rect 23290 11200 23296 11212
rect 23247 11172 23296 11200
rect 23247 11169 23259 11172
rect 23201 11163 23259 11169
rect 23290 11160 23296 11172
rect 23348 11160 23354 11212
rect 23382 11160 23388 11212
rect 23440 11160 23446 11212
rect 23658 11160 23664 11212
rect 23716 11200 23722 11212
rect 24578 11200 24584 11212
rect 23716 11172 24584 11200
rect 23716 11160 23722 11172
rect 24578 11160 24584 11172
rect 24636 11160 24642 11212
rect 24854 11160 24860 11212
rect 24912 11160 24918 11212
rect 27246 11160 27252 11212
rect 27304 11200 27310 11212
rect 27304 11172 28580 11200
rect 27304 11160 27310 11172
rect 17862 11132 17868 11144
rect 17236 11104 17868 11132
rect 17129 11095 17187 11101
rect 17862 11092 17868 11104
rect 17920 11092 17926 11144
rect 18325 11135 18383 11141
rect 18325 11101 18337 11135
rect 18371 11132 18383 11135
rect 19150 11132 19156 11144
rect 18371 11104 19156 11132
rect 18371 11101 18383 11104
rect 18325 11095 18383 11101
rect 19150 11092 19156 11104
rect 19208 11092 19214 11144
rect 21818 11092 21824 11144
rect 21876 11092 21882 11144
rect 23750 11132 23756 11144
rect 22066 11104 23756 11132
rect 11241 11067 11299 11073
rect 11241 11033 11253 11067
rect 11287 11033 11299 11067
rect 11241 11027 11299 11033
rect 11256 10996 11284 11027
rect 12250 11024 12256 11076
rect 12308 11024 12314 11076
rect 17221 11067 17279 11073
rect 17221 11033 17233 11067
rect 17267 11064 17279 11067
rect 18966 11064 18972 11076
rect 17267 11036 18972 11064
rect 17267 11033 17279 11036
rect 17221 11027 17279 11033
rect 18966 11024 18972 11036
rect 19024 11024 19030 11076
rect 20717 11067 20775 11073
rect 20717 11033 20729 11067
rect 20763 11064 20775 11067
rect 22066 11064 22094 11104
rect 23750 11092 23756 11104
rect 23808 11092 23814 11144
rect 26878 11092 26884 11144
rect 26936 11092 26942 11144
rect 20763 11036 21128 11064
rect 20763 11033 20775 11036
rect 20717 11027 20775 11033
rect 12158 10996 12164 11008
rect 11256 10968 12164 10996
rect 12158 10956 12164 10968
rect 12216 10956 12222 11008
rect 13446 10956 13452 11008
rect 13504 10996 13510 11008
rect 18138 10996 18144 11008
rect 13504 10968 18144 10996
rect 13504 10956 13510 10968
rect 18138 10956 18144 10968
rect 18196 10956 18202 11008
rect 18417 10999 18475 11005
rect 18417 10965 18429 10999
rect 18463 10996 18475 10999
rect 18690 10996 18696 11008
rect 18463 10968 18696 10996
rect 18463 10965 18475 10968
rect 18417 10959 18475 10965
rect 18690 10956 18696 10968
rect 18748 10956 18754 11008
rect 21100 10996 21128 11036
rect 22020 11036 22094 11064
rect 23109 11067 23167 11073
rect 22020 10996 22048 11036
rect 23109 11033 23121 11067
rect 23155 11064 23167 11067
rect 23290 11064 23296 11076
rect 23155 11036 23296 11064
rect 23155 11033 23167 11036
rect 23109 11027 23167 11033
rect 23290 11024 23296 11036
rect 23348 11024 23354 11076
rect 25314 11024 25320 11076
rect 25372 11024 25378 11076
rect 28552 11064 28580 11172
rect 28626 11160 28632 11212
rect 28684 11160 28690 11212
rect 28718 11160 28724 11212
rect 28776 11200 28782 11212
rect 30300 11209 30328 11240
rect 32582 11228 32588 11280
rect 32640 11268 32646 11280
rect 32876 11277 32904 11308
rect 32861 11271 32919 11277
rect 32861 11268 32873 11271
rect 32640 11240 32873 11268
rect 32640 11228 32646 11240
rect 32861 11237 32873 11240
rect 32907 11237 32919 11271
rect 32861 11231 32919 11237
rect 33321 11271 33379 11277
rect 33321 11237 33333 11271
rect 33367 11268 33379 11271
rect 33888 11268 33916 11308
rect 33962 11296 33968 11348
rect 34020 11336 34026 11348
rect 38289 11339 38347 11345
rect 34020 11308 37136 11336
rect 34020 11296 34026 11308
rect 33367 11240 33732 11268
rect 33888 11240 34008 11268
rect 33367 11237 33379 11240
rect 33321 11231 33379 11237
rect 30193 11203 30251 11209
rect 30193 11200 30205 11203
rect 28776 11172 30205 11200
rect 28776 11160 28782 11172
rect 30193 11169 30205 11172
rect 30239 11169 30251 11203
rect 30193 11163 30251 11169
rect 30285 11203 30343 11209
rect 30285 11169 30297 11203
rect 30331 11169 30343 11203
rect 30285 11163 30343 11169
rect 31018 11160 31024 11212
rect 31076 11200 31082 11212
rect 31076 11172 32812 11200
rect 31076 11160 31082 11172
rect 29730 11092 29736 11144
rect 29788 11132 29794 11144
rect 31113 11135 31171 11141
rect 31113 11132 31125 11135
rect 29788 11104 31125 11132
rect 29788 11092 29794 11104
rect 31113 11101 31125 11104
rect 31159 11101 31171 11135
rect 32784 11132 32812 11172
rect 33704 11132 33732 11240
rect 33980 11209 34008 11240
rect 33965 11203 34023 11209
rect 33965 11169 33977 11203
rect 34011 11169 34023 11203
rect 33965 11163 34023 11169
rect 36078 11160 36084 11212
rect 36136 11160 36142 11212
rect 37108 11200 37136 11308
rect 38289 11305 38301 11339
rect 38335 11336 38347 11339
rect 42610 11336 42616 11348
rect 38335 11308 42616 11336
rect 38335 11305 38347 11308
rect 38289 11299 38347 11305
rect 42610 11296 42616 11308
rect 42668 11296 42674 11348
rect 40773 11271 40831 11277
rect 40773 11237 40785 11271
rect 40819 11268 40831 11271
rect 40819 11240 41414 11268
rect 40819 11237 40831 11240
rect 40773 11231 40831 11237
rect 41386 11200 41414 11240
rect 42702 11228 42708 11280
rect 42760 11268 42766 11280
rect 42760 11240 47992 11268
rect 42760 11228 42766 11240
rect 37108 11172 38516 11200
rect 41386 11172 45554 11200
rect 34422 11132 34428 11144
rect 32784 11104 33640 11132
rect 33704 11104 34428 11132
rect 31113 11095 31171 11101
rect 30101 11067 30159 11073
rect 30101 11064 30113 11067
rect 28382 11036 28488 11064
rect 28552 11036 30113 11064
rect 21100 10968 22048 10996
rect 28460 10996 28488 11036
rect 30101 11033 30113 11036
rect 30147 11033 30159 11067
rect 30101 11027 30159 11033
rect 31386 11024 31392 11076
rect 31444 11064 31450 11076
rect 31662 11064 31668 11076
rect 31444 11036 31668 11064
rect 31444 11024 31450 11036
rect 31662 11024 31668 11036
rect 31720 11024 31726 11076
rect 32766 11064 32772 11076
rect 32614 11036 32772 11064
rect 32766 11024 32772 11036
rect 32824 11064 32830 11076
rect 33318 11064 33324 11076
rect 32824 11036 33324 11064
rect 32824 11024 32830 11036
rect 33318 11024 33324 11036
rect 33376 11024 33382 11076
rect 33612 11064 33640 11104
rect 34422 11092 34428 11104
rect 34480 11092 34486 11144
rect 34790 11092 34796 11144
rect 34848 11132 34854 11144
rect 38488 11141 38516 11172
rect 35805 11135 35863 11141
rect 35805 11132 35817 11135
rect 34848 11104 35817 11132
rect 34848 11092 34854 11104
rect 35805 11101 35817 11104
rect 35851 11101 35863 11135
rect 38473 11135 38531 11141
rect 35805 11095 35863 11101
rect 37384 11104 37964 11132
rect 33689 11067 33747 11073
rect 33689 11064 33701 11067
rect 33612 11036 33701 11064
rect 33689 11033 33701 11036
rect 33735 11033 33747 11067
rect 33689 11027 33747 11033
rect 33778 11024 33784 11076
rect 33836 11024 33842 11076
rect 35342 11024 35348 11076
rect 35400 11064 35406 11076
rect 36538 11064 36544 11076
rect 35400 11036 36544 11064
rect 35400 11024 35406 11036
rect 36538 11024 36544 11036
rect 36596 11024 36602 11076
rect 28626 10996 28632 11008
rect 28460 10968 28632 10996
rect 28626 10956 28632 10968
rect 28684 10956 28690 11008
rect 30282 10956 30288 11008
rect 30340 10996 30346 11008
rect 31754 10996 31760 11008
rect 30340 10968 31760 10996
rect 30340 10956 30346 10968
rect 31754 10956 31760 10968
rect 31812 10996 31818 11008
rect 35526 10996 35532 11008
rect 31812 10968 35532 10996
rect 31812 10956 31818 10968
rect 35526 10956 35532 10968
rect 35584 10956 35590 11008
rect 36446 10956 36452 11008
rect 36504 10996 36510 11008
rect 37384 10996 37412 11104
rect 37458 11024 37464 11076
rect 37516 11064 37522 11076
rect 37829 11067 37887 11073
rect 37829 11064 37841 11067
rect 37516 11036 37841 11064
rect 37516 11024 37522 11036
rect 37829 11033 37841 11036
rect 37875 11033 37887 11067
rect 37936 11064 37964 11104
rect 38473 11101 38485 11135
rect 38519 11101 38531 11135
rect 38473 11095 38531 11101
rect 40954 11092 40960 11144
rect 41012 11092 41018 11144
rect 45526 11132 45554 11172
rect 47964 11141 47992 11240
rect 49142 11160 49148 11212
rect 49200 11160 49206 11212
rect 45649 11135 45707 11141
rect 45649 11132 45661 11135
rect 45526 11104 45661 11132
rect 45649 11101 45661 11104
rect 45695 11101 45707 11135
rect 45649 11095 45707 11101
rect 47949 11135 48007 11141
rect 47949 11101 47961 11135
rect 47995 11101 48007 11135
rect 47949 11095 48007 11101
rect 40129 11067 40187 11073
rect 40129 11064 40141 11067
rect 37936 11036 40141 11064
rect 37829 11027 37887 11033
rect 40129 11033 40141 11036
rect 40175 11033 40187 11067
rect 40129 11027 40187 11033
rect 40313 11067 40371 11073
rect 40313 11033 40325 11067
rect 40359 11064 40371 11067
rect 45738 11064 45744 11076
rect 40359 11036 45744 11064
rect 40359 11033 40371 11036
rect 40313 11027 40371 11033
rect 45738 11024 45744 11036
rect 45796 11024 45802 11076
rect 45833 11067 45891 11073
rect 45833 11033 45845 11067
rect 45879 11064 45891 11067
rect 46934 11064 46940 11076
rect 45879 11036 46940 11064
rect 45879 11033 45891 11036
rect 45833 11027 45891 11033
rect 46934 11024 46940 11036
rect 46992 11024 46998 11076
rect 36504 10968 37412 10996
rect 36504 10956 36510 10968
rect 1104 10906 49864 10928
rect 1104 10854 7950 10906
rect 8002 10854 8014 10906
rect 8066 10854 8078 10906
rect 8130 10854 8142 10906
rect 8194 10854 8206 10906
rect 8258 10854 17950 10906
rect 18002 10854 18014 10906
rect 18066 10854 18078 10906
rect 18130 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 27950 10906
rect 28002 10854 28014 10906
rect 28066 10854 28078 10906
rect 28130 10854 28142 10906
rect 28194 10854 28206 10906
rect 28258 10854 37950 10906
rect 38002 10854 38014 10906
rect 38066 10854 38078 10906
rect 38130 10854 38142 10906
rect 38194 10854 38206 10906
rect 38258 10854 47950 10906
rect 48002 10854 48014 10906
rect 48066 10854 48078 10906
rect 48130 10854 48142 10906
rect 48194 10854 48206 10906
rect 48258 10854 49864 10906
rect 1104 10832 49864 10854
rect 1765 10795 1823 10801
rect 1765 10761 1777 10795
rect 1811 10792 1823 10795
rect 13173 10795 13231 10801
rect 1811 10764 6914 10792
rect 1811 10761 1823 10764
rect 1765 10755 1823 10761
rect 934 10616 940 10668
rect 992 10656 998 10668
rect 1581 10659 1639 10665
rect 1581 10656 1593 10659
rect 992 10628 1593 10656
rect 992 10616 998 10628
rect 1581 10625 1593 10628
rect 1627 10625 1639 10659
rect 1581 10619 1639 10625
rect 2317 10659 2375 10665
rect 2317 10625 2329 10659
rect 2363 10625 2375 10659
rect 6886 10656 6914 10764
rect 13173 10761 13185 10795
rect 13219 10792 13231 10795
rect 15933 10795 15991 10801
rect 15933 10792 15945 10795
rect 13219 10764 15945 10792
rect 13219 10761 13231 10764
rect 13173 10755 13231 10761
rect 15933 10761 15945 10764
rect 15979 10761 15991 10795
rect 15933 10755 15991 10761
rect 16022 10752 16028 10804
rect 16080 10752 16086 10804
rect 17773 10795 17831 10801
rect 17773 10761 17785 10795
rect 17819 10761 17831 10795
rect 17773 10755 17831 10761
rect 18233 10795 18291 10801
rect 18233 10761 18245 10795
rect 18279 10792 18291 10795
rect 18598 10792 18604 10804
rect 18279 10764 18604 10792
rect 18279 10761 18291 10764
rect 18233 10755 18291 10761
rect 13541 10727 13599 10733
rect 13541 10693 13553 10727
rect 13587 10724 13599 10727
rect 17788 10724 17816 10755
rect 18598 10752 18604 10764
rect 18656 10752 18662 10804
rect 18966 10752 18972 10804
rect 19024 10752 19030 10804
rect 19426 10752 19432 10804
rect 19484 10752 19490 10804
rect 20530 10752 20536 10804
rect 20588 10792 20594 10804
rect 20625 10795 20683 10801
rect 20625 10792 20637 10795
rect 20588 10764 20637 10792
rect 20588 10752 20594 10764
rect 20625 10761 20637 10764
rect 20671 10761 20683 10795
rect 20625 10755 20683 10761
rect 20714 10752 20720 10804
rect 20772 10792 20778 10804
rect 20772 10764 24164 10792
rect 20772 10752 20778 10764
rect 13587 10696 17816 10724
rect 13587 10693 13599 10696
rect 13541 10687 13599 10693
rect 19518 10684 19524 10736
rect 19576 10724 19582 10736
rect 21726 10724 21732 10736
rect 19576 10696 21732 10724
rect 19576 10684 19582 10696
rect 21726 10684 21732 10696
rect 21784 10724 21790 10736
rect 22281 10727 22339 10733
rect 22281 10724 22293 10727
rect 21784 10696 22293 10724
rect 21784 10684 21790 10696
rect 22281 10693 22293 10696
rect 22327 10693 22339 10727
rect 24136 10724 24164 10764
rect 24210 10752 24216 10804
rect 24268 10752 24274 10804
rect 27157 10795 27215 10801
rect 27157 10761 27169 10795
rect 27203 10792 27215 10795
rect 31754 10792 31760 10804
rect 27203 10764 31760 10792
rect 27203 10761 27215 10764
rect 27157 10755 27215 10761
rect 31754 10752 31760 10764
rect 31812 10752 31818 10804
rect 31938 10752 31944 10804
rect 31996 10792 32002 10804
rect 34238 10792 34244 10804
rect 31996 10764 34244 10792
rect 31996 10752 32002 10764
rect 34238 10752 34244 10764
rect 34296 10752 34302 10804
rect 34882 10792 34888 10804
rect 34440 10764 34888 10792
rect 28813 10727 28871 10733
rect 24136 10696 27568 10724
rect 22281 10687 22339 10693
rect 27540 10668 27568 10696
rect 28813 10693 28825 10727
rect 28859 10724 28871 10727
rect 28902 10724 28908 10736
rect 28859 10696 28908 10724
rect 28859 10693 28871 10696
rect 28813 10687 28871 10693
rect 28902 10684 28908 10696
rect 28960 10684 28966 10736
rect 30282 10724 30288 10736
rect 29472 10696 30288 10724
rect 13446 10656 13452 10668
rect 6886 10628 13452 10656
rect 2317 10619 2375 10625
rect 1210 10548 1216 10600
rect 1268 10588 1274 10600
rect 2332 10588 2360 10619
rect 13446 10616 13452 10628
rect 13504 10616 13510 10668
rect 13633 10659 13691 10665
rect 13633 10625 13645 10659
rect 13679 10656 13691 10659
rect 14366 10656 14372 10668
rect 13679 10628 14372 10656
rect 13679 10625 13691 10628
rect 13633 10619 13691 10625
rect 14366 10616 14372 10628
rect 14424 10616 14430 10668
rect 14458 10616 14464 10668
rect 14516 10656 14522 10668
rect 14737 10659 14795 10665
rect 14737 10656 14749 10659
rect 14516 10628 14749 10656
rect 14516 10616 14522 10628
rect 14737 10625 14749 10628
rect 14783 10625 14795 10659
rect 14737 10619 14795 10625
rect 14829 10659 14887 10665
rect 14829 10625 14841 10659
rect 14875 10656 14887 10659
rect 16206 10656 16212 10668
rect 14875 10628 16212 10656
rect 14875 10625 14887 10628
rect 14829 10619 14887 10625
rect 16206 10616 16212 10628
rect 16264 10616 16270 10668
rect 16942 10616 16948 10668
rect 17000 10656 17006 10668
rect 17313 10659 17371 10665
rect 17313 10656 17325 10659
rect 17000 10628 17325 10656
rect 17000 10616 17006 10628
rect 17313 10625 17325 10628
rect 17359 10625 17371 10659
rect 17313 10619 17371 10625
rect 18141 10659 18199 10665
rect 18141 10625 18153 10659
rect 18187 10656 18199 10659
rect 19150 10656 19156 10668
rect 18187 10628 19156 10656
rect 18187 10625 18199 10628
rect 18141 10619 18199 10625
rect 19150 10616 19156 10628
rect 19208 10616 19214 10668
rect 19334 10616 19340 10668
rect 19392 10616 19398 10668
rect 20533 10659 20591 10665
rect 20533 10656 20545 10659
rect 19444 10628 20545 10656
rect 12802 10588 12808 10600
rect 1268 10560 2360 10588
rect 6886 10560 12808 10588
rect 1268 10548 1274 10560
rect 2501 10523 2559 10529
rect 2501 10489 2513 10523
rect 2547 10520 2559 10523
rect 6886 10520 6914 10560
rect 12802 10548 12808 10560
rect 12860 10548 12866 10600
rect 13722 10548 13728 10600
rect 13780 10548 13786 10600
rect 14918 10548 14924 10600
rect 14976 10548 14982 10600
rect 15286 10548 15292 10600
rect 15344 10588 15350 10600
rect 16117 10591 16175 10597
rect 16117 10588 16129 10591
rect 15344 10560 16129 10588
rect 15344 10548 15350 10560
rect 16117 10557 16129 10560
rect 16163 10557 16175 10591
rect 16117 10551 16175 10557
rect 18325 10591 18383 10597
rect 18325 10557 18337 10591
rect 18371 10557 18383 10591
rect 18325 10551 18383 10557
rect 2547 10492 6914 10520
rect 2547 10489 2559 10492
rect 2501 10483 2559 10489
rect 12066 10480 12072 10532
rect 12124 10520 12130 10532
rect 14369 10523 14427 10529
rect 14369 10520 14381 10523
rect 12124 10492 14381 10520
rect 12124 10480 12130 10492
rect 14369 10489 14381 10492
rect 14415 10489 14427 10523
rect 15654 10520 15660 10532
rect 14369 10483 14427 10489
rect 14476 10492 15660 10520
rect 11882 10412 11888 10464
rect 11940 10452 11946 10464
rect 14476 10452 14504 10492
rect 15654 10480 15660 10492
rect 15712 10480 15718 10532
rect 15930 10480 15936 10532
rect 15988 10520 15994 10532
rect 18340 10520 18368 10551
rect 18966 10548 18972 10600
rect 19024 10588 19030 10600
rect 19444 10588 19472 10628
rect 20533 10625 20545 10628
rect 20579 10625 20591 10659
rect 20533 10619 20591 10625
rect 23382 10616 23388 10668
rect 23440 10616 23446 10668
rect 24581 10659 24639 10665
rect 24581 10625 24593 10659
rect 24627 10656 24639 10659
rect 25593 10659 25651 10665
rect 25593 10656 25605 10659
rect 24627 10628 25605 10656
rect 24627 10625 24639 10628
rect 24581 10619 24639 10625
rect 25593 10625 25605 10628
rect 25639 10625 25651 10659
rect 25593 10619 25651 10625
rect 27522 10616 27528 10668
rect 27580 10616 27586 10668
rect 19024 10560 19472 10588
rect 19613 10591 19671 10597
rect 19024 10548 19030 10560
rect 19613 10557 19625 10591
rect 19659 10588 19671 10591
rect 19702 10588 19708 10600
rect 19659 10560 19708 10588
rect 19659 10557 19671 10560
rect 19613 10551 19671 10557
rect 19702 10548 19708 10560
rect 19760 10548 19766 10600
rect 20717 10591 20775 10597
rect 20717 10588 20729 10591
rect 19812 10560 20729 10588
rect 19812 10520 19840 10560
rect 20717 10557 20729 10560
rect 20763 10557 20775 10591
rect 20717 10551 20775 10557
rect 22002 10548 22008 10600
rect 22060 10548 22066 10600
rect 24670 10548 24676 10600
rect 24728 10548 24734 10600
rect 24854 10548 24860 10600
rect 24912 10588 24918 10600
rect 26510 10588 26516 10600
rect 24912 10560 26516 10588
rect 24912 10548 24918 10560
rect 26510 10548 26516 10560
rect 26568 10548 26574 10600
rect 27617 10591 27675 10597
rect 27617 10557 27629 10591
rect 27663 10557 27675 10591
rect 27617 10551 27675 10557
rect 27801 10591 27859 10597
rect 27801 10557 27813 10591
rect 27847 10588 27859 10591
rect 29472 10588 29500 10696
rect 30282 10684 30288 10696
rect 30340 10684 30346 10736
rect 30374 10684 30380 10736
rect 30432 10724 30438 10736
rect 30432 10696 30696 10724
rect 30432 10684 30438 10696
rect 29914 10616 29920 10668
rect 29972 10656 29978 10668
rect 30561 10659 30619 10665
rect 30561 10656 30573 10659
rect 29972 10628 30573 10656
rect 29972 10616 29978 10628
rect 30561 10625 30573 10628
rect 30607 10625 30619 10659
rect 30668 10656 30696 10696
rect 31110 10684 31116 10736
rect 31168 10724 31174 10736
rect 32030 10724 32036 10736
rect 31168 10696 32036 10724
rect 31168 10684 31174 10696
rect 32030 10684 32036 10696
rect 32088 10724 32094 10736
rect 32766 10724 32772 10736
rect 32088 10696 32772 10724
rect 32088 10684 32094 10696
rect 32766 10684 32772 10696
rect 32824 10684 32830 10736
rect 34057 10727 34115 10733
rect 34057 10693 34069 10727
rect 34103 10724 34115 10727
rect 34440 10724 34468 10764
rect 34882 10752 34888 10764
rect 34940 10752 34946 10804
rect 35066 10752 35072 10804
rect 35124 10792 35130 10804
rect 36081 10795 36139 10801
rect 35124 10764 36032 10792
rect 35124 10752 35130 10764
rect 35342 10724 35348 10736
rect 34103 10696 34468 10724
rect 35282 10696 35348 10724
rect 34103 10693 34115 10696
rect 34057 10687 34115 10693
rect 35342 10684 35348 10696
rect 35400 10684 35406 10736
rect 36004 10724 36032 10764
rect 36081 10761 36093 10795
rect 36127 10792 36139 10795
rect 36998 10792 37004 10804
rect 36127 10764 37004 10792
rect 36127 10761 36139 10764
rect 36081 10755 36139 10761
rect 36998 10752 37004 10764
rect 37056 10752 37062 10804
rect 37200 10764 38056 10792
rect 37200 10724 37228 10764
rect 36004 10696 37228 10724
rect 37274 10684 37280 10736
rect 37332 10724 37338 10736
rect 37921 10727 37979 10733
rect 37921 10724 37933 10727
rect 37332 10696 37933 10724
rect 37332 10684 37338 10696
rect 37921 10693 37933 10696
rect 37967 10693 37979 10727
rect 37921 10687 37979 10693
rect 31573 10659 31631 10665
rect 30668 10628 30788 10656
rect 30561 10619 30619 10625
rect 27847 10560 29500 10588
rect 29641 10591 29699 10597
rect 27847 10557 27859 10560
rect 27801 10551 27859 10557
rect 29641 10557 29653 10591
rect 29687 10588 29699 10591
rect 29730 10588 29736 10600
rect 29687 10560 29736 10588
rect 29687 10557 29699 10560
rect 29641 10551 29699 10557
rect 15988 10492 18368 10520
rect 18984 10492 19840 10520
rect 15988 10480 15994 10492
rect 11940 10424 14504 10452
rect 11940 10412 11946 10424
rect 15562 10412 15568 10464
rect 15620 10412 15626 10464
rect 17678 10412 17684 10464
rect 17736 10452 17742 10464
rect 18984 10452 19012 10492
rect 23750 10480 23756 10532
rect 23808 10520 23814 10532
rect 24762 10520 24768 10532
rect 23808 10492 24768 10520
rect 23808 10480 23814 10492
rect 24762 10480 24768 10492
rect 24820 10480 24826 10532
rect 25590 10480 25596 10532
rect 25648 10520 25654 10532
rect 27632 10520 27660 10551
rect 29730 10548 29736 10560
rect 29788 10548 29794 10600
rect 30374 10548 30380 10600
rect 30432 10588 30438 10600
rect 30760 10597 30788 10628
rect 31573 10625 31585 10659
rect 31619 10656 31631 10659
rect 32677 10659 32735 10665
rect 32677 10656 32689 10659
rect 31619 10628 32689 10656
rect 31619 10625 31631 10628
rect 31573 10619 31631 10625
rect 32677 10625 32689 10628
rect 32723 10625 32735 10659
rect 32677 10619 32735 10625
rect 35802 10616 35808 10668
rect 35860 10656 35866 10668
rect 35860 10628 36400 10656
rect 35860 10616 35866 10628
rect 30653 10591 30711 10597
rect 30653 10588 30665 10591
rect 30432 10560 30665 10588
rect 30432 10548 30438 10560
rect 30653 10557 30665 10560
rect 30699 10557 30711 10591
rect 30653 10551 30711 10557
rect 30745 10591 30803 10597
rect 30745 10557 30757 10591
rect 30791 10557 30803 10591
rect 30745 10551 30803 10557
rect 31754 10548 31760 10600
rect 31812 10588 31818 10600
rect 32769 10591 32827 10597
rect 32769 10588 32781 10591
rect 31812 10560 32781 10588
rect 31812 10548 31818 10560
rect 32769 10557 32781 10560
rect 32815 10557 32827 10591
rect 32769 10551 32827 10557
rect 32950 10548 32956 10600
rect 33008 10548 33014 10600
rect 33502 10548 33508 10600
rect 33560 10588 33566 10600
rect 33781 10591 33839 10597
rect 33781 10588 33793 10591
rect 33560 10560 33793 10588
rect 33560 10548 33566 10560
rect 33781 10557 33793 10560
rect 33827 10557 33839 10591
rect 36262 10588 36268 10600
rect 33781 10551 33839 10557
rect 33888 10560 36268 10588
rect 28353 10523 28411 10529
rect 28353 10520 28365 10523
rect 25648 10492 28365 10520
rect 25648 10480 25654 10492
rect 28353 10489 28365 10492
rect 28399 10520 28411 10523
rect 28534 10520 28540 10532
rect 28399 10492 28540 10520
rect 28399 10489 28411 10492
rect 28353 10483 28411 10489
rect 28534 10480 28540 10492
rect 28592 10480 28598 10532
rect 30193 10523 30251 10529
rect 30193 10489 30205 10523
rect 30239 10520 30251 10523
rect 31202 10520 31208 10532
rect 30239 10492 31208 10520
rect 30239 10489 30251 10492
rect 30193 10483 30251 10489
rect 31202 10480 31208 10492
rect 31260 10480 31266 10532
rect 31938 10520 31944 10532
rect 31496 10492 31944 10520
rect 17736 10424 19012 10452
rect 17736 10412 17742 10424
rect 19058 10412 19064 10464
rect 19116 10452 19122 10464
rect 20165 10455 20223 10461
rect 20165 10452 20177 10455
rect 19116 10424 20177 10452
rect 19116 10412 19122 10424
rect 20165 10421 20177 10424
rect 20211 10421 20223 10455
rect 20165 10415 20223 10421
rect 28442 10412 28448 10464
rect 28500 10452 28506 10464
rect 31496 10452 31524 10492
rect 31938 10480 31944 10492
rect 31996 10480 32002 10532
rect 32309 10523 32367 10529
rect 32309 10489 32321 10523
rect 32355 10520 32367 10523
rect 33888 10520 33916 10560
rect 36262 10548 36268 10560
rect 36320 10548 36326 10600
rect 36372 10588 36400 10628
rect 36446 10616 36452 10668
rect 36504 10616 36510 10668
rect 36538 10616 36544 10668
rect 36596 10616 36602 10668
rect 37829 10659 37887 10665
rect 37829 10625 37841 10659
rect 37875 10625 37887 10659
rect 37829 10619 37887 10625
rect 36633 10591 36691 10597
rect 36633 10588 36645 10591
rect 36372 10560 36645 10588
rect 36633 10557 36645 10560
rect 36679 10588 36691 10591
rect 37642 10588 37648 10600
rect 36679 10560 37648 10588
rect 36679 10557 36691 10560
rect 36633 10551 36691 10557
rect 37642 10548 37648 10560
rect 37700 10548 37706 10600
rect 37844 10520 37872 10619
rect 38028 10597 38056 10764
rect 49145 10727 49203 10733
rect 49145 10693 49157 10727
rect 49191 10724 49203 10727
rect 49234 10724 49240 10736
rect 49191 10696 49240 10724
rect 49191 10693 49203 10696
rect 49145 10687 49203 10693
rect 49234 10684 49240 10696
rect 49292 10684 49298 10736
rect 39758 10616 39764 10668
rect 39816 10616 39822 10668
rect 46934 10616 46940 10668
rect 46992 10656 46998 10668
rect 47949 10659 48007 10665
rect 47949 10656 47961 10659
rect 46992 10628 47961 10656
rect 46992 10616 46998 10628
rect 47949 10625 47961 10628
rect 47995 10625 48007 10659
rect 47949 10619 48007 10625
rect 38013 10591 38071 10597
rect 38013 10557 38025 10591
rect 38059 10557 38071 10591
rect 38013 10551 38071 10557
rect 32355 10492 33916 10520
rect 35084 10492 37872 10520
rect 39945 10523 40003 10529
rect 32355 10489 32367 10492
rect 32309 10483 32367 10489
rect 28500 10424 31524 10452
rect 28500 10412 28506 10424
rect 32674 10412 32680 10464
rect 32732 10452 32738 10464
rect 35084 10452 35112 10492
rect 39945 10489 39957 10523
rect 39991 10520 40003 10523
rect 43714 10520 43720 10532
rect 39991 10492 43720 10520
rect 39991 10489 40003 10492
rect 39945 10483 40003 10489
rect 43714 10480 43720 10492
rect 43772 10480 43778 10532
rect 32732 10424 35112 10452
rect 32732 10412 32738 10424
rect 35526 10412 35532 10464
rect 35584 10412 35590 10464
rect 37461 10455 37519 10461
rect 37461 10421 37473 10455
rect 37507 10452 37519 10455
rect 37826 10452 37832 10464
rect 37507 10424 37832 10452
rect 37507 10421 37519 10424
rect 37461 10415 37519 10421
rect 37826 10412 37832 10424
rect 37884 10412 37890 10464
rect 1104 10362 49864 10384
rect 1104 10310 2950 10362
rect 3002 10310 3014 10362
rect 3066 10310 3078 10362
rect 3130 10310 3142 10362
rect 3194 10310 3206 10362
rect 3258 10310 12950 10362
rect 13002 10310 13014 10362
rect 13066 10310 13078 10362
rect 13130 10310 13142 10362
rect 13194 10310 13206 10362
rect 13258 10310 22950 10362
rect 23002 10310 23014 10362
rect 23066 10310 23078 10362
rect 23130 10310 23142 10362
rect 23194 10310 23206 10362
rect 23258 10310 32950 10362
rect 33002 10310 33014 10362
rect 33066 10310 33078 10362
rect 33130 10310 33142 10362
rect 33194 10310 33206 10362
rect 33258 10310 42950 10362
rect 43002 10310 43014 10362
rect 43066 10310 43078 10362
rect 43130 10310 43142 10362
rect 43194 10310 43206 10362
rect 43258 10310 49864 10362
rect 1104 10288 49864 10310
rect 12526 10208 12532 10260
rect 12584 10248 12590 10260
rect 12805 10251 12863 10257
rect 12805 10248 12817 10251
rect 12584 10220 12817 10248
rect 12584 10208 12590 10220
rect 12805 10217 12817 10220
rect 12851 10217 12863 10251
rect 12805 10211 12863 10217
rect 13630 10208 13636 10260
rect 13688 10248 13694 10260
rect 16025 10251 16083 10257
rect 16025 10248 16037 10251
rect 13688 10220 16037 10248
rect 13688 10208 13694 10220
rect 16025 10217 16037 10220
rect 16071 10217 16083 10251
rect 16025 10211 16083 10217
rect 17954 10208 17960 10260
rect 18012 10248 18018 10260
rect 18012 10220 18368 10248
rect 18012 10208 18018 10220
rect 11609 10183 11667 10189
rect 11609 10149 11621 10183
rect 11655 10180 11667 10183
rect 12434 10180 12440 10192
rect 11655 10152 12440 10180
rect 11655 10149 11667 10152
rect 11609 10143 11667 10149
rect 12434 10140 12440 10152
rect 12492 10140 12498 10192
rect 16577 10183 16635 10189
rect 16577 10149 16589 10183
rect 16623 10180 16635 10183
rect 16623 10152 18276 10180
rect 16623 10149 16635 10152
rect 16577 10143 16635 10149
rect 1857 10115 1915 10121
rect 1857 10081 1869 10115
rect 1903 10112 1915 10115
rect 11882 10112 11888 10124
rect 1903 10084 11888 10112
rect 1903 10081 1915 10084
rect 1857 10075 1915 10081
rect 11882 10072 11888 10084
rect 11940 10072 11946 10124
rect 12066 10072 12072 10124
rect 12124 10072 12130 10124
rect 12158 10072 12164 10124
rect 12216 10072 12222 10124
rect 13354 10072 13360 10124
rect 13412 10072 13418 10124
rect 16114 10072 16120 10124
rect 16172 10112 16178 10124
rect 17037 10115 17095 10121
rect 17037 10112 17049 10115
rect 16172 10084 17049 10112
rect 16172 10072 16178 10084
rect 17037 10081 17049 10084
rect 17083 10081 17095 10115
rect 17037 10075 17095 10081
rect 17129 10115 17187 10121
rect 17129 10081 17141 10115
rect 17175 10112 17187 10115
rect 17678 10112 17684 10124
rect 17175 10084 17684 10112
rect 17175 10081 17187 10084
rect 17129 10075 17187 10081
rect 934 10004 940 10056
rect 992 10044 998 10056
rect 1581 10047 1639 10053
rect 1581 10044 1593 10047
rect 992 10016 1593 10044
rect 992 10004 998 10016
rect 1581 10013 1593 10016
rect 1627 10013 1639 10047
rect 1581 10007 1639 10013
rect 11974 10004 11980 10056
rect 12032 10004 12038 10056
rect 13262 10004 13268 10056
rect 13320 10004 13326 10056
rect 13814 10004 13820 10056
rect 13872 10044 13878 10056
rect 14277 10047 14335 10053
rect 14277 10044 14289 10047
rect 13872 10016 14289 10044
rect 13872 10004 13878 10016
rect 14277 10013 14289 10016
rect 14323 10013 14335 10047
rect 16390 10044 16396 10056
rect 14277 10007 14335 10013
rect 16132 10016 16396 10044
rect 16132 9988 16160 10016
rect 16390 10004 16396 10016
rect 16448 10004 16454 10056
rect 16574 10004 16580 10056
rect 16632 10044 16638 10056
rect 17144 10044 17172 10075
rect 17678 10072 17684 10084
rect 17736 10072 17742 10124
rect 18248 10121 18276 10152
rect 18340 10121 18368 10220
rect 19242 10208 19248 10260
rect 19300 10248 19306 10260
rect 19705 10251 19763 10257
rect 19705 10248 19717 10251
rect 19300 10220 19717 10248
rect 19300 10208 19306 10220
rect 19705 10217 19717 10220
rect 19751 10217 19763 10251
rect 20990 10248 20996 10260
rect 19705 10211 19763 10217
rect 20180 10220 20996 10248
rect 18233 10115 18291 10121
rect 18233 10081 18245 10115
rect 18279 10081 18291 10115
rect 18233 10075 18291 10081
rect 18325 10115 18383 10121
rect 18325 10081 18337 10115
rect 18371 10081 18383 10115
rect 18325 10075 18383 10081
rect 18141 10047 18199 10053
rect 16632 10016 17172 10044
rect 17696 10016 18092 10044
rect 16632 10004 16638 10016
rect 13173 9979 13231 9985
rect 13173 9945 13185 9979
rect 13219 9976 13231 9979
rect 13446 9976 13452 9988
rect 13219 9948 13452 9976
rect 13219 9945 13231 9948
rect 13173 9939 13231 9945
rect 13446 9936 13452 9948
rect 13504 9936 13510 9988
rect 14550 9936 14556 9988
rect 14608 9936 14614 9988
rect 16114 9976 16120 9988
rect 15778 9948 16120 9976
rect 16114 9936 16120 9948
rect 16172 9936 16178 9988
rect 16206 9936 16212 9988
rect 16264 9976 16270 9988
rect 17696 9976 17724 10016
rect 16264 9948 17724 9976
rect 16264 9936 16270 9948
rect 14568 9908 14596 9936
rect 15930 9908 15936 9920
rect 14568 9880 15936 9908
rect 15930 9868 15936 9880
rect 15988 9868 15994 9920
rect 16942 9868 16948 9920
rect 17000 9868 17006 9920
rect 17773 9911 17831 9917
rect 17773 9877 17785 9911
rect 17819 9908 17831 9911
rect 17954 9908 17960 9920
rect 17819 9880 17960 9908
rect 17819 9877 17831 9880
rect 17773 9871 17831 9877
rect 17954 9868 17960 9880
rect 18012 9868 18018 9920
rect 18064 9908 18092 10016
rect 18141 10013 18153 10047
rect 18187 10044 18199 10047
rect 19058 10044 19064 10056
rect 18187 10016 19064 10044
rect 18187 10013 18199 10016
rect 18141 10007 18199 10013
rect 19058 10004 19064 10016
rect 19116 10004 19122 10056
rect 20180 9908 20208 10220
rect 20990 10208 20996 10220
rect 21048 10208 21054 10260
rect 21726 10208 21732 10260
rect 21784 10248 21790 10260
rect 22005 10251 22063 10257
rect 22005 10248 22017 10251
rect 21784 10220 22017 10248
rect 21784 10208 21790 10220
rect 22005 10217 22017 10220
rect 22051 10217 22063 10251
rect 22005 10211 22063 10217
rect 23290 10208 23296 10260
rect 23348 10248 23354 10260
rect 24029 10251 24087 10257
rect 24029 10248 24041 10251
rect 23348 10220 24041 10248
rect 23348 10208 23354 10220
rect 24029 10217 24041 10220
rect 24075 10217 24087 10251
rect 24029 10211 24087 10217
rect 24670 10208 24676 10260
rect 24728 10248 24734 10260
rect 28721 10251 28779 10257
rect 24728 10220 28672 10248
rect 24728 10208 24734 10220
rect 28644 10180 28672 10220
rect 28721 10217 28733 10251
rect 28767 10248 28779 10251
rect 29086 10248 29092 10260
rect 28767 10220 29092 10248
rect 28767 10217 28779 10220
rect 28721 10211 28779 10217
rect 29086 10208 29092 10220
rect 29144 10248 29150 10260
rect 30190 10248 30196 10260
rect 29144 10220 30196 10248
rect 29144 10208 29150 10220
rect 30190 10208 30196 10220
rect 30248 10208 30254 10260
rect 30466 10208 30472 10260
rect 30524 10208 30530 10260
rect 31386 10208 31392 10260
rect 31444 10248 31450 10260
rect 32125 10251 32183 10257
rect 32125 10248 32137 10251
rect 31444 10220 32137 10248
rect 31444 10208 31450 10220
rect 32125 10217 32137 10220
rect 32171 10217 32183 10251
rect 32125 10211 32183 10217
rect 34882 10208 34888 10260
rect 34940 10248 34946 10260
rect 36633 10251 36691 10257
rect 36633 10248 36645 10251
rect 34940 10220 36645 10248
rect 34940 10208 34946 10220
rect 36633 10217 36645 10220
rect 36679 10217 36691 10251
rect 36633 10211 36691 10217
rect 37461 10251 37519 10257
rect 37461 10217 37473 10251
rect 37507 10248 37519 10251
rect 40954 10248 40960 10260
rect 37507 10220 40960 10248
rect 37507 10217 37519 10220
rect 37461 10211 37519 10217
rect 30484 10180 30512 10208
rect 28644 10152 30512 10180
rect 31662 10140 31668 10192
rect 31720 10180 31726 10192
rect 32674 10180 32680 10192
rect 31720 10152 32680 10180
rect 31720 10140 31726 10152
rect 32674 10140 32680 10152
rect 32732 10140 32738 10192
rect 32766 10140 32772 10192
rect 32824 10180 32830 10192
rect 33965 10183 34023 10189
rect 33965 10180 33977 10183
rect 32824 10152 33977 10180
rect 32824 10140 32830 10152
rect 33965 10149 33977 10152
rect 34011 10149 34023 10183
rect 36648 10180 36676 10211
rect 40954 10208 40960 10220
rect 41012 10208 41018 10260
rect 36648 10152 38056 10180
rect 33965 10143 34023 10149
rect 20254 10072 20260 10124
rect 20312 10112 20318 10124
rect 22002 10112 22008 10124
rect 20312 10084 22008 10112
rect 20312 10072 20318 10084
rect 22002 10072 22008 10084
rect 22060 10112 22066 10124
rect 23201 10115 23259 10121
rect 23201 10112 23213 10115
rect 22060 10084 23213 10112
rect 22060 10072 22066 10084
rect 23201 10081 23213 10084
rect 23247 10081 23259 10115
rect 23201 10075 23259 10081
rect 24581 10115 24639 10121
rect 24581 10081 24593 10115
rect 24627 10112 24639 10115
rect 30377 10115 30435 10121
rect 24627 10084 27016 10112
rect 24627 10081 24639 10084
rect 24581 10075 24639 10081
rect 26988 10056 27016 10084
rect 30377 10081 30389 10115
rect 30423 10112 30435 10115
rect 30742 10112 30748 10124
rect 30423 10084 30748 10112
rect 30423 10081 30435 10084
rect 30377 10075 30435 10081
rect 30742 10072 30748 10084
rect 30800 10072 30806 10124
rect 31202 10072 31208 10124
rect 31260 10112 31266 10124
rect 32214 10112 32220 10124
rect 31260 10084 32220 10112
rect 31260 10072 31266 10084
rect 32214 10072 32220 10084
rect 32272 10072 32278 10124
rect 32398 10072 32404 10124
rect 32456 10112 32462 10124
rect 33137 10115 33195 10121
rect 33137 10112 33149 10115
rect 32456 10084 33149 10112
rect 32456 10072 32462 10084
rect 33137 10081 33149 10084
rect 33183 10081 33195 10115
rect 33137 10075 33195 10081
rect 33502 10072 33508 10124
rect 33560 10112 33566 10124
rect 34885 10115 34943 10121
rect 34885 10112 34897 10115
rect 33560 10084 34897 10112
rect 33560 10072 33566 10084
rect 34885 10081 34897 10084
rect 34931 10081 34943 10115
rect 34885 10075 34943 10081
rect 37734 10072 37740 10124
rect 37792 10112 37798 10124
rect 38028 10121 38056 10152
rect 37921 10115 37979 10121
rect 37921 10112 37933 10115
rect 37792 10084 37933 10112
rect 37792 10072 37798 10084
rect 37921 10081 37933 10084
rect 37967 10081 37979 10115
rect 37921 10075 37979 10081
rect 38013 10115 38071 10121
rect 38013 10081 38025 10115
rect 38059 10081 38071 10115
rect 38013 10075 38071 10081
rect 40313 10115 40371 10121
rect 40313 10081 40325 10115
rect 40359 10112 40371 10115
rect 40359 10084 41414 10112
rect 40359 10081 40371 10084
rect 40313 10075 40371 10081
rect 22462 10004 22468 10056
rect 22520 10004 22526 10056
rect 26970 10004 26976 10056
rect 27028 10004 27034 10056
rect 29917 10047 29975 10053
rect 29917 10013 29929 10047
rect 29963 10013 29975 10047
rect 29917 10007 29975 10013
rect 33045 10047 33103 10053
rect 33045 10013 33057 10047
rect 33091 10044 33103 10047
rect 33410 10044 33416 10056
rect 33091 10016 33416 10044
rect 33091 10013 33103 10016
rect 33045 10007 33103 10013
rect 20533 9979 20591 9985
rect 20533 9945 20545 9979
rect 20579 9976 20591 9979
rect 20806 9976 20812 9988
rect 20579 9948 20812 9976
rect 20579 9945 20591 9948
rect 20533 9939 20591 9945
rect 20806 9936 20812 9948
rect 20864 9936 20870 9988
rect 21818 9976 21824 9988
rect 21758 9948 21824 9976
rect 21818 9936 21824 9948
rect 21876 9976 21882 9988
rect 23382 9976 23388 9988
rect 21876 9948 23388 9976
rect 21876 9936 21882 9948
rect 23382 9936 23388 9948
rect 23440 9936 23446 9988
rect 24854 9936 24860 9988
rect 24912 9936 24918 9988
rect 25314 9936 25320 9988
rect 25372 9936 25378 9988
rect 26878 9936 26884 9988
rect 26936 9976 26942 9988
rect 27249 9979 27307 9985
rect 27249 9976 27261 9979
rect 26936 9948 27261 9976
rect 26936 9936 26942 9948
rect 27249 9945 27261 9948
rect 27295 9976 27307 9979
rect 27338 9976 27344 9988
rect 27295 9948 27344 9976
rect 27295 9945 27307 9948
rect 27249 9939 27307 9945
rect 27338 9936 27344 9948
rect 27396 9936 27402 9988
rect 28626 9976 28632 9988
rect 28474 9948 28632 9976
rect 28626 9936 28632 9948
rect 28684 9976 28690 9988
rect 28902 9976 28908 9988
rect 28684 9948 28908 9976
rect 28684 9936 28690 9948
rect 28902 9936 28908 9948
rect 28960 9936 28966 9988
rect 29932 9976 29960 10007
rect 33410 10004 33416 10016
rect 33468 10004 33474 10056
rect 37826 10004 37832 10056
rect 37884 10004 37890 10056
rect 38933 10047 38991 10053
rect 38933 10013 38945 10047
rect 38979 10044 38991 10047
rect 38979 10016 40356 10044
rect 38979 10013 38991 10016
rect 38933 10007 38991 10013
rect 30558 9976 30564 9988
rect 29932 9948 30564 9976
rect 30558 9936 30564 9948
rect 30616 9936 30622 9988
rect 30650 9936 30656 9988
rect 30708 9936 30714 9988
rect 32030 9976 32036 9988
rect 31878 9948 32036 9976
rect 32030 9936 32036 9948
rect 32088 9936 32094 9988
rect 34330 9976 34336 9988
rect 32600 9948 34336 9976
rect 18064 9880 20208 9908
rect 23566 9868 23572 9920
rect 23624 9908 23630 9920
rect 26329 9911 26387 9917
rect 26329 9908 26341 9911
rect 23624 9880 26341 9908
rect 23624 9868 23630 9880
rect 26329 9877 26341 9880
rect 26375 9877 26387 9911
rect 26329 9871 26387 9877
rect 28534 9868 28540 9920
rect 28592 9908 28598 9920
rect 31386 9908 31392 9920
rect 28592 9880 31392 9908
rect 28592 9868 28598 9880
rect 31386 9868 31392 9880
rect 31444 9868 31450 9920
rect 32600 9917 32628 9948
rect 34330 9936 34336 9948
rect 34388 9936 34394 9988
rect 35066 9936 35072 9988
rect 35124 9976 35130 9988
rect 35161 9979 35219 9985
rect 35161 9976 35173 9979
rect 35124 9948 35173 9976
rect 35124 9936 35130 9948
rect 35161 9945 35173 9948
rect 35207 9945 35219 9979
rect 35161 9939 35219 9945
rect 35434 9936 35440 9988
rect 35492 9976 35498 9988
rect 35618 9976 35624 9988
rect 35492 9948 35624 9976
rect 35492 9936 35498 9948
rect 35618 9936 35624 9948
rect 35676 9936 35682 9988
rect 38746 9936 38752 9988
rect 38804 9936 38810 9988
rect 40126 9936 40132 9988
rect 40184 9936 40190 9988
rect 32585 9911 32643 9917
rect 32585 9877 32597 9911
rect 32631 9877 32643 9911
rect 32585 9871 32643 9877
rect 32674 9868 32680 9920
rect 32732 9908 32738 9920
rect 32953 9911 33011 9917
rect 32953 9908 32965 9911
rect 32732 9880 32965 9908
rect 32732 9868 32738 9880
rect 32953 9877 32965 9880
rect 32999 9877 33011 9911
rect 32953 9871 33011 9877
rect 34514 9868 34520 9920
rect 34572 9908 34578 9920
rect 35452 9908 35480 9936
rect 34572 9880 35480 9908
rect 40328 9908 40356 10016
rect 41386 9976 41414 10084
rect 49142 10072 49148 10124
rect 49200 10072 49206 10124
rect 42610 10004 42616 10056
rect 42668 10044 42674 10056
rect 44361 10047 44419 10053
rect 44361 10044 44373 10047
rect 42668 10016 44373 10044
rect 42668 10004 42674 10016
rect 44361 10013 44373 10016
rect 44407 10013 44419 10047
rect 44361 10007 44419 10013
rect 45738 10004 45744 10056
rect 45796 10044 45802 10056
rect 46109 10047 46167 10053
rect 46109 10044 46121 10047
rect 45796 10016 46121 10044
rect 45796 10004 45802 10016
rect 46109 10013 46121 10016
rect 46155 10013 46167 10047
rect 46109 10007 46167 10013
rect 46658 10004 46664 10056
rect 46716 10044 46722 10056
rect 47949 10047 48007 10053
rect 47949 10044 47961 10047
rect 46716 10016 47961 10044
rect 46716 10004 46722 10016
rect 47949 10013 47961 10016
rect 47995 10013 48007 10047
rect 47949 10007 48007 10013
rect 42702 9976 42708 9988
rect 41386 9948 42708 9976
rect 42702 9936 42708 9948
rect 42760 9936 42766 9988
rect 44545 9979 44603 9985
rect 44545 9945 44557 9979
rect 44591 9976 44603 9979
rect 46750 9976 46756 9988
rect 44591 9948 46756 9976
rect 44591 9945 44603 9948
rect 44545 9939 44603 9945
rect 46750 9936 46756 9948
rect 46808 9936 46814 9988
rect 47302 9936 47308 9988
rect 47360 9936 47366 9988
rect 42794 9908 42800 9920
rect 40328 9880 42800 9908
rect 34572 9868 34578 9880
rect 42794 9868 42800 9880
rect 42852 9868 42858 9920
rect 1104 9818 49864 9840
rect 1104 9766 7950 9818
rect 8002 9766 8014 9818
rect 8066 9766 8078 9818
rect 8130 9766 8142 9818
rect 8194 9766 8206 9818
rect 8258 9766 17950 9818
rect 18002 9766 18014 9818
rect 18066 9766 18078 9818
rect 18130 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 27950 9818
rect 28002 9766 28014 9818
rect 28066 9766 28078 9818
rect 28130 9766 28142 9818
rect 28194 9766 28206 9818
rect 28258 9766 37950 9818
rect 38002 9766 38014 9818
rect 38066 9766 38078 9818
rect 38130 9766 38142 9818
rect 38194 9766 38206 9818
rect 38258 9766 47950 9818
rect 48002 9766 48014 9818
rect 48066 9766 48078 9818
rect 48130 9766 48142 9818
rect 48194 9766 48206 9818
rect 48258 9766 49864 9818
rect 1104 9744 49864 9766
rect 16114 9664 16120 9716
rect 16172 9664 16178 9716
rect 25590 9704 25596 9716
rect 16776 9676 25596 9704
rect 12434 9596 12440 9648
rect 12492 9596 12498 9648
rect 12529 9639 12587 9645
rect 12529 9605 12541 9639
rect 12575 9636 12587 9639
rect 12618 9636 12624 9648
rect 12575 9608 12624 9636
rect 12575 9605 12587 9608
rect 12529 9599 12587 9605
rect 12618 9596 12624 9608
rect 12676 9596 12682 9648
rect 13814 9636 13820 9648
rect 13280 9608 13820 9636
rect 934 9528 940 9580
rect 992 9568 998 9580
rect 13280 9577 13308 9608
rect 13814 9596 13820 9608
rect 13872 9596 13878 9648
rect 15010 9596 15016 9648
rect 15068 9636 15074 9648
rect 15289 9639 15347 9645
rect 15289 9636 15301 9639
rect 15068 9608 15301 9636
rect 15068 9596 15074 9608
rect 15289 9605 15301 9608
rect 15335 9605 15347 9639
rect 15289 9599 15347 9605
rect 16132 9636 16160 9664
rect 16666 9636 16672 9648
rect 16132 9608 16672 9636
rect 1581 9571 1639 9577
rect 1581 9568 1593 9571
rect 992 9540 1593 9568
rect 992 9528 998 9540
rect 1581 9537 1593 9540
rect 1627 9537 1639 9571
rect 1581 9531 1639 9537
rect 13265 9571 13323 9577
rect 13265 9537 13277 9571
rect 13311 9537 13323 9571
rect 16132 9568 16160 9608
rect 16666 9596 16672 9608
rect 16724 9596 16730 9648
rect 14674 9540 16160 9568
rect 13265 9531 13323 9537
rect 12710 9460 12716 9512
rect 12768 9460 12774 9512
rect 13541 9503 13599 9509
rect 13541 9469 13553 9503
rect 13587 9500 13599 9503
rect 15194 9500 15200 9512
rect 13587 9472 15200 9500
rect 13587 9469 13599 9472
rect 13541 9463 13599 9469
rect 15194 9460 15200 9472
rect 15252 9460 15258 9512
rect 1762 9392 1768 9444
rect 1820 9392 1826 9444
rect 12069 9435 12127 9441
rect 12069 9401 12081 9435
rect 12115 9432 12127 9435
rect 12802 9432 12808 9444
rect 12115 9404 12808 9432
rect 12115 9401 12127 9404
rect 12069 9395 12127 9401
rect 12802 9392 12808 9404
rect 12860 9392 12866 9444
rect 12158 9324 12164 9376
rect 12216 9364 12222 9376
rect 16776 9364 16804 9676
rect 25590 9664 25596 9676
rect 25648 9664 25654 9716
rect 25685 9707 25743 9713
rect 25685 9673 25697 9707
rect 25731 9673 25743 9707
rect 25685 9667 25743 9673
rect 28184 9676 29132 9704
rect 18874 9596 18880 9648
rect 18932 9596 18938 9648
rect 19610 9596 19616 9648
rect 19668 9596 19674 9648
rect 21082 9636 21088 9648
rect 20838 9608 21088 9636
rect 21082 9596 21088 9608
rect 21140 9596 21146 9648
rect 22554 9596 22560 9648
rect 22612 9636 22618 9648
rect 22741 9639 22799 9645
rect 22741 9636 22753 9639
rect 22612 9608 22753 9636
rect 22612 9596 22618 9608
rect 22741 9605 22753 9608
rect 22787 9605 22799 9639
rect 22741 9599 22799 9605
rect 23566 9596 23572 9648
rect 23624 9636 23630 9648
rect 23937 9639 23995 9645
rect 23937 9636 23949 9639
rect 23624 9608 23949 9636
rect 23624 9596 23630 9608
rect 23937 9605 23949 9608
rect 23983 9605 23995 9639
rect 25700 9636 25728 9667
rect 28184 9636 28212 9676
rect 25700 9608 28212 9636
rect 29104 9636 29132 9676
rect 29270 9664 29276 9716
rect 29328 9664 29334 9716
rect 30374 9664 30380 9716
rect 30432 9664 30438 9716
rect 30650 9664 30656 9716
rect 30708 9704 30714 9716
rect 31294 9704 31300 9716
rect 30708 9676 31300 9704
rect 30708 9664 30714 9676
rect 31294 9664 31300 9676
rect 31352 9664 31358 9716
rect 31386 9664 31392 9716
rect 31444 9704 31450 9716
rect 38746 9704 38752 9716
rect 31444 9676 38752 9704
rect 31444 9664 31450 9676
rect 38746 9664 38752 9676
rect 38804 9664 38810 9716
rect 30392 9636 30420 9664
rect 32030 9636 32036 9648
rect 29104 9608 30420 9636
rect 31234 9608 32036 9636
rect 23937 9599 23995 9605
rect 32030 9596 32036 9608
rect 32088 9596 32094 9648
rect 32214 9596 32220 9648
rect 32272 9636 32278 9648
rect 32953 9639 33011 9645
rect 32953 9636 32965 9639
rect 32272 9608 32965 9636
rect 32272 9596 32278 9608
rect 32953 9605 32965 9608
rect 32999 9605 33011 9639
rect 35618 9636 35624 9648
rect 35374 9608 35624 9636
rect 32953 9599 33011 9605
rect 35618 9596 35624 9608
rect 35676 9596 35682 9648
rect 49145 9639 49203 9645
rect 49145 9605 49157 9639
rect 49191 9636 49203 9639
rect 49326 9636 49332 9648
rect 49191 9608 49332 9636
rect 49191 9605 49203 9608
rect 49145 9599 49203 9605
rect 49326 9596 49332 9608
rect 49384 9596 49390 9648
rect 18230 9528 18236 9580
rect 18288 9528 18294 9580
rect 20990 9528 20996 9580
rect 21048 9568 21054 9580
rect 22649 9571 22707 9577
rect 22649 9568 22661 9571
rect 21048 9540 22661 9568
rect 21048 9528 21054 9540
rect 22649 9537 22661 9540
rect 22695 9568 22707 9571
rect 22695 9540 23612 9568
rect 22695 9537 22707 9540
rect 22649 9531 22707 9537
rect 16850 9460 16856 9512
rect 16908 9460 16914 9512
rect 17129 9503 17187 9509
rect 17129 9469 17141 9503
rect 17175 9500 17187 9503
rect 18598 9500 18604 9512
rect 17175 9472 18604 9500
rect 17175 9469 17187 9472
rect 17129 9463 17187 9469
rect 18598 9460 18604 9472
rect 18656 9460 18662 9512
rect 19337 9503 19395 9509
rect 19337 9469 19349 9503
rect 19383 9469 19395 9503
rect 19337 9463 19395 9469
rect 12216 9336 16804 9364
rect 12216 9324 12222 9336
rect 16850 9324 16856 9376
rect 16908 9364 16914 9376
rect 19352 9364 19380 9463
rect 20806 9460 20812 9512
rect 20864 9500 20870 9512
rect 21085 9503 21143 9509
rect 21085 9500 21097 9503
rect 20864 9472 21097 9500
rect 20864 9460 20870 9472
rect 21085 9469 21097 9472
rect 21131 9500 21143 9503
rect 22833 9503 22891 9509
rect 21131 9472 22094 9500
rect 21131 9469 21143 9472
rect 21085 9463 21143 9469
rect 22066 9432 22094 9472
rect 22833 9469 22845 9503
rect 22879 9469 22891 9503
rect 22833 9463 22891 9469
rect 22848 9432 22876 9463
rect 22066 9404 22876 9432
rect 16908 9336 19380 9364
rect 16908 9324 16914 9336
rect 20898 9324 20904 9376
rect 20956 9364 20962 9376
rect 23584 9373 23612 9540
rect 23658 9528 23664 9580
rect 23716 9528 23722 9580
rect 25038 9528 25044 9580
rect 25096 9568 25102 9580
rect 25314 9568 25320 9580
rect 25096 9540 25320 9568
rect 25096 9528 25102 9540
rect 25314 9528 25320 9540
rect 25372 9528 25378 9580
rect 26050 9528 26056 9580
rect 26108 9528 26114 9580
rect 26142 9528 26148 9580
rect 26200 9528 26206 9580
rect 28902 9528 28908 9580
rect 28960 9568 28966 9580
rect 29638 9568 29644 9580
rect 28960 9540 29644 9568
rect 28960 9528 28966 9540
rect 29638 9528 29644 9540
rect 29696 9528 29702 9580
rect 31294 9528 31300 9580
rect 31352 9568 31358 9580
rect 31352 9540 32444 9568
rect 31352 9528 31358 9540
rect 26329 9503 26387 9509
rect 26329 9469 26341 9503
rect 26375 9500 26387 9503
rect 26878 9500 26884 9512
rect 26375 9472 26884 9500
rect 26375 9469 26387 9472
rect 26329 9463 26387 9469
rect 26878 9460 26884 9472
rect 26936 9460 26942 9512
rect 26970 9460 26976 9512
rect 27028 9500 27034 9512
rect 27525 9503 27583 9509
rect 27525 9500 27537 9503
rect 27028 9472 27537 9500
rect 27028 9460 27034 9472
rect 27525 9469 27537 9472
rect 27571 9469 27583 9503
rect 27525 9463 27583 9469
rect 27801 9503 27859 9509
rect 27801 9469 27813 9503
rect 27847 9500 27859 9503
rect 27847 9472 28856 9500
rect 27847 9469 27859 9472
rect 27801 9463 27859 9469
rect 26786 9432 26792 9444
rect 25332 9404 26792 9432
rect 22281 9367 22339 9373
rect 22281 9364 22293 9367
rect 20956 9336 22293 9364
rect 20956 9324 20962 9336
rect 22281 9333 22293 9336
rect 22327 9333 22339 9367
rect 22281 9327 22339 9333
rect 23569 9367 23627 9373
rect 23569 9333 23581 9367
rect 23615 9364 23627 9367
rect 25332 9364 25360 9404
rect 26786 9392 26792 9404
rect 26844 9392 26850 9444
rect 23615 9336 25360 9364
rect 23615 9333 23627 9336
rect 23569 9327 23627 9333
rect 25406 9324 25412 9376
rect 25464 9324 25470 9376
rect 27540 9364 27568 9463
rect 28828 9432 28856 9472
rect 29730 9460 29736 9512
rect 29788 9460 29794 9512
rect 30006 9460 30012 9512
rect 30064 9460 30070 9512
rect 30098 9460 30104 9512
rect 30156 9500 30162 9512
rect 32306 9500 32312 9512
rect 30156 9472 32312 9500
rect 30156 9460 30162 9472
rect 32306 9460 32312 9472
rect 32364 9460 32370 9512
rect 32416 9432 32444 9540
rect 32490 9528 32496 9580
rect 32548 9568 32554 9580
rect 33045 9571 33103 9577
rect 33045 9568 33057 9571
rect 32548 9540 33057 9568
rect 32548 9528 32554 9540
rect 33045 9537 33057 9540
rect 33091 9537 33103 9571
rect 33045 9531 33103 9537
rect 33502 9528 33508 9580
rect 33560 9568 33566 9580
rect 33873 9571 33931 9577
rect 33873 9568 33885 9571
rect 33560 9540 33885 9568
rect 33560 9528 33566 9540
rect 33873 9537 33885 9540
rect 33919 9537 33931 9571
rect 33873 9531 33931 9537
rect 47026 9528 47032 9580
rect 47084 9568 47090 9580
rect 47949 9571 48007 9577
rect 47949 9568 47961 9571
rect 47084 9540 47961 9568
rect 47084 9528 47090 9540
rect 47949 9537 47961 9540
rect 47995 9537 48007 9571
rect 47949 9531 48007 9537
rect 33137 9503 33195 9509
rect 33137 9469 33149 9503
rect 33183 9469 33195 9503
rect 33137 9463 33195 9469
rect 33152 9432 33180 9463
rect 33686 9460 33692 9512
rect 33744 9500 33750 9512
rect 34149 9503 34207 9509
rect 34149 9500 34161 9503
rect 33744 9472 34161 9500
rect 33744 9460 33750 9472
rect 33888 9444 33916 9472
rect 34149 9469 34161 9472
rect 34195 9500 34207 9503
rect 37458 9500 37464 9512
rect 34195 9472 37464 9500
rect 34195 9469 34207 9472
rect 34149 9463 34207 9469
rect 37458 9460 37464 9472
rect 37516 9460 37522 9512
rect 28828 9404 29868 9432
rect 32416 9404 33180 9432
rect 29730 9364 29736 9376
rect 27540 9336 29736 9364
rect 29730 9324 29736 9336
rect 29788 9324 29794 9376
rect 29840 9364 29868 9404
rect 33870 9392 33876 9444
rect 33928 9392 33934 9444
rect 35158 9392 35164 9444
rect 35216 9432 35222 9444
rect 35621 9435 35679 9441
rect 35621 9432 35633 9435
rect 35216 9404 35633 9432
rect 35216 9392 35222 9404
rect 35621 9401 35633 9404
rect 35667 9401 35679 9435
rect 35621 9395 35679 9401
rect 31481 9367 31539 9373
rect 31481 9364 31493 9367
rect 29840 9336 31493 9364
rect 31481 9333 31493 9336
rect 31527 9364 31539 9367
rect 32398 9364 32404 9376
rect 31527 9336 32404 9364
rect 31527 9333 31539 9336
rect 31481 9327 31539 9333
rect 32398 9324 32404 9336
rect 32456 9324 32462 9376
rect 32585 9367 32643 9373
rect 32585 9333 32597 9367
rect 32631 9364 32643 9367
rect 35526 9364 35532 9376
rect 32631 9336 35532 9364
rect 32631 9333 32643 9336
rect 32585 9327 32643 9333
rect 35526 9324 35532 9336
rect 35584 9324 35590 9376
rect 1104 9274 49864 9296
rect 1104 9222 2950 9274
rect 3002 9222 3014 9274
rect 3066 9222 3078 9274
rect 3130 9222 3142 9274
rect 3194 9222 3206 9274
rect 3258 9222 12950 9274
rect 13002 9222 13014 9274
rect 13066 9222 13078 9274
rect 13130 9222 13142 9274
rect 13194 9222 13206 9274
rect 13258 9222 22950 9274
rect 23002 9222 23014 9274
rect 23066 9222 23078 9274
rect 23130 9222 23142 9274
rect 23194 9222 23206 9274
rect 23258 9222 32950 9274
rect 33002 9222 33014 9274
rect 33066 9222 33078 9274
rect 33130 9222 33142 9274
rect 33194 9222 33206 9274
rect 33258 9222 42950 9274
rect 43002 9222 43014 9274
rect 43066 9222 43078 9274
rect 43130 9222 43142 9274
rect 43194 9222 43206 9274
rect 43258 9222 49864 9274
rect 1104 9200 49864 9222
rect 1765 9163 1823 9169
rect 1765 9129 1777 9163
rect 1811 9160 1823 9163
rect 12158 9160 12164 9172
rect 1811 9132 12164 9160
rect 1811 9129 1823 9132
rect 1765 9123 1823 9129
rect 12158 9120 12164 9132
rect 12216 9120 12222 9172
rect 14366 9120 14372 9172
rect 14424 9120 14430 9172
rect 15102 9120 15108 9172
rect 15160 9160 15166 9172
rect 17034 9160 17040 9172
rect 15160 9132 17040 9160
rect 15160 9120 15166 9132
rect 17034 9120 17040 9132
rect 17092 9120 17098 9172
rect 17862 9120 17868 9172
rect 17920 9160 17926 9172
rect 18049 9163 18107 9169
rect 18049 9160 18061 9163
rect 17920 9132 18061 9160
rect 17920 9120 17926 9132
rect 18049 9129 18061 9132
rect 18095 9129 18107 9163
rect 18049 9123 18107 9129
rect 18877 9163 18935 9169
rect 18877 9129 18889 9163
rect 18923 9160 18935 9163
rect 18966 9160 18972 9172
rect 18923 9132 18972 9160
rect 18923 9129 18935 9132
rect 18877 9123 18935 9129
rect 18966 9120 18972 9132
rect 19024 9120 19030 9172
rect 22278 9120 22284 9172
rect 22336 9160 22342 9172
rect 24029 9163 24087 9169
rect 24029 9160 24041 9163
rect 22336 9132 24041 9160
rect 22336 9120 22342 9132
rect 24029 9129 24041 9132
rect 24075 9129 24087 9163
rect 24029 9123 24087 9129
rect 27062 9120 27068 9172
rect 27120 9160 27126 9172
rect 27706 9160 27712 9172
rect 27120 9132 27712 9160
rect 27120 9120 27126 9132
rect 27706 9120 27712 9132
rect 27764 9120 27770 9172
rect 28169 9163 28227 9169
rect 28169 9129 28181 9163
rect 28215 9160 28227 9163
rect 32674 9160 32680 9172
rect 28215 9132 32680 9160
rect 28215 9129 28227 9132
rect 28169 9123 28227 9129
rect 32674 9120 32680 9132
rect 32732 9120 32738 9172
rect 33321 9163 33379 9169
rect 33321 9129 33333 9163
rect 33367 9160 33379 9163
rect 37274 9160 37280 9172
rect 33367 9132 37280 9160
rect 33367 9129 33379 9132
rect 33321 9123 33379 9129
rect 37274 9120 37280 9132
rect 37332 9120 37338 9172
rect 14550 9052 14556 9104
rect 14608 9092 14614 9104
rect 14608 9064 15056 9092
rect 14608 9052 14614 9064
rect 14826 8984 14832 9036
rect 14884 8984 14890 9036
rect 15028 9033 15056 9064
rect 23842 9052 23848 9104
rect 23900 9092 23906 9104
rect 24581 9095 24639 9101
rect 24581 9092 24593 9095
rect 23900 9064 24593 9092
rect 23900 9052 23906 9064
rect 24581 9061 24593 9064
rect 24627 9061 24639 9095
rect 24581 9055 24639 9061
rect 26142 9052 26148 9104
rect 26200 9092 26206 9104
rect 30098 9092 30104 9104
rect 26200 9064 30104 9092
rect 26200 9052 26206 9064
rect 30098 9052 30104 9064
rect 30156 9052 30162 9104
rect 32306 9052 32312 9104
rect 32364 9092 32370 9104
rect 34974 9092 34980 9104
rect 32364 9064 34980 9092
rect 32364 9052 32370 9064
rect 34974 9052 34980 9064
rect 35032 9092 35038 9104
rect 35618 9092 35624 9104
rect 35032 9064 35624 9092
rect 35032 9052 35038 9064
rect 35618 9052 35624 9064
rect 35676 9052 35682 9104
rect 36633 9095 36691 9101
rect 36633 9061 36645 9095
rect 36679 9092 36691 9095
rect 36679 9064 41414 9092
rect 36679 9061 36691 9064
rect 36633 9055 36691 9061
rect 15013 9027 15071 9033
rect 15013 8993 15025 9027
rect 15059 8993 15071 9027
rect 15013 8987 15071 8993
rect 18506 8984 18512 9036
rect 18564 9024 18570 9036
rect 20990 9024 20996 9036
rect 18564 8996 20996 9024
rect 18564 8984 18570 8996
rect 20990 8984 20996 8996
rect 21048 8984 21054 9036
rect 22002 8984 22008 9036
rect 22060 9024 22066 9036
rect 22281 9027 22339 9033
rect 22281 9024 22293 9027
rect 22060 8996 22293 9024
rect 22060 8984 22066 8996
rect 22281 8993 22293 8996
rect 22327 8993 22339 9027
rect 22281 8987 22339 8993
rect 22557 9027 22615 9033
rect 22557 8993 22569 9027
rect 22603 9024 22615 9027
rect 25133 9027 25191 9033
rect 25133 9024 25145 9027
rect 22603 8996 25145 9024
rect 22603 8993 22615 8996
rect 22557 8987 22615 8993
rect 25133 8993 25145 8996
rect 25179 9024 25191 9027
rect 25406 9024 25412 9036
rect 25179 8996 25412 9024
rect 25179 8993 25191 8996
rect 25133 8987 25191 8993
rect 25406 8984 25412 8996
rect 25464 8984 25470 9036
rect 28813 9027 28871 9033
rect 28813 8993 28825 9027
rect 28859 9024 28871 9027
rect 30006 9024 30012 9036
rect 28859 8996 30012 9024
rect 28859 8993 28871 8996
rect 28813 8987 28871 8993
rect 30006 8984 30012 8996
rect 30064 8984 30070 9036
rect 31021 9027 31079 9033
rect 31021 8993 31033 9027
rect 31067 9024 31079 9027
rect 31067 8996 33824 9024
rect 31067 8993 31079 8996
rect 31021 8987 31079 8993
rect 934 8916 940 8968
rect 992 8956 998 8968
rect 1581 8959 1639 8965
rect 1581 8956 1593 8959
rect 992 8928 1593 8956
rect 992 8916 998 8928
rect 1581 8925 1593 8928
rect 1627 8925 1639 8959
rect 1581 8919 1639 8925
rect 2317 8959 2375 8965
rect 2317 8925 2329 8959
rect 2363 8925 2375 8959
rect 2317 8919 2375 8925
rect 1210 8848 1216 8900
rect 1268 8888 1274 8900
rect 2332 8888 2360 8919
rect 13538 8916 13544 8968
rect 13596 8956 13602 8968
rect 13725 8959 13783 8965
rect 13725 8956 13737 8959
rect 13596 8928 13737 8956
rect 13596 8916 13602 8928
rect 13725 8925 13737 8928
rect 13771 8925 13783 8959
rect 13725 8919 13783 8925
rect 13814 8916 13820 8968
rect 13872 8956 13878 8968
rect 16301 8959 16359 8965
rect 16301 8956 16313 8959
rect 13872 8928 16313 8956
rect 13872 8916 13878 8928
rect 16301 8925 16313 8928
rect 16347 8925 16359 8959
rect 16301 8919 16359 8925
rect 16206 8888 16212 8900
rect 1268 8860 2360 8888
rect 12406 8860 16212 8888
rect 1268 8848 1274 8860
rect 2501 8823 2559 8829
rect 2501 8789 2513 8823
rect 2547 8820 2559 8823
rect 12406 8820 12434 8860
rect 16206 8848 16212 8860
rect 16264 8848 16270 8900
rect 2547 8792 12434 8820
rect 13541 8823 13599 8829
rect 2547 8789 2559 8792
rect 2501 8783 2559 8789
rect 13541 8789 13553 8823
rect 13587 8820 13599 8823
rect 14550 8820 14556 8832
rect 13587 8792 14556 8820
rect 13587 8789 13599 8792
rect 13541 8783 13599 8789
rect 14550 8780 14556 8792
rect 14608 8780 14614 8832
rect 14734 8780 14740 8832
rect 14792 8820 14798 8832
rect 15102 8820 15108 8832
rect 14792 8792 15108 8820
rect 14792 8780 14798 8792
rect 15102 8780 15108 8792
rect 15160 8780 15166 8832
rect 16316 8820 16344 8919
rect 19426 8916 19432 8968
rect 19484 8916 19490 8968
rect 21821 8959 21879 8965
rect 21821 8925 21833 8959
rect 21867 8956 21879 8959
rect 22186 8956 22192 8968
rect 21867 8928 22192 8956
rect 21867 8925 21879 8928
rect 21821 8919 21879 8925
rect 22186 8916 22192 8928
rect 22244 8916 22250 8968
rect 28537 8959 28595 8965
rect 28537 8925 28549 8959
rect 28583 8956 28595 8959
rect 29917 8959 29975 8965
rect 29917 8956 29929 8959
rect 28583 8928 29929 8956
rect 28583 8925 28595 8928
rect 28537 8919 28595 8925
rect 29917 8925 29929 8928
rect 29963 8925 29975 8959
rect 29917 8919 29975 8925
rect 30742 8916 30748 8968
rect 30800 8916 30806 8968
rect 32030 8916 32036 8968
rect 32088 8956 32094 8968
rect 32088 8928 32154 8956
rect 32088 8916 32094 8928
rect 33594 8916 33600 8968
rect 33652 8956 33658 8968
rect 33689 8959 33747 8965
rect 33689 8956 33701 8959
rect 33652 8928 33701 8956
rect 33652 8916 33658 8928
rect 33689 8925 33701 8928
rect 33735 8925 33747 8959
rect 33796 8956 33824 8996
rect 33870 8984 33876 9036
rect 33928 8984 33934 9036
rect 34422 8984 34428 9036
rect 34480 9024 34486 9036
rect 35345 9027 35403 9033
rect 35345 9024 35357 9027
rect 34480 8996 35357 9024
rect 34480 8984 34486 8996
rect 35345 8993 35357 8996
rect 35391 8993 35403 9027
rect 35345 8987 35403 8993
rect 35437 9027 35495 9033
rect 35437 8993 35449 9027
rect 35483 8993 35495 9027
rect 35437 8987 35495 8993
rect 34054 8956 34060 8968
rect 33796 8928 34060 8956
rect 33689 8919 33747 8925
rect 34054 8916 34060 8928
rect 34112 8956 34118 8968
rect 35452 8956 35480 8987
rect 35526 8984 35532 9036
rect 35584 9024 35590 9036
rect 39485 9027 39543 9033
rect 35584 8996 37872 9024
rect 35584 8984 35590 8996
rect 37844 8965 37872 8996
rect 39485 8993 39497 9027
rect 39531 9024 39543 9027
rect 39531 8996 40448 9024
rect 39531 8993 39543 8996
rect 39485 8987 39543 8993
rect 34112 8928 35480 8956
rect 36817 8959 36875 8965
rect 34112 8916 34118 8928
rect 36817 8925 36829 8959
rect 36863 8925 36875 8959
rect 36817 8919 36875 8925
rect 37829 8959 37887 8965
rect 37829 8925 37841 8959
rect 37875 8925 37887 8959
rect 37829 8919 37887 8925
rect 16574 8848 16580 8900
rect 16632 8848 16638 8900
rect 16666 8848 16672 8900
rect 16724 8888 16730 8900
rect 18230 8888 18236 8900
rect 16724 8860 16988 8888
rect 17802 8860 18236 8888
rect 16724 8848 16730 8860
rect 16850 8820 16856 8832
rect 16316 8792 16856 8820
rect 16850 8780 16856 8792
rect 16908 8780 16914 8832
rect 16960 8820 16988 8860
rect 17880 8820 17908 8860
rect 18230 8848 18236 8860
rect 18288 8888 18294 8900
rect 18414 8888 18420 8900
rect 18288 8860 18420 8888
rect 18288 8848 18294 8860
rect 18414 8848 18420 8860
rect 18472 8848 18478 8900
rect 19702 8848 19708 8900
rect 19760 8848 19766 8900
rect 21082 8888 21088 8900
rect 20930 8860 21088 8888
rect 21082 8848 21088 8860
rect 21140 8848 21146 8900
rect 23290 8848 23296 8900
rect 23348 8848 23354 8900
rect 25041 8891 25099 8897
rect 25041 8857 25053 8891
rect 25087 8888 25099 8891
rect 25130 8888 25136 8900
rect 25087 8860 25136 8888
rect 25087 8857 25099 8860
rect 25041 8851 25099 8857
rect 25130 8848 25136 8860
rect 25188 8848 25194 8900
rect 32858 8848 32864 8900
rect 32916 8888 32922 8900
rect 36832 8888 36860 8919
rect 39301 8891 39359 8897
rect 39301 8888 39313 8891
rect 32916 8860 36860 8888
rect 36924 8860 39313 8888
rect 32916 8848 32922 8860
rect 16960 8792 17908 8820
rect 19610 8780 19616 8832
rect 19668 8820 19674 8832
rect 21177 8823 21235 8829
rect 21177 8820 21189 8823
rect 19668 8792 21189 8820
rect 19668 8780 19674 8792
rect 21177 8789 21189 8792
rect 21223 8789 21235 8823
rect 21177 8783 21235 8789
rect 24946 8780 24952 8832
rect 25004 8780 25010 8832
rect 27614 8780 27620 8832
rect 27672 8820 27678 8832
rect 28626 8820 28632 8832
rect 27672 8792 28632 8820
rect 27672 8780 27678 8792
rect 28626 8780 28632 8792
rect 28684 8780 28690 8832
rect 30006 8780 30012 8832
rect 30064 8820 30070 8832
rect 32493 8823 32551 8829
rect 32493 8820 32505 8823
rect 30064 8792 32505 8820
rect 30064 8780 30070 8792
rect 32493 8789 32505 8792
rect 32539 8789 32551 8823
rect 32493 8783 32551 8789
rect 33778 8780 33784 8832
rect 33836 8780 33842 8832
rect 34882 8780 34888 8832
rect 34940 8780 34946 8832
rect 35250 8780 35256 8832
rect 35308 8780 35314 8832
rect 35618 8780 35624 8832
rect 35676 8820 35682 8832
rect 36924 8820 36952 8860
rect 39301 8857 39313 8860
rect 39347 8857 39359 8891
rect 40420 8888 40448 8996
rect 41386 8956 41414 9064
rect 49145 9027 49203 9033
rect 49145 8993 49157 9027
rect 49191 9024 49203 9027
rect 49234 9024 49240 9036
rect 49191 8996 49240 9024
rect 49191 8993 49203 8996
rect 49145 8987 49203 8993
rect 49234 8984 49240 8996
rect 49292 8984 49298 9036
rect 43622 8956 43628 8968
rect 41386 8928 43628 8956
rect 43622 8916 43628 8928
rect 43680 8916 43686 8968
rect 44174 8916 44180 8968
rect 44232 8956 44238 8968
rect 47949 8959 48007 8965
rect 47949 8956 47961 8959
rect 44232 8928 47961 8956
rect 44232 8916 44238 8928
rect 47949 8925 47961 8928
rect 47995 8925 48007 8959
rect 47949 8919 48007 8925
rect 46566 8888 46572 8900
rect 40420 8860 46572 8888
rect 39301 8851 39359 8857
rect 46566 8848 46572 8860
rect 46624 8848 46630 8900
rect 35676 8792 36952 8820
rect 37645 8823 37703 8829
rect 35676 8780 35682 8792
rect 37645 8789 37657 8823
rect 37691 8820 37703 8823
rect 44266 8820 44272 8832
rect 37691 8792 44272 8820
rect 37691 8789 37703 8792
rect 37645 8783 37703 8789
rect 44266 8780 44272 8792
rect 44324 8780 44330 8832
rect 1104 8730 49864 8752
rect 1104 8678 7950 8730
rect 8002 8678 8014 8730
rect 8066 8678 8078 8730
rect 8130 8678 8142 8730
rect 8194 8678 8206 8730
rect 8258 8678 17950 8730
rect 18002 8678 18014 8730
rect 18066 8678 18078 8730
rect 18130 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 27950 8730
rect 28002 8678 28014 8730
rect 28066 8678 28078 8730
rect 28130 8678 28142 8730
rect 28194 8678 28206 8730
rect 28258 8678 37950 8730
rect 38002 8678 38014 8730
rect 38066 8678 38078 8730
rect 38130 8678 38142 8730
rect 38194 8678 38206 8730
rect 38258 8678 47950 8730
rect 48002 8678 48014 8730
rect 48066 8678 48078 8730
rect 48130 8678 48142 8730
rect 48194 8678 48206 8730
rect 48258 8678 49864 8730
rect 1104 8656 49864 8678
rect 14642 8576 14648 8628
rect 14700 8616 14706 8628
rect 14700 8588 15240 8616
rect 14700 8576 14706 8588
rect 13814 8548 13820 8560
rect 13556 8520 13820 8548
rect 1854 8440 1860 8492
rect 1912 8440 1918 8492
rect 13556 8489 13584 8520
rect 13814 8508 13820 8520
rect 13872 8508 13878 8560
rect 15212 8548 15240 8588
rect 15286 8576 15292 8628
rect 15344 8576 15350 8628
rect 18506 8616 18512 8628
rect 17512 8588 18512 8616
rect 17512 8548 17540 8588
rect 18506 8576 18512 8588
rect 18564 8576 18570 8628
rect 18598 8576 18604 8628
rect 18656 8576 18662 8628
rect 19978 8576 19984 8628
rect 20036 8616 20042 8628
rect 21453 8619 21511 8625
rect 21453 8616 21465 8619
rect 20036 8588 21465 8616
rect 20036 8576 20042 8588
rect 21453 8585 21465 8588
rect 21499 8585 21511 8619
rect 21453 8579 21511 8585
rect 30561 8619 30619 8625
rect 30561 8585 30573 8619
rect 30607 8616 30619 8619
rect 30650 8616 30656 8628
rect 30607 8588 30656 8616
rect 30607 8585 30619 8588
rect 30561 8579 30619 8585
rect 30650 8576 30656 8588
rect 30708 8576 30714 8628
rect 31021 8619 31079 8625
rect 31021 8585 31033 8619
rect 31067 8616 31079 8619
rect 31662 8616 31668 8628
rect 31067 8588 31668 8616
rect 31067 8585 31079 8588
rect 31021 8579 31079 8585
rect 31662 8576 31668 8588
rect 31720 8576 31726 8628
rect 33502 8616 33508 8628
rect 32324 8588 33508 8616
rect 20254 8548 20260 8560
rect 15212 8520 17540 8548
rect 19720 8520 20260 8548
rect 13541 8483 13599 8489
rect 13541 8449 13553 8483
rect 13587 8449 13599 8483
rect 16666 8480 16672 8492
rect 14950 8452 16672 8480
rect 13541 8443 13599 8449
rect 16666 8440 16672 8452
rect 16724 8440 16730 8492
rect 16850 8440 16856 8492
rect 16908 8440 16914 8492
rect 1578 8372 1584 8424
rect 1636 8372 1642 8424
rect 13817 8415 13875 8421
rect 13817 8412 13829 8415
rect 13556 8384 13829 8412
rect 13556 8356 13584 8384
rect 13817 8381 13829 8384
rect 13863 8381 13875 8415
rect 13817 8375 13875 8381
rect 14550 8372 14556 8424
rect 14608 8412 14614 8424
rect 16390 8412 16396 8424
rect 14608 8384 16396 8412
rect 14608 8372 14614 8384
rect 16390 8372 16396 8384
rect 16448 8372 16454 8424
rect 17129 8415 17187 8421
rect 17129 8381 17141 8415
rect 17175 8412 17187 8415
rect 17862 8412 17868 8424
rect 17175 8384 17868 8412
rect 17175 8381 17187 8384
rect 17129 8375 17187 8381
rect 17862 8372 17868 8384
rect 17920 8372 17926 8424
rect 13538 8304 13544 8356
rect 13596 8304 13602 8356
rect 18248 8344 18276 8466
rect 19150 8440 19156 8492
rect 19208 8480 19214 8492
rect 19245 8483 19303 8489
rect 19245 8480 19257 8483
rect 19208 8452 19257 8480
rect 19208 8440 19214 8452
rect 19245 8449 19257 8452
rect 19291 8449 19303 8483
rect 19245 8443 19303 8449
rect 19426 8440 19432 8492
rect 19484 8480 19490 8492
rect 19720 8489 19748 8520
rect 20254 8508 20260 8520
rect 20312 8508 20318 8560
rect 22278 8508 22284 8560
rect 22336 8508 22342 8560
rect 29086 8508 29092 8560
rect 29144 8508 29150 8560
rect 29638 8508 29644 8560
rect 29696 8508 29702 8560
rect 30742 8508 30748 8560
rect 30800 8548 30806 8560
rect 30800 8520 31754 8548
rect 30800 8508 30806 8520
rect 19705 8483 19763 8489
rect 19705 8480 19717 8483
rect 19484 8452 19717 8480
rect 19484 8440 19490 8452
rect 19705 8449 19717 8452
rect 19751 8449 19763 8483
rect 19705 8443 19763 8449
rect 21082 8440 21088 8492
rect 21140 8440 21146 8492
rect 22002 8440 22008 8492
rect 22060 8440 22066 8492
rect 23382 8440 23388 8492
rect 23440 8480 23446 8492
rect 25038 8480 25044 8492
rect 23440 8452 25044 8480
rect 23440 8440 23446 8452
rect 25038 8440 25044 8452
rect 25096 8440 25102 8492
rect 31386 8440 31392 8492
rect 31444 8440 31450 8492
rect 31726 8480 31754 8520
rect 32324 8489 32352 8588
rect 33502 8576 33508 8588
rect 33560 8576 33566 8628
rect 34054 8576 34060 8628
rect 34112 8576 34118 8628
rect 37461 8619 37519 8625
rect 37461 8585 37473 8619
rect 37507 8616 37519 8619
rect 40218 8616 40224 8628
rect 37507 8588 40224 8616
rect 37507 8585 37519 8588
rect 37461 8579 37519 8585
rect 40218 8576 40224 8588
rect 40276 8576 40282 8628
rect 40405 8619 40463 8625
rect 40405 8585 40417 8619
rect 40451 8616 40463 8619
rect 47670 8616 47676 8628
rect 40451 8588 47676 8616
rect 40451 8585 40463 8588
rect 40405 8579 40463 8585
rect 47670 8576 47676 8588
rect 47728 8576 47734 8628
rect 32582 8508 32588 8560
rect 32640 8508 32646 8560
rect 34514 8548 34520 8560
rect 33810 8520 34520 8548
rect 34514 8508 34520 8520
rect 34572 8508 34578 8560
rect 34882 8508 34888 8560
rect 34940 8548 34946 8560
rect 34940 8520 39160 8548
rect 34940 8508 34946 8520
rect 32309 8483 32367 8489
rect 32309 8480 32321 8483
rect 31726 8452 32321 8480
rect 32309 8449 32321 8452
rect 32355 8449 32367 8483
rect 32309 8443 32367 8449
rect 34330 8440 34336 8492
rect 34388 8480 34394 8492
rect 39132 8489 39160 8520
rect 44266 8508 44272 8560
rect 44324 8508 44330 8560
rect 49142 8508 49148 8560
rect 49200 8508 49206 8560
rect 37645 8483 37703 8489
rect 37645 8480 37657 8483
rect 34388 8452 37657 8480
rect 34388 8440 34394 8452
rect 37645 8449 37657 8452
rect 37691 8449 37703 8483
rect 37645 8443 37703 8449
rect 39117 8483 39175 8489
rect 39117 8449 39129 8483
rect 39163 8449 39175 8483
rect 39117 8443 39175 8449
rect 40313 8483 40371 8489
rect 40313 8449 40325 8483
rect 40359 8449 40371 8483
rect 40313 8443 40371 8449
rect 19981 8415 20039 8421
rect 19981 8381 19993 8415
rect 20027 8412 20039 8415
rect 20027 8384 22094 8412
rect 20027 8381 20039 8384
rect 19981 8375 20039 8381
rect 18414 8344 18420 8356
rect 18248 8316 18420 8344
rect 18414 8304 18420 8316
rect 18472 8344 18478 8356
rect 18472 8316 19472 8344
rect 18472 8304 18478 8316
rect 19444 8276 19472 8316
rect 21082 8276 21088 8288
rect 19444 8248 21088 8276
rect 21082 8236 21088 8248
rect 21140 8236 21146 8288
rect 22066 8276 22094 8384
rect 28810 8372 28816 8424
rect 28868 8412 28874 8424
rect 29730 8412 29736 8424
rect 28868 8384 29736 8412
rect 28868 8372 28874 8384
rect 29730 8372 29736 8384
rect 29788 8372 29794 8424
rect 31481 8415 31539 8421
rect 31481 8381 31493 8415
rect 31527 8381 31539 8415
rect 31481 8375 31539 8381
rect 31665 8415 31723 8421
rect 31665 8381 31677 8415
rect 31711 8412 31723 8415
rect 33870 8412 33876 8424
rect 31711 8384 33876 8412
rect 31711 8381 31723 8384
rect 31665 8375 31723 8381
rect 23753 8347 23811 8353
rect 23753 8344 23765 8347
rect 23308 8316 23765 8344
rect 22646 8276 22652 8288
rect 22066 8248 22652 8276
rect 22646 8236 22652 8248
rect 22704 8276 22710 8288
rect 23308 8276 23336 8316
rect 23753 8313 23765 8316
rect 23799 8313 23811 8347
rect 23753 8307 23811 8313
rect 31496 8288 31524 8375
rect 33870 8372 33876 8384
rect 33928 8372 33934 8424
rect 34698 8372 34704 8424
rect 34756 8412 34762 8424
rect 35526 8412 35532 8424
rect 34756 8384 35532 8412
rect 34756 8372 34762 8384
rect 35526 8372 35532 8384
rect 35584 8412 35590 8424
rect 40328 8412 40356 8443
rect 42702 8440 42708 8492
rect 42760 8480 42766 8492
rect 45833 8483 45891 8489
rect 45833 8480 45845 8483
rect 42760 8452 45845 8480
rect 42760 8440 42766 8452
rect 45833 8449 45845 8452
rect 45879 8449 45891 8483
rect 45833 8443 45891 8449
rect 46750 8440 46756 8492
rect 46808 8480 46814 8492
rect 47949 8483 48007 8489
rect 47949 8480 47961 8483
rect 46808 8452 47961 8480
rect 46808 8440 46814 8452
rect 47949 8449 47961 8452
rect 47995 8449 48007 8483
rect 47949 8443 48007 8449
rect 35584 8384 40356 8412
rect 35584 8372 35590 8384
rect 46842 8372 46848 8424
rect 46900 8372 46906 8424
rect 38933 8347 38991 8353
rect 38933 8313 38945 8347
rect 38979 8344 38991 8347
rect 40126 8344 40132 8356
rect 38979 8316 40132 8344
rect 38979 8313 38991 8316
rect 38933 8307 38991 8313
rect 40126 8304 40132 8316
rect 40184 8304 40190 8356
rect 44453 8347 44511 8353
rect 44453 8313 44465 8347
rect 44499 8344 44511 8347
rect 47854 8344 47860 8356
rect 44499 8316 47860 8344
rect 44499 8313 44511 8316
rect 44453 8307 44511 8313
rect 47854 8304 47860 8316
rect 47912 8304 47918 8356
rect 22704 8248 23336 8276
rect 22704 8236 22710 8248
rect 31478 8236 31484 8288
rect 31536 8276 31542 8288
rect 38470 8276 38476 8288
rect 31536 8248 38476 8276
rect 31536 8236 31542 8248
rect 38470 8236 38476 8248
rect 38528 8236 38534 8288
rect 1104 8186 49864 8208
rect 1104 8134 2950 8186
rect 3002 8134 3014 8186
rect 3066 8134 3078 8186
rect 3130 8134 3142 8186
rect 3194 8134 3206 8186
rect 3258 8134 12950 8186
rect 13002 8134 13014 8186
rect 13066 8134 13078 8186
rect 13130 8134 13142 8186
rect 13194 8134 13206 8186
rect 13258 8134 22950 8186
rect 23002 8134 23014 8186
rect 23066 8134 23078 8186
rect 23130 8134 23142 8186
rect 23194 8134 23206 8186
rect 23258 8134 32950 8186
rect 33002 8134 33014 8186
rect 33066 8134 33078 8186
rect 33130 8134 33142 8186
rect 33194 8134 33206 8186
rect 33258 8134 42950 8186
rect 43002 8134 43014 8186
rect 43066 8134 43078 8186
rect 43130 8134 43142 8186
rect 43194 8134 43206 8186
rect 43258 8134 49864 8186
rect 1104 8112 49864 8134
rect 19702 8032 19708 8084
rect 19760 8072 19766 8084
rect 21177 8075 21235 8081
rect 21177 8072 21189 8075
rect 19760 8044 21189 8072
rect 19760 8032 19766 8044
rect 21177 8041 21189 8044
rect 21223 8041 21235 8075
rect 21177 8035 21235 8041
rect 21910 8032 21916 8084
rect 21968 8072 21974 8084
rect 22005 8075 22063 8081
rect 22005 8072 22017 8075
rect 21968 8044 22017 8072
rect 21968 8032 21974 8044
rect 22005 8041 22017 8044
rect 22051 8041 22063 8075
rect 22005 8035 22063 8041
rect 29914 8032 29920 8084
rect 29972 8032 29978 8084
rect 30561 8075 30619 8081
rect 30561 8041 30573 8075
rect 30607 8072 30619 8075
rect 35250 8072 35256 8084
rect 30607 8044 35256 8072
rect 30607 8041 30619 8044
rect 30561 8035 30619 8041
rect 35250 8032 35256 8044
rect 35308 8032 35314 8084
rect 17681 8007 17739 8013
rect 17681 7973 17693 8007
rect 17727 8004 17739 8007
rect 19242 8004 19248 8016
rect 17727 7976 19248 8004
rect 17727 7973 17739 7976
rect 17681 7967 17739 7973
rect 19242 7964 19248 7976
rect 19300 7964 19306 8016
rect 32309 8007 32367 8013
rect 32309 7973 32321 8007
rect 32355 8004 32367 8007
rect 38378 8004 38384 8016
rect 32355 7976 38384 8004
rect 32355 7973 32367 7976
rect 32309 7967 32367 7973
rect 38378 7964 38384 7976
rect 38436 7964 38442 8016
rect 16482 7896 16488 7948
rect 16540 7936 16546 7948
rect 18141 7939 18199 7945
rect 18141 7936 18153 7939
rect 16540 7908 18153 7936
rect 16540 7896 16546 7908
rect 18141 7905 18153 7908
rect 18187 7905 18199 7939
rect 18141 7899 18199 7905
rect 18233 7939 18291 7945
rect 18233 7905 18245 7939
rect 18279 7936 18291 7939
rect 18598 7936 18604 7948
rect 18279 7908 18604 7936
rect 18279 7905 18291 7908
rect 18233 7899 18291 7905
rect 18598 7896 18604 7908
rect 18656 7896 18662 7948
rect 19426 7896 19432 7948
rect 19484 7896 19490 7948
rect 22649 7939 22707 7945
rect 22649 7905 22661 7939
rect 22695 7936 22707 7939
rect 23750 7936 23756 7948
rect 22695 7908 23756 7936
rect 22695 7905 22707 7908
rect 22649 7899 22707 7905
rect 23750 7896 23756 7908
rect 23808 7896 23814 7948
rect 31205 7939 31263 7945
rect 31205 7905 31217 7939
rect 31251 7936 31263 7939
rect 32582 7936 32588 7948
rect 31251 7908 32588 7936
rect 31251 7905 31263 7908
rect 31205 7899 31263 7905
rect 32582 7896 32588 7908
rect 32640 7896 32646 7948
rect 32953 7939 33011 7945
rect 32953 7905 32965 7939
rect 32999 7936 33011 7939
rect 35802 7936 35808 7948
rect 32999 7908 35808 7936
rect 32999 7905 33011 7908
rect 32953 7899 33011 7905
rect 35802 7896 35808 7908
rect 35860 7896 35866 7948
rect 49145 7939 49203 7945
rect 49145 7905 49157 7939
rect 49191 7936 49203 7939
rect 49234 7936 49240 7948
rect 49191 7908 49240 7936
rect 49191 7905 49203 7908
rect 49145 7899 49203 7905
rect 49234 7896 49240 7908
rect 49292 7896 49298 7948
rect 934 7828 940 7880
rect 992 7868 998 7880
rect 1581 7871 1639 7877
rect 1581 7868 1593 7871
rect 992 7840 1593 7868
rect 992 7828 998 7840
rect 1581 7837 1593 7840
rect 1627 7837 1639 7871
rect 1581 7831 1639 7837
rect 12802 7828 12808 7880
rect 12860 7868 12866 7880
rect 15841 7871 15899 7877
rect 15841 7868 15853 7871
rect 12860 7840 15853 7868
rect 12860 7828 12866 7840
rect 15841 7837 15853 7840
rect 15887 7837 15899 7871
rect 15841 7831 15899 7837
rect 18049 7871 18107 7877
rect 18049 7837 18061 7871
rect 18095 7868 18107 7871
rect 18322 7868 18328 7880
rect 18095 7840 18328 7868
rect 18095 7837 18107 7840
rect 18049 7831 18107 7837
rect 18322 7828 18328 7840
rect 18380 7828 18386 7880
rect 22186 7828 22192 7880
rect 22244 7868 22250 7880
rect 22373 7871 22431 7877
rect 22373 7868 22385 7871
rect 22244 7840 22385 7868
rect 22244 7828 22250 7840
rect 22373 7837 22385 7840
rect 22419 7837 22431 7871
rect 22373 7831 22431 7837
rect 30558 7828 30564 7880
rect 30616 7868 30622 7880
rect 30929 7871 30987 7877
rect 30929 7868 30941 7871
rect 30616 7840 30941 7868
rect 30616 7828 30622 7840
rect 30929 7837 30941 7840
rect 30975 7837 30987 7871
rect 30929 7831 30987 7837
rect 31021 7871 31079 7877
rect 31021 7837 31033 7871
rect 31067 7868 31079 7871
rect 31754 7868 31760 7880
rect 31067 7840 31760 7868
rect 31067 7837 31079 7840
rect 31021 7831 31079 7837
rect 31754 7828 31760 7840
rect 31812 7828 31818 7880
rect 31846 7828 31852 7880
rect 31904 7868 31910 7880
rect 32766 7868 32772 7880
rect 31904 7840 32772 7868
rect 31904 7828 31910 7840
rect 32766 7828 32772 7840
rect 32824 7828 32830 7880
rect 38746 7828 38752 7880
rect 38804 7828 38810 7880
rect 43714 7828 43720 7880
rect 43772 7868 43778 7880
rect 47949 7871 48007 7877
rect 47949 7868 47961 7871
rect 43772 7840 47961 7868
rect 43772 7828 43778 7840
rect 47949 7837 47961 7840
rect 47995 7837 48007 7871
rect 47949 7831 48007 7837
rect 15470 7800 15476 7812
rect 6886 7772 15476 7800
rect 1765 7735 1823 7741
rect 1765 7701 1777 7735
rect 1811 7732 1823 7735
rect 6886 7732 6914 7772
rect 15470 7760 15476 7772
rect 15528 7760 15534 7812
rect 18966 7800 18972 7812
rect 15672 7772 18972 7800
rect 15672 7741 15700 7772
rect 18966 7760 18972 7772
rect 19024 7760 19030 7812
rect 19705 7803 19763 7809
rect 19705 7769 19717 7803
rect 19751 7800 19763 7803
rect 19978 7800 19984 7812
rect 19751 7772 19984 7800
rect 19751 7769 19763 7772
rect 19705 7763 19763 7769
rect 19978 7760 19984 7772
rect 20036 7760 20042 7812
rect 21082 7800 21088 7812
rect 20930 7772 21088 7800
rect 21082 7760 21088 7772
rect 21140 7800 21146 7812
rect 21818 7800 21824 7812
rect 21140 7772 21824 7800
rect 21140 7760 21146 7772
rect 21818 7760 21824 7772
rect 21876 7760 21882 7812
rect 27706 7760 27712 7812
rect 27764 7800 27770 7812
rect 38013 7803 38071 7809
rect 38013 7800 38025 7803
rect 27764 7772 38025 7800
rect 27764 7760 27770 7772
rect 38013 7769 38025 7772
rect 38059 7769 38071 7803
rect 38013 7763 38071 7769
rect 38933 7803 38991 7809
rect 38933 7769 38945 7803
rect 38979 7800 38991 7803
rect 40034 7800 40040 7812
rect 38979 7772 40040 7800
rect 38979 7769 38991 7772
rect 38933 7763 38991 7769
rect 40034 7760 40040 7772
rect 40092 7760 40098 7812
rect 1811 7704 6914 7732
rect 15657 7735 15715 7741
rect 1811 7701 1823 7704
rect 1765 7695 1823 7701
rect 15657 7701 15669 7735
rect 15703 7701 15715 7735
rect 15657 7695 15715 7701
rect 22465 7735 22523 7741
rect 22465 7701 22477 7735
rect 22511 7732 22523 7735
rect 22738 7732 22744 7744
rect 22511 7704 22744 7732
rect 22511 7701 22523 7704
rect 22465 7695 22523 7701
rect 22738 7692 22744 7704
rect 22796 7732 22802 7744
rect 26050 7732 26056 7744
rect 22796 7704 26056 7732
rect 22796 7692 22802 7704
rect 26050 7692 26056 7704
rect 26108 7692 26114 7744
rect 32674 7692 32680 7744
rect 32732 7692 32738 7744
rect 32766 7692 32772 7744
rect 32824 7692 32830 7744
rect 38105 7735 38163 7741
rect 38105 7701 38117 7735
rect 38151 7732 38163 7735
rect 38654 7732 38660 7744
rect 38151 7704 38660 7732
rect 38151 7701 38163 7704
rect 38105 7695 38163 7701
rect 38654 7692 38660 7704
rect 38712 7692 38718 7744
rect 1104 7642 49864 7664
rect 1104 7590 7950 7642
rect 8002 7590 8014 7642
rect 8066 7590 8078 7642
rect 8130 7590 8142 7642
rect 8194 7590 8206 7642
rect 8258 7590 17950 7642
rect 18002 7590 18014 7642
rect 18066 7590 18078 7642
rect 18130 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 27950 7642
rect 28002 7590 28014 7642
rect 28066 7590 28078 7642
rect 28130 7590 28142 7642
rect 28194 7590 28206 7642
rect 28258 7590 37950 7642
rect 38002 7590 38014 7642
rect 38066 7590 38078 7642
rect 38130 7590 38142 7642
rect 38194 7590 38206 7642
rect 38258 7590 47950 7642
rect 48002 7590 48014 7642
rect 48066 7590 48078 7642
rect 48130 7590 48142 7642
rect 48194 7590 48206 7642
rect 48258 7590 49864 7642
rect 1104 7568 49864 7590
rect 1765 7531 1823 7537
rect 1765 7497 1777 7531
rect 1811 7528 1823 7531
rect 1811 7500 6914 7528
rect 1811 7497 1823 7500
rect 1765 7491 1823 7497
rect 6886 7460 6914 7500
rect 21174 7488 21180 7540
rect 21232 7528 21238 7540
rect 22005 7531 22063 7537
rect 22005 7528 22017 7531
rect 21232 7500 22017 7528
rect 21232 7488 21238 7500
rect 22005 7497 22017 7500
rect 22051 7497 22063 7531
rect 22005 7491 22063 7497
rect 22370 7488 22376 7540
rect 22428 7528 22434 7540
rect 22465 7531 22523 7537
rect 22465 7528 22477 7531
rect 22428 7500 22477 7528
rect 22428 7488 22434 7500
rect 22465 7497 22477 7500
rect 22511 7497 22523 7531
rect 22465 7491 22523 7497
rect 23293 7531 23351 7537
rect 23293 7497 23305 7531
rect 23339 7528 23351 7531
rect 31478 7528 31484 7540
rect 23339 7500 31484 7528
rect 23339 7497 23351 7500
rect 23293 7491 23351 7497
rect 18782 7460 18788 7472
rect 6886 7432 18788 7460
rect 18782 7420 18788 7432
rect 18840 7420 18846 7472
rect 934 7352 940 7404
rect 992 7392 998 7404
rect 1581 7395 1639 7401
rect 1581 7392 1593 7395
rect 992 7364 1593 7392
rect 992 7352 998 7364
rect 1581 7361 1593 7364
rect 1627 7361 1639 7395
rect 1581 7355 1639 7361
rect 15562 7352 15568 7404
rect 15620 7392 15626 7404
rect 17865 7395 17923 7401
rect 17865 7392 17877 7395
rect 15620 7364 17877 7392
rect 15620 7352 15626 7364
rect 17865 7361 17877 7364
rect 17911 7361 17923 7395
rect 22373 7395 22431 7401
rect 22373 7392 22385 7395
rect 17865 7355 17923 7361
rect 22066 7364 22385 7392
rect 16942 7284 16948 7336
rect 17000 7324 17006 7336
rect 22066 7324 22094 7364
rect 22373 7361 22385 7364
rect 22419 7392 22431 7395
rect 23308 7392 23336 7491
rect 31478 7488 31484 7500
rect 31536 7488 31542 7540
rect 31846 7528 31852 7540
rect 31588 7500 31852 7528
rect 24946 7420 24952 7472
rect 25004 7460 25010 7472
rect 31588 7460 31616 7500
rect 31846 7488 31852 7500
rect 31904 7488 31910 7540
rect 38654 7488 38660 7540
rect 38712 7528 38718 7540
rect 47578 7528 47584 7540
rect 38712 7500 47584 7528
rect 38712 7488 38718 7500
rect 47578 7488 47584 7500
rect 47636 7488 47642 7540
rect 37829 7463 37887 7469
rect 37829 7460 37841 7463
rect 25004 7432 31616 7460
rect 31726 7432 37841 7460
rect 25004 7420 25010 7432
rect 22419 7364 23336 7392
rect 31113 7395 31171 7401
rect 22419 7361 22431 7364
rect 22373 7355 22431 7361
rect 31113 7361 31125 7395
rect 31159 7392 31171 7395
rect 31386 7392 31392 7404
rect 31159 7364 31392 7392
rect 31159 7361 31171 7364
rect 31113 7355 31171 7361
rect 31386 7352 31392 7364
rect 31444 7352 31450 7404
rect 31726 7392 31754 7432
rect 37829 7429 37841 7432
rect 37875 7429 37887 7463
rect 37829 7423 37887 7429
rect 40126 7420 40132 7472
rect 40184 7460 40190 7472
rect 44913 7463 44971 7469
rect 44913 7460 44925 7463
rect 40184 7432 44925 7460
rect 40184 7420 40190 7432
rect 44913 7429 44925 7432
rect 44959 7429 44971 7463
rect 44913 7423 44971 7429
rect 49145 7463 49203 7469
rect 49145 7429 49157 7463
rect 49191 7460 49203 7463
rect 49326 7460 49332 7472
rect 49191 7432 49332 7460
rect 49191 7429 49203 7432
rect 49145 7423 49203 7429
rect 49326 7420 49332 7432
rect 49384 7420 49390 7472
rect 31496 7364 31754 7392
rect 17000 7296 22094 7324
rect 17000 7284 17006 7296
rect 22646 7284 22652 7336
rect 22704 7284 22710 7336
rect 27798 7284 27804 7336
rect 27856 7324 27862 7336
rect 31496 7324 31524 7364
rect 34238 7352 34244 7404
rect 34296 7392 34302 7404
rect 38565 7395 38623 7401
rect 38565 7392 38577 7395
rect 34296 7364 38577 7392
rect 34296 7352 34302 7364
rect 38565 7361 38577 7364
rect 38611 7361 38623 7395
rect 38565 7355 38623 7361
rect 42794 7352 42800 7404
rect 42852 7392 42858 7404
rect 47949 7395 48007 7401
rect 47949 7392 47961 7395
rect 42852 7364 47961 7392
rect 42852 7352 42858 7364
rect 47949 7361 47961 7364
rect 47995 7361 48007 7395
rect 47949 7355 48007 7361
rect 27856 7296 31524 7324
rect 27856 7284 27862 7296
rect 31754 7284 31760 7336
rect 31812 7324 31818 7336
rect 35526 7324 35532 7336
rect 31812 7296 35532 7324
rect 31812 7284 31818 7296
rect 35526 7284 35532 7296
rect 35584 7284 35590 7336
rect 38749 7259 38807 7265
rect 38749 7225 38761 7259
rect 38795 7256 38807 7259
rect 45738 7256 45744 7268
rect 38795 7228 45744 7256
rect 38795 7225 38807 7228
rect 38749 7219 38807 7225
rect 45738 7216 45744 7228
rect 45796 7216 45802 7268
rect 17681 7191 17739 7197
rect 17681 7157 17693 7191
rect 17727 7188 17739 7191
rect 20438 7188 20444 7200
rect 17727 7160 20444 7188
rect 17727 7157 17739 7160
rect 17681 7151 17739 7157
rect 20438 7148 20444 7160
rect 20496 7148 20502 7200
rect 37918 7148 37924 7200
rect 37976 7148 37982 7200
rect 45005 7191 45063 7197
rect 45005 7157 45017 7191
rect 45051 7188 45063 7191
rect 47762 7188 47768 7200
rect 45051 7160 47768 7188
rect 45051 7157 45063 7160
rect 45005 7151 45063 7157
rect 47762 7148 47768 7160
rect 47820 7148 47826 7200
rect 1104 7098 49864 7120
rect 1104 7046 2950 7098
rect 3002 7046 3014 7098
rect 3066 7046 3078 7098
rect 3130 7046 3142 7098
rect 3194 7046 3206 7098
rect 3258 7046 12950 7098
rect 13002 7046 13014 7098
rect 13066 7046 13078 7098
rect 13130 7046 13142 7098
rect 13194 7046 13206 7098
rect 13258 7046 22950 7098
rect 23002 7046 23014 7098
rect 23066 7046 23078 7098
rect 23130 7046 23142 7098
rect 23194 7046 23206 7098
rect 23258 7046 32950 7098
rect 33002 7046 33014 7098
rect 33066 7046 33078 7098
rect 33130 7046 33142 7098
rect 33194 7046 33206 7098
rect 33258 7046 42950 7098
rect 43002 7046 43014 7098
rect 43066 7046 43078 7098
rect 43130 7046 43142 7098
rect 43194 7046 43206 7098
rect 43258 7046 49864 7098
rect 1104 7024 49864 7046
rect 37918 6876 37924 6928
rect 37976 6916 37982 6928
rect 46934 6916 46940 6928
rect 37976 6888 46940 6916
rect 37976 6876 37982 6888
rect 46934 6876 46940 6888
rect 46992 6876 46998 6928
rect 32766 6808 32772 6860
rect 32824 6848 32830 6860
rect 37734 6848 37740 6860
rect 32824 6820 37740 6848
rect 32824 6808 32830 6820
rect 37734 6808 37740 6820
rect 37792 6808 37798 6860
rect 49142 6808 49148 6860
rect 49200 6808 49206 6860
rect 934 6740 940 6792
rect 992 6780 998 6792
rect 1673 6783 1731 6789
rect 1673 6780 1685 6783
rect 992 6752 1685 6780
rect 992 6740 998 6752
rect 1673 6749 1685 6752
rect 1719 6749 1731 6783
rect 2501 6783 2559 6789
rect 2501 6780 2513 6783
rect 1673 6743 1731 6749
rect 1780 6752 2513 6780
rect 1302 6672 1308 6724
rect 1360 6712 1366 6724
rect 1780 6712 1808 6752
rect 2501 6749 2513 6752
rect 2547 6749 2559 6783
rect 2501 6743 2559 6749
rect 19242 6740 19248 6792
rect 19300 6780 19306 6792
rect 19889 6783 19947 6789
rect 19889 6780 19901 6783
rect 19300 6752 19901 6780
rect 19300 6740 19306 6752
rect 19889 6749 19901 6752
rect 19935 6749 19947 6783
rect 19889 6743 19947 6749
rect 40034 6740 40040 6792
rect 40092 6780 40098 6792
rect 46109 6783 46167 6789
rect 46109 6780 46121 6783
rect 40092 6752 46121 6780
rect 40092 6740 40098 6752
rect 46109 6749 46121 6752
rect 46155 6749 46167 6783
rect 46109 6743 46167 6749
rect 47854 6740 47860 6792
rect 47912 6780 47918 6792
rect 47949 6783 48007 6789
rect 47949 6780 47961 6783
rect 47912 6752 47961 6780
rect 47912 6740 47918 6752
rect 47949 6749 47961 6752
rect 47995 6749 48007 6783
rect 47949 6743 48007 6749
rect 1360 6684 1808 6712
rect 1857 6715 1915 6721
rect 1360 6672 1366 6684
rect 1857 6681 1869 6715
rect 1903 6712 1915 6715
rect 27614 6712 27620 6724
rect 1903 6684 27620 6712
rect 1903 6681 1915 6684
rect 1857 6675 1915 6681
rect 27614 6672 27620 6684
rect 27672 6672 27678 6724
rect 47305 6715 47363 6721
rect 47305 6681 47317 6715
rect 47351 6712 47363 6715
rect 48866 6712 48872 6724
rect 47351 6684 48872 6712
rect 47351 6681 47363 6684
rect 47305 6675 47363 6681
rect 48866 6672 48872 6684
rect 48924 6672 48930 6724
rect 2314 6604 2320 6656
rect 2372 6604 2378 6656
rect 19705 6647 19763 6653
rect 19705 6613 19717 6647
rect 19751 6644 19763 6647
rect 21910 6644 21916 6656
rect 19751 6616 21916 6644
rect 19751 6613 19763 6616
rect 19705 6607 19763 6613
rect 21910 6604 21916 6616
rect 21968 6604 21974 6656
rect 1104 6554 49864 6576
rect 1104 6502 7950 6554
rect 8002 6502 8014 6554
rect 8066 6502 8078 6554
rect 8130 6502 8142 6554
rect 8194 6502 8206 6554
rect 8258 6502 17950 6554
rect 18002 6502 18014 6554
rect 18066 6502 18078 6554
rect 18130 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 27950 6554
rect 28002 6502 28014 6554
rect 28066 6502 28078 6554
rect 28130 6502 28142 6554
rect 28194 6502 28206 6554
rect 28258 6502 37950 6554
rect 38002 6502 38014 6554
rect 38066 6502 38078 6554
rect 38130 6502 38142 6554
rect 38194 6502 38206 6554
rect 38258 6502 47950 6554
rect 48002 6502 48014 6554
rect 48066 6502 48078 6554
rect 48130 6502 48142 6554
rect 48194 6502 48206 6554
rect 48258 6502 49864 6554
rect 1104 6480 49864 6502
rect 30466 6332 30472 6384
rect 30524 6372 30530 6384
rect 37553 6375 37611 6381
rect 37553 6372 37565 6375
rect 30524 6344 37565 6372
rect 30524 6332 30530 6344
rect 37553 6341 37565 6344
rect 37599 6341 37611 6375
rect 37553 6335 37611 6341
rect 40218 6332 40224 6384
rect 40276 6372 40282 6384
rect 43993 6375 44051 6381
rect 43993 6372 44005 6375
rect 40276 6344 44005 6372
rect 40276 6332 40282 6344
rect 43993 6341 44005 6344
rect 44039 6341 44051 6375
rect 43993 6335 44051 6341
rect 49145 6375 49203 6381
rect 49145 6341 49157 6375
rect 49191 6372 49203 6375
rect 49234 6372 49240 6384
rect 49191 6344 49240 6372
rect 49191 6341 49203 6344
rect 49145 6335 49203 6341
rect 49234 6332 49240 6344
rect 49292 6332 49298 6384
rect 934 6264 940 6316
rect 992 6304 998 6316
rect 1581 6307 1639 6313
rect 1581 6304 1593 6307
rect 992 6276 1593 6304
rect 992 6264 998 6276
rect 1581 6273 1593 6276
rect 1627 6273 1639 6307
rect 1581 6267 1639 6273
rect 16390 6264 16396 6316
rect 16448 6304 16454 6316
rect 18049 6307 18107 6313
rect 18049 6304 18061 6307
rect 16448 6276 18061 6304
rect 16448 6264 16454 6276
rect 18049 6273 18061 6276
rect 18095 6273 18107 6307
rect 18049 6267 18107 6273
rect 46566 6264 46572 6316
rect 46624 6304 46630 6316
rect 47949 6307 48007 6313
rect 47949 6304 47961 6307
rect 46624 6276 47961 6304
rect 46624 6264 46630 6276
rect 47949 6273 47961 6276
rect 47995 6273 48007 6307
rect 47949 6267 48007 6273
rect 18233 6239 18291 6245
rect 18233 6205 18245 6239
rect 18279 6236 18291 6239
rect 18322 6236 18328 6248
rect 18279 6208 18328 6236
rect 18279 6205 18291 6208
rect 18233 6199 18291 6205
rect 18322 6196 18328 6208
rect 18380 6196 18386 6248
rect 1854 6128 1860 6180
rect 1912 6168 1918 6180
rect 24946 6168 24952 6180
rect 1912 6140 24952 6168
rect 1912 6128 1918 6140
rect 24946 6128 24952 6140
rect 25004 6128 25010 6180
rect 32122 6128 32128 6180
rect 32180 6168 32186 6180
rect 44177 6171 44235 6177
rect 32180 6140 41414 6168
rect 32180 6128 32186 6140
rect 1765 6103 1823 6109
rect 1765 6069 1777 6103
rect 1811 6100 1823 6103
rect 16298 6100 16304 6112
rect 1811 6072 16304 6100
rect 1811 6069 1823 6072
rect 1765 6063 1823 6069
rect 16298 6060 16304 6072
rect 16356 6060 16362 6112
rect 18693 6103 18751 6109
rect 18693 6069 18705 6103
rect 18739 6100 18751 6103
rect 19610 6100 19616 6112
rect 18739 6072 19616 6100
rect 18739 6069 18751 6072
rect 18693 6063 18751 6069
rect 19610 6060 19616 6072
rect 19668 6060 19674 6112
rect 37642 6060 37648 6112
rect 37700 6060 37706 6112
rect 41386 6100 41414 6140
rect 44177 6137 44189 6171
rect 44223 6168 44235 6171
rect 47026 6168 47032 6180
rect 44223 6140 47032 6168
rect 44223 6137 44235 6140
rect 44177 6131 44235 6137
rect 47026 6128 47032 6140
rect 47084 6128 47090 6180
rect 45554 6100 45560 6112
rect 41386 6072 45560 6100
rect 45554 6060 45560 6072
rect 45612 6060 45618 6112
rect 1104 6010 49864 6032
rect 1104 5958 2950 6010
rect 3002 5958 3014 6010
rect 3066 5958 3078 6010
rect 3130 5958 3142 6010
rect 3194 5958 3206 6010
rect 3258 5958 12950 6010
rect 13002 5958 13014 6010
rect 13066 5958 13078 6010
rect 13130 5958 13142 6010
rect 13194 5958 13206 6010
rect 13258 5958 22950 6010
rect 23002 5958 23014 6010
rect 23066 5958 23078 6010
rect 23130 5958 23142 6010
rect 23194 5958 23206 6010
rect 23258 5958 32950 6010
rect 33002 5958 33014 6010
rect 33066 5958 33078 6010
rect 33130 5958 33142 6010
rect 33194 5958 33206 6010
rect 33258 5958 42950 6010
rect 43002 5958 43014 6010
rect 43066 5958 43078 6010
rect 43130 5958 43142 6010
rect 43194 5958 43206 6010
rect 43258 5958 49864 6010
rect 1104 5936 49864 5958
rect 37642 5856 37648 5908
rect 37700 5896 37706 5908
rect 47210 5896 47216 5908
rect 37700 5868 47216 5896
rect 37700 5856 37706 5868
rect 47210 5856 47216 5868
rect 47268 5856 47274 5908
rect 2501 5831 2559 5837
rect 2501 5797 2513 5831
rect 2547 5828 2559 5831
rect 17218 5828 17224 5840
rect 2547 5800 17224 5828
rect 2547 5797 2559 5800
rect 2501 5791 2559 5797
rect 17218 5788 17224 5800
rect 17276 5788 17282 5840
rect 49145 5763 49203 5769
rect 49145 5729 49157 5763
rect 49191 5760 49203 5763
rect 49418 5760 49424 5772
rect 49191 5732 49424 5760
rect 49191 5729 49203 5732
rect 49145 5723 49203 5729
rect 49418 5720 49424 5732
rect 49476 5720 49482 5772
rect 934 5652 940 5704
rect 992 5692 998 5704
rect 1581 5695 1639 5701
rect 1581 5692 1593 5695
rect 992 5664 1593 5692
rect 992 5652 998 5664
rect 1581 5661 1593 5664
rect 1627 5661 1639 5695
rect 1581 5655 1639 5661
rect 2314 5652 2320 5704
rect 2372 5652 2378 5704
rect 43714 5652 43720 5704
rect 43772 5652 43778 5704
rect 47670 5652 47676 5704
rect 47728 5692 47734 5704
rect 47949 5695 48007 5701
rect 47949 5692 47961 5695
rect 47728 5664 47961 5692
rect 47728 5652 47734 5664
rect 47949 5661 47961 5664
rect 47995 5661 48007 5695
rect 47949 5655 48007 5661
rect 43901 5627 43959 5633
rect 1780 5596 6914 5624
rect 1780 5565 1808 5596
rect 1765 5559 1823 5565
rect 1765 5525 1777 5559
rect 1811 5525 1823 5559
rect 6886 5556 6914 5596
rect 43901 5593 43913 5627
rect 43947 5624 43959 5627
rect 45830 5624 45836 5636
rect 43947 5596 45836 5624
rect 43947 5593 43959 5596
rect 43901 5587 43959 5593
rect 45830 5584 45836 5596
rect 45888 5584 45894 5636
rect 18690 5556 18696 5568
rect 6886 5528 18696 5556
rect 1765 5519 1823 5525
rect 18690 5516 18696 5528
rect 18748 5516 18754 5568
rect 1104 5466 49864 5488
rect 1104 5414 7950 5466
rect 8002 5414 8014 5466
rect 8066 5414 8078 5466
rect 8130 5414 8142 5466
rect 8194 5414 8206 5466
rect 8258 5414 17950 5466
rect 18002 5414 18014 5466
rect 18066 5414 18078 5466
rect 18130 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 27950 5466
rect 28002 5414 28014 5466
rect 28066 5414 28078 5466
rect 28130 5414 28142 5466
rect 28194 5414 28206 5466
rect 28258 5414 37950 5466
rect 38002 5414 38014 5466
rect 38066 5414 38078 5466
rect 38130 5414 38142 5466
rect 38194 5414 38206 5466
rect 38258 5414 47950 5466
rect 48002 5414 48014 5466
rect 48066 5414 48078 5466
rect 48130 5414 48142 5466
rect 48194 5414 48206 5466
rect 48258 5414 49864 5466
rect 1104 5392 49864 5414
rect 37734 5244 37740 5296
rect 37792 5244 37798 5296
rect 38470 5244 38476 5296
rect 38528 5244 38534 5296
rect 49142 5244 49148 5296
rect 49200 5244 49206 5296
rect 18966 5176 18972 5228
rect 19024 5176 19030 5228
rect 22716 5219 22774 5225
rect 22716 5216 22728 5219
rect 22066 5188 22728 5216
rect 934 5108 940 5160
rect 992 5148 998 5160
rect 1581 5151 1639 5157
rect 1581 5148 1593 5151
rect 992 5120 1593 5148
rect 992 5108 998 5120
rect 1581 5117 1593 5120
rect 1627 5117 1639 5151
rect 1581 5111 1639 5117
rect 1857 5151 1915 5157
rect 1857 5117 1869 5151
rect 1903 5148 1915 5151
rect 15746 5148 15752 5160
rect 1903 5120 15752 5148
rect 1903 5117 1915 5120
rect 1857 5111 1915 5117
rect 15746 5108 15752 5120
rect 15804 5108 15810 5160
rect 19150 5108 19156 5160
rect 19208 5148 19214 5160
rect 22066 5148 22094 5188
rect 22716 5185 22728 5188
rect 22762 5216 22774 5219
rect 24026 5216 24032 5228
rect 22762 5188 24032 5216
rect 22762 5185 22774 5188
rect 22716 5179 22774 5185
rect 24026 5176 24032 5188
rect 24084 5176 24090 5228
rect 45738 5176 45744 5228
rect 45796 5216 45802 5228
rect 45833 5219 45891 5225
rect 45833 5216 45845 5219
rect 45796 5188 45845 5216
rect 45796 5176 45802 5188
rect 45833 5185 45845 5188
rect 45879 5185 45891 5219
rect 45833 5179 45891 5185
rect 47762 5176 47768 5228
rect 47820 5216 47826 5228
rect 47949 5219 48007 5225
rect 47949 5216 47961 5219
rect 47820 5188 47961 5216
rect 47820 5176 47826 5188
rect 47949 5185 47961 5188
rect 47995 5185 48007 5219
rect 47949 5179 48007 5185
rect 19208 5120 22094 5148
rect 46845 5151 46903 5157
rect 19208 5108 19214 5120
rect 46845 5117 46857 5151
rect 46891 5148 46903 5151
rect 48314 5148 48320 5160
rect 46891 5120 48320 5148
rect 46891 5117 46903 5120
rect 46845 5111 46903 5117
rect 48314 5108 48320 5120
rect 48372 5108 48378 5160
rect 38657 5083 38715 5089
rect 38657 5049 38669 5083
rect 38703 5080 38715 5083
rect 40034 5080 40040 5092
rect 38703 5052 40040 5080
rect 38703 5049 38715 5052
rect 38657 5043 38715 5049
rect 40034 5040 40040 5052
rect 40092 5040 40098 5092
rect 19613 5015 19671 5021
rect 19613 4981 19625 5015
rect 19659 5012 19671 5015
rect 20806 5012 20812 5024
rect 19659 4984 20812 5012
rect 19659 4981 19671 4984
rect 19613 4975 19671 4981
rect 20806 4972 20812 4984
rect 20864 4972 20870 5024
rect 22787 5015 22845 5021
rect 22787 4981 22799 5015
rect 22833 5012 22845 5015
rect 24302 5012 24308 5024
rect 22833 4984 24308 5012
rect 22833 4981 22845 4984
rect 22787 4975 22845 4981
rect 24302 4972 24308 4984
rect 24360 4972 24366 5024
rect 26786 4972 26792 5024
rect 26844 5012 26850 5024
rect 37274 5012 37280 5024
rect 26844 4984 37280 5012
rect 26844 4972 26850 4984
rect 37274 4972 37280 4984
rect 37332 4972 37338 5024
rect 37826 4972 37832 5024
rect 37884 4972 37890 5024
rect 1104 4922 49864 4944
rect 1104 4870 2950 4922
rect 3002 4870 3014 4922
rect 3066 4870 3078 4922
rect 3130 4870 3142 4922
rect 3194 4870 3206 4922
rect 3258 4870 12950 4922
rect 13002 4870 13014 4922
rect 13066 4870 13078 4922
rect 13130 4870 13142 4922
rect 13194 4870 13206 4922
rect 13258 4870 22950 4922
rect 23002 4870 23014 4922
rect 23066 4870 23078 4922
rect 23130 4870 23142 4922
rect 23194 4870 23206 4922
rect 23258 4870 32950 4922
rect 33002 4870 33014 4922
rect 33066 4870 33078 4922
rect 33130 4870 33142 4922
rect 33194 4870 33206 4922
rect 33258 4870 42950 4922
rect 43002 4870 43014 4922
rect 43066 4870 43078 4922
rect 43130 4870 43142 4922
rect 43194 4870 43206 4922
rect 43258 4870 49864 4922
rect 1104 4848 49864 4870
rect 37826 4768 37832 4820
rect 37884 4808 37890 4820
rect 47118 4808 47124 4820
rect 37884 4780 47124 4808
rect 37884 4768 37890 4780
rect 47118 4768 47124 4780
rect 47176 4768 47182 4820
rect 24670 4740 24676 4752
rect 6886 4712 24676 4740
rect 1857 4675 1915 4681
rect 1857 4641 1869 4675
rect 1903 4672 1915 4675
rect 6886 4672 6914 4712
rect 24670 4700 24676 4712
rect 24728 4700 24734 4752
rect 28718 4740 28724 4752
rect 25148 4712 28724 4740
rect 1903 4644 6914 4672
rect 1903 4641 1915 4644
rect 1857 4635 1915 4641
rect 20438 4632 20444 4684
rect 20496 4632 20502 4684
rect 21910 4632 21916 4684
rect 21968 4632 21974 4684
rect 25148 4681 25176 4712
rect 28718 4700 28724 4712
rect 28776 4700 28782 4752
rect 33778 4700 33784 4752
rect 33836 4740 33842 4752
rect 46753 4743 46811 4749
rect 46753 4740 46765 4743
rect 33836 4712 46765 4740
rect 33836 4700 33842 4712
rect 46753 4709 46765 4712
rect 46799 4709 46811 4743
rect 46753 4703 46811 4709
rect 25133 4675 25191 4681
rect 25133 4641 25145 4675
rect 25179 4641 25191 4675
rect 25133 4635 25191 4641
rect 25590 4632 25596 4684
rect 25648 4632 25654 4684
rect 36538 4632 36544 4684
rect 36596 4672 36602 4684
rect 47489 4675 47547 4681
rect 47489 4672 47501 4675
rect 36596 4644 47501 4672
rect 36596 4632 36602 4644
rect 47489 4641 47501 4644
rect 47535 4641 47547 4675
rect 47489 4635 47547 4641
rect 49145 4675 49203 4681
rect 49145 4641 49157 4675
rect 49191 4672 49203 4675
rect 49418 4672 49424 4684
rect 49191 4644 49424 4672
rect 49191 4641 49203 4644
rect 49145 4635 49203 4641
rect 49418 4632 49424 4644
rect 49476 4632 49482 4684
rect 19518 4564 19524 4616
rect 19576 4604 19582 4616
rect 20625 4607 20683 4613
rect 20625 4604 20637 4607
rect 19576 4576 20637 4604
rect 19576 4564 19582 4576
rect 20625 4573 20637 4576
rect 20671 4573 20683 4607
rect 20625 4567 20683 4573
rect 934 4496 940 4548
rect 992 4536 998 4548
rect 1673 4539 1731 4545
rect 1673 4536 1685 4539
rect 992 4508 1685 4536
rect 992 4496 998 4508
rect 1673 4505 1685 4508
rect 1719 4505 1731 4539
rect 20640 4536 20668 4567
rect 22094 4564 22100 4616
rect 22152 4564 22158 4616
rect 23436 4607 23494 4613
rect 23436 4604 23448 4607
rect 23032 4576 23448 4604
rect 23032 4536 23060 4576
rect 23436 4573 23448 4576
rect 23482 4604 23494 4607
rect 23658 4604 23664 4616
rect 23482 4576 23664 4604
rect 23482 4573 23494 4576
rect 23436 4567 23494 4573
rect 23658 4564 23664 4576
rect 23716 4564 23722 4616
rect 27522 4564 27528 4616
rect 27580 4604 27586 4616
rect 38013 4607 38071 4613
rect 38013 4604 38025 4607
rect 27580 4576 38025 4604
rect 27580 4564 27586 4576
rect 38013 4573 38025 4576
rect 38059 4573 38071 4607
rect 38013 4567 38071 4573
rect 47578 4564 47584 4616
rect 47636 4604 47642 4616
rect 47949 4607 48007 4613
rect 47949 4604 47961 4607
rect 47636 4576 47961 4604
rect 47636 4564 47642 4576
rect 47949 4573 47961 4576
rect 47995 4573 48007 4607
rect 47949 4567 48007 4573
rect 20640 4508 23060 4536
rect 23523 4539 23581 4545
rect 1673 4499 1731 4505
rect 23523 4505 23535 4539
rect 23569 4536 23581 4539
rect 25317 4539 25375 4545
rect 25317 4536 25329 4539
rect 23569 4508 25329 4536
rect 23569 4505 23581 4508
rect 23523 4499 23581 4505
rect 25317 4505 25329 4508
rect 25363 4505 25375 4539
rect 25317 4499 25375 4505
rect 37274 4496 37280 4548
rect 37332 4496 37338 4548
rect 37461 4539 37519 4545
rect 37461 4505 37473 4539
rect 37507 4536 37519 4539
rect 39850 4536 39856 4548
rect 37507 4508 39856 4536
rect 37507 4505 37519 4508
rect 37461 4499 37519 4505
rect 39850 4496 39856 4508
rect 39908 4496 39914 4548
rect 46569 4539 46627 4545
rect 46569 4505 46581 4539
rect 46615 4505 46627 4539
rect 46569 4499 46627 4505
rect 47305 4539 47363 4545
rect 47305 4505 47317 4539
rect 47351 4536 47363 4539
rect 47670 4536 47676 4548
rect 47351 4508 47676 4536
rect 47351 4505 47363 4508
rect 47305 4499 47363 4505
rect 21085 4471 21143 4477
rect 21085 4437 21097 4471
rect 21131 4468 21143 4471
rect 21450 4468 21456 4480
rect 21131 4440 21456 4468
rect 21131 4437 21143 4440
rect 21085 4431 21143 4437
rect 21450 4428 21456 4440
rect 21508 4428 21514 4480
rect 22557 4471 22615 4477
rect 22557 4437 22569 4471
rect 22603 4468 22615 4471
rect 26142 4468 26148 4480
rect 22603 4440 26148 4468
rect 22603 4437 22615 4440
rect 22557 4431 22615 4437
rect 26142 4428 26148 4440
rect 26200 4428 26206 4480
rect 38105 4471 38163 4477
rect 38105 4437 38117 4471
rect 38151 4468 38163 4471
rect 44634 4468 44640 4480
rect 38151 4440 44640 4468
rect 38151 4437 38163 4440
rect 38105 4431 38163 4437
rect 44634 4428 44640 4440
rect 44692 4428 44698 4480
rect 46584 4468 46612 4499
rect 47670 4496 47676 4508
rect 47728 4496 47734 4548
rect 49786 4468 49792 4480
rect 46584 4440 49792 4468
rect 49786 4428 49792 4440
rect 49844 4428 49850 4480
rect 1104 4378 49864 4400
rect 1104 4326 7950 4378
rect 8002 4326 8014 4378
rect 8066 4326 8078 4378
rect 8130 4326 8142 4378
rect 8194 4326 8206 4378
rect 8258 4326 17950 4378
rect 18002 4326 18014 4378
rect 18066 4326 18078 4378
rect 18130 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 27950 4378
rect 28002 4326 28014 4378
rect 28066 4326 28078 4378
rect 28130 4326 28142 4378
rect 28194 4326 28206 4378
rect 28258 4326 37950 4378
rect 38002 4326 38014 4378
rect 38066 4326 38078 4378
rect 38130 4326 38142 4378
rect 38194 4326 38206 4378
rect 38258 4326 47950 4378
rect 48002 4326 48014 4378
rect 48066 4326 48078 4378
rect 48130 4326 48142 4378
rect 48194 4326 48206 4378
rect 48258 4326 49864 4378
rect 1104 4304 49864 4326
rect 20714 4224 20720 4276
rect 20772 4264 20778 4276
rect 21634 4264 21640 4276
rect 20772 4236 21640 4264
rect 20772 4224 20778 4236
rect 21634 4224 21640 4236
rect 21692 4264 21698 4276
rect 25590 4264 25596 4276
rect 21692 4236 25596 4264
rect 21692 4224 21698 4236
rect 25590 4224 25596 4236
rect 25648 4224 25654 4276
rect 1670 4156 1676 4208
rect 1728 4156 1734 4208
rect 27341 4199 27399 4205
rect 27341 4196 27353 4199
rect 26896 4168 27353 4196
rect 934 4088 940 4140
rect 992 4128 998 4140
rect 2317 4131 2375 4137
rect 2317 4128 2329 4131
rect 992 4100 2329 4128
rect 992 4088 998 4100
rect 2317 4097 2329 4100
rect 2363 4097 2375 4131
rect 2317 4091 2375 4097
rect 18322 4088 18328 4140
rect 18380 4128 18386 4140
rect 22646 4137 22652 4140
rect 22624 4131 22652 4137
rect 22624 4128 22636 4131
rect 18380 4100 22636 4128
rect 18380 4088 18386 4100
rect 22624 4097 22636 4100
rect 22624 4091 22652 4097
rect 22646 4088 22652 4091
rect 22704 4088 22710 4140
rect 23512 4131 23570 4137
rect 23512 4128 23524 4131
rect 22756 4100 23524 4128
rect 1854 4020 1860 4072
rect 1912 4020 1918 4072
rect 22094 4020 22100 4072
rect 22152 4060 22158 4072
rect 22756 4060 22784 4100
rect 23512 4097 23524 4100
rect 23558 4097 23570 4131
rect 26896 4128 26924 4168
rect 27341 4165 27353 4168
rect 27387 4165 27399 4199
rect 27341 4159 27399 4165
rect 27157 4131 27215 4137
rect 27157 4128 27169 4131
rect 23512 4091 23570 4097
rect 25516 4100 26924 4128
rect 26988 4100 27169 4128
rect 22152 4032 22784 4060
rect 22152 4020 22158 4032
rect 24118 4020 24124 4072
rect 24176 4020 24182 4072
rect 24302 4020 24308 4072
rect 24360 4020 24366 4072
rect 24394 4020 24400 4072
rect 24452 4060 24458 4072
rect 24581 4063 24639 4069
rect 24581 4060 24593 4063
rect 24452 4032 24593 4060
rect 24452 4020 24458 4032
rect 24581 4029 24593 4032
rect 24627 4029 24639 4063
rect 24581 4023 24639 4029
rect 23615 3995 23673 4001
rect 23615 3961 23627 3995
rect 23661 3992 23673 3995
rect 25516 3992 25544 4100
rect 23661 3964 25544 3992
rect 23661 3961 23673 3964
rect 23615 3955 23673 3961
rect 2501 3927 2559 3933
rect 2501 3893 2513 3927
rect 2547 3924 2559 3927
rect 16942 3924 16948 3936
rect 2547 3896 16948 3924
rect 2547 3893 2559 3896
rect 2501 3887 2559 3893
rect 16942 3884 16948 3896
rect 17000 3884 17006 3936
rect 22695 3927 22753 3933
rect 22695 3893 22707 3927
rect 22741 3924 22753 3927
rect 24762 3924 24768 3936
rect 22741 3896 24768 3924
rect 22741 3893 22753 3896
rect 22695 3887 22753 3893
rect 24762 3884 24768 3896
rect 24820 3884 24826 3936
rect 26988 3924 27016 4100
rect 27157 4097 27169 4100
rect 27203 4097 27215 4131
rect 27157 4091 27215 4097
rect 36538 4088 36544 4140
rect 36596 4128 36602 4140
rect 45833 4131 45891 4137
rect 45833 4128 45845 4131
rect 36596 4100 45845 4128
rect 36596 4088 36602 4100
rect 45833 4097 45845 4100
rect 45879 4097 45891 4131
rect 45833 4091 45891 4097
rect 46934 4088 46940 4140
rect 46992 4128 46998 4140
rect 47949 4131 48007 4137
rect 47949 4128 47961 4131
rect 46992 4100 47961 4128
rect 46992 4088 46998 4100
rect 47949 4097 47961 4100
rect 47995 4097 48007 4131
rect 47949 4091 48007 4097
rect 49145 4131 49203 4137
rect 49145 4097 49157 4131
rect 49191 4128 49203 4131
rect 49326 4128 49332 4140
rect 49191 4100 49332 4128
rect 49191 4097 49203 4100
rect 49145 4091 49203 4097
rect 49326 4088 49332 4100
rect 49384 4088 49390 4140
rect 27614 4020 27620 4072
rect 27672 4020 27678 4072
rect 46658 4020 46664 4072
rect 46716 4020 46722 4072
rect 34422 3924 34428 3936
rect 26988 3896 34428 3924
rect 34422 3884 34428 3896
rect 34480 3884 34486 3936
rect 1104 3834 49864 3856
rect 1104 3782 2950 3834
rect 3002 3782 3014 3834
rect 3066 3782 3078 3834
rect 3130 3782 3142 3834
rect 3194 3782 3206 3834
rect 3258 3782 12950 3834
rect 13002 3782 13014 3834
rect 13066 3782 13078 3834
rect 13130 3782 13142 3834
rect 13194 3782 13206 3834
rect 13258 3782 22950 3834
rect 23002 3782 23014 3834
rect 23066 3782 23078 3834
rect 23130 3782 23142 3834
rect 23194 3782 23206 3834
rect 23258 3782 32950 3834
rect 33002 3782 33014 3834
rect 33066 3782 33078 3834
rect 33130 3782 33142 3834
rect 33194 3782 33206 3834
rect 33258 3782 42950 3834
rect 43002 3782 43014 3834
rect 43066 3782 43078 3834
rect 43130 3782 43142 3834
rect 43194 3782 43206 3834
rect 43258 3782 49864 3834
rect 1104 3760 49864 3782
rect 23845 3723 23903 3729
rect 23845 3689 23857 3723
rect 23891 3720 23903 3723
rect 25866 3720 25872 3732
rect 23891 3692 25872 3720
rect 23891 3689 23903 3692
rect 23845 3683 23903 3689
rect 25866 3680 25872 3692
rect 25924 3680 25930 3732
rect 36538 3680 36544 3732
rect 36596 3680 36602 3732
rect 45554 3680 45560 3732
rect 45612 3680 45618 3732
rect 23382 3652 23388 3664
rect 22480 3624 23388 3652
rect 3326 3544 3332 3596
rect 3384 3584 3390 3596
rect 20714 3584 20720 3596
rect 3384 3556 20720 3584
rect 3384 3544 3390 3556
rect 20714 3544 20720 3556
rect 20772 3544 20778 3596
rect 21910 3584 21916 3596
rect 20824 3556 21916 3584
rect 934 3476 940 3528
rect 992 3516 998 3528
rect 1581 3519 1639 3525
rect 1581 3516 1593 3519
rect 992 3488 1593 3516
rect 992 3476 998 3488
rect 1581 3485 1593 3488
rect 1627 3485 1639 3519
rect 1581 3479 1639 3485
rect 1857 3519 1915 3525
rect 1857 3485 1869 3519
rect 1903 3516 1915 3519
rect 14734 3516 14740 3528
rect 1903 3488 14740 3516
rect 1903 3485 1915 3488
rect 1857 3479 1915 3485
rect 14734 3476 14740 3488
rect 14792 3476 14798 3528
rect 16485 3519 16543 3525
rect 16485 3485 16497 3519
rect 16531 3516 16543 3519
rect 18322 3516 18328 3528
rect 16531 3488 18328 3516
rect 16531 3485 16543 3488
rect 16485 3479 16543 3485
rect 18322 3476 18328 3488
rect 18380 3476 18386 3528
rect 18414 3476 18420 3528
rect 18472 3516 18478 3528
rect 20824 3516 20852 3556
rect 21910 3544 21916 3556
rect 21968 3584 21974 3596
rect 22480 3584 22508 3624
rect 23382 3612 23388 3624
rect 23440 3652 23446 3664
rect 24302 3652 24308 3664
rect 23440 3624 24308 3652
rect 23440 3612 23446 3624
rect 24302 3612 24308 3624
rect 24360 3612 24366 3664
rect 28902 3652 28908 3664
rect 24596 3624 28908 3652
rect 21968 3556 22508 3584
rect 22572 3556 23980 3584
rect 21968 3544 21974 3556
rect 18472 3488 20852 3516
rect 18472 3476 18478 3488
rect 20898 3476 20904 3528
rect 20956 3476 20962 3528
rect 17862 3408 17868 3460
rect 17920 3448 17926 3460
rect 21174 3448 21180 3460
rect 17920 3420 21180 3448
rect 17920 3408 17926 3420
rect 21174 3408 21180 3420
rect 21232 3408 21238 3460
rect 21910 3408 21916 3460
rect 21968 3408 21974 3460
rect 12526 3340 12532 3392
rect 12584 3380 12590 3392
rect 16577 3383 16635 3389
rect 16577 3380 16589 3383
rect 12584 3352 16589 3380
rect 12584 3340 12590 3352
rect 16577 3349 16589 3352
rect 16623 3349 16635 3383
rect 16577 3343 16635 3349
rect 17218 3340 17224 3392
rect 17276 3380 17282 3392
rect 22572 3380 22600 3556
rect 22646 3476 22652 3528
rect 22704 3476 22710 3528
rect 23566 3476 23572 3528
rect 23624 3476 23630 3528
rect 23952 3516 23980 3556
rect 24026 3544 24032 3596
rect 24084 3544 24090 3596
rect 24596 3593 24624 3624
rect 28902 3612 28908 3624
rect 28960 3612 28966 3664
rect 24581 3587 24639 3593
rect 24581 3553 24593 3587
rect 24627 3553 24639 3587
rect 24581 3547 24639 3553
rect 24762 3544 24768 3596
rect 24820 3544 24826 3596
rect 24854 3544 24860 3596
rect 24912 3584 24918 3596
rect 25041 3587 25099 3593
rect 25041 3584 25053 3587
rect 24912 3556 25053 3584
rect 24912 3544 24918 3556
rect 25041 3553 25053 3556
rect 25087 3584 25099 3587
rect 25682 3584 25688 3596
rect 25087 3556 25688 3584
rect 25087 3553 25099 3556
rect 25041 3547 25099 3553
rect 25682 3544 25688 3556
rect 25740 3544 25746 3596
rect 31726 3556 36492 3584
rect 24486 3516 24492 3528
rect 23952 3488 24492 3516
rect 24486 3476 24492 3488
rect 24544 3476 24550 3528
rect 27798 3516 27804 3528
rect 25976 3488 27804 3516
rect 22664 3448 22692 3476
rect 25976 3448 26004 3488
rect 27798 3476 27804 3488
rect 27856 3476 27862 3528
rect 31726 3448 31754 3556
rect 36464 3457 36492 3556
rect 40034 3544 40040 3596
rect 40092 3584 40098 3596
rect 40092 3556 46152 3584
rect 40092 3544 40098 3556
rect 45465 3519 45523 3525
rect 45465 3485 45477 3519
rect 45511 3516 45523 3519
rect 45554 3516 45560 3528
rect 45511 3488 45560 3516
rect 45511 3485 45523 3488
rect 45465 3479 45523 3485
rect 45554 3476 45560 3488
rect 45612 3476 45618 3528
rect 46124 3525 46152 3556
rect 49142 3544 49148 3596
rect 49200 3544 49206 3596
rect 46109 3519 46167 3525
rect 46109 3485 46121 3519
rect 46155 3485 46167 3519
rect 46109 3479 46167 3485
rect 47026 3476 47032 3528
rect 47084 3516 47090 3528
rect 47949 3519 48007 3525
rect 47949 3516 47961 3519
rect 47084 3488 47961 3516
rect 47084 3476 47090 3488
rect 47949 3485 47961 3488
rect 47995 3485 48007 3519
rect 47949 3479 48007 3485
rect 22664 3420 26004 3448
rect 26528 3420 31754 3448
rect 36449 3451 36507 3457
rect 17276 3352 22600 3380
rect 22649 3383 22707 3389
rect 17276 3340 17282 3352
rect 22649 3349 22661 3383
rect 22695 3380 22707 3383
rect 23290 3380 23296 3392
rect 22695 3352 23296 3380
rect 22695 3349 22707 3352
rect 22649 3343 22707 3349
rect 23290 3340 23296 3352
rect 23348 3340 23354 3392
rect 23382 3340 23388 3392
rect 23440 3380 23446 3392
rect 26528 3380 26556 3420
rect 36449 3417 36461 3451
rect 36495 3417 36507 3451
rect 36449 3411 36507 3417
rect 47305 3451 47363 3457
rect 47305 3417 47317 3451
rect 47351 3448 47363 3451
rect 48682 3448 48688 3460
rect 47351 3420 48688 3448
rect 47351 3417 47363 3420
rect 47305 3411 47363 3417
rect 48682 3408 48688 3420
rect 48740 3408 48746 3460
rect 23440 3352 26556 3380
rect 23440 3340 23446 3352
rect 27154 3340 27160 3392
rect 27212 3380 27218 3392
rect 39206 3380 39212 3392
rect 27212 3352 39212 3380
rect 27212 3340 27218 3352
rect 39206 3340 39212 3352
rect 39264 3340 39270 3392
rect 1104 3290 49864 3312
rect 1104 3238 7950 3290
rect 8002 3238 8014 3290
rect 8066 3238 8078 3290
rect 8130 3238 8142 3290
rect 8194 3238 8206 3290
rect 8258 3238 17950 3290
rect 18002 3238 18014 3290
rect 18066 3238 18078 3290
rect 18130 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 27950 3290
rect 28002 3238 28014 3290
rect 28066 3238 28078 3290
rect 28130 3238 28142 3290
rect 28194 3238 28206 3290
rect 28258 3238 37950 3290
rect 38002 3238 38014 3290
rect 38066 3238 38078 3290
rect 38130 3238 38142 3290
rect 38194 3238 38206 3290
rect 38258 3238 47950 3290
rect 48002 3238 48014 3290
rect 48066 3238 48078 3290
rect 48130 3238 48142 3290
rect 48194 3238 48206 3290
rect 48258 3238 49864 3290
rect 1104 3216 49864 3238
rect 7466 3136 7472 3188
rect 7524 3176 7530 3188
rect 17218 3176 17224 3188
rect 7524 3148 17224 3176
rect 7524 3136 7530 3148
rect 17218 3136 17224 3148
rect 17276 3136 17282 3188
rect 18414 3176 18420 3188
rect 17512 3148 18420 3176
rect 17512 3108 17540 3148
rect 18414 3136 18420 3148
rect 18472 3136 18478 3188
rect 21269 3179 21327 3185
rect 21269 3145 21281 3179
rect 21315 3176 21327 3179
rect 23106 3176 23112 3188
rect 21315 3148 23112 3176
rect 21315 3145 21327 3148
rect 21269 3139 21327 3145
rect 23106 3136 23112 3148
rect 23164 3136 23170 3188
rect 23566 3176 23572 3188
rect 23216 3148 23572 3176
rect 19150 3108 19156 3120
rect 16054 3080 17540 3108
rect 17604 3080 19156 3108
rect 934 3000 940 3052
rect 992 3040 998 3052
rect 1581 3043 1639 3049
rect 1581 3040 1593 3043
rect 992 3012 1593 3040
rect 992 3000 998 3012
rect 1581 3009 1593 3012
rect 1627 3009 1639 3043
rect 1581 3003 1639 3009
rect 13814 3000 13820 3052
rect 13872 3040 13878 3052
rect 17604 3049 17632 3080
rect 19150 3068 19156 3080
rect 19208 3068 19214 3120
rect 22094 3108 22100 3120
rect 20180 3080 22100 3108
rect 20180 3049 20208 3080
rect 22094 3068 22100 3080
rect 22152 3108 22158 3120
rect 22646 3108 22652 3120
rect 22152 3080 22652 3108
rect 22152 3068 22158 3080
rect 22646 3068 22652 3080
rect 22704 3068 22710 3120
rect 14553 3043 14611 3049
rect 14553 3040 14565 3043
rect 13872 3012 14565 3040
rect 13872 3000 13878 3012
rect 14553 3009 14565 3012
rect 14599 3009 14611 3043
rect 14553 3003 14611 3009
rect 17589 3043 17647 3049
rect 17589 3009 17601 3043
rect 17635 3009 17647 3043
rect 17589 3003 17647 3009
rect 18325 3043 18383 3049
rect 18325 3009 18337 3043
rect 18371 3009 18383 3043
rect 18325 3003 18383 3009
rect 20165 3043 20223 3049
rect 20165 3009 20177 3043
rect 20211 3009 20223 3043
rect 20165 3003 20223 3009
rect 11054 2932 11060 2984
rect 11112 2972 11118 2984
rect 14829 2975 14887 2981
rect 14829 2972 14841 2975
rect 11112 2944 14841 2972
rect 11112 2932 11118 2944
rect 14829 2941 14841 2944
rect 14875 2941 14887 2975
rect 14829 2935 14887 2941
rect 16301 2975 16359 2981
rect 16301 2941 16313 2975
rect 16347 2972 16359 2975
rect 17862 2972 17868 2984
rect 16347 2944 17868 2972
rect 16347 2941 16359 2944
rect 16301 2935 16359 2941
rect 17862 2932 17868 2944
rect 17920 2932 17926 2984
rect 1765 2907 1823 2913
rect 1765 2873 1777 2907
rect 1811 2904 1823 2907
rect 14458 2904 14464 2916
rect 1811 2876 14464 2904
rect 1811 2873 1823 2876
rect 1765 2867 1823 2873
rect 14458 2864 14464 2876
rect 14516 2864 14522 2916
rect 18340 2904 18368 3003
rect 20806 3000 20812 3052
rect 20864 3000 20870 3052
rect 21450 3000 21456 3052
rect 21508 3000 21514 3052
rect 23216 3049 23244 3148
rect 23566 3136 23572 3148
rect 23624 3176 23630 3188
rect 36814 3176 36820 3188
rect 23624 3148 36820 3176
rect 23624 3136 23630 3148
rect 23290 3068 23296 3120
rect 23348 3108 23354 3120
rect 24397 3111 24455 3117
rect 24397 3108 24409 3111
rect 23348 3080 24409 3108
rect 23348 3068 23354 3080
rect 24397 3077 24409 3080
rect 24443 3077 24455 3111
rect 24397 3071 24455 3077
rect 24486 3068 24492 3120
rect 24544 3108 24550 3120
rect 24544 3080 24886 3108
rect 24544 3068 24550 3080
rect 22189 3043 22247 3049
rect 22189 3009 22201 3043
rect 22235 3040 22247 3043
rect 23201 3043 23259 3049
rect 23201 3040 23213 3043
rect 22235 3012 23213 3040
rect 22235 3009 22247 3012
rect 22189 3003 22247 3009
rect 23201 3009 23213 3012
rect 23247 3009 23259 3043
rect 23201 3003 23259 3009
rect 26142 3000 26148 3052
rect 26200 3040 26206 3052
rect 26513 3043 26571 3049
rect 26513 3040 26525 3043
rect 26200 3012 26525 3040
rect 26200 3000 26206 3012
rect 26513 3009 26525 3012
rect 26559 3009 26571 3043
rect 27356 3040 27384 3148
rect 36814 3136 36820 3148
rect 36872 3136 36878 3188
rect 27522 3068 27528 3120
rect 27580 3108 27586 3120
rect 29638 3108 29644 3120
rect 27580 3080 29644 3108
rect 27580 3068 27586 3080
rect 29638 3068 29644 3080
rect 29696 3068 29702 3120
rect 49145 3111 49203 3117
rect 49145 3077 49157 3111
rect 49191 3108 49203 3111
rect 49234 3108 49240 3120
rect 49191 3080 49240 3108
rect 49191 3077 49203 3080
rect 49145 3071 49203 3077
rect 49234 3068 49240 3080
rect 49292 3068 49298 3120
rect 27433 3043 27491 3049
rect 27433 3040 27445 3043
rect 27356 3012 27445 3040
rect 26513 3003 26571 3009
rect 27433 3009 27445 3012
rect 27479 3009 27491 3043
rect 27433 3003 27491 3009
rect 28810 3000 28816 3052
rect 28868 3040 28874 3052
rect 28905 3043 28963 3049
rect 28905 3040 28917 3043
rect 28868 3012 28917 3040
rect 28868 3000 28874 3012
rect 28905 3009 28917 3012
rect 28951 3009 28963 3043
rect 28905 3003 28963 3009
rect 39850 3000 39856 3052
rect 39908 3040 39914 3052
rect 43993 3043 44051 3049
rect 43993 3040 44005 3043
rect 39908 3012 44005 3040
rect 39908 3000 39914 3012
rect 43993 3009 44005 3012
rect 44039 3009 44051 3043
rect 43993 3003 44051 3009
rect 45830 3000 45836 3052
rect 45888 3000 45894 3052
rect 47210 3000 47216 3052
rect 47268 3040 47274 3052
rect 47949 3043 48007 3049
rect 47949 3040 47961 3043
rect 47268 3012 47961 3040
rect 47268 3000 47274 3012
rect 47949 3009 47961 3012
rect 47995 3009 48007 3043
rect 47949 3003 48007 3009
rect 18414 2932 18420 2984
rect 18472 2972 18478 2984
rect 18601 2975 18659 2981
rect 18601 2972 18613 2975
rect 18472 2944 18613 2972
rect 18472 2932 18478 2944
rect 18601 2941 18613 2944
rect 18647 2941 18659 2975
rect 18601 2935 18659 2941
rect 20898 2932 20904 2984
rect 20956 2972 20962 2984
rect 22002 2972 22008 2984
rect 20956 2944 22008 2972
rect 20956 2932 20962 2944
rect 22002 2932 22008 2944
rect 22060 2972 22066 2984
rect 24121 2975 24179 2981
rect 24121 2972 24133 2975
rect 22060 2944 24133 2972
rect 22060 2932 22066 2944
rect 24121 2941 24133 2944
rect 24167 2941 24179 2975
rect 24121 2935 24179 2941
rect 24486 2932 24492 2984
rect 24544 2972 24550 2984
rect 24544 2944 25820 2972
rect 24544 2932 24550 2944
rect 19981 2907 20039 2913
rect 19981 2904 19993 2907
rect 18340 2876 19993 2904
rect 19981 2873 19993 2876
rect 20027 2873 20039 2907
rect 19981 2867 20039 2873
rect 20625 2907 20683 2913
rect 20625 2873 20637 2907
rect 20671 2904 20683 2907
rect 22370 2904 22376 2916
rect 20671 2876 22376 2904
rect 20671 2873 20683 2876
rect 20625 2867 20683 2873
rect 22370 2864 22376 2876
rect 22428 2864 22434 2916
rect 22646 2864 22652 2916
rect 22704 2864 22710 2916
rect 23106 2864 23112 2916
rect 23164 2904 23170 2916
rect 25792 2904 25820 2944
rect 25866 2932 25872 2984
rect 25924 2972 25930 2984
rect 29181 2975 29239 2981
rect 29181 2972 29193 2975
rect 25924 2944 29193 2972
rect 25924 2932 25930 2944
rect 29181 2941 29193 2944
rect 29227 2941 29239 2975
rect 29181 2935 29239 2941
rect 45189 2975 45247 2981
rect 45189 2941 45201 2975
rect 45235 2972 45247 2975
rect 46750 2972 46756 2984
rect 45235 2944 46756 2972
rect 45235 2941 45247 2944
rect 45189 2935 45247 2941
rect 46750 2932 46756 2944
rect 46808 2932 46814 2984
rect 46842 2932 46848 2984
rect 46900 2932 46906 2984
rect 27522 2904 27528 2916
rect 23164 2876 23796 2904
rect 25792 2876 27528 2904
rect 23164 2864 23170 2876
rect 16390 2796 16396 2848
rect 16448 2836 16454 2848
rect 17405 2839 17463 2845
rect 17405 2836 17417 2839
rect 16448 2808 17417 2836
rect 16448 2796 16454 2808
rect 17405 2805 17417 2808
rect 17451 2805 17463 2839
rect 17405 2799 17463 2805
rect 21174 2796 21180 2848
rect 21232 2836 21238 2848
rect 22281 2839 22339 2845
rect 22281 2836 22293 2839
rect 21232 2808 22293 2836
rect 21232 2796 21238 2808
rect 22281 2805 22293 2808
rect 22327 2805 22339 2839
rect 22281 2799 22339 2805
rect 23290 2796 23296 2848
rect 23348 2796 23354 2848
rect 23658 2796 23664 2848
rect 23716 2796 23722 2848
rect 23768 2836 23796 2876
rect 27522 2864 27528 2876
rect 27580 2864 27586 2916
rect 27724 2876 29040 2904
rect 24578 2836 24584 2848
rect 23768 2808 24584 2836
rect 24578 2796 24584 2808
rect 24636 2796 24642 2848
rect 26329 2839 26387 2845
rect 26329 2805 26341 2839
rect 26375 2836 26387 2839
rect 27154 2836 27160 2848
rect 26375 2808 27160 2836
rect 26375 2805 26387 2808
rect 26329 2799 26387 2805
rect 27154 2796 27160 2808
rect 27212 2796 27218 2848
rect 27724 2845 27752 2876
rect 27709 2839 27767 2845
rect 27709 2805 27721 2839
rect 27755 2805 27767 2839
rect 27709 2799 27767 2805
rect 27798 2796 27804 2848
rect 27856 2836 27862 2848
rect 27893 2839 27951 2845
rect 27893 2836 27905 2839
rect 27856 2808 27905 2836
rect 27856 2796 27862 2808
rect 27893 2805 27905 2808
rect 27939 2805 27951 2839
rect 29012 2836 29040 2876
rect 30653 2839 30711 2845
rect 30653 2836 30665 2839
rect 29012 2808 30665 2836
rect 27893 2799 27951 2805
rect 30653 2805 30665 2808
rect 30699 2836 30711 2839
rect 38102 2836 38108 2848
rect 30699 2808 38108 2836
rect 30699 2805 30711 2808
rect 30653 2799 30711 2805
rect 38102 2796 38108 2808
rect 38160 2796 38166 2848
rect 1104 2746 49864 2768
rect 1104 2694 2950 2746
rect 3002 2694 3014 2746
rect 3066 2694 3078 2746
rect 3130 2694 3142 2746
rect 3194 2694 3206 2746
rect 3258 2694 12950 2746
rect 13002 2694 13014 2746
rect 13066 2694 13078 2746
rect 13130 2694 13142 2746
rect 13194 2694 13206 2746
rect 13258 2694 22950 2746
rect 23002 2694 23014 2746
rect 23066 2694 23078 2746
rect 23130 2694 23142 2746
rect 23194 2694 23206 2746
rect 23258 2694 32950 2746
rect 33002 2694 33014 2746
rect 33066 2694 33078 2746
rect 33130 2694 33142 2746
rect 33194 2694 33206 2746
rect 33258 2694 42950 2746
rect 43002 2694 43014 2746
rect 43066 2694 43078 2746
rect 43130 2694 43142 2746
rect 43194 2694 43206 2746
rect 43258 2694 49864 2746
rect 1104 2672 49864 2694
rect 2501 2635 2559 2641
rect 2501 2601 2513 2635
rect 2547 2632 2559 2635
rect 22462 2632 22468 2644
rect 2547 2604 22468 2632
rect 2547 2601 2559 2604
rect 2501 2595 2559 2601
rect 22462 2592 22468 2604
rect 22520 2592 22526 2644
rect 28902 2592 28908 2644
rect 28960 2632 28966 2644
rect 28997 2635 29055 2641
rect 28997 2632 29009 2635
rect 28960 2604 29009 2632
rect 28960 2592 28966 2604
rect 28997 2601 29009 2604
rect 29043 2601 29055 2635
rect 28997 2595 29055 2601
rect 34422 2592 34428 2644
rect 34480 2632 34486 2644
rect 35069 2635 35127 2641
rect 35069 2632 35081 2635
rect 34480 2604 35081 2632
rect 34480 2592 34486 2604
rect 35069 2601 35081 2604
rect 35115 2601 35127 2635
rect 35069 2595 35127 2601
rect 1765 2567 1823 2573
rect 1765 2533 1777 2567
rect 1811 2533 1823 2567
rect 1765 2527 1823 2533
rect 3053 2567 3111 2573
rect 3053 2533 3065 2567
rect 3099 2564 3111 2567
rect 9677 2567 9735 2573
rect 3099 2536 6914 2564
rect 3099 2533 3111 2536
rect 3053 2527 3111 2533
rect 1780 2496 1808 2527
rect 6886 2496 6914 2536
rect 9677 2533 9689 2567
rect 9723 2564 9735 2567
rect 11054 2564 11060 2576
rect 9723 2536 11060 2564
rect 9723 2533 9735 2536
rect 9677 2527 9735 2533
rect 11054 2524 11060 2536
rect 11112 2524 11118 2576
rect 13446 2564 13452 2576
rect 11164 2536 13452 2564
rect 11164 2496 11192 2536
rect 13446 2524 13452 2536
rect 13504 2524 13510 2576
rect 19429 2567 19487 2573
rect 19429 2533 19441 2567
rect 19475 2564 19487 2567
rect 19475 2536 20116 2564
rect 19475 2533 19487 2536
rect 19429 2527 19487 2533
rect 1780 2468 4384 2496
rect 6886 2468 11192 2496
rect 934 2388 940 2440
rect 992 2428 998 2440
rect 1581 2431 1639 2437
rect 1581 2428 1593 2431
rect 992 2400 1593 2428
rect 992 2388 998 2400
rect 1581 2397 1593 2400
rect 1627 2397 1639 2431
rect 1581 2391 1639 2397
rect 3237 2431 3295 2437
rect 3237 2397 3249 2431
rect 3283 2397 3295 2431
rect 3237 2391 3295 2397
rect 1210 2320 1216 2372
rect 1268 2360 1274 2372
rect 2409 2363 2467 2369
rect 2409 2360 2421 2363
rect 1268 2332 2421 2360
rect 1268 2320 1274 2332
rect 2409 2329 2421 2332
rect 2455 2329 2467 2363
rect 2409 2323 2467 2329
rect 1302 2252 1308 2304
rect 1360 2292 1366 2304
rect 3252 2292 3280 2391
rect 4356 2360 4384 2468
rect 11698 2456 11704 2508
rect 11756 2496 11762 2508
rect 12253 2499 12311 2505
rect 12253 2496 12265 2499
rect 11756 2468 12265 2496
rect 11756 2456 11762 2468
rect 12253 2465 12265 2468
rect 12299 2465 12311 2499
rect 12253 2459 12311 2465
rect 13814 2456 13820 2508
rect 13872 2496 13878 2508
rect 14737 2499 14795 2505
rect 14737 2496 14749 2499
rect 13872 2468 14749 2496
rect 13872 2456 13878 2468
rect 14737 2465 14749 2468
rect 14783 2465 14795 2499
rect 14737 2459 14795 2465
rect 15930 2456 15936 2508
rect 15988 2496 15994 2508
rect 17313 2499 17371 2505
rect 17313 2496 17325 2499
rect 15988 2468 17325 2496
rect 15988 2456 15994 2468
rect 17313 2465 17325 2468
rect 17359 2465 17371 2499
rect 17313 2459 17371 2465
rect 9582 2388 9588 2440
rect 9640 2428 9646 2440
rect 9861 2431 9919 2437
rect 9861 2428 9873 2431
rect 9640 2400 9873 2428
rect 9640 2388 9646 2400
rect 9861 2397 9873 2400
rect 9907 2397 9919 2431
rect 9861 2391 9919 2397
rect 11977 2431 12035 2437
rect 11977 2397 11989 2431
rect 12023 2428 12035 2431
rect 12526 2428 12532 2440
rect 12023 2400 12532 2428
rect 12023 2397 12035 2400
rect 11977 2391 12035 2397
rect 12526 2388 12532 2400
rect 12584 2388 12590 2440
rect 14461 2431 14519 2437
rect 14461 2397 14473 2431
rect 14507 2428 14519 2431
rect 16390 2428 16396 2440
rect 14507 2400 16396 2428
rect 14507 2397 14519 2400
rect 14461 2391 14519 2397
rect 16390 2388 16396 2400
rect 16448 2388 16454 2440
rect 17037 2431 17095 2437
rect 17037 2397 17049 2431
rect 17083 2428 17095 2431
rect 18877 2431 18935 2437
rect 17083 2400 18736 2428
rect 17083 2397 17095 2400
rect 17037 2391 17095 2397
rect 14642 2360 14648 2372
rect 4356 2332 14648 2360
rect 14642 2320 14648 2332
rect 14700 2320 14706 2372
rect 18708 2301 18736 2400
rect 18877 2397 18889 2431
rect 18923 2428 18935 2431
rect 19518 2428 19524 2440
rect 18923 2400 19524 2428
rect 18923 2397 18935 2400
rect 18877 2391 18935 2397
rect 19518 2388 19524 2400
rect 19576 2388 19582 2440
rect 19610 2388 19616 2440
rect 19668 2388 19674 2440
rect 20088 2437 20116 2536
rect 24118 2524 24124 2576
rect 24176 2564 24182 2576
rect 30837 2567 30895 2573
rect 30837 2564 30849 2567
rect 24176 2536 30849 2564
rect 24176 2524 24182 2536
rect 30837 2533 30849 2536
rect 30883 2533 30895 2567
rect 30837 2527 30895 2533
rect 34330 2524 34336 2576
rect 34388 2564 34394 2576
rect 34388 2536 43852 2564
rect 34388 2524 34394 2536
rect 20162 2456 20168 2508
rect 20220 2496 20226 2508
rect 20533 2499 20591 2505
rect 20533 2496 20545 2499
rect 20220 2468 20545 2496
rect 20220 2456 20226 2468
rect 20533 2465 20545 2468
rect 20579 2465 20591 2499
rect 20533 2459 20591 2465
rect 22278 2456 22284 2508
rect 22336 2496 22342 2508
rect 22833 2499 22891 2505
rect 22833 2496 22845 2499
rect 22336 2468 22845 2496
rect 22336 2456 22342 2468
rect 22833 2465 22845 2468
rect 22879 2465 22891 2499
rect 22833 2459 22891 2465
rect 24394 2456 24400 2508
rect 24452 2496 24458 2508
rect 25041 2499 25099 2505
rect 25041 2496 25053 2499
rect 24452 2468 25053 2496
rect 24452 2456 24458 2468
rect 25041 2465 25053 2468
rect 25087 2465 25099 2499
rect 25041 2459 25099 2465
rect 26510 2456 26516 2508
rect 26568 2496 26574 2508
rect 27617 2499 27675 2505
rect 27617 2496 27629 2499
rect 26568 2468 27629 2496
rect 26568 2456 26574 2468
rect 27617 2465 27629 2468
rect 27663 2465 27675 2499
rect 27617 2459 27675 2465
rect 36814 2456 36820 2508
rect 36872 2496 36878 2508
rect 37737 2499 37795 2505
rect 37737 2496 37749 2499
rect 36872 2468 37749 2496
rect 36872 2456 36878 2468
rect 37737 2465 37749 2468
rect 37783 2465 37795 2499
rect 37737 2459 37795 2465
rect 41322 2456 41328 2508
rect 41380 2496 41386 2508
rect 43824 2505 43852 2536
rect 41417 2499 41475 2505
rect 41417 2496 41429 2499
rect 41380 2468 41429 2496
rect 41380 2456 41386 2468
rect 41417 2465 41429 2468
rect 41463 2465 41475 2499
rect 41417 2459 41475 2465
rect 43809 2499 43867 2505
rect 43809 2465 43821 2499
rect 43855 2465 43867 2499
rect 43809 2459 43867 2465
rect 49142 2456 49148 2508
rect 49200 2456 49206 2508
rect 20073 2431 20131 2437
rect 20073 2397 20085 2431
rect 20119 2397 20131 2431
rect 20073 2391 20131 2397
rect 22370 2388 22376 2440
rect 22428 2388 22434 2440
rect 24578 2388 24584 2440
rect 24636 2388 24642 2440
rect 27154 2388 27160 2440
rect 27212 2388 27218 2440
rect 28626 2388 28632 2440
rect 28684 2428 28690 2440
rect 29181 2431 29239 2437
rect 29181 2428 29193 2431
rect 28684 2400 29193 2428
rect 28684 2388 28690 2400
rect 29181 2397 29193 2400
rect 29227 2397 29239 2431
rect 29181 2391 29239 2397
rect 30742 2388 30748 2440
rect 30800 2428 30806 2440
rect 31021 2431 31079 2437
rect 31021 2428 31033 2431
rect 30800 2400 31033 2428
rect 30800 2388 30806 2400
rect 31021 2397 31033 2400
rect 31067 2397 31079 2431
rect 31021 2391 31079 2397
rect 32858 2388 32864 2440
rect 32916 2428 32922 2440
rect 33137 2431 33195 2437
rect 33137 2428 33149 2431
rect 32916 2400 33149 2428
rect 32916 2388 32922 2400
rect 33137 2397 33149 2400
rect 33183 2397 33195 2431
rect 33137 2391 33195 2397
rect 34974 2388 34980 2440
rect 35032 2428 35038 2440
rect 35253 2431 35311 2437
rect 35253 2428 35265 2431
rect 35032 2400 35265 2428
rect 35032 2388 35038 2400
rect 35253 2397 35265 2400
rect 35299 2397 35311 2431
rect 35253 2391 35311 2397
rect 37090 2388 37096 2440
rect 37148 2428 37154 2440
rect 37461 2431 37519 2437
rect 37461 2428 37473 2431
rect 37148 2400 37473 2428
rect 37148 2388 37154 2400
rect 37461 2397 37473 2400
rect 37507 2397 37519 2431
rect 37461 2391 37519 2397
rect 38102 2388 38108 2440
rect 38160 2428 38166 2440
rect 40681 2431 40739 2437
rect 40681 2428 40693 2431
rect 38160 2400 40693 2428
rect 38160 2388 38166 2400
rect 40681 2397 40693 2400
rect 40727 2397 40739 2431
rect 40681 2391 40739 2397
rect 43438 2388 43444 2440
rect 43496 2428 43502 2440
rect 43533 2431 43591 2437
rect 43533 2428 43545 2431
rect 43496 2400 43545 2428
rect 43496 2388 43502 2400
rect 43533 2397 43545 2400
rect 43579 2397 43591 2431
rect 43533 2391 43591 2397
rect 44634 2388 44640 2440
rect 44692 2428 44698 2440
rect 45833 2431 45891 2437
rect 45833 2428 45845 2431
rect 44692 2400 45845 2428
rect 44692 2388 44698 2400
rect 45833 2397 45845 2400
rect 45879 2397 45891 2431
rect 45833 2391 45891 2397
rect 47118 2388 47124 2440
rect 47176 2428 47182 2440
rect 47949 2431 48007 2437
rect 47949 2428 47961 2431
rect 47176 2400 47961 2428
rect 47176 2388 47182 2400
rect 47949 2397 47961 2400
rect 47995 2397 48007 2431
rect 47949 2391 48007 2397
rect 47029 2363 47087 2369
rect 47029 2329 47041 2363
rect 47075 2360 47087 2363
rect 48498 2360 48504 2372
rect 47075 2332 48504 2360
rect 47075 2329 47087 2332
rect 47029 2323 47087 2329
rect 48498 2320 48504 2332
rect 48556 2320 48562 2372
rect 1360 2264 3280 2292
rect 18693 2295 18751 2301
rect 1360 2252 1366 2264
rect 18693 2261 18705 2295
rect 18739 2261 18751 2295
rect 18693 2255 18751 2261
rect 28718 2252 28724 2304
rect 28776 2292 28782 2304
rect 32953 2295 33011 2301
rect 32953 2292 32965 2295
rect 28776 2264 32965 2292
rect 28776 2252 28782 2264
rect 32953 2261 32965 2264
rect 32999 2261 33011 2295
rect 32953 2255 33011 2261
rect 1104 2202 49864 2224
rect 1104 2150 7950 2202
rect 8002 2150 8014 2202
rect 8066 2150 8078 2202
rect 8130 2150 8142 2202
rect 8194 2150 8206 2202
rect 8258 2150 17950 2202
rect 18002 2150 18014 2202
rect 18066 2150 18078 2202
rect 18130 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 27950 2202
rect 28002 2150 28014 2202
rect 28066 2150 28078 2202
rect 28130 2150 28142 2202
rect 28194 2150 28206 2202
rect 28258 2150 37950 2202
rect 38002 2150 38014 2202
rect 38066 2150 38078 2202
rect 38130 2150 38142 2202
rect 38194 2150 38206 2202
rect 38258 2150 47950 2202
rect 48002 2150 48014 2202
rect 48066 2150 48078 2202
rect 48130 2150 48142 2202
rect 48194 2150 48206 2202
rect 48258 2150 49864 2202
rect 1104 2128 49864 2150
<< via1 >>
rect 3424 25168 3476 25220
rect 9220 25168 9272 25220
rect 3332 25032 3384 25084
rect 8852 25032 8904 25084
rect 32128 24896 32180 24948
rect 39212 24896 39264 24948
rect 28816 24828 28868 24880
rect 48688 24828 48740 24880
rect 24032 24760 24084 24812
rect 27804 24760 27856 24812
rect 32864 24760 32916 24812
rect 36544 24760 36596 24812
rect 38936 24760 38988 24812
rect 41788 24760 41840 24812
rect 19064 24692 19116 24744
rect 22100 24692 22152 24744
rect 17592 24624 17644 24676
rect 27436 24692 27488 24744
rect 36268 24692 36320 24744
rect 40684 24692 40736 24744
rect 3148 24556 3200 24608
rect 5724 24556 5776 24608
rect 17776 24556 17828 24608
rect 20076 24556 20128 24608
rect 21456 24556 21508 24608
rect 29092 24624 29144 24676
rect 29276 24624 29328 24676
rect 35072 24624 35124 24676
rect 35716 24624 35768 24676
rect 43536 24624 43588 24676
rect 24768 24556 24820 24608
rect 31208 24556 31260 24608
rect 34980 24556 35032 24608
rect 40040 24556 40092 24608
rect 2950 24454 3002 24506
rect 3014 24454 3066 24506
rect 3078 24454 3130 24506
rect 3142 24454 3194 24506
rect 3206 24454 3258 24506
rect 12950 24454 13002 24506
rect 13014 24454 13066 24506
rect 13078 24454 13130 24506
rect 13142 24454 13194 24506
rect 13206 24454 13258 24506
rect 22950 24454 23002 24506
rect 23014 24454 23066 24506
rect 23078 24454 23130 24506
rect 23142 24454 23194 24506
rect 23206 24454 23258 24506
rect 32950 24454 33002 24506
rect 33014 24454 33066 24506
rect 33078 24454 33130 24506
rect 33142 24454 33194 24506
rect 33206 24454 33258 24506
rect 42950 24454 43002 24506
rect 43014 24454 43066 24506
rect 43078 24454 43130 24506
rect 43142 24454 43194 24506
rect 43206 24454 43258 24506
rect 2780 24352 2832 24404
rect 6276 24352 6328 24404
rect 6736 24284 6788 24336
rect 3516 24216 3568 24268
rect 8668 24216 8720 24268
rect 11888 24284 11940 24336
rect 16028 24284 16080 24336
rect 19432 24284 19484 24336
rect 2320 24148 2372 24200
rect 4712 24148 4764 24200
rect 6552 24148 6604 24200
rect 7472 24148 7524 24200
rect 9680 24148 9732 24200
rect 13820 24216 13872 24268
rect 17684 24216 17736 24268
rect 19524 24216 19576 24268
rect 10324 24080 10376 24132
rect 12624 24148 12676 24200
rect 14464 24191 14516 24200
rect 14464 24157 14473 24191
rect 14473 24157 14507 24191
rect 14507 24157 14516 24191
rect 14464 24148 14516 24157
rect 16580 24148 16632 24200
rect 17592 24191 17644 24200
rect 17592 24157 17601 24191
rect 17601 24157 17635 24191
rect 17635 24157 17644 24191
rect 17592 24148 17644 24157
rect 24032 24352 24084 24404
rect 24124 24352 24176 24404
rect 20536 24284 20588 24336
rect 13636 24080 13688 24132
rect 13728 24080 13780 24132
rect 4620 24012 4672 24064
rect 7472 24012 7524 24064
rect 9128 24055 9180 24064
rect 9128 24021 9137 24055
rect 9137 24021 9171 24055
rect 9171 24021 9180 24055
rect 9128 24012 9180 24021
rect 13452 24012 13504 24064
rect 20904 24259 20956 24268
rect 20904 24225 20913 24259
rect 20913 24225 20947 24259
rect 20947 24225 20956 24259
rect 20904 24216 20956 24225
rect 23572 24284 23624 24336
rect 24952 24284 25004 24336
rect 26148 24284 26200 24336
rect 28724 24284 28776 24336
rect 28908 24284 28960 24336
rect 25136 24259 25188 24268
rect 25136 24225 25145 24259
rect 25145 24225 25179 24259
rect 25179 24225 25188 24259
rect 25136 24216 25188 24225
rect 26332 24259 26384 24268
rect 26332 24225 26341 24259
rect 26341 24225 26375 24259
rect 26375 24225 26384 24259
rect 26332 24216 26384 24225
rect 27988 24216 28040 24268
rect 22192 24191 22244 24200
rect 22192 24157 22201 24191
rect 22201 24157 22235 24191
rect 22235 24157 22244 24191
rect 22192 24148 22244 24157
rect 25412 24148 25464 24200
rect 26056 24148 26108 24200
rect 26700 24148 26752 24200
rect 28724 24191 28776 24200
rect 28724 24157 28733 24191
rect 28733 24157 28767 24191
rect 28767 24157 28776 24191
rect 28724 24148 28776 24157
rect 26424 24080 26476 24132
rect 27252 24123 27304 24132
rect 27252 24089 27261 24123
rect 27261 24089 27295 24123
rect 27295 24089 27304 24123
rect 27252 24080 27304 24089
rect 29092 24080 29144 24132
rect 31208 24191 31260 24200
rect 31208 24157 31217 24191
rect 31217 24157 31251 24191
rect 31251 24157 31260 24191
rect 31208 24148 31260 24157
rect 31484 24352 31536 24404
rect 31852 24284 31904 24336
rect 37556 24352 37608 24404
rect 38568 24352 38620 24404
rect 39212 24395 39264 24404
rect 39212 24361 39221 24395
rect 39221 24361 39255 24395
rect 39255 24361 39264 24395
rect 39212 24352 39264 24361
rect 40040 24395 40092 24404
rect 40040 24361 40049 24395
rect 40049 24361 40083 24395
rect 40083 24361 40092 24395
rect 40040 24352 40092 24361
rect 40684 24395 40736 24404
rect 40684 24361 40693 24395
rect 40693 24361 40727 24395
rect 40727 24361 40736 24395
rect 40684 24352 40736 24361
rect 48320 24395 48372 24404
rect 48320 24361 48329 24395
rect 48329 24361 48363 24395
rect 48363 24361 48372 24395
rect 48320 24352 48372 24361
rect 39672 24284 39724 24336
rect 39948 24284 40000 24336
rect 40960 24284 41012 24336
rect 35072 24191 35124 24200
rect 35072 24157 35081 24191
rect 35081 24157 35115 24191
rect 35115 24157 35124 24191
rect 35072 24148 35124 24157
rect 36360 24191 36412 24200
rect 36360 24157 36369 24191
rect 36369 24157 36403 24191
rect 36403 24157 36412 24191
rect 36360 24148 36412 24157
rect 36544 24259 36596 24268
rect 36544 24225 36553 24259
rect 36553 24225 36587 24259
rect 36587 24225 36596 24259
rect 36544 24216 36596 24225
rect 37556 24216 37608 24268
rect 37924 24259 37976 24268
rect 37924 24225 37933 24259
rect 37933 24225 37967 24259
rect 37967 24225 37976 24259
rect 37924 24216 37976 24225
rect 38384 24216 38436 24268
rect 38660 24216 38712 24268
rect 26240 24012 26292 24064
rect 27712 24012 27764 24064
rect 28448 24012 28500 24064
rect 29184 24012 29236 24064
rect 30472 24012 30524 24064
rect 31944 24012 31996 24064
rect 39120 24148 39172 24200
rect 39212 24148 39264 24200
rect 48228 24216 48280 24268
rect 33968 24055 34020 24064
rect 33968 24021 33977 24055
rect 33977 24021 34011 24055
rect 34011 24021 34020 24055
rect 33968 24012 34020 24021
rect 34888 24055 34940 24064
rect 34888 24021 34897 24055
rect 34897 24021 34931 24055
rect 34931 24021 34940 24055
rect 34888 24012 34940 24021
rect 35624 24012 35676 24064
rect 37464 24055 37516 24064
rect 37464 24021 37473 24055
rect 37473 24021 37507 24055
rect 37507 24021 37516 24055
rect 37464 24012 37516 24021
rect 37740 24080 37792 24132
rect 42156 24148 42208 24200
rect 44732 24148 44784 24200
rect 45560 24148 45612 24200
rect 46020 24148 46072 24200
rect 47308 24148 47360 24200
rect 48596 24148 48648 24200
rect 40960 24080 41012 24132
rect 41144 24080 41196 24132
rect 46940 24123 46992 24132
rect 46940 24089 46949 24123
rect 46949 24089 46983 24123
rect 46983 24089 46992 24123
rect 46940 24080 46992 24089
rect 39856 24012 39908 24064
rect 40776 24012 40828 24064
rect 43352 24012 43404 24064
rect 46112 24055 46164 24064
rect 46112 24021 46121 24055
rect 46121 24021 46155 24055
rect 46155 24021 46164 24055
rect 46112 24012 46164 24021
rect 7950 23910 8002 23962
rect 8014 23910 8066 23962
rect 8078 23910 8130 23962
rect 8142 23910 8194 23962
rect 8206 23910 8258 23962
rect 17950 23910 18002 23962
rect 18014 23910 18066 23962
rect 18078 23910 18130 23962
rect 18142 23910 18194 23962
rect 18206 23910 18258 23962
rect 27950 23910 28002 23962
rect 28014 23910 28066 23962
rect 28078 23910 28130 23962
rect 28142 23910 28194 23962
rect 28206 23910 28258 23962
rect 37950 23910 38002 23962
rect 38014 23910 38066 23962
rect 38078 23910 38130 23962
rect 38142 23910 38194 23962
rect 38206 23910 38258 23962
rect 47950 23910 48002 23962
rect 48014 23910 48066 23962
rect 48078 23910 48130 23962
rect 48142 23910 48194 23962
rect 48206 23910 48258 23962
rect 6552 23851 6604 23860
rect 6552 23817 6561 23851
rect 6561 23817 6595 23851
rect 6595 23817 6604 23851
rect 6552 23808 6604 23817
rect 4160 23740 4212 23792
rect 3516 23672 3568 23724
rect 4620 23715 4672 23724
rect 4620 23681 4629 23715
rect 4629 23681 4663 23715
rect 4663 23681 4672 23715
rect 4620 23672 4672 23681
rect 7288 23672 7340 23724
rect 12716 23808 12768 23860
rect 9312 23740 9364 23792
rect 10600 23740 10652 23792
rect 14372 23783 14424 23792
rect 14372 23749 14381 23783
rect 14381 23749 14415 23783
rect 14415 23749 14424 23783
rect 14372 23740 14424 23749
rect 16120 23783 16172 23792
rect 16120 23749 16129 23783
rect 16129 23749 16163 23783
rect 16163 23749 16172 23783
rect 16120 23740 16172 23749
rect 18328 23740 18380 23792
rect 5448 23647 5500 23656
rect 5448 23613 5457 23647
rect 5457 23613 5491 23647
rect 5491 23613 5500 23647
rect 5448 23604 5500 23613
rect 9588 23604 9640 23656
rect 3424 23536 3476 23588
rect 5540 23536 5592 23588
rect 12072 23647 12124 23656
rect 12072 23613 12081 23647
rect 12081 23613 12115 23647
rect 12115 23613 12124 23647
rect 12072 23604 12124 23613
rect 12440 23536 12492 23588
rect 13452 23715 13504 23724
rect 13452 23681 13461 23715
rect 13461 23681 13495 23715
rect 13495 23681 13504 23715
rect 13452 23672 13504 23681
rect 19064 23783 19116 23792
rect 19064 23749 19073 23783
rect 19073 23749 19107 23783
rect 19107 23749 19116 23783
rect 19064 23740 19116 23749
rect 20444 23808 20496 23860
rect 23480 23808 23532 23860
rect 18788 23715 18840 23724
rect 18788 23681 18797 23715
rect 18797 23681 18831 23715
rect 18831 23681 18840 23715
rect 18788 23672 18840 23681
rect 20168 23672 20220 23724
rect 17960 23604 18012 23656
rect 20260 23604 20312 23656
rect 20536 23740 20588 23792
rect 27804 23808 27856 23860
rect 25228 23740 25280 23792
rect 26424 23740 26476 23792
rect 27344 23740 27396 23792
rect 21456 23715 21508 23724
rect 21456 23681 21465 23715
rect 21465 23681 21499 23715
rect 21499 23681 21508 23715
rect 21456 23672 21508 23681
rect 23480 23672 23532 23724
rect 27160 23672 27212 23724
rect 27436 23715 27488 23724
rect 27436 23681 27445 23715
rect 27445 23681 27479 23715
rect 27479 23681 27488 23715
rect 27436 23672 27488 23681
rect 33968 23808 34020 23860
rect 37464 23808 37516 23860
rect 39856 23851 39908 23860
rect 39856 23817 39865 23851
rect 39865 23817 39899 23851
rect 39899 23817 39908 23851
rect 39856 23808 39908 23817
rect 30748 23740 30800 23792
rect 34152 23740 34204 23792
rect 34336 23740 34388 23792
rect 35256 23740 35308 23792
rect 20076 23536 20128 23588
rect 4804 23468 4856 23520
rect 9680 23468 9732 23520
rect 16580 23468 16632 23520
rect 18788 23468 18840 23520
rect 20352 23468 20404 23520
rect 20536 23511 20588 23520
rect 20536 23477 20545 23511
rect 20545 23477 20579 23511
rect 20579 23477 20588 23511
rect 20536 23468 20588 23477
rect 21272 23511 21324 23520
rect 21272 23477 21281 23511
rect 21281 23477 21315 23511
rect 21315 23477 21324 23511
rect 21272 23468 21324 23477
rect 23296 23604 23348 23656
rect 24860 23647 24912 23656
rect 24860 23613 24869 23647
rect 24869 23613 24903 23647
rect 24903 23613 24912 23647
rect 24860 23604 24912 23613
rect 27620 23604 27672 23656
rect 32680 23715 32732 23724
rect 32680 23681 32689 23715
rect 32689 23681 32723 23715
rect 32723 23681 32732 23715
rect 32680 23672 32732 23681
rect 37372 23672 37424 23724
rect 37832 23715 37884 23724
rect 37832 23681 37841 23715
rect 37841 23681 37875 23715
rect 37875 23681 37884 23715
rect 37832 23672 37884 23681
rect 38752 23672 38804 23724
rect 29736 23604 29788 23656
rect 30012 23647 30064 23656
rect 30012 23613 30021 23647
rect 30021 23613 30055 23647
rect 30055 23613 30064 23647
rect 30012 23604 30064 23613
rect 24768 23536 24820 23588
rect 25136 23468 25188 23520
rect 25228 23468 25280 23520
rect 29276 23536 29328 23588
rect 29368 23536 29420 23588
rect 32404 23604 32456 23656
rect 32864 23604 32916 23656
rect 26608 23511 26660 23520
rect 26608 23477 26617 23511
rect 26617 23477 26651 23511
rect 26651 23477 26660 23511
rect 26608 23468 26660 23477
rect 28632 23468 28684 23520
rect 29000 23468 29052 23520
rect 30288 23468 30340 23520
rect 31484 23468 31536 23520
rect 31668 23468 31720 23520
rect 33324 23604 33376 23656
rect 33876 23647 33928 23656
rect 33876 23613 33885 23647
rect 33885 23613 33919 23647
rect 33919 23613 33928 23647
rect 33876 23604 33928 23613
rect 34244 23604 34296 23656
rect 34888 23536 34940 23588
rect 35624 23536 35676 23588
rect 36544 23647 36596 23656
rect 36544 23613 36553 23647
rect 36553 23613 36587 23647
rect 36587 23613 36596 23647
rect 36544 23604 36596 23613
rect 36728 23647 36780 23656
rect 36728 23613 36737 23647
rect 36737 23613 36771 23647
rect 36771 23613 36780 23647
rect 36728 23604 36780 23613
rect 38292 23604 38344 23656
rect 40040 23740 40092 23792
rect 35348 23511 35400 23520
rect 35348 23477 35357 23511
rect 35357 23477 35391 23511
rect 35391 23477 35400 23511
rect 35348 23468 35400 23477
rect 35440 23468 35492 23520
rect 38568 23468 38620 23520
rect 39948 23647 40000 23656
rect 39948 23613 39957 23647
rect 39957 23613 39991 23647
rect 39991 23613 40000 23647
rect 39948 23604 40000 23613
rect 39764 23536 39816 23588
rect 41236 23808 41288 23860
rect 41328 23740 41380 23792
rect 41420 23740 41472 23792
rect 46848 23783 46900 23792
rect 46848 23749 46857 23783
rect 46857 23749 46891 23783
rect 46891 23749 46900 23783
rect 46848 23740 46900 23749
rect 47860 23740 47912 23792
rect 45468 23715 45520 23724
rect 45468 23681 45477 23715
rect 45477 23681 45511 23715
rect 45511 23681 45520 23715
rect 45468 23672 45520 23681
rect 48780 23715 48832 23724
rect 48780 23681 48789 23715
rect 48789 23681 48823 23715
rect 48823 23681 48832 23715
rect 48780 23672 48832 23681
rect 41236 23604 41288 23656
rect 43536 23647 43588 23656
rect 43536 23613 43545 23647
rect 43545 23613 43579 23647
rect 43579 23613 43588 23647
rect 43536 23604 43588 23613
rect 40500 23468 40552 23520
rect 42800 23468 42852 23520
rect 47124 23468 47176 23520
rect 2950 23366 3002 23418
rect 3014 23366 3066 23418
rect 3078 23366 3130 23418
rect 3142 23366 3194 23418
rect 3206 23366 3258 23418
rect 12950 23366 13002 23418
rect 13014 23366 13066 23418
rect 13078 23366 13130 23418
rect 13142 23366 13194 23418
rect 13206 23366 13258 23418
rect 22950 23366 23002 23418
rect 23014 23366 23066 23418
rect 23078 23366 23130 23418
rect 23142 23366 23194 23418
rect 23206 23366 23258 23418
rect 32950 23366 33002 23418
rect 33014 23366 33066 23418
rect 33078 23366 33130 23418
rect 33142 23366 33194 23418
rect 33206 23366 33258 23418
rect 42950 23366 43002 23418
rect 43014 23366 43066 23418
rect 43078 23366 43130 23418
rect 43142 23366 43194 23418
rect 43206 23366 43258 23418
rect 1584 23196 1636 23248
rect 4344 23196 4396 23248
rect 7748 23196 7800 23248
rect 4436 23060 4488 23112
rect 5264 23060 5316 23112
rect 6092 23171 6144 23180
rect 6092 23137 6101 23171
rect 6101 23137 6135 23171
rect 6135 23137 6144 23171
rect 6092 23128 6144 23137
rect 7840 23171 7892 23180
rect 7840 23137 7849 23171
rect 7849 23137 7883 23171
rect 7883 23137 7892 23171
rect 7840 23128 7892 23137
rect 2780 23035 2832 23044
rect 2780 23001 2789 23035
rect 2789 23001 2823 23035
rect 2823 23001 2832 23035
rect 2780 22992 2832 23001
rect 2872 22992 2924 23044
rect 4160 22992 4212 23044
rect 3608 22924 3660 22976
rect 7104 23060 7156 23112
rect 8300 23060 8352 23112
rect 9128 23060 9180 23112
rect 17592 23264 17644 23316
rect 17960 23264 18012 23316
rect 13820 23196 13872 23248
rect 11244 23171 11296 23180
rect 11244 23137 11253 23171
rect 11253 23137 11287 23171
rect 11287 23137 11296 23171
rect 11244 23128 11296 23137
rect 13360 23171 13412 23180
rect 13360 23137 13369 23171
rect 13369 23137 13403 23171
rect 13403 23137 13412 23171
rect 13360 23128 13412 23137
rect 15752 23171 15804 23180
rect 15752 23137 15761 23171
rect 15761 23137 15795 23171
rect 15795 23137 15804 23171
rect 15752 23128 15804 23137
rect 22008 23264 22060 23316
rect 22192 23264 22244 23316
rect 22836 23264 22888 23316
rect 23388 23264 23440 23316
rect 22100 23196 22152 23248
rect 23296 23196 23348 23248
rect 20352 23171 20404 23180
rect 20352 23137 20361 23171
rect 20361 23137 20395 23171
rect 20395 23137 20404 23171
rect 20352 23128 20404 23137
rect 20720 23128 20772 23180
rect 10692 23103 10744 23112
rect 10692 23069 10701 23103
rect 10701 23069 10735 23103
rect 10735 23069 10744 23103
rect 10692 23060 10744 23069
rect 14372 23060 14424 23112
rect 15108 23060 15160 23112
rect 5448 22992 5500 23044
rect 7656 22992 7708 23044
rect 17040 23060 17092 23112
rect 22744 23128 22796 23180
rect 27804 23264 27856 23316
rect 27896 23307 27948 23316
rect 27896 23273 27905 23307
rect 27905 23273 27939 23307
rect 27939 23273 27948 23307
rect 27896 23264 27948 23273
rect 29736 23307 29788 23316
rect 29736 23273 29745 23307
rect 29745 23273 29779 23307
rect 29779 23273 29788 23307
rect 29736 23264 29788 23273
rect 30564 23264 30616 23316
rect 25136 23196 25188 23248
rect 26608 23128 26660 23180
rect 26976 23128 27028 23180
rect 21916 23060 21968 23112
rect 17316 22992 17368 23044
rect 17500 22992 17552 23044
rect 18696 22992 18748 23044
rect 9312 22967 9364 22976
rect 9312 22933 9321 22967
rect 9321 22933 9355 22967
rect 9355 22933 9364 22967
rect 9312 22924 9364 22933
rect 12808 22924 12860 22976
rect 19064 22924 19116 22976
rect 20628 23035 20680 23044
rect 20628 23001 20637 23035
rect 20637 23001 20671 23035
rect 20671 23001 20680 23035
rect 20628 22992 20680 23001
rect 22008 22992 22060 23044
rect 22284 22992 22336 23044
rect 24952 23060 25004 23112
rect 25688 23103 25740 23112
rect 25688 23069 25697 23103
rect 25697 23069 25731 23103
rect 25731 23069 25740 23103
rect 25688 23060 25740 23069
rect 30656 23196 30708 23248
rect 30288 23128 30340 23180
rect 31668 23171 31720 23180
rect 31668 23137 31677 23171
rect 31677 23137 31711 23171
rect 31711 23137 31720 23171
rect 31668 23128 31720 23137
rect 30012 23060 30064 23112
rect 33048 23264 33100 23316
rect 34704 23264 34756 23316
rect 35164 23264 35216 23316
rect 38568 23264 38620 23316
rect 38660 23264 38712 23316
rect 40040 23307 40092 23316
rect 40040 23273 40049 23307
rect 40049 23273 40083 23307
rect 40083 23273 40092 23307
rect 40040 23264 40092 23273
rect 40224 23264 40276 23316
rect 41604 23264 41656 23316
rect 32956 23196 33008 23248
rect 38844 23196 38896 23248
rect 43352 23264 43404 23316
rect 33324 23128 33376 23180
rect 34612 23128 34664 23180
rect 21916 22924 21968 22976
rect 22100 22967 22152 22976
rect 22100 22933 22109 22967
rect 22109 22933 22143 22967
rect 22143 22933 22152 22967
rect 22100 22924 22152 22933
rect 22192 22924 22244 22976
rect 23664 22967 23716 22976
rect 23664 22933 23673 22967
rect 23673 22933 23707 22967
rect 23707 22933 23716 22967
rect 23664 22924 23716 22933
rect 24676 23035 24728 23044
rect 24676 23001 24685 23035
rect 24685 23001 24719 23035
rect 24719 23001 24728 23035
rect 24676 22992 24728 23001
rect 25320 22992 25372 23044
rect 26424 22992 26476 23044
rect 25136 22924 25188 22976
rect 30840 22992 30892 23044
rect 37280 23103 37332 23112
rect 37280 23069 37289 23103
rect 37289 23069 37323 23103
rect 37323 23069 37332 23103
rect 37280 23060 37332 23069
rect 40592 23171 40644 23180
rect 40592 23137 40601 23171
rect 40601 23137 40635 23171
rect 40635 23137 40644 23171
rect 40592 23128 40644 23137
rect 31576 22992 31628 23044
rect 28356 22967 28408 22976
rect 28356 22933 28365 22967
rect 28365 22933 28399 22967
rect 28399 22933 28408 22967
rect 28356 22924 28408 22933
rect 30104 22967 30156 22976
rect 30104 22933 30113 22967
rect 30113 22933 30147 22967
rect 30147 22933 30156 22967
rect 30104 22924 30156 22933
rect 30748 22924 30800 22976
rect 31208 22924 31260 22976
rect 32128 22992 32180 23044
rect 35348 23035 35400 23044
rect 35348 23001 35357 23035
rect 35357 23001 35391 23035
rect 35391 23001 35400 23035
rect 35348 22992 35400 23001
rect 35808 22992 35860 23044
rect 36728 22992 36780 23044
rect 37188 22992 37240 23044
rect 38844 22992 38896 23044
rect 39580 22992 39632 23044
rect 40316 22992 40368 23044
rect 42156 22992 42208 23044
rect 43352 22992 43404 23044
rect 43628 23035 43680 23044
rect 43628 23001 43637 23035
rect 43637 23001 43671 23035
rect 43671 23001 43680 23035
rect 43628 22992 43680 23001
rect 31760 22924 31812 22976
rect 33048 22924 33100 22976
rect 33324 22924 33376 22976
rect 35072 22924 35124 22976
rect 35164 22924 35216 22976
rect 38568 22924 38620 22976
rect 40224 22924 40276 22976
rect 41420 22924 41472 22976
rect 41604 22924 41656 22976
rect 42616 22924 42668 22976
rect 42800 22924 42852 22976
rect 43996 23103 44048 23112
rect 43996 23069 44005 23103
rect 44005 23069 44039 23103
rect 44039 23069 44048 23103
rect 43996 23060 44048 23069
rect 44088 23060 44140 23112
rect 43812 22992 43864 23044
rect 46296 23103 46348 23112
rect 46296 23069 46305 23103
rect 46305 23069 46339 23103
rect 46339 23069 46348 23103
rect 46296 23060 46348 23069
rect 49240 23128 49292 23180
rect 47860 23103 47912 23112
rect 47860 23069 47869 23103
rect 47869 23069 47903 23103
rect 47903 23069 47912 23103
rect 47860 23060 47912 23069
rect 48320 23103 48372 23112
rect 48320 23069 48329 23103
rect 48329 23069 48363 23103
rect 48363 23069 48372 23103
rect 48320 23060 48372 23069
rect 49148 23060 49200 23112
rect 46848 22992 46900 23044
rect 45192 22967 45244 22976
rect 45192 22933 45201 22967
rect 45201 22933 45235 22967
rect 45235 22933 45244 22967
rect 45192 22924 45244 22933
rect 45376 22967 45428 22976
rect 45376 22933 45385 22967
rect 45385 22933 45419 22967
rect 45419 22933 45428 22967
rect 45376 22924 45428 22933
rect 45468 22924 45520 22976
rect 47676 22967 47728 22976
rect 47676 22933 47685 22967
rect 47685 22933 47719 22967
rect 47719 22933 47728 22967
rect 47676 22924 47728 22933
rect 48504 22967 48556 22976
rect 48504 22933 48513 22967
rect 48513 22933 48547 22967
rect 48547 22933 48556 22967
rect 48504 22924 48556 22933
rect 7950 22822 8002 22874
rect 8014 22822 8066 22874
rect 8078 22822 8130 22874
rect 8142 22822 8194 22874
rect 8206 22822 8258 22874
rect 17950 22822 18002 22874
rect 18014 22822 18066 22874
rect 18078 22822 18130 22874
rect 18142 22822 18194 22874
rect 18206 22822 18258 22874
rect 27950 22822 28002 22874
rect 28014 22822 28066 22874
rect 28078 22822 28130 22874
rect 28142 22822 28194 22874
rect 28206 22822 28258 22874
rect 37950 22822 38002 22874
rect 38014 22822 38066 22874
rect 38078 22822 38130 22874
rect 38142 22822 38194 22874
rect 38206 22822 38258 22874
rect 47950 22822 48002 22874
rect 48014 22822 48066 22874
rect 48078 22822 48130 22874
rect 48142 22822 48194 22874
rect 48206 22822 48258 22874
rect 3332 22720 3384 22772
rect 6736 22720 6788 22772
rect 2872 22652 2924 22704
rect 13360 22720 13412 22772
rect 4804 22627 4856 22636
rect 4804 22593 4813 22627
rect 4813 22593 4847 22627
rect 4847 22593 4856 22627
rect 4804 22584 4856 22593
rect 5080 22559 5132 22568
rect 5080 22525 5089 22559
rect 5089 22525 5123 22559
rect 5123 22525 5132 22559
rect 5080 22516 5132 22525
rect 7564 22652 7616 22704
rect 7472 22627 7524 22636
rect 7472 22593 7481 22627
rect 7481 22593 7515 22627
rect 7515 22593 7524 22627
rect 7472 22584 7524 22593
rect 7380 22516 7432 22568
rect 10048 22516 10100 22568
rect 6460 22380 6512 22432
rect 9128 22380 9180 22432
rect 12808 22627 12860 22636
rect 12808 22593 12817 22627
rect 12817 22593 12851 22627
rect 12851 22593 12860 22627
rect 12808 22584 12860 22593
rect 17408 22720 17460 22772
rect 20628 22720 20680 22772
rect 22652 22720 22704 22772
rect 24768 22720 24820 22772
rect 24860 22720 24912 22772
rect 17040 22652 17092 22704
rect 18696 22652 18748 22704
rect 18880 22652 18932 22704
rect 20168 22652 20220 22704
rect 22284 22695 22336 22704
rect 22284 22661 22293 22695
rect 22293 22661 22327 22695
rect 22327 22661 22336 22695
rect 22284 22652 22336 22661
rect 22744 22652 22796 22704
rect 25044 22652 25096 22704
rect 25136 22695 25188 22704
rect 25136 22661 25145 22695
rect 25145 22661 25179 22695
rect 25179 22661 25188 22695
rect 25136 22652 25188 22661
rect 26424 22652 26476 22704
rect 27436 22652 27488 22704
rect 27620 22652 27672 22704
rect 27896 22652 27948 22704
rect 12532 22516 12584 22568
rect 15016 22516 15068 22568
rect 17132 22559 17184 22568
rect 17132 22525 17141 22559
rect 17141 22525 17175 22559
rect 17175 22525 17184 22559
rect 17132 22516 17184 22525
rect 18604 22516 18656 22568
rect 22008 22559 22060 22568
rect 22008 22525 22017 22559
rect 22017 22525 22051 22559
rect 22051 22525 22060 22559
rect 22008 22516 22060 22525
rect 14740 22448 14792 22500
rect 15660 22380 15712 22432
rect 17500 22380 17552 22432
rect 24860 22627 24912 22636
rect 24860 22593 24869 22627
rect 24869 22593 24903 22627
rect 24903 22593 24912 22627
rect 24860 22584 24912 22593
rect 27344 22627 27396 22636
rect 27344 22593 27353 22627
rect 27353 22593 27387 22627
rect 27387 22593 27396 22627
rect 27344 22584 27396 22593
rect 30012 22720 30064 22772
rect 30748 22652 30800 22704
rect 32496 22720 32548 22772
rect 32588 22652 32640 22704
rect 33324 22652 33376 22704
rect 33692 22652 33744 22704
rect 36360 22720 36412 22772
rect 37188 22720 37240 22772
rect 37740 22652 37792 22704
rect 23664 22516 23716 22568
rect 27620 22516 27672 22568
rect 29000 22516 29052 22568
rect 30748 22559 30800 22568
rect 30748 22525 30757 22559
rect 30757 22525 30791 22559
rect 30791 22525 30800 22559
rect 30748 22516 30800 22525
rect 30840 22559 30892 22568
rect 30840 22525 30849 22559
rect 30849 22525 30883 22559
rect 30883 22525 30892 22559
rect 30840 22516 30892 22525
rect 31668 22627 31720 22636
rect 31668 22593 31677 22627
rect 31677 22593 31711 22627
rect 31711 22593 31720 22627
rect 31668 22584 31720 22593
rect 26148 22448 26200 22500
rect 26976 22448 27028 22500
rect 27160 22491 27212 22500
rect 27160 22457 27169 22491
rect 27169 22457 27203 22491
rect 27203 22457 27212 22491
rect 27160 22448 27212 22457
rect 30380 22448 30432 22500
rect 23664 22380 23716 22432
rect 26608 22423 26660 22432
rect 26608 22389 26617 22423
rect 26617 22389 26651 22423
rect 26651 22389 26660 22423
rect 26608 22380 26660 22389
rect 28908 22380 28960 22432
rect 30288 22423 30340 22432
rect 30288 22389 30297 22423
rect 30297 22389 30331 22423
rect 30331 22389 30340 22423
rect 30288 22380 30340 22389
rect 31484 22423 31536 22432
rect 31484 22389 31493 22423
rect 31493 22389 31527 22423
rect 31527 22389 31536 22423
rect 31484 22380 31536 22389
rect 33140 22627 33192 22636
rect 33140 22593 33149 22627
rect 33149 22593 33183 22627
rect 33183 22593 33192 22627
rect 33140 22584 33192 22593
rect 36084 22584 36136 22636
rect 38844 22584 38896 22636
rect 33048 22516 33100 22568
rect 33876 22516 33928 22568
rect 35256 22516 35308 22568
rect 36176 22516 36228 22568
rect 36452 22559 36504 22568
rect 36452 22525 36461 22559
rect 36461 22525 36495 22559
rect 36495 22525 36504 22559
rect 36452 22516 36504 22525
rect 37280 22516 37332 22568
rect 37740 22559 37792 22568
rect 37740 22525 37749 22559
rect 37749 22525 37783 22559
rect 37783 22525 37792 22559
rect 37740 22516 37792 22525
rect 39672 22763 39724 22772
rect 39672 22729 39681 22763
rect 39681 22729 39715 22763
rect 39715 22729 39724 22763
rect 39672 22720 39724 22729
rect 40132 22763 40184 22772
rect 40132 22729 40141 22763
rect 40141 22729 40175 22763
rect 40175 22729 40184 22763
rect 40132 22720 40184 22729
rect 48688 22720 48740 22772
rect 40316 22652 40368 22704
rect 40040 22627 40092 22636
rect 40040 22593 40049 22627
rect 40049 22593 40083 22627
rect 40083 22593 40092 22627
rect 40040 22584 40092 22593
rect 41512 22627 41564 22636
rect 41512 22593 41521 22627
rect 41521 22593 41555 22627
rect 41555 22593 41564 22627
rect 41512 22584 41564 22593
rect 41788 22627 41840 22636
rect 41788 22593 41797 22627
rect 41797 22593 41831 22627
rect 41831 22593 41840 22627
rect 41788 22584 41840 22593
rect 41880 22584 41932 22636
rect 43444 22584 43496 22636
rect 46756 22584 46808 22636
rect 48412 22584 48464 22636
rect 49056 22627 49108 22636
rect 49056 22593 49065 22627
rect 49065 22593 49099 22627
rect 49099 22593 49108 22627
rect 49056 22584 49108 22593
rect 40960 22559 41012 22568
rect 40960 22525 40969 22559
rect 40969 22525 41003 22559
rect 41003 22525 41012 22559
rect 40960 22516 41012 22525
rect 41052 22559 41104 22568
rect 41052 22525 41061 22559
rect 41061 22525 41095 22559
rect 41095 22525 41104 22559
rect 41052 22516 41104 22525
rect 43536 22559 43588 22568
rect 43536 22525 43545 22559
rect 43545 22525 43579 22559
rect 43579 22525 43588 22559
rect 43536 22516 43588 22525
rect 35256 22380 35308 22432
rect 37004 22380 37056 22432
rect 39028 22448 39080 22500
rect 39120 22448 39172 22500
rect 47308 22448 47360 22500
rect 41328 22423 41380 22432
rect 41328 22389 41337 22423
rect 41337 22389 41371 22423
rect 41371 22389 41380 22423
rect 41328 22380 41380 22389
rect 41604 22423 41656 22432
rect 41604 22389 41613 22423
rect 41613 22389 41647 22423
rect 41647 22389 41656 22423
rect 41604 22380 41656 22389
rect 41696 22380 41748 22432
rect 44732 22423 44784 22432
rect 44732 22389 44741 22423
rect 44741 22389 44775 22423
rect 44775 22389 44784 22423
rect 44732 22380 44784 22389
rect 2950 22278 3002 22330
rect 3014 22278 3066 22330
rect 3078 22278 3130 22330
rect 3142 22278 3194 22330
rect 3206 22278 3258 22330
rect 12950 22278 13002 22330
rect 13014 22278 13066 22330
rect 13078 22278 13130 22330
rect 13142 22278 13194 22330
rect 13206 22278 13258 22330
rect 22950 22278 23002 22330
rect 23014 22278 23066 22330
rect 23078 22278 23130 22330
rect 23142 22278 23194 22330
rect 23206 22278 23258 22330
rect 32950 22278 33002 22330
rect 33014 22278 33066 22330
rect 33078 22278 33130 22330
rect 33142 22278 33194 22330
rect 33206 22278 33258 22330
rect 42950 22278 43002 22330
rect 43014 22278 43066 22330
rect 43078 22278 43130 22330
rect 43142 22278 43194 22330
rect 43206 22278 43258 22330
rect 2228 22176 2280 22228
rect 4896 22176 4948 22228
rect 7104 22176 7156 22228
rect 17132 22176 17184 22228
rect 17408 22176 17460 22228
rect 20996 22176 21048 22228
rect 22376 22176 22428 22228
rect 23204 22176 23256 22228
rect 3424 22108 3476 22160
rect 1308 22040 1360 22092
rect 3792 22040 3844 22092
rect 10508 22108 10560 22160
rect 13728 22108 13780 22160
rect 17224 22108 17276 22160
rect 9220 22040 9272 22092
rect 13820 22040 13872 22092
rect 18972 22108 19024 22160
rect 21732 22108 21784 22160
rect 4068 22015 4120 22024
rect 4068 21981 4077 22015
rect 4077 21981 4111 22015
rect 4111 21981 4120 22015
rect 4068 21972 4120 21981
rect 6000 22015 6052 22024
rect 6000 21981 6009 22015
rect 6009 21981 6043 22015
rect 6043 21981 6052 22015
rect 6000 21972 6052 21981
rect 7748 22015 7800 22024
rect 7748 21981 7757 22015
rect 7757 21981 7791 22015
rect 7791 21981 7800 22015
rect 7748 21972 7800 21981
rect 9128 22015 9180 22024
rect 9128 21981 9137 22015
rect 9137 21981 9171 22015
rect 9171 21981 9180 22015
rect 9128 21972 9180 21981
rect 11980 21972 12032 22024
rect 12072 22015 12124 22024
rect 12072 21981 12081 22015
rect 12081 21981 12115 22015
rect 12115 21981 12124 22015
rect 12072 21972 12124 21981
rect 12440 21972 12492 22024
rect 14004 21972 14056 22024
rect 4712 21836 4764 21888
rect 12808 21904 12860 21956
rect 14924 21904 14976 21956
rect 21272 21972 21324 22024
rect 23204 22083 23256 22092
rect 23204 22049 23213 22083
rect 23213 22049 23247 22083
rect 23247 22049 23256 22083
rect 23204 22040 23256 22049
rect 23388 22108 23440 22160
rect 25504 22108 25556 22160
rect 27804 22176 27856 22228
rect 29276 22176 29328 22228
rect 31300 22176 31352 22228
rect 32220 22176 32272 22228
rect 35808 22176 35860 22228
rect 38844 22176 38896 22228
rect 40040 22176 40092 22228
rect 42156 22176 42208 22228
rect 24584 22040 24636 22092
rect 24768 22040 24820 22092
rect 26148 22040 26200 22092
rect 26424 22083 26476 22092
rect 26424 22049 26433 22083
rect 26433 22049 26467 22083
rect 26467 22049 26476 22083
rect 26424 22040 26476 22049
rect 26608 22108 26660 22160
rect 27068 22040 27120 22092
rect 27896 22040 27948 22092
rect 28908 22040 28960 22092
rect 29552 22040 29604 22092
rect 30472 22040 30524 22092
rect 31576 22040 31628 22092
rect 32404 22040 32456 22092
rect 33876 22108 33928 22160
rect 38568 22108 38620 22160
rect 35900 22083 35952 22092
rect 35900 22049 35909 22083
rect 35909 22049 35943 22083
rect 35943 22049 35952 22083
rect 35900 22040 35952 22049
rect 37556 22083 37608 22092
rect 37556 22049 37565 22083
rect 37565 22049 37599 22083
rect 37599 22049 37608 22083
rect 37556 22040 37608 22049
rect 37648 22040 37700 22092
rect 40776 22108 40828 22160
rect 23940 21972 23992 22024
rect 11428 21836 11480 21888
rect 11612 21879 11664 21888
rect 11612 21845 11621 21879
rect 11621 21845 11655 21879
rect 11655 21845 11664 21879
rect 11612 21836 11664 21845
rect 12440 21836 12492 21888
rect 12624 21836 12676 21888
rect 16304 21836 16356 21888
rect 16488 21836 16540 21888
rect 20444 21904 20496 21956
rect 22284 21904 22336 21956
rect 25228 21904 25280 21956
rect 18696 21836 18748 21888
rect 19248 21836 19300 21888
rect 21548 21836 21600 21888
rect 22836 21836 22888 21888
rect 23112 21879 23164 21888
rect 23112 21845 23121 21879
rect 23121 21845 23155 21879
rect 23155 21845 23164 21879
rect 23112 21836 23164 21845
rect 23480 21836 23532 21888
rect 24952 21879 25004 21888
rect 24952 21845 24961 21879
rect 24961 21845 24995 21879
rect 24995 21845 25004 21879
rect 24952 21836 25004 21845
rect 25136 21836 25188 21888
rect 25872 21879 25924 21888
rect 25872 21845 25881 21879
rect 25881 21845 25915 21879
rect 25915 21845 25924 21879
rect 25872 21836 25924 21845
rect 27712 21972 27764 22024
rect 29828 21972 29880 22024
rect 30380 21904 30432 21956
rect 26240 21836 26292 21888
rect 26516 21836 26568 21888
rect 26608 21836 26660 21888
rect 27160 21836 27212 21888
rect 27436 21836 27488 21888
rect 28540 21836 28592 21888
rect 29552 21836 29604 21888
rect 34152 21972 34204 22024
rect 37280 22015 37332 22024
rect 37280 21981 37289 22015
rect 37289 21981 37323 22015
rect 37323 21981 37332 22015
rect 37280 21972 37332 21981
rect 38844 21972 38896 22024
rect 39028 21972 39080 22024
rect 31116 21947 31168 21956
rect 31116 21913 31125 21947
rect 31125 21913 31159 21947
rect 31159 21913 31168 21947
rect 31116 21904 31168 21913
rect 31208 21904 31260 21956
rect 31300 21836 31352 21888
rect 31392 21836 31444 21888
rect 42616 22040 42668 22092
rect 45468 22040 45520 22092
rect 46756 21972 46808 22024
rect 48596 22015 48648 22024
rect 48596 21981 48605 22015
rect 48605 21981 48639 22015
rect 48639 21981 48648 22015
rect 48596 21972 48648 21981
rect 32680 21836 32732 21888
rect 33416 21879 33468 21888
rect 33416 21845 33425 21879
rect 33425 21845 33459 21879
rect 33459 21845 33468 21879
rect 33416 21836 33468 21845
rect 34796 21836 34848 21888
rect 35808 21879 35860 21888
rect 35808 21845 35817 21879
rect 35817 21845 35851 21879
rect 35851 21845 35860 21879
rect 35808 21836 35860 21845
rect 36544 21879 36596 21888
rect 36544 21845 36553 21879
rect 36553 21845 36587 21879
rect 36587 21845 36596 21879
rect 36544 21836 36596 21845
rect 39120 21836 39172 21888
rect 39764 21836 39816 21888
rect 41512 21904 41564 21956
rect 47676 21904 47728 21956
rect 49148 21947 49200 21956
rect 49148 21913 49157 21947
rect 49157 21913 49191 21947
rect 49191 21913 49200 21947
rect 49148 21904 49200 21913
rect 40592 21836 40644 21888
rect 40960 21836 41012 21888
rect 41144 21836 41196 21888
rect 43260 21879 43312 21888
rect 43260 21845 43269 21879
rect 43269 21845 43303 21879
rect 43303 21845 43312 21879
rect 43260 21836 43312 21845
rect 48412 21879 48464 21888
rect 48412 21845 48421 21879
rect 48421 21845 48455 21879
rect 48455 21845 48464 21879
rect 48412 21836 48464 21845
rect 48688 21836 48740 21888
rect 7950 21734 8002 21786
rect 8014 21734 8066 21786
rect 8078 21734 8130 21786
rect 8142 21734 8194 21786
rect 8206 21734 8258 21786
rect 17950 21734 18002 21786
rect 18014 21734 18066 21786
rect 18078 21734 18130 21786
rect 18142 21734 18194 21786
rect 18206 21734 18258 21786
rect 27950 21734 28002 21786
rect 28014 21734 28066 21786
rect 28078 21734 28130 21786
rect 28142 21734 28194 21786
rect 28206 21734 28258 21786
rect 37950 21734 38002 21786
rect 38014 21734 38066 21786
rect 38078 21734 38130 21786
rect 38142 21734 38194 21786
rect 38206 21734 38258 21786
rect 47950 21734 48002 21786
rect 48014 21734 48066 21786
rect 48078 21734 48130 21786
rect 48142 21734 48194 21786
rect 48206 21734 48258 21786
rect 4068 21632 4120 21684
rect 9680 21632 9732 21684
rect 10324 21675 10376 21684
rect 10324 21641 10333 21675
rect 10333 21641 10367 21675
rect 10367 21641 10376 21675
rect 10324 21632 10376 21641
rect 10692 21632 10744 21684
rect 5632 21564 5684 21616
rect 3608 21539 3660 21548
rect 3608 21505 3617 21539
rect 3617 21505 3651 21539
rect 3651 21505 3660 21539
rect 3608 21496 3660 21505
rect 10416 21564 10468 21616
rect 6552 21539 6604 21548
rect 6552 21505 6561 21539
rect 6561 21505 6595 21539
rect 6595 21505 6604 21539
rect 6552 21496 6604 21505
rect 12164 21564 12216 21616
rect 13728 21632 13780 21684
rect 12348 21564 12400 21616
rect 13452 21564 13504 21616
rect 3332 21428 3384 21480
rect 4160 21471 4212 21480
rect 4160 21437 4169 21471
rect 4169 21437 4203 21471
rect 4203 21437 4212 21471
rect 4160 21428 4212 21437
rect 5540 21428 5592 21480
rect 8852 21471 8904 21480
rect 8852 21437 8861 21471
rect 8861 21437 8895 21471
rect 8895 21437 8904 21471
rect 8852 21428 8904 21437
rect 9864 21428 9916 21480
rect 11612 21428 11664 21480
rect 12624 21496 12676 21548
rect 17132 21632 17184 21684
rect 17408 21675 17460 21684
rect 17408 21641 17417 21675
rect 17417 21641 17451 21675
rect 17451 21641 17460 21675
rect 17408 21632 17460 21641
rect 17776 21632 17828 21684
rect 14832 21607 14884 21616
rect 14832 21573 14841 21607
rect 14841 21573 14875 21607
rect 14875 21573 14884 21607
rect 14832 21564 14884 21573
rect 16120 21564 16172 21616
rect 16488 21564 16540 21616
rect 12532 21428 12584 21480
rect 17776 21539 17828 21548
rect 17776 21505 17785 21539
rect 17785 21505 17819 21539
rect 17819 21505 17828 21539
rect 17776 21496 17828 21505
rect 11244 21360 11296 21412
rect 13728 21428 13780 21480
rect 14556 21471 14608 21480
rect 14556 21437 14565 21471
rect 14565 21437 14599 21471
rect 14599 21437 14608 21471
rect 14556 21428 14608 21437
rect 16396 21428 16448 21480
rect 20536 21632 20588 21684
rect 20996 21675 21048 21684
rect 20996 21641 21005 21675
rect 21005 21641 21039 21675
rect 21039 21641 21048 21675
rect 20996 21632 21048 21641
rect 22560 21632 22612 21684
rect 23112 21632 23164 21684
rect 24768 21675 24820 21684
rect 24768 21641 24777 21675
rect 24777 21641 24811 21675
rect 24811 21641 24820 21675
rect 24768 21632 24820 21641
rect 27252 21632 27304 21684
rect 27712 21632 27764 21684
rect 27804 21632 27856 21684
rect 28448 21632 28500 21684
rect 31116 21632 31168 21684
rect 18788 21564 18840 21616
rect 20352 21564 20404 21616
rect 22284 21564 22336 21616
rect 22744 21564 22796 21616
rect 21640 21496 21692 21548
rect 27436 21564 27488 21616
rect 29092 21564 29144 21616
rect 32496 21564 32548 21616
rect 18604 21471 18656 21480
rect 18604 21437 18613 21471
rect 18613 21437 18647 21471
rect 18647 21437 18656 21471
rect 18604 21428 18656 21437
rect 20720 21428 20772 21480
rect 22008 21428 22060 21480
rect 17040 21360 17092 21412
rect 23388 21428 23440 21480
rect 25136 21539 25188 21548
rect 25136 21505 25145 21539
rect 25145 21505 25179 21539
rect 25179 21505 25188 21539
rect 25136 21496 25188 21505
rect 24216 21471 24268 21480
rect 24216 21437 24225 21471
rect 24225 21437 24259 21471
rect 24259 21437 24268 21471
rect 24216 21428 24268 21437
rect 25412 21471 25464 21480
rect 25412 21437 25421 21471
rect 25421 21437 25455 21471
rect 25455 21437 25464 21471
rect 25412 21428 25464 21437
rect 4068 21292 4120 21344
rect 13544 21292 13596 21344
rect 15476 21292 15528 21344
rect 16304 21335 16356 21344
rect 16304 21301 16313 21335
rect 16313 21301 16347 21335
rect 16347 21301 16356 21335
rect 16304 21292 16356 21301
rect 19064 21292 19116 21344
rect 23756 21360 23808 21412
rect 27896 21496 27948 21548
rect 28264 21428 28316 21480
rect 28908 21471 28960 21480
rect 28908 21437 28917 21471
rect 28917 21437 28951 21471
rect 28951 21437 28960 21471
rect 28908 21428 28960 21437
rect 29736 21360 29788 21412
rect 30472 21496 30524 21548
rect 31024 21496 31076 21548
rect 33416 21564 33468 21616
rect 33692 21564 33744 21616
rect 33876 21564 33928 21616
rect 34888 21675 34940 21684
rect 34888 21641 34897 21675
rect 34897 21641 34931 21675
rect 34931 21641 34940 21675
rect 34888 21632 34940 21641
rect 37740 21632 37792 21684
rect 40132 21632 40184 21684
rect 40592 21632 40644 21684
rect 46848 21632 46900 21684
rect 36268 21564 36320 21616
rect 39028 21564 39080 21616
rect 39488 21564 39540 21616
rect 41144 21564 41196 21616
rect 41328 21564 41380 21616
rect 47124 21564 47176 21616
rect 34704 21496 34756 21548
rect 37096 21496 37148 21548
rect 37280 21496 37332 21548
rect 39672 21496 39724 21548
rect 46940 21496 46992 21548
rect 49056 21539 49108 21548
rect 49056 21505 49065 21539
rect 49065 21505 49099 21539
rect 49099 21505 49108 21539
rect 49056 21496 49108 21505
rect 30012 21428 30064 21480
rect 31208 21471 31260 21480
rect 31208 21437 31217 21471
rect 31217 21437 31251 21471
rect 31251 21437 31260 21471
rect 31208 21428 31260 21437
rect 31484 21428 31536 21480
rect 31576 21428 31628 21480
rect 33416 21471 33468 21480
rect 33416 21437 33425 21471
rect 33425 21437 33459 21471
rect 33459 21437 33468 21471
rect 33416 21428 33468 21437
rect 36176 21471 36228 21480
rect 36176 21437 36185 21471
rect 36185 21437 36219 21471
rect 36219 21437 36228 21471
rect 36176 21428 36228 21437
rect 36912 21428 36964 21480
rect 32680 21360 32732 21412
rect 32864 21360 32916 21412
rect 20260 21292 20312 21344
rect 21916 21292 21968 21344
rect 26148 21292 26200 21344
rect 26240 21292 26292 21344
rect 28632 21292 28684 21344
rect 28908 21292 28960 21344
rect 29092 21292 29144 21344
rect 29276 21292 29328 21344
rect 29552 21335 29604 21344
rect 29552 21301 29561 21335
rect 29561 21301 29595 21335
rect 29595 21301 29604 21335
rect 29552 21292 29604 21301
rect 30380 21292 30432 21344
rect 30840 21292 30892 21344
rect 36544 21360 36596 21412
rect 39120 21428 39172 21480
rect 40408 21428 40460 21480
rect 40684 21471 40736 21480
rect 40684 21437 40693 21471
rect 40693 21437 40727 21471
rect 40727 21437 40736 21471
rect 40684 21428 40736 21437
rect 40776 21471 40828 21480
rect 40776 21437 40785 21471
rect 40785 21437 40819 21471
rect 40819 21437 40828 21471
rect 40776 21428 40828 21437
rect 35624 21292 35676 21344
rect 36176 21292 36228 21344
rect 37924 21292 37976 21344
rect 43260 21360 43312 21412
rect 43628 21360 43680 21412
rect 48964 21360 49016 21412
rect 39212 21335 39264 21344
rect 39212 21301 39221 21335
rect 39221 21301 39255 21335
rect 39255 21301 39264 21335
rect 39212 21292 39264 21301
rect 39672 21335 39724 21344
rect 39672 21301 39681 21335
rect 39681 21301 39715 21335
rect 39715 21301 39724 21335
rect 39672 21292 39724 21301
rect 41604 21292 41656 21344
rect 2950 21190 3002 21242
rect 3014 21190 3066 21242
rect 3078 21190 3130 21242
rect 3142 21190 3194 21242
rect 3206 21190 3258 21242
rect 12950 21190 13002 21242
rect 13014 21190 13066 21242
rect 13078 21190 13130 21242
rect 13142 21190 13194 21242
rect 13206 21190 13258 21242
rect 22950 21190 23002 21242
rect 23014 21190 23066 21242
rect 23078 21190 23130 21242
rect 23142 21190 23194 21242
rect 23206 21190 23258 21242
rect 32950 21190 33002 21242
rect 33014 21190 33066 21242
rect 33078 21190 33130 21242
rect 33142 21190 33194 21242
rect 33206 21190 33258 21242
rect 42950 21190 43002 21242
rect 43014 21190 43066 21242
rect 43078 21190 43130 21242
rect 43142 21190 43194 21242
rect 43206 21190 43258 21242
rect 6000 21088 6052 21140
rect 4252 20952 4304 21004
rect 2780 20859 2832 20868
rect 2780 20825 2789 20859
rect 2789 20825 2823 20859
rect 2823 20825 2832 20859
rect 2780 20816 2832 20825
rect 4068 20927 4120 20936
rect 4068 20893 4077 20927
rect 4077 20893 4111 20927
rect 4111 20893 4120 20927
rect 4068 20884 4120 20893
rect 12624 21088 12676 21140
rect 12716 21088 12768 21140
rect 13636 21131 13688 21140
rect 13636 21097 13645 21131
rect 13645 21097 13679 21131
rect 13679 21097 13688 21131
rect 13636 21088 13688 21097
rect 6736 20995 6788 21004
rect 6736 20961 6745 20995
rect 6745 20961 6779 20995
rect 6779 20961 6788 20995
rect 6736 20952 6788 20961
rect 13636 20952 13688 21004
rect 10968 20884 11020 20936
rect 11152 20927 11204 20936
rect 11152 20893 11161 20927
rect 11161 20893 11195 20927
rect 11195 20893 11204 20927
rect 11152 20884 11204 20893
rect 15292 21088 15344 21140
rect 17776 21088 17828 21140
rect 13912 21020 13964 21072
rect 14188 21020 14240 21072
rect 18880 21131 18932 21140
rect 18880 21097 18889 21131
rect 18889 21097 18923 21131
rect 18923 21097 18932 21131
rect 18880 21088 18932 21097
rect 22376 21088 22428 21140
rect 14556 20952 14608 21004
rect 17040 20952 17092 21004
rect 20996 21020 21048 21072
rect 22468 21020 22520 21072
rect 22100 20952 22152 21004
rect 22376 20952 22428 21004
rect 22560 20952 22612 21004
rect 27804 21088 27856 21140
rect 27896 21131 27948 21140
rect 27896 21097 27905 21131
rect 27905 21097 27939 21131
rect 27939 21097 27948 21131
rect 27896 21088 27948 21097
rect 30104 21088 30156 21140
rect 30288 21088 30340 21140
rect 31208 21088 31260 21140
rect 33140 21088 33192 21140
rect 36268 21088 36320 21140
rect 37372 21088 37424 21140
rect 38752 21088 38804 21140
rect 40316 21088 40368 21140
rect 43628 21088 43680 21140
rect 48964 21088 49016 21140
rect 26148 21020 26200 21072
rect 14004 20884 14056 20936
rect 11520 20816 11572 20868
rect 7840 20748 7892 20800
rect 13544 20859 13596 20868
rect 13544 20825 13553 20859
rect 13553 20825 13587 20859
rect 13587 20825 13596 20859
rect 13544 20816 13596 20825
rect 13912 20816 13964 20868
rect 15844 20816 15896 20868
rect 16120 20816 16172 20868
rect 14648 20748 14700 20800
rect 14832 20748 14884 20800
rect 16488 20791 16540 20800
rect 16488 20757 16497 20791
rect 16497 20757 16531 20791
rect 16531 20757 16540 20791
rect 16488 20748 16540 20757
rect 19524 20884 19576 20936
rect 20720 20884 20772 20936
rect 18696 20816 18748 20868
rect 20812 20816 20864 20868
rect 21824 20816 21876 20868
rect 22008 20748 22060 20800
rect 22100 20748 22152 20800
rect 26332 20952 26384 21004
rect 27804 20952 27856 21004
rect 28448 20952 28500 21004
rect 29368 20952 29420 21004
rect 34796 21020 34848 21072
rect 33416 20952 33468 21004
rect 33692 20952 33744 21004
rect 34612 20952 34664 21004
rect 35164 20995 35216 21004
rect 35164 20961 35173 20995
rect 35173 20961 35207 20995
rect 35207 20961 35216 20995
rect 35164 20952 35216 20961
rect 35900 20952 35952 21004
rect 37280 20952 37332 21004
rect 37740 20995 37792 21004
rect 37740 20961 37749 20995
rect 37749 20961 37783 20995
rect 37783 20961 37792 20995
rect 37740 20952 37792 20961
rect 39212 20952 39264 21004
rect 40500 20995 40552 21004
rect 40500 20961 40509 20995
rect 40509 20961 40543 20995
rect 40543 20961 40552 20995
rect 40500 20952 40552 20961
rect 40592 20995 40644 21004
rect 40592 20961 40601 20995
rect 40601 20961 40635 20995
rect 40635 20961 40644 20995
rect 40592 20952 40644 20961
rect 24768 20884 24820 20936
rect 25044 20927 25096 20936
rect 25044 20893 25053 20927
rect 25053 20893 25087 20927
rect 25087 20893 25096 20927
rect 25044 20884 25096 20893
rect 25320 20884 25372 20936
rect 30288 20884 30340 20936
rect 32220 20927 32272 20936
rect 32220 20893 32229 20927
rect 32229 20893 32263 20927
rect 32263 20893 32272 20927
rect 32220 20884 32272 20893
rect 34704 20884 34756 20936
rect 39488 20884 39540 20936
rect 39764 20884 39816 20936
rect 23756 20859 23808 20868
rect 23756 20825 23765 20859
rect 23765 20825 23799 20859
rect 23799 20825 23808 20859
rect 23756 20816 23808 20825
rect 23296 20791 23348 20800
rect 23296 20757 23305 20791
rect 23305 20757 23339 20791
rect 23339 20757 23348 20791
rect 23296 20748 23348 20757
rect 29368 20816 29420 20868
rect 31484 20816 31536 20868
rect 33140 20816 33192 20868
rect 24952 20791 25004 20800
rect 24952 20757 24961 20791
rect 24961 20757 24995 20791
rect 24995 20757 25004 20791
rect 24952 20748 25004 20757
rect 25320 20748 25372 20800
rect 26240 20791 26292 20800
rect 26240 20757 26249 20791
rect 26249 20757 26283 20791
rect 26283 20757 26292 20791
rect 26240 20748 26292 20757
rect 26424 20748 26476 20800
rect 26884 20748 26936 20800
rect 27620 20748 27672 20800
rect 28632 20748 28684 20800
rect 28724 20791 28776 20800
rect 28724 20757 28733 20791
rect 28733 20757 28767 20791
rect 28767 20757 28776 20791
rect 28724 20748 28776 20757
rect 31208 20791 31260 20800
rect 31208 20757 31217 20791
rect 31217 20757 31251 20791
rect 31251 20757 31260 20791
rect 31208 20748 31260 20757
rect 32036 20791 32088 20800
rect 32036 20757 32045 20791
rect 32045 20757 32079 20791
rect 32079 20757 32088 20791
rect 32036 20748 32088 20757
rect 32496 20748 32548 20800
rect 32864 20748 32916 20800
rect 34428 20816 34480 20868
rect 37924 20816 37976 20868
rect 39948 20816 40000 20868
rect 49056 20927 49108 20936
rect 49056 20893 49065 20927
rect 49065 20893 49099 20927
rect 49099 20893 49108 20927
rect 49056 20884 49108 20893
rect 48412 20816 48464 20868
rect 38292 20748 38344 20800
rect 7950 20646 8002 20698
rect 8014 20646 8066 20698
rect 8078 20646 8130 20698
rect 8142 20646 8194 20698
rect 8206 20646 8258 20698
rect 17950 20646 18002 20698
rect 18014 20646 18066 20698
rect 18078 20646 18130 20698
rect 18142 20646 18194 20698
rect 18206 20646 18258 20698
rect 27950 20646 28002 20698
rect 28014 20646 28066 20698
rect 28078 20646 28130 20698
rect 28142 20646 28194 20698
rect 28206 20646 28258 20698
rect 37950 20646 38002 20698
rect 38014 20646 38066 20698
rect 38078 20646 38130 20698
rect 38142 20646 38194 20698
rect 38206 20646 38258 20698
rect 47950 20646 48002 20698
rect 48014 20646 48066 20698
rect 48078 20646 48130 20698
rect 48142 20646 48194 20698
rect 48206 20646 48258 20698
rect 6552 20544 6604 20596
rect 8300 20544 8352 20596
rect 9588 20544 9640 20596
rect 10416 20544 10468 20596
rect 10692 20544 10744 20596
rect 11336 20544 11388 20596
rect 1768 20451 1820 20460
rect 1768 20417 1777 20451
rect 1777 20417 1811 20451
rect 1811 20417 1820 20451
rect 1768 20408 1820 20417
rect 3608 20451 3660 20460
rect 3608 20417 3617 20451
rect 3617 20417 3651 20451
rect 3651 20417 3660 20451
rect 3608 20408 3660 20417
rect 6368 20408 6420 20460
rect 6460 20408 6512 20460
rect 2872 20340 2924 20392
rect 3884 20383 3936 20392
rect 3884 20349 3893 20383
rect 3893 20349 3927 20383
rect 3927 20349 3936 20383
rect 3884 20340 3936 20349
rect 5724 20340 5776 20392
rect 10048 20408 10100 20460
rect 11244 20476 11296 20528
rect 11428 20476 11480 20528
rect 13636 20544 13688 20596
rect 14372 20544 14424 20596
rect 9772 20340 9824 20392
rect 7656 20272 7708 20324
rect 11888 20408 11940 20460
rect 13636 20408 13688 20460
rect 9680 20204 9732 20256
rect 11980 20204 12032 20256
rect 14832 20340 14884 20392
rect 15384 20451 15436 20460
rect 15384 20417 15393 20451
rect 15393 20417 15427 20451
rect 15427 20417 15436 20451
rect 15384 20408 15436 20417
rect 15660 20476 15712 20528
rect 19156 20544 19208 20596
rect 18696 20476 18748 20528
rect 19432 20476 19484 20528
rect 16120 20451 16172 20460
rect 16120 20417 16129 20451
rect 16129 20417 16163 20451
rect 16163 20417 16172 20451
rect 16120 20408 16172 20417
rect 17040 20451 17092 20460
rect 17040 20417 17049 20451
rect 17049 20417 17083 20451
rect 17083 20417 17092 20451
rect 17040 20408 17092 20417
rect 16764 20340 16816 20392
rect 16856 20272 16908 20324
rect 19616 20340 19668 20392
rect 20628 20544 20680 20596
rect 20996 20544 21048 20596
rect 22100 20544 22152 20596
rect 21272 20476 21324 20528
rect 21824 20476 21876 20528
rect 25412 20544 25464 20596
rect 26608 20544 26660 20596
rect 27160 20544 27212 20596
rect 22560 20476 22612 20528
rect 23664 20476 23716 20528
rect 24124 20476 24176 20528
rect 27436 20476 27488 20528
rect 27712 20544 27764 20596
rect 28540 20544 28592 20596
rect 21364 20340 21416 20392
rect 23756 20408 23808 20460
rect 25504 20408 25556 20460
rect 29000 20587 29052 20596
rect 29000 20553 29009 20587
rect 29009 20553 29043 20587
rect 29043 20553 29052 20587
rect 29000 20544 29052 20553
rect 30840 20544 30892 20596
rect 31116 20587 31168 20596
rect 31116 20553 31125 20587
rect 31125 20553 31159 20587
rect 31159 20553 31168 20587
rect 31116 20544 31168 20553
rect 33416 20544 33468 20596
rect 35808 20544 35860 20596
rect 40408 20587 40460 20596
rect 40408 20553 40417 20587
rect 40417 20553 40451 20587
rect 40451 20553 40460 20587
rect 40408 20544 40460 20553
rect 32496 20476 32548 20528
rect 33876 20476 33928 20528
rect 34428 20476 34480 20528
rect 34612 20476 34664 20528
rect 35900 20476 35952 20528
rect 29644 20408 29696 20460
rect 29828 20408 29880 20460
rect 34520 20408 34572 20460
rect 22376 20272 22428 20324
rect 23388 20340 23440 20392
rect 24124 20383 24176 20392
rect 24124 20349 24133 20383
rect 24133 20349 24167 20383
rect 24167 20349 24176 20383
rect 24124 20340 24176 20349
rect 25596 20340 25648 20392
rect 26976 20340 27028 20392
rect 25228 20272 25280 20324
rect 26056 20315 26108 20324
rect 26056 20281 26065 20315
rect 26065 20281 26099 20315
rect 26099 20281 26108 20315
rect 26056 20272 26108 20281
rect 12716 20204 12768 20256
rect 18420 20204 18472 20256
rect 18788 20247 18840 20256
rect 18788 20213 18797 20247
rect 18797 20213 18831 20247
rect 18831 20213 18840 20247
rect 18788 20204 18840 20213
rect 18972 20204 19024 20256
rect 21732 20204 21784 20256
rect 21916 20204 21968 20256
rect 23664 20204 23716 20256
rect 25596 20247 25648 20256
rect 25596 20213 25605 20247
rect 25605 20213 25639 20247
rect 25639 20213 25648 20247
rect 25596 20204 25648 20213
rect 27896 20340 27948 20392
rect 29368 20340 29420 20392
rect 29920 20383 29972 20392
rect 29920 20349 29929 20383
rect 29929 20349 29963 20383
rect 29963 20349 29972 20383
rect 29920 20340 29972 20349
rect 30104 20383 30156 20392
rect 30104 20349 30113 20383
rect 30113 20349 30147 20383
rect 30147 20349 30156 20383
rect 30104 20340 30156 20349
rect 30196 20340 30248 20392
rect 31576 20340 31628 20392
rect 32588 20340 32640 20392
rect 33600 20340 33652 20392
rect 35348 20408 35400 20460
rect 37924 20476 37976 20528
rect 38292 20476 38344 20528
rect 39488 20476 39540 20528
rect 36084 20408 36136 20460
rect 37556 20408 37608 20460
rect 37740 20451 37792 20460
rect 37740 20417 37749 20451
rect 37749 20417 37783 20451
rect 37783 20417 37792 20451
rect 37740 20408 37792 20417
rect 40316 20451 40368 20460
rect 40316 20417 40325 20451
rect 40325 20417 40359 20451
rect 40359 20417 40368 20451
rect 40316 20408 40368 20417
rect 35164 20383 35216 20392
rect 35164 20349 35173 20383
rect 35173 20349 35207 20383
rect 35207 20349 35216 20383
rect 35164 20340 35216 20349
rect 37648 20340 37700 20392
rect 45376 20408 45428 20460
rect 48596 20451 48648 20460
rect 48596 20417 48605 20451
rect 48605 20417 48639 20451
rect 48639 20417 48648 20451
rect 48596 20408 48648 20417
rect 49056 20451 49108 20460
rect 49056 20417 49065 20451
rect 49065 20417 49099 20451
rect 49099 20417 49108 20451
rect 49056 20408 49108 20417
rect 30564 20204 30616 20256
rect 31116 20204 31168 20256
rect 31300 20204 31352 20256
rect 34060 20204 34112 20256
rect 40500 20383 40552 20392
rect 40500 20349 40509 20383
rect 40509 20349 40543 20383
rect 40543 20349 40552 20383
rect 40500 20340 40552 20349
rect 38660 20204 38712 20256
rect 40132 20272 40184 20324
rect 40408 20272 40460 20324
rect 40868 20204 40920 20256
rect 48412 20247 48464 20256
rect 48412 20213 48421 20247
rect 48421 20213 48455 20247
rect 48455 20213 48464 20247
rect 48412 20204 48464 20213
rect 2950 20102 3002 20154
rect 3014 20102 3066 20154
rect 3078 20102 3130 20154
rect 3142 20102 3194 20154
rect 3206 20102 3258 20154
rect 12950 20102 13002 20154
rect 13014 20102 13066 20154
rect 13078 20102 13130 20154
rect 13142 20102 13194 20154
rect 13206 20102 13258 20154
rect 22950 20102 23002 20154
rect 23014 20102 23066 20154
rect 23078 20102 23130 20154
rect 23142 20102 23194 20154
rect 23206 20102 23258 20154
rect 32950 20102 33002 20154
rect 33014 20102 33066 20154
rect 33078 20102 33130 20154
rect 33142 20102 33194 20154
rect 33206 20102 33258 20154
rect 42950 20102 43002 20154
rect 43014 20102 43066 20154
rect 43078 20102 43130 20154
rect 43142 20102 43194 20154
rect 43206 20102 43258 20154
rect 3608 19932 3660 19984
rect 13360 19932 13412 19984
rect 13544 19932 13596 19984
rect 14740 20043 14792 20052
rect 14740 20009 14749 20043
rect 14749 20009 14783 20043
rect 14783 20009 14792 20043
rect 14740 20000 14792 20009
rect 16396 20000 16448 20052
rect 17316 19932 17368 19984
rect 4896 19907 4948 19916
rect 4896 19873 4905 19907
rect 4905 19873 4939 19907
rect 4939 19873 4948 19907
rect 4896 19864 4948 19873
rect 6276 19907 6328 19916
rect 6276 19873 6285 19907
rect 6285 19873 6319 19907
rect 6319 19873 6328 19907
rect 6276 19864 6328 19873
rect 9312 19864 9364 19916
rect 16304 19864 16356 19916
rect 2780 19771 2832 19780
rect 2780 19737 2789 19771
rect 2789 19737 2823 19771
rect 2823 19737 2832 19771
rect 2780 19728 2832 19737
rect 9496 19796 9548 19848
rect 7288 19728 7340 19780
rect 11060 19839 11112 19848
rect 11060 19805 11069 19839
rect 11069 19805 11103 19839
rect 11103 19805 11112 19839
rect 11060 19796 11112 19805
rect 11336 19839 11388 19848
rect 11336 19805 11345 19839
rect 11345 19805 11379 19839
rect 11379 19805 11388 19839
rect 11336 19796 11388 19805
rect 11980 19839 12032 19848
rect 11980 19805 11989 19839
rect 11989 19805 12023 19839
rect 12023 19805 12032 19839
rect 11980 19796 12032 19805
rect 14280 19796 14332 19848
rect 14648 19796 14700 19848
rect 23296 20000 23348 20052
rect 24124 20000 24176 20052
rect 21824 19932 21876 19984
rect 22836 19932 22888 19984
rect 18880 19864 18932 19916
rect 12164 19728 12216 19780
rect 12256 19771 12308 19780
rect 12256 19737 12265 19771
rect 12265 19737 12299 19771
rect 12299 19737 12308 19771
rect 12256 19728 12308 19737
rect 12072 19660 12124 19712
rect 12624 19660 12676 19712
rect 13268 19660 13320 19712
rect 14740 19728 14792 19780
rect 13820 19660 13872 19712
rect 16672 19771 16724 19780
rect 16672 19737 16681 19771
rect 16681 19737 16715 19771
rect 16715 19737 16724 19771
rect 16672 19728 16724 19737
rect 16948 19728 17000 19780
rect 20536 19839 20588 19848
rect 20536 19805 20545 19839
rect 20545 19805 20579 19839
rect 20579 19805 20588 19839
rect 20536 19796 20588 19805
rect 25136 19864 25188 19916
rect 25596 19864 25648 19916
rect 30012 20000 30064 20052
rect 31392 20000 31444 20052
rect 34704 20000 34756 20052
rect 36728 20000 36780 20052
rect 37832 20000 37884 20052
rect 40132 20000 40184 20052
rect 27160 19932 27212 19984
rect 29000 19932 29052 19984
rect 33508 19932 33560 19984
rect 27528 19864 27580 19916
rect 27896 19907 27948 19916
rect 27896 19873 27905 19907
rect 27905 19873 27939 19907
rect 27939 19873 27948 19907
rect 27896 19864 27948 19873
rect 28540 19907 28592 19916
rect 28540 19873 28549 19907
rect 28549 19873 28583 19907
rect 28583 19873 28592 19907
rect 28540 19864 28592 19873
rect 28632 19907 28684 19916
rect 28632 19873 28641 19907
rect 28641 19873 28675 19907
rect 28675 19873 28684 19907
rect 28632 19864 28684 19873
rect 23848 19796 23900 19848
rect 29552 19864 29604 19916
rect 31760 19864 31812 19916
rect 32128 19907 32180 19916
rect 32128 19873 32137 19907
rect 32137 19873 32171 19907
rect 32171 19873 32180 19907
rect 32128 19864 32180 19873
rect 33416 19864 33468 19916
rect 35256 19864 35308 19916
rect 35440 19907 35492 19916
rect 35440 19873 35449 19907
rect 35449 19873 35483 19907
rect 35483 19873 35492 19907
rect 35440 19864 35492 19873
rect 37280 19864 37332 19916
rect 37924 19864 37976 19916
rect 38384 19864 38436 19916
rect 38568 19864 38620 19916
rect 40592 19907 40644 19916
rect 40592 19873 40601 19907
rect 40601 19873 40635 19907
rect 40635 19873 40644 19907
rect 40592 19864 40644 19873
rect 41604 19864 41656 19916
rect 41880 19864 41932 19916
rect 28816 19796 28868 19848
rect 30288 19796 30340 19848
rect 17224 19660 17276 19712
rect 17408 19703 17460 19712
rect 17408 19669 17417 19703
rect 17417 19669 17451 19703
rect 17451 19669 17460 19703
rect 17408 19660 17460 19669
rect 18328 19660 18380 19712
rect 18512 19703 18564 19712
rect 18512 19669 18521 19703
rect 18521 19669 18555 19703
rect 18555 19669 18564 19703
rect 18512 19660 18564 19669
rect 21272 19728 21324 19780
rect 21456 19660 21508 19712
rect 22744 19703 22796 19712
rect 22744 19669 22753 19703
rect 22753 19669 22787 19703
rect 22787 19669 22796 19703
rect 22744 19660 22796 19669
rect 22836 19660 22888 19712
rect 26792 19771 26844 19780
rect 26792 19737 26801 19771
rect 26801 19737 26835 19771
rect 26835 19737 26844 19771
rect 26792 19728 26844 19737
rect 27620 19771 27672 19780
rect 27620 19737 27629 19771
rect 27629 19737 27663 19771
rect 27663 19737 27672 19771
rect 27620 19728 27672 19737
rect 30932 19728 30984 19780
rect 32036 19796 32088 19848
rect 34060 19796 34112 19848
rect 37372 19796 37424 19848
rect 39120 19796 39172 19848
rect 26976 19660 27028 19712
rect 27252 19703 27304 19712
rect 27252 19669 27261 19703
rect 27261 19669 27295 19703
rect 27295 19669 27304 19703
rect 27252 19660 27304 19669
rect 28908 19660 28960 19712
rect 30656 19660 30708 19712
rect 30840 19703 30892 19712
rect 30840 19669 30849 19703
rect 30849 19669 30883 19703
rect 30883 19669 30892 19703
rect 30840 19660 30892 19669
rect 34060 19660 34112 19712
rect 35072 19728 35124 19780
rect 39948 19728 40000 19780
rect 48412 19728 48464 19780
rect 49332 19728 49384 19780
rect 35900 19660 35952 19712
rect 35992 19660 36044 19712
rect 36544 19703 36596 19712
rect 36544 19669 36553 19703
rect 36553 19669 36587 19703
rect 36587 19669 36596 19703
rect 36544 19660 36596 19669
rect 40960 19660 41012 19712
rect 41144 19660 41196 19712
rect 7950 19558 8002 19610
rect 8014 19558 8066 19610
rect 8078 19558 8130 19610
rect 8142 19558 8194 19610
rect 8206 19558 8258 19610
rect 17950 19558 18002 19610
rect 18014 19558 18066 19610
rect 18078 19558 18130 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 27950 19558 28002 19610
rect 28014 19558 28066 19610
rect 28078 19558 28130 19610
rect 28142 19558 28194 19610
rect 28206 19558 28258 19610
rect 37950 19558 38002 19610
rect 38014 19558 38066 19610
rect 38078 19558 38130 19610
rect 38142 19558 38194 19610
rect 38206 19558 38258 19610
rect 47950 19558 48002 19610
rect 48014 19558 48066 19610
rect 48078 19558 48130 19610
rect 48142 19558 48194 19610
rect 48206 19558 48258 19610
rect 9312 19456 9364 19508
rect 4344 19431 4396 19440
rect 4344 19397 4353 19431
rect 4353 19397 4387 19431
rect 4387 19397 4396 19431
rect 4344 19388 4396 19397
rect 2872 19320 2924 19372
rect 10876 19388 10928 19440
rect 5356 19363 5408 19372
rect 5356 19329 5365 19363
rect 5365 19329 5399 19363
rect 5399 19329 5408 19363
rect 5356 19320 5408 19329
rect 7564 19320 7616 19372
rect 11060 19456 11112 19508
rect 12624 19456 12676 19508
rect 13360 19456 13412 19508
rect 15292 19456 15344 19508
rect 16856 19499 16908 19508
rect 16856 19465 16865 19499
rect 16865 19465 16899 19499
rect 16899 19465 16908 19499
rect 16856 19456 16908 19465
rect 19248 19456 19300 19508
rect 20812 19456 20864 19508
rect 23940 19456 23992 19508
rect 25136 19499 25188 19508
rect 25136 19465 25145 19499
rect 25145 19465 25179 19499
rect 25179 19465 25188 19499
rect 25136 19456 25188 19465
rect 13268 19388 13320 19440
rect 14280 19388 14332 19440
rect 15752 19388 15804 19440
rect 17040 19388 17092 19440
rect 12072 19363 12124 19372
rect 12072 19329 12081 19363
rect 12081 19329 12115 19363
rect 12115 19329 12124 19363
rect 12072 19320 12124 19329
rect 15844 19320 15896 19372
rect 16488 19320 16540 19372
rect 17224 19363 17276 19372
rect 17224 19329 17233 19363
rect 17233 19329 17267 19363
rect 17267 19329 17276 19363
rect 17224 19320 17276 19329
rect 18604 19388 18656 19440
rect 19616 19388 19668 19440
rect 26608 19456 26660 19508
rect 27528 19456 27580 19508
rect 27988 19456 28040 19508
rect 28724 19456 28776 19508
rect 28816 19499 28868 19508
rect 28816 19465 28825 19499
rect 28825 19465 28859 19499
rect 28859 19465 28868 19499
rect 28816 19456 28868 19465
rect 29644 19499 29696 19508
rect 29644 19465 29653 19499
rect 29653 19465 29687 19499
rect 29687 19465 29696 19499
rect 29644 19456 29696 19465
rect 31760 19456 31812 19508
rect 32588 19456 32640 19508
rect 32680 19499 32732 19508
rect 32680 19465 32689 19499
rect 32689 19465 32723 19499
rect 32723 19465 32732 19499
rect 32680 19456 32732 19465
rect 32864 19456 32916 19508
rect 33508 19499 33560 19508
rect 33508 19465 33517 19499
rect 33517 19465 33551 19499
rect 33551 19465 33560 19499
rect 33508 19456 33560 19465
rect 34336 19456 34388 19508
rect 36544 19456 36596 19508
rect 40408 19456 40460 19508
rect 41052 19456 41104 19508
rect 19432 19320 19484 19372
rect 19892 19320 19944 19372
rect 20352 19320 20404 19372
rect 21548 19320 21600 19372
rect 26148 19431 26200 19440
rect 26148 19397 26157 19431
rect 26157 19397 26191 19431
rect 26191 19397 26200 19431
rect 26148 19388 26200 19397
rect 26240 19388 26292 19440
rect 27160 19388 27212 19440
rect 27712 19388 27764 19440
rect 29920 19388 29972 19440
rect 30196 19388 30248 19440
rect 30656 19388 30708 19440
rect 31300 19388 31352 19440
rect 31576 19431 31628 19440
rect 31576 19397 31585 19431
rect 31585 19397 31619 19431
rect 31619 19397 31628 19431
rect 31576 19388 31628 19397
rect 35256 19388 35308 19440
rect 9128 19252 9180 19304
rect 15936 19252 15988 19304
rect 11612 19184 11664 19236
rect 11980 19184 12032 19236
rect 2320 19116 2372 19168
rect 10416 19116 10468 19168
rect 11336 19116 11388 19168
rect 11520 19116 11572 19168
rect 12716 19184 12768 19236
rect 14004 19116 14056 19168
rect 16212 19159 16264 19168
rect 16212 19125 16221 19159
rect 16221 19125 16255 19159
rect 16255 19125 16264 19159
rect 16212 19116 16264 19125
rect 23388 19363 23440 19372
rect 23388 19329 23397 19363
rect 23397 19329 23431 19363
rect 23431 19329 23440 19363
rect 23388 19320 23440 19329
rect 25872 19320 25924 19372
rect 23296 19252 23348 19304
rect 23664 19295 23716 19304
rect 23664 19261 23673 19295
rect 23673 19261 23707 19295
rect 23707 19261 23716 19295
rect 23664 19252 23716 19261
rect 28632 19320 28684 19372
rect 22468 19184 22520 19236
rect 27804 19252 27856 19304
rect 30012 19363 30064 19372
rect 30012 19329 30021 19363
rect 30021 19329 30055 19363
rect 30055 19329 30064 19363
rect 30012 19320 30064 19329
rect 30840 19363 30892 19372
rect 30840 19329 30849 19363
rect 30849 19329 30883 19363
rect 30883 19329 30892 19363
rect 30840 19320 30892 19329
rect 30932 19320 30984 19372
rect 31944 19320 31996 19372
rect 32404 19320 32456 19372
rect 34612 19320 34664 19372
rect 35072 19363 35124 19372
rect 26884 19184 26936 19236
rect 27528 19184 27580 19236
rect 32128 19252 32180 19304
rect 32864 19295 32916 19304
rect 32864 19261 32873 19295
rect 32873 19261 32907 19295
rect 32907 19261 32916 19295
rect 32864 19252 32916 19261
rect 33968 19295 34020 19304
rect 33968 19261 33977 19295
rect 33977 19261 34011 19295
rect 34011 19261 34020 19295
rect 33968 19252 34020 19261
rect 34520 19252 34572 19304
rect 35072 19329 35081 19363
rect 35081 19329 35115 19363
rect 35115 19329 35124 19363
rect 35072 19320 35124 19329
rect 35164 19363 35216 19372
rect 35164 19329 35173 19363
rect 35173 19329 35207 19363
rect 35207 19329 35216 19363
rect 35164 19320 35216 19329
rect 36176 19388 36228 19440
rect 36636 19388 36688 19440
rect 39488 19388 39540 19440
rect 39948 19388 40000 19440
rect 41144 19388 41196 19440
rect 35900 19320 35952 19372
rect 37188 19320 37240 19372
rect 37740 19320 37792 19372
rect 49148 19363 49200 19372
rect 49148 19329 49157 19363
rect 49157 19329 49191 19363
rect 49191 19329 49200 19363
rect 49148 19320 49200 19329
rect 18788 19116 18840 19168
rect 21088 19116 21140 19168
rect 23480 19116 23532 19168
rect 25780 19159 25832 19168
rect 25780 19125 25789 19159
rect 25789 19125 25823 19159
rect 25823 19125 25832 19159
rect 25780 19116 25832 19125
rect 26516 19116 26568 19168
rect 33324 19116 33376 19168
rect 37832 19252 37884 19304
rect 36176 19184 36228 19236
rect 38660 19252 38712 19304
rect 39212 19252 39264 19304
rect 37004 19116 37056 19168
rect 40500 19184 40552 19236
rect 41788 19184 41840 19236
rect 39672 19159 39724 19168
rect 39672 19125 39681 19159
rect 39681 19125 39715 19159
rect 39715 19125 39724 19159
rect 39672 19116 39724 19125
rect 40132 19159 40184 19168
rect 40132 19125 40141 19159
rect 40141 19125 40175 19159
rect 40175 19125 40184 19159
rect 40132 19116 40184 19125
rect 47400 19116 47452 19168
rect 2950 19014 3002 19066
rect 3014 19014 3066 19066
rect 3078 19014 3130 19066
rect 3142 19014 3194 19066
rect 3206 19014 3258 19066
rect 12950 19014 13002 19066
rect 13014 19014 13066 19066
rect 13078 19014 13130 19066
rect 13142 19014 13194 19066
rect 13206 19014 13258 19066
rect 22950 19014 23002 19066
rect 23014 19014 23066 19066
rect 23078 19014 23130 19066
rect 23142 19014 23194 19066
rect 23206 19014 23258 19066
rect 32950 19014 33002 19066
rect 33014 19014 33066 19066
rect 33078 19014 33130 19066
rect 33142 19014 33194 19066
rect 33206 19014 33258 19066
rect 42950 19014 43002 19066
rect 43014 19014 43066 19066
rect 43078 19014 43130 19066
rect 43142 19014 43194 19066
rect 43206 19014 43258 19066
rect 2780 18683 2832 18692
rect 2780 18649 2789 18683
rect 2789 18649 2823 18683
rect 2823 18649 2832 18683
rect 2780 18640 2832 18649
rect 3700 18776 3752 18828
rect 9864 18912 9916 18964
rect 10876 18955 10928 18964
rect 10876 18921 10885 18955
rect 10885 18921 10919 18955
rect 10919 18921 10928 18955
rect 10876 18912 10928 18921
rect 10968 18912 11020 18964
rect 11980 18912 12032 18964
rect 9128 18819 9180 18828
rect 9128 18785 9137 18819
rect 9137 18785 9171 18819
rect 9171 18785 9180 18819
rect 9128 18776 9180 18785
rect 11060 18776 11112 18828
rect 7840 18708 7892 18760
rect 12164 18844 12216 18896
rect 13084 18776 13136 18828
rect 13360 18776 13412 18828
rect 13728 18776 13780 18828
rect 15200 18776 15252 18828
rect 15292 18776 15344 18828
rect 15752 18776 15804 18828
rect 8300 18615 8352 18624
rect 8300 18581 8309 18615
rect 8309 18581 8343 18615
rect 8343 18581 8352 18615
rect 8300 18572 8352 18581
rect 11244 18640 11296 18692
rect 11336 18640 11388 18692
rect 11520 18572 11572 18624
rect 12164 18572 12216 18624
rect 14832 18640 14884 18692
rect 15936 18912 15988 18964
rect 16580 18912 16632 18964
rect 17224 18912 17276 18964
rect 18512 18912 18564 18964
rect 21088 18844 21140 18896
rect 16028 18708 16080 18760
rect 17408 18776 17460 18828
rect 18972 18776 19024 18828
rect 20996 18776 21048 18828
rect 21824 18844 21876 18896
rect 24584 18955 24636 18964
rect 24584 18921 24593 18955
rect 24593 18921 24627 18955
rect 24627 18921 24636 18955
rect 24584 18912 24636 18921
rect 24676 18912 24728 18964
rect 29736 18912 29788 18964
rect 25320 18844 25372 18896
rect 22192 18776 22244 18828
rect 24492 18776 24544 18828
rect 25044 18819 25096 18828
rect 25044 18785 25053 18819
rect 25053 18785 25087 18819
rect 25087 18785 25096 18819
rect 25044 18776 25096 18785
rect 18144 18640 18196 18692
rect 22284 18751 22336 18760
rect 22284 18717 22293 18751
rect 22293 18717 22327 18751
rect 22327 18717 22336 18751
rect 22284 18708 22336 18717
rect 25688 18776 25740 18828
rect 27160 18844 27212 18896
rect 27528 18887 27580 18896
rect 27528 18853 27537 18887
rect 27537 18853 27571 18887
rect 27571 18853 27580 18887
rect 27528 18844 27580 18853
rect 32496 18912 32548 18964
rect 32772 18912 32824 18964
rect 32956 18912 33008 18964
rect 35992 18912 36044 18964
rect 37004 18955 37056 18964
rect 37004 18921 37013 18955
rect 37013 18921 37047 18955
rect 37047 18921 37056 18955
rect 37004 18912 37056 18921
rect 27068 18776 27120 18828
rect 30196 18819 30248 18828
rect 30196 18785 30205 18819
rect 30205 18785 30239 18819
rect 30239 18785 30248 18819
rect 30196 18776 30248 18785
rect 30288 18819 30340 18828
rect 30288 18785 30297 18819
rect 30297 18785 30331 18819
rect 30331 18785 30340 18819
rect 30288 18776 30340 18785
rect 19064 18640 19116 18692
rect 21272 18640 21324 18692
rect 23020 18640 23072 18692
rect 13084 18572 13136 18624
rect 15568 18572 15620 18624
rect 18328 18615 18380 18624
rect 18328 18581 18337 18615
rect 18337 18581 18371 18615
rect 18371 18581 18380 18615
rect 18328 18572 18380 18581
rect 19248 18572 19300 18624
rect 20444 18572 20496 18624
rect 20720 18572 20772 18624
rect 21548 18572 21600 18624
rect 23848 18572 23900 18624
rect 30472 18708 30524 18760
rect 25136 18640 25188 18692
rect 26608 18640 26660 18692
rect 29276 18640 29328 18692
rect 32956 18776 33008 18828
rect 33048 18776 33100 18828
rect 32496 18708 32548 18760
rect 34888 18776 34940 18828
rect 35256 18819 35308 18828
rect 35256 18785 35265 18819
rect 35265 18785 35299 18819
rect 35299 18785 35308 18819
rect 35256 18776 35308 18785
rect 41328 18912 41380 18964
rect 41788 18955 41840 18964
rect 41788 18921 41797 18955
rect 41797 18921 41831 18955
rect 41831 18921 41840 18955
rect 41788 18912 41840 18921
rect 40040 18844 40092 18896
rect 38292 18776 38344 18828
rect 39488 18776 39540 18828
rect 37464 18751 37516 18760
rect 37464 18717 37473 18751
rect 37473 18717 37507 18751
rect 37507 18717 37516 18751
rect 37464 18708 37516 18717
rect 38660 18708 38712 18760
rect 36544 18640 36596 18692
rect 37648 18640 37700 18692
rect 39856 18640 39908 18692
rect 48596 18751 48648 18760
rect 48596 18717 48605 18751
rect 48605 18717 48639 18751
rect 48639 18717 48648 18751
rect 48596 18708 48648 18717
rect 49148 18708 49200 18760
rect 24860 18572 24912 18624
rect 27620 18572 27672 18624
rect 29184 18572 29236 18624
rect 29828 18572 29880 18624
rect 31852 18615 31904 18624
rect 31852 18581 31861 18615
rect 31861 18581 31895 18615
rect 31895 18581 31904 18615
rect 31852 18572 31904 18581
rect 32496 18572 32548 18624
rect 33416 18572 33468 18624
rect 33692 18572 33744 18624
rect 35348 18572 35400 18624
rect 38384 18615 38436 18624
rect 38384 18581 38393 18615
rect 38393 18581 38427 18615
rect 38427 18581 38436 18615
rect 38384 18572 38436 18581
rect 47400 18572 47452 18624
rect 48412 18615 48464 18624
rect 48412 18581 48421 18615
rect 48421 18581 48455 18615
rect 48455 18581 48464 18615
rect 48412 18572 48464 18581
rect 49240 18615 49292 18624
rect 49240 18581 49249 18615
rect 49249 18581 49283 18615
rect 49283 18581 49292 18615
rect 49240 18572 49292 18581
rect 7950 18470 8002 18522
rect 8014 18470 8066 18522
rect 8078 18470 8130 18522
rect 8142 18470 8194 18522
rect 8206 18470 8258 18522
rect 17950 18470 18002 18522
rect 18014 18470 18066 18522
rect 18078 18470 18130 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 27950 18470 28002 18522
rect 28014 18470 28066 18522
rect 28078 18470 28130 18522
rect 28142 18470 28194 18522
rect 28206 18470 28258 18522
rect 37950 18470 38002 18522
rect 38014 18470 38066 18522
rect 38078 18470 38130 18522
rect 38142 18470 38194 18522
rect 38206 18470 38258 18522
rect 47950 18470 48002 18522
rect 48014 18470 48066 18522
rect 48078 18470 48130 18522
rect 48142 18470 48194 18522
rect 48206 18470 48258 18522
rect 5632 18368 5684 18420
rect 9772 18411 9824 18420
rect 9772 18377 9781 18411
rect 9781 18377 9815 18411
rect 9815 18377 9824 18411
rect 9772 18368 9824 18377
rect 10416 18368 10468 18420
rect 11152 18368 11204 18420
rect 11244 18368 11296 18420
rect 11980 18368 12032 18420
rect 3516 18232 3568 18284
rect 9864 18232 9916 18284
rect 2780 18207 2832 18216
rect 2780 18173 2789 18207
rect 2789 18173 2823 18207
rect 2823 18173 2832 18207
rect 2780 18164 2832 18173
rect 4160 18207 4212 18216
rect 4160 18173 4169 18207
rect 4169 18173 4203 18207
rect 4203 18173 4212 18207
rect 4160 18164 4212 18173
rect 12256 18300 12308 18352
rect 12624 18368 12676 18420
rect 14832 18368 14884 18420
rect 15384 18368 15436 18420
rect 15476 18411 15528 18420
rect 15476 18377 15485 18411
rect 15485 18377 15519 18411
rect 15519 18377 15528 18411
rect 15476 18368 15528 18377
rect 16120 18411 16172 18420
rect 16120 18377 16129 18411
rect 16129 18377 16163 18411
rect 16163 18377 16172 18411
rect 16120 18368 16172 18377
rect 16764 18368 16816 18420
rect 17316 18368 17368 18420
rect 18604 18368 18656 18420
rect 25780 18368 25832 18420
rect 27252 18368 27304 18420
rect 27620 18368 27672 18420
rect 29644 18368 29696 18420
rect 31208 18368 31260 18420
rect 36268 18411 36320 18420
rect 36268 18377 36277 18411
rect 36277 18377 36311 18411
rect 36311 18377 36320 18411
rect 36268 18368 36320 18377
rect 37556 18368 37608 18420
rect 13820 18300 13872 18352
rect 10048 18096 10100 18148
rect 11612 18164 11664 18216
rect 13360 18164 13412 18216
rect 13452 18164 13504 18216
rect 11428 18096 11480 18148
rect 15200 18164 15252 18216
rect 16028 18164 16080 18216
rect 16396 18164 16448 18216
rect 16488 18164 16540 18216
rect 18972 18300 19024 18352
rect 19524 18232 19576 18284
rect 22284 18300 22336 18352
rect 22744 18300 22796 18352
rect 25688 18300 25740 18352
rect 20996 18232 21048 18284
rect 21364 18232 21416 18284
rect 22376 18275 22428 18284
rect 22376 18241 22385 18275
rect 22385 18241 22419 18275
rect 22419 18241 22428 18275
rect 22376 18232 22428 18241
rect 23296 18275 23348 18284
rect 23296 18241 23305 18275
rect 23305 18241 23339 18275
rect 23339 18241 23348 18275
rect 23296 18232 23348 18241
rect 26240 18232 26292 18284
rect 26792 18232 26844 18284
rect 27528 18232 27580 18284
rect 29000 18343 29052 18352
rect 29000 18309 29009 18343
rect 29009 18309 29043 18343
rect 29043 18309 29052 18343
rect 29000 18300 29052 18309
rect 30748 18300 30800 18352
rect 31576 18300 31628 18352
rect 16764 18096 16816 18148
rect 20904 18164 20956 18216
rect 21548 18164 21600 18216
rect 11244 18028 11296 18080
rect 12716 18028 12768 18080
rect 18236 18071 18288 18080
rect 18236 18037 18245 18071
rect 18245 18037 18279 18071
rect 18279 18037 18288 18071
rect 18236 18028 18288 18037
rect 21180 18028 21232 18080
rect 21456 18028 21508 18080
rect 22008 18071 22060 18080
rect 22008 18037 22017 18071
rect 22017 18037 22051 18071
rect 22051 18037 22060 18071
rect 22008 18028 22060 18037
rect 22468 18207 22520 18216
rect 22468 18173 22477 18207
rect 22477 18173 22511 18207
rect 22511 18173 22520 18207
rect 22468 18164 22520 18173
rect 22652 18207 22704 18216
rect 22652 18173 22661 18207
rect 22661 18173 22695 18207
rect 22695 18173 22704 18207
rect 22652 18164 22704 18173
rect 25504 18164 25556 18216
rect 25964 18164 26016 18216
rect 26516 18164 26568 18216
rect 23020 18096 23072 18148
rect 23480 18096 23532 18148
rect 23756 18096 23808 18148
rect 23848 18028 23900 18080
rect 23940 18028 23992 18080
rect 26056 18028 26108 18080
rect 27620 18028 27672 18080
rect 27804 18028 27856 18080
rect 30380 18232 30432 18284
rect 32036 18232 32088 18284
rect 28816 18164 28868 18216
rect 32404 18164 32456 18216
rect 28908 18096 28960 18148
rect 33416 18164 33468 18216
rect 35256 18300 35308 18352
rect 35716 18300 35768 18352
rect 33600 18207 33652 18216
rect 33600 18173 33609 18207
rect 33609 18173 33643 18207
rect 33643 18173 33652 18207
rect 33600 18164 33652 18173
rect 37280 18232 37332 18284
rect 38660 18300 38712 18352
rect 39856 18411 39908 18420
rect 39856 18377 39865 18411
rect 39865 18377 39899 18411
rect 39899 18377 39908 18411
rect 39856 18368 39908 18377
rect 40868 18411 40920 18420
rect 40868 18377 40877 18411
rect 40877 18377 40911 18411
rect 40911 18377 40920 18411
rect 40868 18368 40920 18377
rect 41420 18368 41472 18420
rect 49240 18368 49292 18420
rect 48412 18300 48464 18352
rect 39488 18232 39540 18284
rect 49056 18275 49108 18284
rect 49056 18241 49065 18275
rect 49065 18241 49099 18275
rect 49099 18241 49108 18275
rect 49056 18232 49108 18241
rect 35348 18207 35400 18216
rect 35348 18173 35357 18207
rect 35357 18173 35391 18207
rect 35391 18173 35400 18207
rect 35348 18164 35400 18173
rect 36360 18207 36412 18216
rect 36360 18173 36369 18207
rect 36369 18173 36403 18207
rect 36403 18173 36412 18207
rect 36360 18164 36412 18173
rect 37556 18164 37608 18216
rect 39672 18164 39724 18216
rect 30196 18028 30248 18080
rect 30472 18028 30524 18080
rect 36452 18096 36504 18148
rect 38476 18028 38528 18080
rect 45560 18028 45612 18080
rect 2950 17926 3002 17978
rect 3014 17926 3066 17978
rect 3078 17926 3130 17978
rect 3142 17926 3194 17978
rect 3206 17926 3258 17978
rect 12950 17926 13002 17978
rect 13014 17926 13066 17978
rect 13078 17926 13130 17978
rect 13142 17926 13194 17978
rect 13206 17926 13258 17978
rect 22950 17926 23002 17978
rect 23014 17926 23066 17978
rect 23078 17926 23130 17978
rect 23142 17926 23194 17978
rect 23206 17926 23258 17978
rect 32950 17926 33002 17978
rect 33014 17926 33066 17978
rect 33078 17926 33130 17978
rect 33142 17926 33194 17978
rect 33206 17926 33258 17978
rect 42950 17926 43002 17978
rect 43014 17926 43066 17978
rect 43078 17926 43130 17978
rect 43142 17926 43194 17978
rect 43206 17926 43258 17978
rect 12256 17824 12308 17876
rect 12808 17824 12860 17876
rect 15108 17824 15160 17876
rect 12532 17756 12584 17808
rect 16028 17867 16080 17876
rect 16028 17833 16037 17867
rect 16037 17833 16071 17867
rect 16071 17833 16080 17867
rect 16028 17824 16080 17833
rect 18328 17824 18380 17876
rect 1216 17688 1268 17740
rect 11612 17688 11664 17740
rect 13820 17688 13872 17740
rect 14004 17688 14056 17740
rect 10508 17620 10560 17672
rect 10600 17663 10652 17672
rect 10600 17629 10609 17663
rect 10609 17629 10643 17663
rect 10643 17629 10652 17663
rect 10600 17620 10652 17629
rect 11980 17620 12032 17672
rect 12164 17484 12216 17536
rect 12716 17484 12768 17536
rect 13636 17620 13688 17672
rect 17132 17688 17184 17740
rect 18972 17688 19024 17740
rect 14556 17595 14608 17604
rect 14556 17561 14565 17595
rect 14565 17561 14599 17595
rect 14599 17561 14608 17595
rect 14556 17552 14608 17561
rect 15292 17552 15344 17604
rect 16672 17484 16724 17536
rect 17224 17484 17276 17536
rect 17776 17552 17828 17604
rect 18696 17552 18748 17604
rect 21916 17824 21968 17876
rect 22836 17824 22888 17876
rect 23848 17824 23900 17876
rect 21640 17756 21692 17808
rect 20536 17688 20588 17740
rect 23664 17688 23716 17740
rect 30104 17824 30156 17876
rect 30380 17824 30432 17876
rect 32772 17824 32824 17876
rect 28356 17756 28408 17808
rect 32680 17756 32732 17808
rect 22652 17663 22704 17672
rect 22652 17629 22661 17663
rect 22661 17629 22695 17663
rect 22695 17629 22704 17663
rect 22652 17620 22704 17629
rect 26332 17688 26384 17740
rect 25412 17620 25464 17672
rect 28540 17688 28592 17740
rect 30932 17731 30984 17740
rect 30932 17697 30941 17731
rect 30941 17697 30975 17731
rect 30975 17697 30984 17731
rect 30932 17688 30984 17697
rect 31668 17688 31720 17740
rect 34612 17824 34664 17876
rect 30840 17620 30892 17672
rect 20260 17552 20312 17604
rect 20628 17552 20680 17604
rect 20996 17552 21048 17604
rect 22192 17552 22244 17604
rect 23112 17552 23164 17604
rect 25688 17595 25740 17604
rect 25688 17561 25697 17595
rect 25697 17561 25731 17595
rect 25731 17561 25740 17595
rect 25688 17552 25740 17561
rect 26792 17552 26844 17604
rect 27804 17552 27856 17604
rect 28632 17552 28684 17604
rect 21916 17484 21968 17536
rect 22468 17527 22520 17536
rect 22468 17493 22477 17527
rect 22477 17493 22511 17527
rect 22511 17493 22520 17527
rect 22468 17484 22520 17493
rect 23664 17527 23716 17536
rect 23664 17493 23673 17527
rect 23673 17493 23707 17527
rect 23707 17493 23716 17527
rect 23664 17484 23716 17493
rect 23756 17527 23808 17536
rect 23756 17493 23765 17527
rect 23765 17493 23799 17527
rect 23799 17493 23808 17527
rect 23756 17484 23808 17493
rect 25596 17527 25648 17536
rect 25596 17493 25605 17527
rect 25605 17493 25639 17527
rect 25639 17493 25648 17527
rect 25596 17484 25648 17493
rect 25872 17484 25924 17536
rect 28816 17527 28868 17536
rect 28816 17493 28825 17527
rect 28825 17493 28859 17527
rect 28859 17493 28868 17527
rect 28816 17484 28868 17493
rect 28908 17484 28960 17536
rect 30380 17484 30432 17536
rect 31484 17484 31536 17536
rect 31944 17595 31996 17604
rect 31944 17561 31953 17595
rect 31953 17561 31987 17595
rect 31987 17561 31996 17595
rect 31944 17552 31996 17561
rect 32220 17552 32272 17604
rect 34888 17756 34940 17808
rect 33232 17731 33284 17740
rect 33232 17697 33241 17731
rect 33241 17697 33275 17731
rect 33275 17697 33284 17731
rect 33232 17688 33284 17697
rect 36820 17824 36872 17876
rect 37188 17824 37240 17876
rect 37280 17756 37332 17808
rect 40868 17756 40920 17808
rect 35716 17688 35768 17740
rect 36176 17688 36228 17740
rect 38476 17731 38528 17740
rect 38476 17697 38485 17731
rect 38485 17697 38519 17731
rect 38519 17697 38528 17731
rect 38476 17688 38528 17697
rect 35072 17663 35124 17672
rect 35072 17629 35081 17663
rect 35081 17629 35115 17663
rect 35115 17629 35124 17663
rect 35072 17620 35124 17629
rect 37372 17620 37424 17672
rect 40132 17688 40184 17740
rect 40684 17620 40736 17672
rect 49056 17663 49108 17672
rect 49056 17629 49065 17663
rect 49065 17629 49099 17663
rect 49099 17629 49108 17663
rect 49056 17620 49108 17629
rect 35992 17552 36044 17604
rect 36544 17552 36596 17604
rect 34244 17484 34296 17536
rect 34520 17484 34572 17536
rect 48412 17552 48464 17604
rect 47400 17484 47452 17536
rect 7950 17382 8002 17434
rect 8014 17382 8066 17434
rect 8078 17382 8130 17434
rect 8142 17382 8194 17434
rect 8206 17382 8258 17434
rect 17950 17382 18002 17434
rect 18014 17382 18066 17434
rect 18078 17382 18130 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 27950 17382 28002 17434
rect 28014 17382 28066 17434
rect 28078 17382 28130 17434
rect 28142 17382 28194 17434
rect 28206 17382 28258 17434
rect 37950 17382 38002 17434
rect 38014 17382 38066 17434
rect 38078 17382 38130 17434
rect 38142 17382 38194 17434
rect 38206 17382 38258 17434
rect 47950 17382 48002 17434
rect 48014 17382 48066 17434
rect 48078 17382 48130 17434
rect 48142 17382 48194 17434
rect 48206 17382 48258 17434
rect 12624 17280 12676 17332
rect 13360 17280 13412 17332
rect 15568 17323 15620 17332
rect 15568 17289 15577 17323
rect 15577 17289 15611 17323
rect 15611 17289 15620 17323
rect 15568 17280 15620 17289
rect 18788 17280 18840 17332
rect 5356 17212 5408 17264
rect 14188 17255 14240 17264
rect 14188 17221 14197 17255
rect 14197 17221 14231 17255
rect 14231 17221 14240 17255
rect 14188 17212 14240 17221
rect 14464 17212 14516 17264
rect 8300 17144 8352 17196
rect 10692 17144 10744 17196
rect 11520 17144 11572 17196
rect 1308 17076 1360 17128
rect 10232 17076 10284 17128
rect 10416 17076 10468 17128
rect 10968 17119 11020 17128
rect 10968 17085 10977 17119
rect 10977 17085 11011 17119
rect 11011 17085 11020 17119
rect 10968 17076 11020 17085
rect 12072 17144 12124 17196
rect 12440 17144 12492 17196
rect 15660 17144 15712 17196
rect 15752 17144 15804 17196
rect 12256 17076 12308 17128
rect 15016 17076 15068 17128
rect 16580 17144 16632 17196
rect 19156 17212 19208 17264
rect 6828 17008 6880 17060
rect 15292 17008 15344 17060
rect 9864 16940 9916 16992
rect 15476 16940 15528 16992
rect 15936 17008 15988 17060
rect 17776 17144 17828 17196
rect 19616 17212 19668 17264
rect 19984 17212 20036 17264
rect 20904 17280 20956 17332
rect 22652 17280 22704 17332
rect 27436 17280 27488 17332
rect 28908 17280 28960 17332
rect 29092 17323 29144 17332
rect 29092 17289 29101 17323
rect 29101 17289 29135 17323
rect 29135 17289 29144 17323
rect 29092 17280 29144 17289
rect 29460 17280 29512 17332
rect 32036 17280 32088 17332
rect 23112 17212 23164 17264
rect 23480 17212 23532 17264
rect 24308 17212 24360 17264
rect 22744 17187 22796 17196
rect 22744 17153 22753 17187
rect 22753 17153 22787 17187
rect 22787 17153 22796 17187
rect 22744 17144 22796 17153
rect 25320 17187 25372 17196
rect 25320 17153 25329 17187
rect 25329 17153 25363 17187
rect 25363 17153 25372 17187
rect 25320 17144 25372 17153
rect 18696 17119 18748 17128
rect 18696 17085 18705 17119
rect 18705 17085 18739 17119
rect 18739 17085 18748 17119
rect 18696 17076 18748 17085
rect 20076 17076 20128 17128
rect 24492 17119 24544 17128
rect 24492 17085 24501 17119
rect 24501 17085 24535 17119
rect 24535 17085 24544 17119
rect 24492 17076 24544 17085
rect 25228 17076 25280 17128
rect 26148 17212 26200 17264
rect 30932 17212 30984 17264
rect 33600 17280 33652 17332
rect 35072 17280 35124 17332
rect 36452 17280 36504 17332
rect 48412 17323 48464 17332
rect 48412 17289 48421 17323
rect 48421 17289 48455 17323
rect 48455 17289 48464 17323
rect 48412 17280 48464 17289
rect 34428 17212 34480 17264
rect 34612 17255 34664 17264
rect 34612 17221 34621 17255
rect 34621 17221 34655 17255
rect 34655 17221 34664 17255
rect 34612 17212 34664 17221
rect 38384 17212 38436 17264
rect 39212 17255 39264 17264
rect 39212 17221 39221 17255
rect 39221 17221 39255 17255
rect 39255 17221 39264 17255
rect 39212 17212 39264 17221
rect 39672 17212 39724 17264
rect 48228 17212 48280 17264
rect 26976 17144 27028 17196
rect 27436 17144 27488 17196
rect 27712 17187 27764 17196
rect 27712 17153 27721 17187
rect 27721 17153 27755 17187
rect 27755 17153 27764 17187
rect 27712 17144 27764 17153
rect 28632 17144 28684 17196
rect 29552 17144 29604 17196
rect 31300 17144 31352 17196
rect 27804 17119 27856 17128
rect 27804 17085 27813 17119
rect 27813 17085 27847 17119
rect 27847 17085 27856 17119
rect 27804 17076 27856 17085
rect 27988 17119 28040 17128
rect 27988 17085 27997 17119
rect 27997 17085 28031 17119
rect 28031 17085 28040 17119
rect 27988 17076 28040 17085
rect 22008 16940 22060 16992
rect 22744 16940 22796 16992
rect 23388 16940 23440 16992
rect 23572 16940 23624 16992
rect 25780 17008 25832 17060
rect 29092 17008 29144 17060
rect 29920 17076 29972 17128
rect 30564 17076 30616 17128
rect 30472 17008 30524 17060
rect 25596 16940 25648 16992
rect 28356 16940 28408 16992
rect 28724 16983 28776 16992
rect 28724 16949 28733 16983
rect 28733 16949 28767 16983
rect 28767 16949 28776 16983
rect 28724 16940 28776 16949
rect 30932 16940 30984 16992
rect 31024 16983 31076 16992
rect 31024 16949 31033 16983
rect 31033 16949 31067 16983
rect 31067 16949 31076 16983
rect 31024 16940 31076 16949
rect 32312 17187 32364 17196
rect 32312 17153 32321 17187
rect 32321 17153 32355 17187
rect 32355 17153 32364 17187
rect 32312 17144 32364 17153
rect 38844 17144 38896 17196
rect 48596 17187 48648 17196
rect 48596 17153 48605 17187
rect 48605 17153 48639 17187
rect 48639 17153 48648 17187
rect 48596 17144 48648 17153
rect 32220 17076 32272 17128
rect 32680 17076 32732 17128
rect 34796 17076 34848 17128
rect 34888 17076 34940 17128
rect 36176 17076 36228 17128
rect 37556 17076 37608 17128
rect 37648 17076 37700 17128
rect 36084 17008 36136 17060
rect 37740 17008 37792 17060
rect 33876 16940 33928 16992
rect 34060 16983 34112 16992
rect 34060 16949 34069 16983
rect 34069 16949 34103 16983
rect 34103 16949 34112 16983
rect 34060 16940 34112 16949
rect 37556 16940 37608 16992
rect 47400 17008 47452 17060
rect 40684 16983 40736 16992
rect 40684 16949 40693 16983
rect 40693 16949 40727 16983
rect 40727 16949 40736 16983
rect 40684 16940 40736 16949
rect 49240 16983 49292 16992
rect 49240 16949 49249 16983
rect 49249 16949 49283 16983
rect 49283 16949 49292 16983
rect 49240 16940 49292 16949
rect 2950 16838 3002 16890
rect 3014 16838 3066 16890
rect 3078 16838 3130 16890
rect 3142 16838 3194 16890
rect 3206 16838 3258 16890
rect 12950 16838 13002 16890
rect 13014 16838 13066 16890
rect 13078 16838 13130 16890
rect 13142 16838 13194 16890
rect 13206 16838 13258 16890
rect 22950 16838 23002 16890
rect 23014 16838 23066 16890
rect 23078 16838 23130 16890
rect 23142 16838 23194 16890
rect 23206 16838 23258 16890
rect 32950 16838 33002 16890
rect 33014 16838 33066 16890
rect 33078 16838 33130 16890
rect 33142 16838 33194 16890
rect 33206 16838 33258 16890
rect 42950 16838 43002 16890
rect 43014 16838 43066 16890
rect 43078 16838 43130 16890
rect 43142 16838 43194 16890
rect 43206 16838 43258 16890
rect 10508 16779 10560 16788
rect 10508 16745 10517 16779
rect 10517 16745 10551 16779
rect 10551 16745 10560 16779
rect 10508 16736 10560 16745
rect 11888 16736 11940 16788
rect 16028 16736 16080 16788
rect 16120 16736 16172 16788
rect 17224 16736 17276 16788
rect 18512 16736 18564 16788
rect 21916 16736 21968 16788
rect 22008 16736 22060 16788
rect 22468 16736 22520 16788
rect 23664 16736 23716 16788
rect 27344 16779 27396 16788
rect 10968 16668 11020 16720
rect 12256 16668 12308 16720
rect 12532 16668 12584 16720
rect 4436 16600 4488 16652
rect 5448 16600 5500 16652
rect 8576 16600 8628 16652
rect 10876 16600 10928 16652
rect 13912 16600 13964 16652
rect 14832 16600 14884 16652
rect 15108 16643 15160 16652
rect 15108 16609 15117 16643
rect 15117 16609 15151 16643
rect 15151 16609 15160 16643
rect 15108 16600 15160 16609
rect 15844 16600 15896 16652
rect 16948 16668 17000 16720
rect 16304 16643 16356 16652
rect 16304 16609 16313 16643
rect 16313 16609 16347 16643
rect 16347 16609 16356 16643
rect 16304 16600 16356 16609
rect 17132 16643 17184 16652
rect 17132 16609 17141 16643
rect 17141 16609 17175 16643
rect 17175 16609 17184 16643
rect 17132 16600 17184 16609
rect 18696 16600 18748 16652
rect 19616 16643 19668 16652
rect 19616 16609 19625 16643
rect 19625 16609 19659 16643
rect 19659 16609 19668 16643
rect 19616 16600 19668 16609
rect 20536 16600 20588 16652
rect 22468 16600 22520 16652
rect 23572 16600 23624 16652
rect 23940 16668 23992 16720
rect 27344 16745 27353 16779
rect 27353 16745 27387 16779
rect 27387 16745 27396 16779
rect 27344 16736 27396 16745
rect 27620 16736 27672 16788
rect 27988 16736 28040 16788
rect 29276 16736 29328 16788
rect 25412 16600 25464 16652
rect 25872 16643 25924 16652
rect 25872 16609 25881 16643
rect 25881 16609 25915 16643
rect 25915 16609 25924 16643
rect 25872 16600 25924 16609
rect 26240 16600 26292 16652
rect 30656 16668 30708 16720
rect 31024 16736 31076 16788
rect 33968 16736 34020 16788
rect 34796 16736 34848 16788
rect 49240 16736 49292 16788
rect 30012 16600 30064 16652
rect 31392 16643 31444 16652
rect 31392 16609 31401 16643
rect 31401 16609 31435 16643
rect 31435 16609 31444 16643
rect 31392 16600 31444 16609
rect 31576 16643 31628 16652
rect 31576 16609 31585 16643
rect 31585 16609 31619 16643
rect 31619 16609 31628 16643
rect 31576 16600 31628 16609
rect 32312 16643 32364 16652
rect 32312 16609 32321 16643
rect 32321 16609 32355 16643
rect 32355 16609 32364 16643
rect 32312 16600 32364 16609
rect 35624 16668 35676 16720
rect 33324 16600 33376 16652
rect 34060 16600 34112 16652
rect 35716 16643 35768 16652
rect 35716 16609 35725 16643
rect 35725 16609 35759 16643
rect 35759 16609 35768 16643
rect 35716 16600 35768 16609
rect 36820 16643 36872 16652
rect 36820 16609 36829 16643
rect 36829 16609 36863 16643
rect 36863 16609 36872 16643
rect 36820 16600 36872 16609
rect 37188 16600 37240 16652
rect 40684 16600 40736 16652
rect 6828 16532 6880 16584
rect 7564 16532 7616 16584
rect 11060 16532 11112 16584
rect 12440 16532 12492 16584
rect 1308 16464 1360 16516
rect 9588 16464 9640 16516
rect 11336 16464 11388 16516
rect 12624 16464 12676 16516
rect 13544 16464 13596 16516
rect 15660 16532 15712 16584
rect 16028 16575 16080 16584
rect 16028 16541 16037 16575
rect 16037 16541 16071 16575
rect 16071 16541 16080 16575
rect 16028 16532 16080 16541
rect 11060 16439 11112 16448
rect 11060 16405 11069 16439
rect 11069 16405 11103 16439
rect 11103 16405 11112 16439
rect 11060 16396 11112 16405
rect 11520 16439 11572 16448
rect 11520 16405 11529 16439
rect 11529 16405 11563 16439
rect 11563 16405 11572 16439
rect 11520 16396 11572 16405
rect 12072 16396 12124 16448
rect 13268 16396 13320 16448
rect 14464 16439 14516 16448
rect 14464 16405 14473 16439
rect 14473 16405 14507 16439
rect 14507 16405 14516 16439
rect 14464 16396 14516 16405
rect 16120 16396 16172 16448
rect 17684 16464 17736 16516
rect 20260 16575 20312 16584
rect 20260 16541 20269 16575
rect 20269 16541 20303 16575
rect 20303 16541 20312 16575
rect 20260 16532 20312 16541
rect 20720 16464 20772 16516
rect 20996 16464 21048 16516
rect 25504 16532 25556 16584
rect 18328 16396 18380 16448
rect 18696 16396 18748 16448
rect 18788 16396 18840 16448
rect 18880 16439 18932 16448
rect 18880 16405 18889 16439
rect 18889 16405 18923 16439
rect 18923 16405 18932 16439
rect 18880 16396 18932 16405
rect 19800 16396 19852 16448
rect 20168 16396 20220 16448
rect 25136 16464 25188 16516
rect 26608 16464 26660 16516
rect 29184 16464 29236 16516
rect 30196 16507 30248 16516
rect 30196 16473 30205 16507
rect 30205 16473 30239 16507
rect 30239 16473 30248 16507
rect 30196 16464 30248 16473
rect 22836 16396 22888 16448
rect 23388 16396 23440 16448
rect 25964 16396 26016 16448
rect 31852 16464 31904 16516
rect 31300 16439 31352 16448
rect 31300 16405 31309 16439
rect 31309 16405 31343 16439
rect 31343 16405 31352 16439
rect 31300 16396 31352 16405
rect 34612 16532 34664 16584
rect 35992 16532 36044 16584
rect 37740 16575 37792 16584
rect 37740 16541 37749 16575
rect 37749 16541 37783 16575
rect 37783 16541 37792 16575
rect 37740 16532 37792 16541
rect 49148 16532 49200 16584
rect 34428 16464 34480 16516
rect 39580 16464 39632 16516
rect 33600 16396 33652 16448
rect 34060 16439 34112 16448
rect 34060 16405 34069 16439
rect 34069 16405 34103 16439
rect 34103 16405 34112 16439
rect 34060 16396 34112 16405
rect 36268 16439 36320 16448
rect 36268 16405 36277 16439
rect 36277 16405 36311 16439
rect 36311 16405 36320 16439
rect 36268 16396 36320 16405
rect 37832 16396 37884 16448
rect 49240 16439 49292 16448
rect 49240 16405 49249 16439
rect 49249 16405 49283 16439
rect 49283 16405 49292 16439
rect 49240 16396 49292 16405
rect 7950 16294 8002 16346
rect 8014 16294 8066 16346
rect 8078 16294 8130 16346
rect 8142 16294 8194 16346
rect 8206 16294 8258 16346
rect 17950 16294 18002 16346
rect 18014 16294 18066 16346
rect 18078 16294 18130 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 27950 16294 28002 16346
rect 28014 16294 28066 16346
rect 28078 16294 28130 16346
rect 28142 16294 28194 16346
rect 28206 16294 28258 16346
rect 37950 16294 38002 16346
rect 38014 16294 38066 16346
rect 38078 16294 38130 16346
rect 38142 16294 38194 16346
rect 38206 16294 38258 16346
rect 47950 16294 48002 16346
rect 48014 16294 48066 16346
rect 48078 16294 48130 16346
rect 48142 16294 48194 16346
rect 48206 16294 48258 16346
rect 6368 16192 6420 16244
rect 1768 16099 1820 16108
rect 1768 16065 1777 16099
rect 1777 16065 1811 16099
rect 1811 16065 1820 16099
rect 1768 16056 1820 16065
rect 9312 16235 9364 16244
rect 9312 16201 9321 16235
rect 9321 16201 9355 16235
rect 9355 16201 9364 16235
rect 9312 16192 9364 16201
rect 11152 16192 11204 16244
rect 11520 16192 11572 16244
rect 13360 16192 13412 16244
rect 15384 16192 15436 16244
rect 12348 16124 12400 16176
rect 12716 16124 12768 16176
rect 14372 16124 14424 16176
rect 15292 16124 15344 16176
rect 16488 16192 16540 16244
rect 19800 16192 19852 16244
rect 20260 16192 20312 16244
rect 16856 16124 16908 16176
rect 17868 16124 17920 16176
rect 1308 15988 1360 16040
rect 4160 15988 4212 16040
rect 8576 16031 8628 16040
rect 8576 15997 8585 16031
rect 8585 15997 8619 16031
rect 8619 15997 8628 16031
rect 8576 15988 8628 15997
rect 11704 16056 11756 16108
rect 13728 16056 13780 16108
rect 14004 16056 14056 16108
rect 12072 15988 12124 16040
rect 12256 16031 12308 16040
rect 12256 15997 12265 16031
rect 12265 15997 12299 16031
rect 12299 15997 12308 16031
rect 12256 15988 12308 15997
rect 12440 16031 12492 16040
rect 12440 15997 12449 16031
rect 12449 15997 12483 16031
rect 12483 15997 12492 16031
rect 12440 15988 12492 15997
rect 12808 15988 12860 16040
rect 14096 15988 14148 16040
rect 14832 16031 14884 16040
rect 14832 15997 14841 16031
rect 14841 15997 14875 16031
rect 14875 15997 14884 16031
rect 14832 15988 14884 15997
rect 16304 16056 16356 16108
rect 15108 15988 15160 16040
rect 16120 16031 16172 16040
rect 16120 15997 16129 16031
rect 16129 15997 16163 16031
rect 16163 15997 16172 16031
rect 16120 15988 16172 15997
rect 18788 16124 18840 16176
rect 18880 16124 18932 16176
rect 19892 16124 19944 16176
rect 23388 16099 23440 16108
rect 23388 16065 23397 16099
rect 23397 16065 23431 16099
rect 23431 16065 23440 16099
rect 23388 16056 23440 16065
rect 25412 16192 25464 16244
rect 25964 16192 26016 16244
rect 26332 16235 26384 16244
rect 26332 16201 26341 16235
rect 26341 16201 26375 16235
rect 26375 16201 26384 16235
rect 26332 16192 26384 16201
rect 27160 16192 27212 16244
rect 30472 16192 30524 16244
rect 30932 16192 30984 16244
rect 31116 16235 31168 16244
rect 31116 16201 31125 16235
rect 31125 16201 31159 16235
rect 31159 16201 31168 16235
rect 31116 16192 31168 16201
rect 31760 16192 31812 16244
rect 32404 16192 32456 16244
rect 32772 16235 32824 16244
rect 32772 16201 32781 16235
rect 32781 16201 32815 16235
rect 32815 16201 32824 16235
rect 32772 16192 32824 16201
rect 33968 16235 34020 16244
rect 33968 16201 33977 16235
rect 33977 16201 34011 16235
rect 34011 16201 34020 16235
rect 33968 16192 34020 16201
rect 24492 16124 24544 16176
rect 25780 16124 25832 16176
rect 26608 16124 26660 16176
rect 28816 16167 28868 16176
rect 28816 16133 28825 16167
rect 28825 16133 28859 16167
rect 28859 16133 28868 16167
rect 28816 16124 28868 16133
rect 30656 16124 30708 16176
rect 37556 16192 37608 16244
rect 38844 16192 38896 16244
rect 40960 16235 41012 16244
rect 40960 16201 40969 16235
rect 40969 16201 41003 16235
rect 41003 16201 41012 16235
rect 40960 16192 41012 16201
rect 26148 16056 26200 16108
rect 18696 15988 18748 16040
rect 20720 15988 20772 16040
rect 23480 16031 23532 16040
rect 23480 15997 23489 16031
rect 23489 15997 23523 16031
rect 23523 15997 23532 16031
rect 23480 15988 23532 15997
rect 25044 15988 25096 16040
rect 28540 16099 28592 16108
rect 28540 16065 28549 16099
rect 28549 16065 28583 16099
rect 28583 16065 28592 16099
rect 28540 16056 28592 16065
rect 37832 16124 37884 16176
rect 9496 15920 9548 15972
rect 11888 15920 11940 15972
rect 14464 15920 14516 15972
rect 15384 15920 15436 15972
rect 17592 15920 17644 15972
rect 9220 15852 9272 15904
rect 12716 15852 12768 15904
rect 14372 15895 14424 15904
rect 14372 15861 14381 15895
rect 14381 15861 14415 15895
rect 14415 15861 14424 15895
rect 14372 15852 14424 15861
rect 14740 15852 14792 15904
rect 17684 15852 17736 15904
rect 19892 15852 19944 15904
rect 20904 15895 20956 15904
rect 20904 15861 20913 15895
rect 20913 15861 20947 15895
rect 20947 15861 20956 15895
rect 20904 15852 20956 15861
rect 23848 15852 23900 15904
rect 26792 15920 26844 15972
rect 31208 16031 31260 16040
rect 31208 15997 31217 16031
rect 31217 15997 31251 16031
rect 31251 15997 31260 16031
rect 31208 15988 31260 15997
rect 31944 15988 31996 16040
rect 32864 16031 32916 16040
rect 32864 15997 32873 16031
rect 32873 15997 32907 16031
rect 32907 15997 32916 16031
rect 32864 15988 32916 15997
rect 33324 16056 33376 16108
rect 36452 16056 36504 16108
rect 39580 16056 39632 16108
rect 48964 16056 49016 16108
rect 49056 16099 49108 16108
rect 49056 16065 49065 16099
rect 49065 16065 49099 16099
rect 49099 16065 49108 16099
rect 49056 16056 49108 16065
rect 33784 15988 33836 16040
rect 29920 15920 29972 15972
rect 30196 15920 30248 15972
rect 32220 15920 32272 15972
rect 34888 15988 34940 16040
rect 37372 15988 37424 16040
rect 37740 15988 37792 16040
rect 32128 15852 32180 15904
rect 32312 15895 32364 15904
rect 32312 15861 32321 15895
rect 32321 15861 32355 15895
rect 32355 15861 32364 15895
rect 32312 15852 32364 15861
rect 35808 15852 35860 15904
rect 35900 15852 35952 15904
rect 36912 15920 36964 15972
rect 38016 15920 38068 15972
rect 41788 15988 41840 16040
rect 38660 15852 38712 15904
rect 39948 15895 40000 15904
rect 39948 15861 39957 15895
rect 39957 15861 39991 15895
rect 39991 15861 40000 15895
rect 39948 15852 40000 15861
rect 48688 15852 48740 15904
rect 2950 15750 3002 15802
rect 3014 15750 3066 15802
rect 3078 15750 3130 15802
rect 3142 15750 3194 15802
rect 3206 15750 3258 15802
rect 12950 15750 13002 15802
rect 13014 15750 13066 15802
rect 13078 15750 13130 15802
rect 13142 15750 13194 15802
rect 13206 15750 13258 15802
rect 22950 15750 23002 15802
rect 23014 15750 23066 15802
rect 23078 15750 23130 15802
rect 23142 15750 23194 15802
rect 23206 15750 23258 15802
rect 32950 15750 33002 15802
rect 33014 15750 33066 15802
rect 33078 15750 33130 15802
rect 33142 15750 33194 15802
rect 33206 15750 33258 15802
rect 42950 15750 43002 15802
rect 43014 15750 43066 15802
rect 43078 15750 43130 15802
rect 43142 15750 43194 15802
rect 43206 15750 43258 15802
rect 1768 15648 1820 15700
rect 1308 15512 1360 15564
rect 10600 15512 10652 15564
rect 11060 15648 11112 15700
rect 12256 15648 12308 15700
rect 13268 15648 13320 15700
rect 13452 15580 13504 15632
rect 15568 15691 15620 15700
rect 15568 15657 15577 15691
rect 15577 15657 15611 15691
rect 15611 15657 15620 15691
rect 15568 15648 15620 15657
rect 16764 15691 16816 15700
rect 16764 15657 16773 15691
rect 16773 15657 16807 15691
rect 16807 15657 16816 15691
rect 16764 15648 16816 15657
rect 16948 15648 17000 15700
rect 11060 15512 11112 15564
rect 13360 15512 13412 15564
rect 14556 15580 14608 15632
rect 18420 15648 18472 15700
rect 19156 15648 19208 15700
rect 20444 15648 20496 15700
rect 23480 15648 23532 15700
rect 15016 15512 15068 15564
rect 16120 15555 16172 15564
rect 16120 15521 16129 15555
rect 16129 15521 16163 15555
rect 16163 15521 16172 15555
rect 16120 15512 16172 15521
rect 16304 15512 16356 15564
rect 21640 15580 21692 15632
rect 18328 15512 18380 15564
rect 19064 15512 19116 15564
rect 21364 15512 21416 15564
rect 21456 15512 21508 15564
rect 23664 15555 23716 15564
rect 23664 15521 23673 15555
rect 23673 15521 23707 15555
rect 23707 15521 23716 15555
rect 23664 15512 23716 15521
rect 24860 15512 24912 15564
rect 26516 15648 26568 15700
rect 31300 15648 31352 15700
rect 32220 15691 32272 15700
rect 32220 15657 32229 15691
rect 32229 15657 32263 15691
rect 32263 15657 32272 15691
rect 32220 15648 32272 15657
rect 34060 15648 34112 15700
rect 36360 15648 36412 15700
rect 37372 15648 37424 15700
rect 37648 15648 37700 15700
rect 41788 15691 41840 15700
rect 41788 15657 41797 15691
rect 41797 15657 41831 15691
rect 41831 15657 41840 15691
rect 41788 15648 41840 15657
rect 48964 15648 49016 15700
rect 10416 15444 10468 15496
rect 12348 15444 12400 15496
rect 10968 15376 11020 15428
rect 6644 15351 6696 15360
rect 6644 15317 6653 15351
rect 6653 15317 6687 15351
rect 6687 15317 6696 15351
rect 6644 15308 6696 15317
rect 12072 15376 12124 15428
rect 13268 15376 13320 15428
rect 14372 15444 14424 15496
rect 15292 15444 15344 15496
rect 18420 15444 18472 15496
rect 22836 15444 22888 15496
rect 24676 15444 24728 15496
rect 26056 15444 26108 15496
rect 26240 15487 26292 15496
rect 26240 15453 26249 15487
rect 26249 15453 26283 15487
rect 26283 15453 26292 15487
rect 26240 15444 26292 15453
rect 16120 15376 16172 15428
rect 12440 15308 12492 15360
rect 13544 15308 13596 15360
rect 14832 15308 14884 15360
rect 16948 15308 17000 15360
rect 17040 15308 17092 15360
rect 19984 15308 20036 15360
rect 21548 15351 21600 15360
rect 21548 15317 21557 15351
rect 21557 15317 21591 15351
rect 21591 15317 21600 15351
rect 21548 15308 21600 15317
rect 21732 15308 21784 15360
rect 25412 15376 25464 15428
rect 26148 15376 26200 15428
rect 29736 15580 29788 15632
rect 34796 15580 34848 15632
rect 26424 15555 26476 15564
rect 26424 15521 26433 15555
rect 26433 15521 26467 15555
rect 26467 15521 26476 15555
rect 26424 15512 26476 15521
rect 26516 15512 26568 15564
rect 28540 15512 28592 15564
rect 32404 15512 32456 15564
rect 33508 15512 33560 15564
rect 35164 15512 35216 15564
rect 28356 15444 28408 15496
rect 30012 15487 30064 15496
rect 30012 15453 30021 15487
rect 30021 15453 30055 15487
rect 30055 15453 30064 15487
rect 30012 15444 30064 15453
rect 34060 15487 34112 15496
rect 34060 15453 34069 15487
rect 34069 15453 34103 15487
rect 34103 15453 34112 15487
rect 34060 15444 34112 15453
rect 34888 15487 34940 15496
rect 34888 15453 34897 15487
rect 34897 15453 34931 15487
rect 34931 15453 34940 15487
rect 34888 15444 34940 15453
rect 37096 15444 37148 15496
rect 37740 15487 37792 15496
rect 37740 15453 37749 15487
rect 37749 15453 37783 15487
rect 37783 15453 37792 15487
rect 37740 15444 37792 15453
rect 49332 15487 49384 15496
rect 49332 15453 49341 15487
rect 49341 15453 49375 15487
rect 49375 15453 49384 15487
rect 49332 15444 49384 15453
rect 28448 15376 28500 15428
rect 30288 15376 30340 15428
rect 30472 15376 30524 15428
rect 34428 15376 34480 15428
rect 36452 15376 36504 15428
rect 37556 15376 37608 15428
rect 38016 15419 38068 15428
rect 38016 15385 38025 15419
rect 38025 15385 38059 15419
rect 38059 15385 38068 15419
rect 38016 15376 38068 15385
rect 26608 15308 26660 15360
rect 29644 15308 29696 15360
rect 30380 15308 30432 15360
rect 31116 15308 31168 15360
rect 31760 15308 31812 15360
rect 32036 15308 32088 15360
rect 32404 15308 32456 15360
rect 33692 15308 33744 15360
rect 34520 15308 34572 15360
rect 35256 15308 35308 15360
rect 35900 15308 35952 15360
rect 39948 15376 40000 15428
rect 39580 15308 39632 15360
rect 7950 15206 8002 15258
rect 8014 15206 8066 15258
rect 8078 15206 8130 15258
rect 8142 15206 8194 15258
rect 8206 15206 8258 15258
rect 17950 15206 18002 15258
rect 18014 15206 18066 15258
rect 18078 15206 18130 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 27950 15206 28002 15258
rect 28014 15206 28066 15258
rect 28078 15206 28130 15258
rect 28142 15206 28194 15258
rect 28206 15206 28258 15258
rect 37950 15206 38002 15258
rect 38014 15206 38066 15258
rect 38078 15206 38130 15258
rect 38142 15206 38194 15258
rect 38206 15206 38258 15258
rect 47950 15206 48002 15258
rect 48014 15206 48066 15258
rect 48078 15206 48130 15258
rect 48142 15206 48194 15258
rect 48206 15206 48258 15258
rect 9220 15104 9272 15156
rect 11060 15147 11112 15156
rect 11060 15113 11069 15147
rect 11069 15113 11103 15147
rect 11103 15113 11112 15147
rect 11060 15104 11112 15113
rect 11428 15104 11480 15156
rect 12256 15147 12308 15156
rect 12256 15113 12265 15147
rect 12265 15113 12299 15147
rect 12299 15113 12308 15147
rect 12256 15104 12308 15113
rect 9588 15036 9640 15088
rect 6644 14968 6696 15020
rect 11060 14968 11112 15020
rect 11796 14968 11848 15020
rect 12164 14968 12216 15020
rect 1308 14900 1360 14952
rect 10784 14900 10836 14952
rect 13728 15104 13780 15156
rect 15660 15104 15712 15156
rect 18880 15104 18932 15156
rect 13176 15011 13228 15020
rect 13176 14977 13185 15011
rect 13185 14977 13219 15011
rect 13219 14977 13228 15011
rect 13176 14968 13228 14977
rect 13820 15036 13872 15088
rect 14188 15036 14240 15088
rect 18052 15036 18104 15088
rect 18696 15079 18748 15088
rect 18696 15045 18705 15079
rect 18705 15045 18739 15079
rect 18739 15045 18748 15079
rect 18696 15036 18748 15045
rect 19524 15147 19576 15156
rect 19524 15113 19533 15147
rect 19533 15113 19567 15147
rect 19567 15113 19576 15147
rect 19524 15104 19576 15113
rect 20352 15104 20404 15156
rect 20444 15104 20496 15156
rect 21732 15104 21784 15156
rect 22560 15104 22612 15156
rect 23756 15104 23808 15156
rect 25136 15147 25188 15156
rect 25136 15113 25145 15147
rect 25145 15113 25179 15147
rect 25179 15113 25188 15147
rect 25136 15104 25188 15113
rect 20812 15036 20864 15088
rect 21088 15079 21140 15088
rect 21088 15045 21097 15079
rect 21097 15045 21131 15079
rect 21131 15045 21140 15079
rect 21088 15036 21140 15045
rect 21180 15036 21232 15088
rect 2320 14832 2372 14884
rect 12256 14832 12308 14884
rect 15016 14943 15068 14952
rect 15016 14909 15025 14943
rect 15025 14909 15059 14943
rect 15059 14909 15068 14943
rect 15016 14900 15068 14909
rect 13176 14832 13228 14884
rect 16948 14832 17000 14884
rect 18236 14968 18288 15020
rect 18328 14968 18380 15020
rect 17316 14943 17368 14952
rect 17316 14909 17325 14943
rect 17325 14909 17359 14943
rect 17359 14909 17368 14943
rect 17316 14900 17368 14909
rect 17408 14943 17460 14952
rect 17408 14909 17417 14943
rect 17417 14909 17451 14943
rect 17451 14909 17460 14943
rect 17408 14900 17460 14909
rect 18420 14900 18472 14952
rect 18788 15011 18840 15020
rect 18788 14977 18797 15011
rect 18797 14977 18831 15011
rect 18831 14977 18840 15011
rect 18788 14968 18840 14977
rect 20904 14968 20956 15020
rect 22100 14968 22152 15020
rect 24400 14968 24452 15020
rect 24860 15036 24912 15088
rect 25688 15036 25740 15088
rect 26700 15104 26752 15156
rect 20076 14943 20128 14952
rect 20076 14909 20085 14943
rect 20085 14909 20119 14943
rect 20119 14909 20128 14943
rect 20076 14900 20128 14909
rect 20352 14900 20404 14952
rect 17224 14832 17276 14884
rect 17500 14832 17552 14884
rect 20996 14900 21048 14952
rect 22652 14900 22704 14952
rect 22744 14832 22796 14884
rect 24124 14900 24176 14952
rect 25504 15011 25556 15020
rect 25504 14977 25513 15011
rect 25513 14977 25547 15011
rect 25547 14977 25556 15011
rect 25504 14968 25556 14977
rect 27528 15011 27580 15020
rect 27528 14977 27537 15011
rect 27537 14977 27571 15011
rect 27571 14977 27580 15011
rect 27528 14968 27580 14977
rect 31116 15104 31168 15156
rect 32036 15104 32088 15156
rect 32312 15104 32364 15156
rect 33692 15104 33744 15156
rect 34060 15104 34112 15156
rect 35164 15104 35216 15156
rect 25872 14900 25924 14952
rect 26148 14900 26200 14952
rect 28356 14968 28408 15020
rect 30748 15036 30800 15088
rect 29736 14968 29788 15020
rect 31760 14968 31812 15020
rect 24768 14832 24820 14884
rect 29276 14900 29328 14952
rect 29552 14943 29604 14952
rect 29552 14909 29561 14943
rect 29561 14909 29595 14943
rect 29595 14909 29604 14943
rect 29552 14900 29604 14909
rect 29460 14832 29512 14884
rect 30380 14900 30432 14952
rect 31116 14900 31168 14952
rect 32588 15036 32640 15088
rect 40040 15104 40092 15156
rect 36728 15036 36780 15088
rect 37648 15036 37700 15088
rect 37832 15036 37884 15088
rect 33416 14968 33468 15020
rect 32680 14900 32732 14952
rect 32772 14900 32824 14952
rect 10876 14764 10928 14816
rect 13728 14764 13780 14816
rect 15936 14764 15988 14816
rect 18052 14764 18104 14816
rect 18420 14764 18472 14816
rect 19248 14764 19300 14816
rect 20628 14764 20680 14816
rect 24860 14764 24912 14816
rect 24952 14764 25004 14816
rect 25136 14764 25188 14816
rect 25412 14764 25464 14816
rect 26332 14764 26384 14816
rect 27436 14764 27488 14816
rect 32220 14832 32272 14884
rect 34152 14943 34204 14952
rect 34152 14909 34161 14943
rect 34161 14909 34195 14943
rect 34195 14909 34204 14943
rect 34152 14900 34204 14909
rect 34980 14900 35032 14952
rect 37188 14968 37240 15020
rect 36452 14943 36504 14952
rect 36452 14909 36461 14943
rect 36461 14909 36495 14943
rect 36495 14909 36504 14943
rect 36452 14900 36504 14909
rect 37096 14900 37148 14952
rect 38292 14900 38344 14952
rect 39304 14900 39356 14952
rect 40868 14968 40920 15020
rect 49056 15011 49108 15020
rect 49056 14977 49065 15011
rect 49065 14977 49099 15011
rect 49099 14977 49108 15011
rect 49056 14968 49108 14977
rect 48412 14900 48464 14952
rect 36636 14832 36688 14884
rect 48320 14832 48372 14884
rect 30104 14764 30156 14816
rect 31300 14764 31352 14816
rect 31668 14764 31720 14816
rect 35716 14764 35768 14816
rect 37280 14764 37332 14816
rect 38476 14764 38528 14816
rect 39304 14764 39356 14816
rect 45836 14764 45888 14816
rect 2950 14662 3002 14714
rect 3014 14662 3066 14714
rect 3078 14662 3130 14714
rect 3142 14662 3194 14714
rect 3206 14662 3258 14714
rect 12950 14662 13002 14714
rect 13014 14662 13066 14714
rect 13078 14662 13130 14714
rect 13142 14662 13194 14714
rect 13206 14662 13258 14714
rect 22950 14662 23002 14714
rect 23014 14662 23066 14714
rect 23078 14662 23130 14714
rect 23142 14662 23194 14714
rect 23206 14662 23258 14714
rect 32950 14662 33002 14714
rect 33014 14662 33066 14714
rect 33078 14662 33130 14714
rect 33142 14662 33194 14714
rect 33206 14662 33258 14714
rect 42950 14662 43002 14714
rect 43014 14662 43066 14714
rect 43078 14662 43130 14714
rect 43142 14662 43194 14714
rect 43206 14662 43258 14714
rect 10416 14603 10468 14612
rect 10416 14569 10425 14603
rect 10425 14569 10459 14603
rect 10459 14569 10468 14603
rect 10416 14560 10468 14569
rect 11244 14560 11296 14612
rect 12256 14560 12308 14612
rect 3608 14492 3660 14544
rect 12532 14492 12584 14544
rect 12624 14492 12676 14544
rect 16856 14560 16908 14612
rect 17224 14560 17276 14612
rect 20536 14560 20588 14612
rect 1308 14424 1360 14476
rect 11704 14424 11756 14476
rect 13176 14424 13228 14476
rect 13544 14467 13596 14476
rect 13544 14433 13553 14467
rect 13553 14433 13587 14467
rect 13587 14433 13596 14467
rect 13544 14424 13596 14433
rect 14924 14467 14976 14476
rect 14924 14433 14933 14467
rect 14933 14433 14967 14467
rect 14967 14433 14976 14467
rect 14924 14424 14976 14433
rect 16212 14424 16264 14476
rect 16948 14467 17000 14476
rect 16948 14433 16957 14467
rect 16957 14433 16991 14467
rect 16991 14433 17000 14467
rect 16948 14424 17000 14433
rect 19432 14492 19484 14544
rect 20444 14492 20496 14544
rect 22468 14492 22520 14544
rect 25504 14560 25556 14612
rect 26056 14560 26108 14612
rect 27804 14560 27856 14612
rect 28264 14560 28316 14612
rect 28448 14560 28500 14612
rect 33324 14560 33376 14612
rect 33416 14603 33468 14612
rect 33416 14569 33425 14603
rect 33425 14569 33459 14603
rect 33459 14569 33468 14603
rect 33416 14560 33468 14569
rect 24952 14492 25004 14544
rect 26884 14492 26936 14544
rect 10140 14288 10192 14340
rect 10324 14331 10376 14340
rect 10324 14297 10333 14331
rect 10333 14297 10367 14331
rect 10367 14297 10376 14331
rect 10324 14288 10376 14297
rect 11152 14331 11204 14340
rect 11152 14297 11161 14331
rect 11161 14297 11195 14331
rect 11195 14297 11204 14331
rect 11152 14288 11204 14297
rect 12624 14288 12676 14340
rect 15476 14399 15528 14408
rect 15476 14365 15485 14399
rect 15485 14365 15519 14399
rect 15519 14365 15528 14399
rect 15476 14356 15528 14365
rect 11244 14263 11296 14272
rect 11244 14229 11253 14263
rect 11253 14229 11287 14263
rect 11287 14229 11296 14263
rect 11244 14220 11296 14229
rect 12532 14220 12584 14272
rect 13728 14220 13780 14272
rect 15660 14220 15712 14272
rect 16764 14220 16816 14272
rect 17960 14356 18012 14408
rect 19248 14424 19300 14476
rect 20720 14424 20772 14476
rect 21364 14467 21416 14476
rect 21364 14433 21373 14467
rect 21373 14433 21407 14467
rect 21407 14433 21416 14467
rect 21364 14424 21416 14433
rect 21456 14424 21508 14476
rect 24400 14424 24452 14476
rect 25412 14424 25464 14476
rect 28264 14467 28316 14476
rect 28264 14433 28273 14467
rect 28273 14433 28307 14467
rect 28307 14433 28316 14467
rect 28264 14424 28316 14433
rect 28816 14424 28868 14476
rect 19892 14356 19944 14408
rect 20628 14356 20680 14408
rect 24952 14399 25004 14408
rect 24952 14365 24961 14399
rect 24961 14365 24995 14399
rect 24995 14365 25004 14399
rect 24952 14356 25004 14365
rect 18604 14331 18656 14340
rect 17408 14220 17460 14272
rect 18604 14297 18613 14331
rect 18613 14297 18647 14331
rect 18647 14297 18656 14331
rect 18604 14288 18656 14297
rect 19340 14288 19392 14340
rect 19800 14288 19852 14340
rect 21456 14288 21508 14340
rect 22744 14288 22796 14340
rect 23572 14288 23624 14340
rect 24860 14288 24912 14340
rect 27712 14356 27764 14408
rect 30012 14356 30064 14408
rect 30380 14492 30432 14544
rect 31668 14492 31720 14544
rect 30288 14467 30340 14476
rect 30288 14433 30297 14467
rect 30297 14433 30331 14467
rect 30331 14433 30340 14467
rect 30288 14424 30340 14433
rect 31300 14424 31352 14476
rect 18696 14220 18748 14272
rect 19524 14263 19576 14272
rect 19524 14229 19533 14263
rect 19533 14229 19567 14263
rect 19567 14229 19576 14263
rect 19524 14220 19576 14229
rect 19708 14220 19760 14272
rect 25596 14288 25648 14340
rect 25780 14288 25832 14340
rect 26700 14220 26752 14272
rect 30932 14356 30984 14408
rect 31116 14356 31168 14408
rect 34060 14492 34112 14544
rect 32312 14424 32364 14476
rect 32864 14467 32916 14476
rect 32864 14433 32873 14467
rect 32873 14433 32907 14467
rect 32907 14433 32916 14467
rect 32864 14424 32916 14433
rect 33416 14424 33468 14476
rect 33600 14424 33652 14476
rect 35348 14560 35400 14612
rect 35808 14560 35860 14612
rect 36820 14560 36872 14612
rect 39304 14492 39356 14544
rect 34888 14467 34940 14476
rect 34888 14433 34897 14467
rect 34897 14433 34931 14467
rect 34931 14433 34940 14467
rect 37096 14467 37148 14476
rect 34888 14424 34940 14433
rect 37096 14433 37105 14467
rect 37105 14433 37139 14467
rect 37139 14433 37148 14467
rect 37096 14424 37148 14433
rect 38108 14424 38160 14476
rect 32220 14356 32272 14408
rect 49056 14399 49108 14408
rect 49056 14365 49065 14399
rect 49065 14365 49099 14399
rect 49099 14365 49108 14399
rect 49056 14356 49108 14365
rect 31024 14263 31076 14272
rect 31024 14229 31033 14263
rect 31033 14229 31067 14263
rect 31067 14229 31076 14263
rect 31024 14220 31076 14229
rect 31668 14288 31720 14340
rect 33784 14331 33836 14340
rect 33784 14297 33793 14331
rect 33793 14297 33827 14331
rect 33827 14297 33836 14331
rect 33784 14288 33836 14297
rect 34520 14288 34572 14340
rect 35256 14288 35308 14340
rect 36544 14288 36596 14340
rect 32036 14220 32088 14272
rect 32496 14220 32548 14272
rect 32680 14220 32732 14272
rect 34244 14220 34296 14272
rect 37832 14288 37884 14340
rect 45008 14220 45060 14272
rect 49240 14263 49292 14272
rect 49240 14229 49249 14263
rect 49249 14229 49283 14263
rect 49283 14229 49292 14263
rect 49240 14220 49292 14229
rect 7950 14118 8002 14170
rect 8014 14118 8066 14170
rect 8078 14118 8130 14170
rect 8142 14118 8194 14170
rect 8206 14118 8258 14170
rect 17950 14118 18002 14170
rect 18014 14118 18066 14170
rect 18078 14118 18130 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 27950 14118 28002 14170
rect 28014 14118 28066 14170
rect 28078 14118 28130 14170
rect 28142 14118 28194 14170
rect 28206 14118 28258 14170
rect 37950 14118 38002 14170
rect 38014 14118 38066 14170
rect 38078 14118 38130 14170
rect 38142 14118 38194 14170
rect 38206 14118 38258 14170
rect 47950 14118 48002 14170
rect 48014 14118 48066 14170
rect 48078 14118 48130 14170
rect 48142 14118 48194 14170
rect 48206 14118 48258 14170
rect 3608 14059 3660 14068
rect 3608 14025 3617 14059
rect 3617 14025 3651 14059
rect 3651 14025 3660 14059
rect 3608 14016 3660 14025
rect 11980 14016 12032 14068
rect 14556 14016 14608 14068
rect 15292 14016 15344 14068
rect 15936 14059 15988 14068
rect 15936 14025 15945 14059
rect 15945 14025 15979 14059
rect 15979 14025 15988 14059
rect 15936 14016 15988 14025
rect 16764 14016 16816 14068
rect 17500 14059 17552 14068
rect 17500 14025 17509 14059
rect 17509 14025 17543 14059
rect 17543 14025 17552 14059
rect 17500 14016 17552 14025
rect 17592 14059 17644 14068
rect 17592 14025 17601 14059
rect 17601 14025 17635 14059
rect 17635 14025 17644 14059
rect 17592 14016 17644 14025
rect 17868 14016 17920 14068
rect 19616 14016 19668 14068
rect 21364 14016 21416 14068
rect 21640 14016 21692 14068
rect 26056 14016 26108 14068
rect 26424 14016 26476 14068
rect 27620 14016 27672 14068
rect 31300 14016 31352 14068
rect 31668 14016 31720 14068
rect 11244 13948 11296 14000
rect 14188 13948 14240 14000
rect 19524 13948 19576 14000
rect 20076 13948 20128 14000
rect 22744 13948 22796 14000
rect 23572 13948 23624 14000
rect 24676 13948 24728 14000
rect 25228 13948 25280 14000
rect 25412 13948 25464 14000
rect 25780 13948 25832 14000
rect 26700 13948 26752 14000
rect 3516 13923 3568 13932
rect 3516 13889 3525 13923
rect 3525 13889 3559 13923
rect 3559 13889 3568 13923
rect 3516 13880 3568 13889
rect 19340 13880 19392 13932
rect 24860 13923 24912 13932
rect 24860 13889 24869 13923
rect 24869 13889 24903 13923
rect 24903 13889 24912 13923
rect 24860 13880 24912 13889
rect 27160 13923 27212 13932
rect 27160 13889 27169 13923
rect 27169 13889 27203 13923
rect 27203 13889 27212 13923
rect 27160 13880 27212 13889
rect 30656 13948 30708 14000
rect 32036 13948 32088 14000
rect 32680 13948 32732 14000
rect 34060 14059 34112 14068
rect 34060 14025 34069 14059
rect 34069 14025 34103 14059
rect 34103 14025 34112 14059
rect 34060 14016 34112 14025
rect 34796 14016 34848 14068
rect 36268 13948 36320 14000
rect 33692 13880 33744 13932
rect 34428 13880 34480 13932
rect 1308 13812 1360 13864
rect 11796 13812 11848 13864
rect 12808 13812 12860 13864
rect 13176 13855 13228 13864
rect 13176 13821 13185 13855
rect 13185 13821 13219 13855
rect 13219 13821 13228 13855
rect 13176 13812 13228 13821
rect 13636 13812 13688 13864
rect 12440 13744 12492 13796
rect 16580 13812 16632 13864
rect 17316 13812 17368 13864
rect 12900 13676 12952 13728
rect 15936 13676 15988 13728
rect 17684 13744 17736 13796
rect 18512 13744 18564 13796
rect 18972 13812 19024 13864
rect 16488 13676 16540 13728
rect 22008 13855 22060 13864
rect 22008 13821 22017 13855
rect 22017 13821 22051 13855
rect 22051 13821 22060 13855
rect 22008 13812 22060 13821
rect 22284 13855 22336 13864
rect 22284 13821 22293 13855
rect 22293 13821 22327 13855
rect 22327 13821 22336 13855
rect 22284 13812 22336 13821
rect 23664 13812 23716 13864
rect 25504 13812 25556 13864
rect 27620 13812 27672 13864
rect 28908 13855 28960 13864
rect 28908 13821 28917 13855
rect 28917 13821 28951 13855
rect 28951 13821 28960 13855
rect 28908 13812 28960 13821
rect 30840 13812 30892 13864
rect 32220 13812 32272 13864
rect 23756 13787 23808 13796
rect 23756 13753 23765 13787
rect 23765 13753 23799 13787
rect 23799 13753 23808 13787
rect 23756 13744 23808 13753
rect 31760 13744 31812 13796
rect 32588 13855 32640 13864
rect 32588 13821 32597 13855
rect 32597 13821 32631 13855
rect 32631 13821 32640 13855
rect 32588 13812 32640 13821
rect 32680 13812 32732 13864
rect 33600 13812 33652 13864
rect 37372 13880 37424 13932
rect 41512 14016 41564 14068
rect 47032 14016 47084 14068
rect 48412 14059 48464 14068
rect 48412 14025 48421 14059
rect 48421 14025 48455 14059
rect 48455 14025 48464 14059
rect 48412 14016 48464 14025
rect 48504 14016 48556 14068
rect 45008 13991 45060 14000
rect 45008 13957 45017 13991
rect 45017 13957 45051 13991
rect 45051 13957 45060 13991
rect 45008 13948 45060 13957
rect 46848 13948 46900 14000
rect 48688 13948 48740 14000
rect 49148 13991 49200 14000
rect 49148 13957 49157 13991
rect 49157 13957 49191 13991
rect 49191 13957 49200 13991
rect 49148 13948 49200 13957
rect 34704 13812 34756 13864
rect 35992 13812 36044 13864
rect 36636 13812 36688 13864
rect 36820 13812 36872 13864
rect 45836 13923 45888 13932
rect 45836 13889 45845 13923
rect 45845 13889 45879 13923
rect 45879 13889 45888 13923
rect 45836 13880 45888 13889
rect 48228 13880 48280 13932
rect 37832 13744 37884 13796
rect 46296 13812 46348 13864
rect 22836 13676 22888 13728
rect 23940 13676 23992 13728
rect 26240 13676 26292 13728
rect 30932 13676 30984 13728
rect 31116 13676 31168 13728
rect 34796 13676 34848 13728
rect 35072 13676 35124 13728
rect 35532 13676 35584 13728
rect 37556 13676 37608 13728
rect 38844 13719 38896 13728
rect 38844 13685 38853 13719
rect 38853 13685 38887 13719
rect 38887 13685 38896 13719
rect 38844 13676 38896 13685
rect 2950 13574 3002 13626
rect 3014 13574 3066 13626
rect 3078 13574 3130 13626
rect 3142 13574 3194 13626
rect 3206 13574 3258 13626
rect 12950 13574 13002 13626
rect 13014 13574 13066 13626
rect 13078 13574 13130 13626
rect 13142 13574 13194 13626
rect 13206 13574 13258 13626
rect 22950 13574 23002 13626
rect 23014 13574 23066 13626
rect 23078 13574 23130 13626
rect 23142 13574 23194 13626
rect 23206 13574 23258 13626
rect 32950 13574 33002 13626
rect 33014 13574 33066 13626
rect 33078 13574 33130 13626
rect 33142 13574 33194 13626
rect 33206 13574 33258 13626
rect 42950 13574 43002 13626
rect 43014 13574 43066 13626
rect 43078 13574 43130 13626
rect 43142 13574 43194 13626
rect 43206 13574 43258 13626
rect 12624 13472 12676 13524
rect 2780 13311 2832 13320
rect 2780 13277 2789 13311
rect 2789 13277 2823 13311
rect 2823 13277 2832 13311
rect 2780 13268 2832 13277
rect 10508 13268 10560 13320
rect 12808 13336 12860 13388
rect 12164 13268 12216 13320
rect 12900 13268 12952 13320
rect 15108 13336 15160 13388
rect 15384 13336 15436 13388
rect 17684 13472 17736 13524
rect 20904 13515 20956 13524
rect 20904 13481 20913 13515
rect 20913 13481 20947 13515
rect 20947 13481 20956 13515
rect 20904 13472 20956 13481
rect 22192 13472 22244 13524
rect 22836 13472 22888 13524
rect 25320 13472 25372 13524
rect 27804 13472 27856 13524
rect 8576 13200 8628 13252
rect 11060 13243 11112 13252
rect 11060 13209 11069 13243
rect 11069 13209 11103 13243
rect 11103 13209 11112 13243
rect 11060 13200 11112 13209
rect 14556 13268 14608 13320
rect 18972 13336 19024 13388
rect 21456 13379 21508 13388
rect 21456 13345 21465 13379
rect 21465 13345 21499 13379
rect 21499 13345 21508 13379
rect 21456 13336 21508 13345
rect 22468 13336 22520 13388
rect 26608 13404 26660 13456
rect 23572 13336 23624 13388
rect 23848 13336 23900 13388
rect 24860 13336 24912 13388
rect 25504 13379 25556 13388
rect 25504 13345 25513 13379
rect 25513 13345 25547 13379
rect 25547 13345 25556 13379
rect 25504 13336 25556 13345
rect 26700 13336 26752 13388
rect 28632 13336 28684 13388
rect 32036 13472 32088 13524
rect 33876 13472 33928 13524
rect 38384 13472 38436 13524
rect 29000 13404 29052 13456
rect 30104 13404 30156 13456
rect 29828 13336 29880 13388
rect 30288 13379 30340 13388
rect 30288 13345 30297 13379
rect 30297 13345 30331 13379
rect 30331 13345 30340 13379
rect 30288 13336 30340 13345
rect 31760 13336 31812 13388
rect 31852 13336 31904 13388
rect 10784 13132 10836 13184
rect 12440 13132 12492 13184
rect 14924 13132 14976 13184
rect 15200 13175 15252 13184
rect 15200 13141 15209 13175
rect 15209 13141 15243 13175
rect 15243 13141 15252 13175
rect 15200 13132 15252 13141
rect 15568 13243 15620 13252
rect 15568 13209 15577 13243
rect 15577 13209 15611 13243
rect 15611 13209 15620 13243
rect 15568 13200 15620 13209
rect 15660 13200 15712 13252
rect 15844 13200 15896 13252
rect 16304 13200 16356 13252
rect 17408 13132 17460 13184
rect 17592 13132 17644 13184
rect 20076 13268 20128 13320
rect 21272 13311 21324 13320
rect 21272 13277 21281 13311
rect 21281 13277 21315 13311
rect 21315 13277 21324 13311
rect 21272 13268 21324 13277
rect 21640 13268 21692 13320
rect 23204 13268 23256 13320
rect 17960 13132 18012 13184
rect 18604 13132 18656 13184
rect 24216 13200 24268 13252
rect 24952 13268 25004 13320
rect 25596 13268 25648 13320
rect 28448 13268 28500 13320
rect 22376 13132 22428 13184
rect 23480 13132 23532 13184
rect 25320 13175 25372 13184
rect 25320 13141 25329 13175
rect 25329 13141 25363 13175
rect 25363 13141 25372 13175
rect 25320 13132 25372 13141
rect 29552 13200 29604 13252
rect 27804 13132 27856 13184
rect 29736 13268 29788 13320
rect 33692 13404 33744 13456
rect 33784 13379 33836 13388
rect 33784 13345 33793 13379
rect 33793 13345 33827 13379
rect 33827 13345 33836 13379
rect 33784 13336 33836 13345
rect 33876 13379 33928 13388
rect 33876 13345 33885 13379
rect 33885 13345 33919 13379
rect 33919 13345 33928 13379
rect 33876 13336 33928 13345
rect 34060 13336 34112 13388
rect 35164 13336 35216 13388
rect 35532 13379 35584 13388
rect 35532 13345 35541 13379
rect 35541 13345 35575 13379
rect 35575 13345 35584 13379
rect 35532 13336 35584 13345
rect 38844 13404 38896 13456
rect 33600 13268 33652 13320
rect 34152 13268 34204 13320
rect 37832 13336 37884 13388
rect 35808 13268 35860 13320
rect 41512 13311 41564 13320
rect 41512 13277 41521 13311
rect 41521 13277 41555 13311
rect 41555 13277 41564 13311
rect 41512 13268 41564 13277
rect 46296 13268 46348 13320
rect 49148 13311 49200 13320
rect 49148 13277 49157 13311
rect 49157 13277 49191 13311
rect 49191 13277 49200 13311
rect 49148 13268 49200 13277
rect 30196 13200 30248 13252
rect 30656 13200 30708 13252
rect 31116 13132 31168 13184
rect 33876 13200 33928 13252
rect 34704 13200 34756 13252
rect 36636 13243 36688 13252
rect 36636 13209 36645 13243
rect 36645 13209 36679 13243
rect 36679 13209 36688 13243
rect 36636 13200 36688 13209
rect 36360 13132 36412 13184
rect 36544 13132 36596 13184
rect 46112 13132 46164 13184
rect 7950 13030 8002 13082
rect 8014 13030 8066 13082
rect 8078 13030 8130 13082
rect 8142 13030 8194 13082
rect 8206 13030 8258 13082
rect 17950 13030 18002 13082
rect 18014 13030 18066 13082
rect 18078 13030 18130 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 27950 13030 28002 13082
rect 28014 13030 28066 13082
rect 28078 13030 28130 13082
rect 28142 13030 28194 13082
rect 28206 13030 28258 13082
rect 37950 13030 38002 13082
rect 38014 13030 38066 13082
rect 38078 13030 38130 13082
rect 38142 13030 38194 13082
rect 38206 13030 38258 13082
rect 47950 13030 48002 13082
rect 48014 13030 48066 13082
rect 48078 13030 48130 13082
rect 48142 13030 48194 13082
rect 48206 13030 48258 13082
rect 5448 12928 5500 12980
rect 10876 12928 10928 12980
rect 12256 12928 12308 12980
rect 14188 12928 14240 12980
rect 940 12860 992 12912
rect 10232 12860 10284 12912
rect 1308 12792 1360 12844
rect 16120 12928 16172 12980
rect 14648 12860 14700 12912
rect 19984 12928 20036 12980
rect 20076 12971 20128 12980
rect 20076 12937 20085 12971
rect 20085 12937 20119 12971
rect 20119 12937 20128 12971
rect 20076 12928 20128 12937
rect 23940 12971 23992 12980
rect 15384 12792 15436 12844
rect 15844 12792 15896 12844
rect 12164 12724 12216 12776
rect 12440 12724 12492 12776
rect 12808 12724 12860 12776
rect 12624 12588 12676 12640
rect 13360 12724 13412 12776
rect 13636 12724 13688 12776
rect 16488 12792 16540 12844
rect 16212 12724 16264 12776
rect 17776 12792 17828 12844
rect 18972 12860 19024 12912
rect 23940 12937 23949 12971
rect 23949 12937 23983 12971
rect 23983 12937 23992 12971
rect 23940 12928 23992 12937
rect 25044 12928 25096 12980
rect 27620 12928 27672 12980
rect 31944 12928 31996 12980
rect 16856 12724 16908 12776
rect 14280 12588 14332 12640
rect 16120 12588 16172 12640
rect 18236 12588 18288 12640
rect 19248 12835 19300 12844
rect 19248 12801 19257 12835
rect 19257 12801 19291 12835
rect 19291 12801 19300 12835
rect 19248 12792 19300 12801
rect 20720 12792 20772 12844
rect 19524 12767 19576 12776
rect 19524 12733 19533 12767
rect 19533 12733 19567 12767
rect 19567 12733 19576 12767
rect 19524 12724 19576 12733
rect 20168 12767 20220 12776
rect 20168 12733 20177 12767
rect 20177 12733 20211 12767
rect 20211 12733 20220 12767
rect 20168 12724 20220 12733
rect 20260 12767 20312 12776
rect 20260 12733 20269 12767
rect 20269 12733 20303 12767
rect 20303 12733 20312 12767
rect 20260 12724 20312 12733
rect 29552 12860 29604 12912
rect 30196 12860 30248 12912
rect 21916 12792 21968 12844
rect 22836 12792 22888 12844
rect 25412 12792 25464 12844
rect 25780 12792 25832 12844
rect 26700 12792 26752 12844
rect 27988 12835 28040 12844
rect 27988 12801 27997 12835
rect 27997 12801 28031 12835
rect 28031 12801 28040 12835
rect 27988 12792 28040 12801
rect 30104 12792 30156 12844
rect 31852 12860 31904 12912
rect 32772 12928 32824 12980
rect 35716 12928 35768 12980
rect 21272 12767 21324 12776
rect 21272 12733 21281 12767
rect 21281 12733 21315 12767
rect 21315 12733 21324 12767
rect 21272 12724 21324 12733
rect 22560 12724 22612 12776
rect 23204 12767 23256 12776
rect 23204 12733 23213 12767
rect 23213 12733 23247 12767
rect 23247 12733 23256 12767
rect 23204 12724 23256 12733
rect 23940 12724 23992 12776
rect 24308 12767 24360 12776
rect 24308 12733 24317 12767
rect 24317 12733 24351 12767
rect 24351 12733 24360 12767
rect 24308 12724 24360 12733
rect 26424 12724 26476 12776
rect 27804 12724 27856 12776
rect 29000 12724 29052 12776
rect 30656 12792 30708 12844
rect 31116 12792 31168 12844
rect 31576 12792 31628 12844
rect 31760 12792 31812 12844
rect 34612 12860 34664 12912
rect 34888 12860 34940 12912
rect 39948 12860 40000 12912
rect 22192 12631 22244 12640
rect 22192 12597 22201 12631
rect 22201 12597 22235 12631
rect 22235 12597 22244 12631
rect 22192 12588 22244 12597
rect 22652 12631 22704 12640
rect 22652 12597 22661 12631
rect 22661 12597 22695 12631
rect 22695 12597 22704 12631
rect 22652 12588 22704 12597
rect 26332 12588 26384 12640
rect 30380 12656 30432 12708
rect 30012 12588 30064 12640
rect 31208 12724 31260 12776
rect 33692 12792 33744 12844
rect 36268 12835 36320 12844
rect 36268 12801 36277 12835
rect 36277 12801 36311 12835
rect 36311 12801 36320 12835
rect 36268 12792 36320 12801
rect 34888 12724 34940 12776
rect 36360 12724 36412 12776
rect 32128 12588 32180 12640
rect 39304 12656 39356 12708
rect 34796 12588 34848 12640
rect 46112 12835 46164 12844
rect 46112 12801 46121 12835
rect 46121 12801 46155 12835
rect 46155 12801 46164 12835
rect 46112 12792 46164 12801
rect 47032 12792 47084 12844
rect 49148 12835 49200 12844
rect 49148 12801 49157 12835
rect 49157 12801 49191 12835
rect 49191 12801 49200 12835
rect 49148 12792 49200 12801
rect 42708 12588 42760 12640
rect 47952 12588 48004 12640
rect 2950 12486 3002 12538
rect 3014 12486 3066 12538
rect 3078 12486 3130 12538
rect 3142 12486 3194 12538
rect 3206 12486 3258 12538
rect 12950 12486 13002 12538
rect 13014 12486 13066 12538
rect 13078 12486 13130 12538
rect 13142 12486 13194 12538
rect 13206 12486 13258 12538
rect 22950 12486 23002 12538
rect 23014 12486 23066 12538
rect 23078 12486 23130 12538
rect 23142 12486 23194 12538
rect 23206 12486 23258 12538
rect 32950 12486 33002 12538
rect 33014 12486 33066 12538
rect 33078 12486 33130 12538
rect 33142 12486 33194 12538
rect 33206 12486 33258 12538
rect 42950 12486 43002 12538
rect 43014 12486 43066 12538
rect 43078 12486 43130 12538
rect 43142 12486 43194 12538
rect 43206 12486 43258 12538
rect 16028 12384 16080 12436
rect 16396 12384 16448 12436
rect 20628 12384 20680 12436
rect 20812 12427 20864 12436
rect 20812 12393 20821 12427
rect 20821 12393 20855 12427
rect 20855 12393 20864 12427
rect 20812 12384 20864 12393
rect 22100 12427 22152 12436
rect 22100 12393 22109 12427
rect 22109 12393 22143 12427
rect 22143 12393 22152 12427
rect 22100 12384 22152 12393
rect 23204 12384 23256 12436
rect 25872 12384 25924 12436
rect 26332 12427 26384 12436
rect 26332 12393 26341 12427
rect 26341 12393 26375 12427
rect 26375 12393 26384 12427
rect 26332 12384 26384 12393
rect 26792 12384 26844 12436
rect 28816 12384 28868 12436
rect 29552 12384 29604 12436
rect 31760 12384 31812 12436
rect 32864 12384 32916 12436
rect 33876 12427 33928 12436
rect 33876 12393 33885 12427
rect 33885 12393 33919 12427
rect 33919 12393 33928 12427
rect 33876 12384 33928 12393
rect 15568 12316 15620 12368
rect 5356 12248 5408 12300
rect 10508 12291 10560 12300
rect 10508 12257 10517 12291
rect 10517 12257 10551 12291
rect 10551 12257 10560 12291
rect 10508 12248 10560 12257
rect 10784 12291 10836 12300
rect 10784 12257 10793 12291
rect 10793 12257 10827 12291
rect 10827 12257 10836 12291
rect 10784 12248 10836 12257
rect 12716 12248 12768 12300
rect 13636 12291 13688 12300
rect 13636 12257 13645 12291
rect 13645 12257 13679 12291
rect 13679 12257 13688 12291
rect 13636 12248 13688 12257
rect 14280 12291 14332 12300
rect 14280 12257 14289 12291
rect 14289 12257 14323 12291
rect 14323 12257 14332 12291
rect 14280 12248 14332 12257
rect 14556 12248 14608 12300
rect 16856 12248 16908 12300
rect 940 12180 992 12232
rect 12256 12180 12308 12232
rect 13360 12180 13412 12232
rect 17224 12291 17276 12300
rect 17224 12257 17233 12291
rect 17233 12257 17267 12291
rect 17267 12257 17276 12291
rect 17224 12248 17276 12257
rect 18696 12248 18748 12300
rect 19984 12291 20036 12300
rect 19984 12257 19993 12291
rect 19993 12257 20027 12291
rect 20027 12257 20036 12291
rect 19984 12248 20036 12257
rect 21456 12291 21508 12300
rect 21456 12257 21465 12291
rect 21465 12257 21499 12291
rect 21499 12257 21508 12291
rect 21456 12248 21508 12257
rect 22560 12248 22612 12300
rect 23296 12316 23348 12368
rect 23756 12248 23808 12300
rect 13452 12112 13504 12164
rect 17776 12180 17828 12232
rect 18236 12180 18288 12232
rect 22192 12180 22244 12232
rect 23664 12223 23716 12232
rect 23664 12189 23673 12223
rect 23673 12189 23707 12223
rect 23707 12189 23716 12223
rect 23664 12180 23716 12189
rect 24308 12180 24360 12232
rect 24584 12223 24636 12232
rect 24584 12189 24593 12223
rect 24593 12189 24627 12223
rect 24627 12189 24636 12223
rect 24584 12180 24636 12189
rect 27528 12291 27580 12300
rect 27528 12257 27537 12291
rect 27537 12257 27571 12291
rect 27571 12257 27580 12291
rect 27528 12248 27580 12257
rect 30012 12291 30064 12300
rect 30012 12257 30021 12291
rect 30021 12257 30055 12291
rect 30055 12257 30064 12291
rect 30012 12248 30064 12257
rect 30748 12248 30800 12300
rect 31208 12248 31260 12300
rect 39396 12384 39448 12436
rect 34888 12291 34940 12300
rect 34888 12257 34897 12291
rect 34897 12257 34931 12291
rect 34931 12257 34940 12291
rect 34888 12248 34940 12257
rect 35808 12248 35860 12300
rect 37832 12248 37884 12300
rect 38292 12248 38344 12300
rect 14464 12112 14516 12164
rect 14648 12112 14700 12164
rect 12164 12044 12216 12096
rect 15292 12044 15344 12096
rect 15384 12044 15436 12096
rect 16396 12112 16448 12164
rect 16856 12112 16908 12164
rect 15936 12044 15988 12096
rect 16212 12044 16264 12096
rect 17224 12044 17276 12096
rect 21180 12044 21232 12096
rect 23204 12044 23256 12096
rect 23388 12044 23440 12096
rect 23756 12087 23808 12096
rect 23756 12053 23765 12087
rect 23765 12053 23799 12087
rect 23799 12053 23808 12087
rect 23756 12044 23808 12053
rect 24952 12112 25004 12164
rect 25412 12112 25464 12164
rect 26240 12112 26292 12164
rect 27068 12112 27120 12164
rect 28908 12112 28960 12164
rect 31116 12180 31168 12232
rect 31576 12180 31628 12232
rect 39304 12180 39356 12232
rect 25596 12044 25648 12096
rect 27252 12044 27304 12096
rect 27344 12087 27396 12096
rect 27344 12053 27353 12087
rect 27353 12053 27387 12087
rect 27387 12053 27396 12087
rect 27344 12044 27396 12053
rect 27988 12044 28040 12096
rect 28448 12044 28500 12096
rect 32496 12112 32548 12164
rect 33692 12112 33744 12164
rect 31392 12044 31444 12096
rect 34520 12044 34572 12096
rect 36544 12112 36596 12164
rect 39948 12223 40000 12232
rect 39948 12189 39957 12223
rect 39957 12189 39991 12223
rect 39991 12189 40000 12223
rect 39948 12180 40000 12189
rect 49148 12291 49200 12300
rect 49148 12257 49157 12291
rect 49157 12257 49191 12291
rect 49191 12257 49200 12291
rect 49148 12248 49200 12257
rect 47952 12223 48004 12232
rect 47952 12189 47961 12223
rect 47961 12189 47995 12223
rect 47995 12189 48004 12223
rect 47952 12180 48004 12189
rect 35440 12044 35492 12096
rect 35808 12044 35860 12096
rect 36452 12044 36504 12096
rect 36728 12044 36780 12096
rect 37648 12044 37700 12096
rect 47032 12112 47084 12164
rect 40224 12087 40276 12096
rect 40224 12053 40233 12087
rect 40233 12053 40267 12087
rect 40267 12053 40276 12087
rect 40224 12044 40276 12053
rect 45928 12087 45980 12096
rect 45928 12053 45937 12087
rect 45937 12053 45971 12087
rect 45971 12053 45980 12087
rect 45928 12044 45980 12053
rect 7950 11942 8002 11994
rect 8014 11942 8066 11994
rect 8078 11942 8130 11994
rect 8142 11942 8194 11994
rect 8206 11942 8258 11994
rect 17950 11942 18002 11994
rect 18014 11942 18066 11994
rect 18078 11942 18130 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 27950 11942 28002 11994
rect 28014 11942 28066 11994
rect 28078 11942 28130 11994
rect 28142 11942 28194 11994
rect 28206 11942 28258 11994
rect 37950 11942 38002 11994
rect 38014 11942 38066 11994
rect 38078 11942 38130 11994
rect 38142 11942 38194 11994
rect 38206 11942 38258 11994
rect 47950 11942 48002 11994
rect 48014 11942 48066 11994
rect 48078 11942 48130 11994
rect 48142 11942 48194 11994
rect 48206 11942 48258 11994
rect 1860 11840 1912 11892
rect 1032 11704 1084 11756
rect 12348 11772 12400 11824
rect 14556 11840 14608 11892
rect 19800 11840 19852 11892
rect 16580 11772 16632 11824
rect 940 11636 992 11688
rect 13452 11704 13504 11756
rect 13820 11704 13872 11756
rect 12716 11636 12768 11688
rect 4160 11500 4212 11552
rect 15292 11568 15344 11620
rect 15476 11747 15528 11756
rect 15476 11713 15485 11747
rect 15485 11713 15519 11747
rect 15519 11713 15528 11747
rect 15476 11704 15528 11713
rect 15844 11704 15896 11756
rect 16396 11704 16448 11756
rect 17592 11772 17644 11824
rect 16856 11679 16908 11688
rect 16856 11645 16865 11679
rect 16865 11645 16899 11679
rect 16899 11645 16908 11679
rect 16856 11636 16908 11645
rect 19800 11636 19852 11688
rect 22284 11772 22336 11824
rect 22468 11772 22520 11824
rect 23296 11772 23348 11824
rect 23388 11772 23440 11824
rect 26332 11840 26384 11892
rect 27620 11840 27672 11892
rect 28908 11840 28960 11892
rect 26792 11772 26844 11824
rect 28816 11772 28868 11824
rect 20168 11704 20220 11756
rect 23848 11704 23900 11756
rect 25320 11704 25372 11756
rect 27344 11704 27396 11756
rect 28448 11747 28500 11756
rect 28448 11713 28457 11747
rect 28457 11713 28491 11747
rect 28491 11713 28500 11747
rect 28448 11704 28500 11713
rect 14096 11500 14148 11552
rect 14832 11500 14884 11552
rect 18144 11568 18196 11620
rect 19892 11568 19944 11620
rect 21456 11636 21508 11688
rect 22008 11636 22060 11688
rect 23664 11636 23716 11688
rect 23940 11679 23992 11688
rect 23940 11645 23949 11679
rect 23949 11645 23983 11679
rect 23983 11645 23992 11679
rect 23940 11636 23992 11645
rect 24860 11636 24912 11688
rect 27436 11636 27488 11688
rect 27804 11679 27856 11688
rect 27804 11645 27813 11679
rect 27813 11645 27847 11679
rect 27847 11645 27856 11679
rect 27804 11636 27856 11645
rect 31760 11772 31812 11824
rect 32128 11772 32180 11824
rect 34612 11772 34664 11824
rect 37280 11772 37332 11824
rect 30472 11704 30524 11756
rect 31208 11747 31260 11756
rect 31208 11713 31217 11747
rect 31217 11713 31251 11747
rect 31251 11713 31260 11747
rect 31208 11704 31260 11713
rect 34888 11704 34940 11756
rect 36544 11704 36596 11756
rect 36728 11704 36780 11756
rect 38384 11704 38436 11756
rect 39396 11815 39448 11824
rect 39396 11781 39405 11815
rect 39405 11781 39439 11815
rect 39439 11781 39448 11815
rect 39396 11772 39448 11781
rect 40224 11772 40276 11824
rect 49148 11815 49200 11824
rect 49148 11781 49157 11815
rect 49157 11781 49191 11815
rect 49191 11781 49200 11815
rect 49148 11772 49200 11781
rect 31392 11679 31444 11688
rect 31392 11645 31401 11679
rect 31401 11645 31435 11679
rect 31435 11645 31444 11679
rect 31392 11636 31444 11645
rect 31944 11636 31996 11688
rect 18328 11500 18380 11552
rect 20076 11500 20128 11552
rect 20628 11500 20680 11552
rect 22284 11568 22336 11620
rect 21548 11500 21600 11552
rect 22100 11500 22152 11552
rect 22836 11500 22888 11552
rect 23296 11500 23348 11552
rect 28356 11568 28408 11620
rect 32220 11568 32272 11620
rect 32588 11568 32640 11620
rect 33508 11636 33560 11688
rect 34796 11636 34848 11688
rect 45928 11704 45980 11756
rect 32956 11568 33008 11620
rect 33968 11568 34020 11620
rect 27344 11500 27396 11552
rect 29736 11500 29788 11552
rect 35992 11500 36044 11552
rect 36084 11500 36136 11552
rect 37004 11568 37056 11620
rect 44180 11568 44232 11620
rect 46664 11568 46716 11620
rect 38292 11500 38344 11552
rect 2950 11398 3002 11450
rect 3014 11398 3066 11450
rect 3078 11398 3130 11450
rect 3142 11398 3194 11450
rect 3206 11398 3258 11450
rect 12950 11398 13002 11450
rect 13014 11398 13066 11450
rect 13078 11398 13130 11450
rect 13142 11398 13194 11450
rect 13206 11398 13258 11450
rect 22950 11398 23002 11450
rect 23014 11398 23066 11450
rect 23078 11398 23130 11450
rect 23142 11398 23194 11450
rect 23206 11398 23258 11450
rect 32950 11398 33002 11450
rect 33014 11398 33066 11450
rect 33078 11398 33130 11450
rect 33142 11398 33194 11450
rect 33206 11398 33258 11450
rect 42950 11398 43002 11450
rect 43014 11398 43066 11450
rect 43078 11398 43130 11450
rect 43142 11398 43194 11450
rect 43206 11398 43258 11450
rect 12716 11271 12768 11280
rect 12716 11237 12725 11271
rect 12725 11237 12759 11271
rect 12759 11237 12768 11271
rect 12716 11228 12768 11237
rect 13728 11296 13780 11348
rect 16672 11296 16724 11348
rect 13912 11228 13964 11280
rect 16488 11228 16540 11280
rect 13820 11160 13872 11212
rect 14832 11203 14884 11212
rect 14832 11169 14841 11203
rect 14841 11169 14875 11203
rect 14875 11169 14884 11203
rect 14832 11160 14884 11169
rect 15108 11160 15160 11212
rect 15200 11160 15252 11212
rect 19616 11296 19668 11348
rect 20168 11296 20220 11348
rect 18420 11228 18472 11280
rect 19800 11228 19852 11280
rect 21272 11296 21324 11348
rect 23480 11296 23532 11348
rect 26516 11296 26568 11348
rect 27528 11296 27580 11348
rect 29092 11296 29144 11348
rect 29276 11296 29328 11348
rect 32772 11296 32824 11348
rect 1584 11135 1636 11144
rect 1584 11101 1593 11135
rect 1593 11101 1627 11135
rect 1627 11101 1636 11135
rect 1584 11092 1636 11101
rect 14740 11135 14792 11144
rect 14740 11101 14749 11135
rect 14749 11101 14783 11135
rect 14783 11101 14792 11135
rect 14740 11092 14792 11101
rect 16764 11092 16816 11144
rect 16948 11092 17000 11144
rect 18512 11160 18564 11212
rect 18880 11160 18932 11212
rect 21456 11160 21508 11212
rect 23296 11160 23348 11212
rect 23388 11203 23440 11212
rect 23388 11169 23397 11203
rect 23397 11169 23431 11203
rect 23431 11169 23440 11203
rect 23388 11160 23440 11169
rect 23664 11160 23716 11212
rect 24584 11203 24636 11212
rect 24584 11169 24593 11203
rect 24593 11169 24627 11203
rect 24627 11169 24636 11203
rect 24584 11160 24636 11169
rect 24860 11203 24912 11212
rect 24860 11169 24869 11203
rect 24869 11169 24903 11203
rect 24903 11169 24912 11203
rect 24860 11160 24912 11169
rect 27252 11160 27304 11212
rect 17868 11092 17920 11144
rect 19156 11092 19208 11144
rect 21824 11092 21876 11144
rect 12256 11024 12308 11076
rect 18972 11024 19024 11076
rect 23756 11092 23808 11144
rect 26884 11135 26936 11144
rect 26884 11101 26893 11135
rect 26893 11101 26927 11135
rect 26927 11101 26936 11135
rect 26884 11092 26936 11101
rect 12164 10956 12216 11008
rect 13452 10956 13504 11008
rect 18144 10956 18196 11008
rect 18696 10956 18748 11008
rect 23296 11024 23348 11076
rect 25320 11024 25372 11076
rect 28632 11203 28684 11212
rect 28632 11169 28641 11203
rect 28641 11169 28675 11203
rect 28675 11169 28684 11203
rect 28632 11160 28684 11169
rect 28724 11160 28776 11212
rect 32588 11228 32640 11280
rect 33968 11296 34020 11348
rect 31024 11160 31076 11212
rect 29736 11092 29788 11144
rect 36084 11203 36136 11212
rect 36084 11169 36093 11203
rect 36093 11169 36127 11203
rect 36127 11169 36136 11203
rect 36084 11160 36136 11169
rect 42616 11296 42668 11348
rect 42708 11228 42760 11280
rect 31392 11067 31444 11076
rect 31392 11033 31401 11067
rect 31401 11033 31435 11067
rect 31435 11033 31444 11067
rect 31392 11024 31444 11033
rect 31668 11024 31720 11076
rect 32772 11024 32824 11076
rect 33324 11024 33376 11076
rect 34428 11092 34480 11144
rect 34796 11092 34848 11144
rect 33784 11067 33836 11076
rect 33784 11033 33793 11067
rect 33793 11033 33827 11067
rect 33827 11033 33836 11067
rect 33784 11024 33836 11033
rect 35348 11024 35400 11076
rect 36544 11024 36596 11076
rect 28632 10956 28684 11008
rect 30288 10956 30340 11008
rect 31760 10956 31812 11008
rect 35532 10956 35584 11008
rect 36452 10956 36504 11008
rect 37464 11024 37516 11076
rect 40960 11135 41012 11144
rect 40960 11101 40969 11135
rect 40969 11101 41003 11135
rect 41003 11101 41012 11135
rect 40960 11092 41012 11101
rect 49148 11203 49200 11212
rect 49148 11169 49157 11203
rect 49157 11169 49191 11203
rect 49191 11169 49200 11203
rect 49148 11160 49200 11169
rect 45744 11024 45796 11076
rect 46940 11024 46992 11076
rect 7950 10854 8002 10906
rect 8014 10854 8066 10906
rect 8078 10854 8130 10906
rect 8142 10854 8194 10906
rect 8206 10854 8258 10906
rect 17950 10854 18002 10906
rect 18014 10854 18066 10906
rect 18078 10854 18130 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 27950 10854 28002 10906
rect 28014 10854 28066 10906
rect 28078 10854 28130 10906
rect 28142 10854 28194 10906
rect 28206 10854 28258 10906
rect 37950 10854 38002 10906
rect 38014 10854 38066 10906
rect 38078 10854 38130 10906
rect 38142 10854 38194 10906
rect 38206 10854 38258 10906
rect 47950 10854 48002 10906
rect 48014 10854 48066 10906
rect 48078 10854 48130 10906
rect 48142 10854 48194 10906
rect 48206 10854 48258 10906
rect 940 10616 992 10668
rect 16028 10795 16080 10804
rect 16028 10761 16037 10795
rect 16037 10761 16071 10795
rect 16071 10761 16080 10795
rect 16028 10752 16080 10761
rect 18604 10752 18656 10804
rect 18972 10795 19024 10804
rect 18972 10761 18981 10795
rect 18981 10761 19015 10795
rect 19015 10761 19024 10795
rect 18972 10752 19024 10761
rect 19432 10795 19484 10804
rect 19432 10761 19441 10795
rect 19441 10761 19475 10795
rect 19475 10761 19484 10795
rect 19432 10752 19484 10761
rect 20536 10752 20588 10804
rect 20720 10752 20772 10804
rect 19524 10684 19576 10736
rect 21732 10684 21784 10736
rect 24216 10795 24268 10804
rect 24216 10761 24225 10795
rect 24225 10761 24259 10795
rect 24259 10761 24268 10795
rect 24216 10752 24268 10761
rect 31760 10752 31812 10804
rect 31944 10752 31996 10804
rect 34244 10752 34296 10804
rect 28908 10684 28960 10736
rect 1216 10548 1268 10600
rect 13452 10616 13504 10668
rect 14372 10616 14424 10668
rect 14464 10616 14516 10668
rect 16212 10616 16264 10668
rect 16948 10616 17000 10668
rect 19156 10616 19208 10668
rect 19340 10659 19392 10668
rect 19340 10625 19349 10659
rect 19349 10625 19383 10659
rect 19383 10625 19392 10659
rect 19340 10616 19392 10625
rect 12808 10548 12860 10600
rect 13728 10591 13780 10600
rect 13728 10557 13737 10591
rect 13737 10557 13771 10591
rect 13771 10557 13780 10591
rect 13728 10548 13780 10557
rect 14924 10591 14976 10600
rect 14924 10557 14933 10591
rect 14933 10557 14967 10591
rect 14967 10557 14976 10591
rect 14924 10548 14976 10557
rect 15292 10548 15344 10600
rect 12072 10480 12124 10532
rect 11888 10412 11940 10464
rect 15660 10480 15712 10532
rect 15936 10480 15988 10532
rect 18972 10548 19024 10600
rect 23388 10616 23440 10668
rect 27528 10659 27580 10668
rect 27528 10625 27537 10659
rect 27537 10625 27571 10659
rect 27571 10625 27580 10659
rect 27528 10616 27580 10625
rect 19708 10548 19760 10600
rect 22008 10591 22060 10600
rect 22008 10557 22017 10591
rect 22017 10557 22051 10591
rect 22051 10557 22060 10591
rect 22008 10548 22060 10557
rect 24676 10591 24728 10600
rect 24676 10557 24685 10591
rect 24685 10557 24719 10591
rect 24719 10557 24728 10591
rect 24676 10548 24728 10557
rect 24860 10591 24912 10600
rect 24860 10557 24869 10591
rect 24869 10557 24903 10591
rect 24903 10557 24912 10591
rect 24860 10548 24912 10557
rect 26516 10548 26568 10600
rect 30288 10684 30340 10736
rect 30380 10684 30432 10736
rect 29920 10616 29972 10668
rect 31116 10684 31168 10736
rect 32036 10684 32088 10736
rect 32772 10684 32824 10736
rect 34888 10752 34940 10804
rect 35072 10752 35124 10804
rect 35348 10684 35400 10736
rect 37004 10752 37056 10804
rect 37280 10684 37332 10736
rect 15568 10455 15620 10464
rect 15568 10421 15577 10455
rect 15577 10421 15611 10455
rect 15611 10421 15620 10455
rect 15568 10412 15620 10421
rect 17684 10412 17736 10464
rect 23756 10523 23808 10532
rect 23756 10489 23765 10523
rect 23765 10489 23799 10523
rect 23799 10489 23808 10523
rect 23756 10480 23808 10489
rect 24768 10480 24820 10532
rect 25596 10480 25648 10532
rect 29736 10548 29788 10600
rect 30380 10548 30432 10600
rect 35808 10616 35860 10668
rect 31760 10548 31812 10600
rect 32956 10591 33008 10600
rect 32956 10557 32965 10591
rect 32965 10557 32999 10591
rect 32999 10557 33008 10591
rect 32956 10548 33008 10557
rect 33508 10548 33560 10600
rect 28540 10480 28592 10532
rect 31208 10480 31260 10532
rect 19064 10412 19116 10464
rect 28448 10412 28500 10464
rect 31944 10480 31996 10532
rect 36268 10548 36320 10600
rect 36452 10659 36504 10668
rect 36452 10625 36461 10659
rect 36461 10625 36495 10659
rect 36495 10625 36504 10659
rect 36452 10616 36504 10625
rect 36544 10659 36596 10668
rect 36544 10625 36553 10659
rect 36553 10625 36587 10659
rect 36587 10625 36596 10659
rect 36544 10616 36596 10625
rect 37648 10548 37700 10600
rect 49240 10684 49292 10736
rect 39764 10659 39816 10668
rect 39764 10625 39773 10659
rect 39773 10625 39807 10659
rect 39807 10625 39816 10659
rect 39764 10616 39816 10625
rect 46940 10616 46992 10668
rect 32680 10412 32732 10464
rect 43720 10480 43772 10532
rect 35532 10455 35584 10464
rect 35532 10421 35541 10455
rect 35541 10421 35575 10455
rect 35575 10421 35584 10455
rect 35532 10412 35584 10421
rect 37832 10412 37884 10464
rect 2950 10310 3002 10362
rect 3014 10310 3066 10362
rect 3078 10310 3130 10362
rect 3142 10310 3194 10362
rect 3206 10310 3258 10362
rect 12950 10310 13002 10362
rect 13014 10310 13066 10362
rect 13078 10310 13130 10362
rect 13142 10310 13194 10362
rect 13206 10310 13258 10362
rect 22950 10310 23002 10362
rect 23014 10310 23066 10362
rect 23078 10310 23130 10362
rect 23142 10310 23194 10362
rect 23206 10310 23258 10362
rect 32950 10310 33002 10362
rect 33014 10310 33066 10362
rect 33078 10310 33130 10362
rect 33142 10310 33194 10362
rect 33206 10310 33258 10362
rect 42950 10310 43002 10362
rect 43014 10310 43066 10362
rect 43078 10310 43130 10362
rect 43142 10310 43194 10362
rect 43206 10310 43258 10362
rect 12532 10208 12584 10260
rect 13636 10208 13688 10260
rect 17960 10208 18012 10260
rect 12440 10140 12492 10192
rect 11888 10072 11940 10124
rect 12072 10115 12124 10124
rect 12072 10081 12081 10115
rect 12081 10081 12115 10115
rect 12115 10081 12124 10115
rect 12072 10072 12124 10081
rect 12164 10115 12216 10124
rect 12164 10081 12173 10115
rect 12173 10081 12207 10115
rect 12207 10081 12216 10115
rect 12164 10072 12216 10081
rect 13360 10115 13412 10124
rect 13360 10081 13369 10115
rect 13369 10081 13403 10115
rect 13403 10081 13412 10115
rect 13360 10072 13412 10081
rect 16120 10072 16172 10124
rect 940 10004 992 10056
rect 11980 10047 12032 10056
rect 11980 10013 11989 10047
rect 11989 10013 12023 10047
rect 12023 10013 12032 10047
rect 11980 10004 12032 10013
rect 13268 10047 13320 10056
rect 13268 10013 13277 10047
rect 13277 10013 13311 10047
rect 13311 10013 13320 10047
rect 13268 10004 13320 10013
rect 13820 10004 13872 10056
rect 16396 10004 16448 10056
rect 16580 10004 16632 10056
rect 17684 10072 17736 10124
rect 19248 10208 19300 10260
rect 13452 9936 13504 9988
rect 14556 9979 14608 9988
rect 14556 9945 14565 9979
rect 14565 9945 14599 9979
rect 14599 9945 14608 9979
rect 14556 9936 14608 9945
rect 16120 9936 16172 9988
rect 16212 9936 16264 9988
rect 15936 9868 15988 9920
rect 16948 9911 17000 9920
rect 16948 9877 16957 9911
rect 16957 9877 16991 9911
rect 16991 9877 17000 9911
rect 16948 9868 17000 9877
rect 17960 9868 18012 9920
rect 19064 10004 19116 10056
rect 20996 10208 21048 10260
rect 21732 10208 21784 10260
rect 23296 10208 23348 10260
rect 24676 10208 24728 10260
rect 29092 10208 29144 10260
rect 30196 10208 30248 10260
rect 30472 10208 30524 10260
rect 31392 10208 31444 10260
rect 34888 10208 34940 10260
rect 31668 10140 31720 10192
rect 32680 10140 32732 10192
rect 32772 10140 32824 10192
rect 40960 10208 41012 10260
rect 20260 10115 20312 10124
rect 20260 10081 20269 10115
rect 20269 10081 20303 10115
rect 20303 10081 20312 10115
rect 20260 10072 20312 10081
rect 22008 10072 22060 10124
rect 30748 10072 30800 10124
rect 31208 10072 31260 10124
rect 32220 10072 32272 10124
rect 32404 10072 32456 10124
rect 33508 10072 33560 10124
rect 37740 10072 37792 10124
rect 22468 10047 22520 10056
rect 22468 10013 22477 10047
rect 22477 10013 22511 10047
rect 22511 10013 22520 10047
rect 22468 10004 22520 10013
rect 26976 10047 27028 10056
rect 26976 10013 26985 10047
rect 26985 10013 27019 10047
rect 27019 10013 27028 10047
rect 26976 10004 27028 10013
rect 20812 9936 20864 9988
rect 21824 9936 21876 9988
rect 23388 9936 23440 9988
rect 24860 9979 24912 9988
rect 24860 9945 24869 9979
rect 24869 9945 24903 9979
rect 24903 9945 24912 9979
rect 24860 9936 24912 9945
rect 25320 9936 25372 9988
rect 26884 9936 26936 9988
rect 27344 9936 27396 9988
rect 28632 9936 28684 9988
rect 28908 9936 28960 9988
rect 33416 10004 33468 10056
rect 37832 10047 37884 10056
rect 37832 10013 37841 10047
rect 37841 10013 37875 10047
rect 37875 10013 37884 10047
rect 37832 10004 37884 10013
rect 30564 9936 30616 9988
rect 30656 9979 30708 9988
rect 30656 9945 30665 9979
rect 30665 9945 30699 9979
rect 30699 9945 30708 9979
rect 30656 9936 30708 9945
rect 32036 9936 32088 9988
rect 23572 9868 23624 9920
rect 28540 9868 28592 9920
rect 31392 9868 31444 9920
rect 34336 9936 34388 9988
rect 35072 9936 35124 9988
rect 35440 9936 35492 9988
rect 35624 9936 35676 9988
rect 38752 9979 38804 9988
rect 38752 9945 38761 9979
rect 38761 9945 38795 9979
rect 38795 9945 38804 9979
rect 38752 9936 38804 9945
rect 40132 9979 40184 9988
rect 40132 9945 40141 9979
rect 40141 9945 40175 9979
rect 40175 9945 40184 9979
rect 40132 9936 40184 9945
rect 32680 9868 32732 9920
rect 34520 9868 34572 9920
rect 49148 10115 49200 10124
rect 49148 10081 49157 10115
rect 49157 10081 49191 10115
rect 49191 10081 49200 10115
rect 49148 10072 49200 10081
rect 42616 10004 42668 10056
rect 45744 10004 45796 10056
rect 46664 10004 46716 10056
rect 42708 9936 42760 9988
rect 46756 9936 46808 9988
rect 47308 9979 47360 9988
rect 47308 9945 47317 9979
rect 47317 9945 47351 9979
rect 47351 9945 47360 9979
rect 47308 9936 47360 9945
rect 42800 9868 42852 9920
rect 7950 9766 8002 9818
rect 8014 9766 8066 9818
rect 8078 9766 8130 9818
rect 8142 9766 8194 9818
rect 8206 9766 8258 9818
rect 17950 9766 18002 9818
rect 18014 9766 18066 9818
rect 18078 9766 18130 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 27950 9766 28002 9818
rect 28014 9766 28066 9818
rect 28078 9766 28130 9818
rect 28142 9766 28194 9818
rect 28206 9766 28258 9818
rect 37950 9766 38002 9818
rect 38014 9766 38066 9818
rect 38078 9766 38130 9818
rect 38142 9766 38194 9818
rect 38206 9766 38258 9818
rect 47950 9766 48002 9818
rect 48014 9766 48066 9818
rect 48078 9766 48130 9818
rect 48142 9766 48194 9818
rect 48206 9766 48258 9818
rect 16120 9664 16172 9716
rect 12440 9639 12492 9648
rect 12440 9605 12449 9639
rect 12449 9605 12483 9639
rect 12483 9605 12492 9639
rect 12440 9596 12492 9605
rect 12624 9596 12676 9648
rect 940 9528 992 9580
rect 13820 9596 13872 9648
rect 15016 9596 15068 9648
rect 16672 9596 16724 9648
rect 12716 9503 12768 9512
rect 12716 9469 12725 9503
rect 12725 9469 12759 9503
rect 12759 9469 12768 9503
rect 12716 9460 12768 9469
rect 15200 9460 15252 9512
rect 1768 9435 1820 9444
rect 1768 9401 1777 9435
rect 1777 9401 1811 9435
rect 1811 9401 1820 9435
rect 1768 9392 1820 9401
rect 12808 9392 12860 9444
rect 12164 9324 12216 9376
rect 25596 9664 25648 9716
rect 18880 9639 18932 9648
rect 18880 9605 18889 9639
rect 18889 9605 18923 9639
rect 18923 9605 18932 9639
rect 18880 9596 18932 9605
rect 19616 9639 19668 9648
rect 19616 9605 19625 9639
rect 19625 9605 19659 9639
rect 19659 9605 19668 9639
rect 19616 9596 19668 9605
rect 21088 9596 21140 9648
rect 22560 9596 22612 9648
rect 23572 9596 23624 9648
rect 29276 9707 29328 9716
rect 29276 9673 29285 9707
rect 29285 9673 29319 9707
rect 29319 9673 29328 9707
rect 29276 9664 29328 9673
rect 30380 9664 30432 9716
rect 30656 9664 30708 9716
rect 31300 9664 31352 9716
rect 31392 9664 31444 9716
rect 38752 9664 38804 9716
rect 32036 9596 32088 9648
rect 32220 9596 32272 9648
rect 35624 9596 35676 9648
rect 49332 9596 49384 9648
rect 18236 9528 18288 9580
rect 20996 9528 21048 9580
rect 16856 9503 16908 9512
rect 16856 9469 16865 9503
rect 16865 9469 16899 9503
rect 16899 9469 16908 9503
rect 16856 9460 16908 9469
rect 18604 9460 18656 9512
rect 16856 9324 16908 9376
rect 20812 9460 20864 9512
rect 20904 9324 20956 9376
rect 23664 9571 23716 9580
rect 23664 9537 23673 9571
rect 23673 9537 23707 9571
rect 23707 9537 23716 9571
rect 23664 9528 23716 9537
rect 25044 9528 25096 9580
rect 25320 9528 25372 9580
rect 26056 9571 26108 9580
rect 26056 9537 26065 9571
rect 26065 9537 26099 9571
rect 26099 9537 26108 9571
rect 26056 9528 26108 9537
rect 26148 9571 26200 9580
rect 26148 9537 26157 9571
rect 26157 9537 26191 9571
rect 26191 9537 26200 9571
rect 26148 9528 26200 9537
rect 28908 9528 28960 9580
rect 29644 9528 29696 9580
rect 31300 9528 31352 9580
rect 26884 9460 26936 9512
rect 26976 9460 27028 9512
rect 26792 9392 26844 9444
rect 25412 9367 25464 9376
rect 25412 9333 25421 9367
rect 25421 9333 25455 9367
rect 25455 9333 25464 9367
rect 25412 9324 25464 9333
rect 29736 9503 29788 9512
rect 29736 9469 29745 9503
rect 29745 9469 29779 9503
rect 29779 9469 29788 9503
rect 29736 9460 29788 9469
rect 30012 9503 30064 9512
rect 30012 9469 30021 9503
rect 30021 9469 30055 9503
rect 30055 9469 30064 9503
rect 30012 9460 30064 9469
rect 30104 9460 30156 9512
rect 32312 9460 32364 9512
rect 32496 9528 32548 9580
rect 33508 9528 33560 9580
rect 47032 9528 47084 9580
rect 33692 9460 33744 9512
rect 37464 9460 37516 9512
rect 29736 9324 29788 9376
rect 33876 9392 33928 9444
rect 35164 9392 35216 9444
rect 32404 9324 32456 9376
rect 35532 9324 35584 9376
rect 2950 9222 3002 9274
rect 3014 9222 3066 9274
rect 3078 9222 3130 9274
rect 3142 9222 3194 9274
rect 3206 9222 3258 9274
rect 12950 9222 13002 9274
rect 13014 9222 13066 9274
rect 13078 9222 13130 9274
rect 13142 9222 13194 9274
rect 13206 9222 13258 9274
rect 22950 9222 23002 9274
rect 23014 9222 23066 9274
rect 23078 9222 23130 9274
rect 23142 9222 23194 9274
rect 23206 9222 23258 9274
rect 32950 9222 33002 9274
rect 33014 9222 33066 9274
rect 33078 9222 33130 9274
rect 33142 9222 33194 9274
rect 33206 9222 33258 9274
rect 42950 9222 43002 9274
rect 43014 9222 43066 9274
rect 43078 9222 43130 9274
rect 43142 9222 43194 9274
rect 43206 9222 43258 9274
rect 12164 9120 12216 9172
rect 14372 9163 14424 9172
rect 14372 9129 14381 9163
rect 14381 9129 14415 9163
rect 14415 9129 14424 9163
rect 14372 9120 14424 9129
rect 15108 9120 15160 9172
rect 17040 9120 17092 9172
rect 17868 9120 17920 9172
rect 18972 9120 19024 9172
rect 22284 9120 22336 9172
rect 27068 9120 27120 9172
rect 27712 9120 27764 9172
rect 32680 9120 32732 9172
rect 37280 9120 37332 9172
rect 14556 9052 14608 9104
rect 14832 9027 14884 9036
rect 14832 8993 14841 9027
rect 14841 8993 14875 9027
rect 14875 8993 14884 9027
rect 14832 8984 14884 8993
rect 23848 9052 23900 9104
rect 26148 9052 26200 9104
rect 30104 9052 30156 9104
rect 32312 9052 32364 9104
rect 34980 9052 35032 9104
rect 35624 9052 35676 9104
rect 18512 8984 18564 9036
rect 20996 8984 21048 9036
rect 22008 8984 22060 9036
rect 25412 8984 25464 9036
rect 30012 8984 30064 9036
rect 940 8916 992 8968
rect 1216 8848 1268 8900
rect 13544 8916 13596 8968
rect 13820 8916 13872 8968
rect 16212 8848 16264 8900
rect 14556 8780 14608 8832
rect 14740 8823 14792 8832
rect 14740 8789 14749 8823
rect 14749 8789 14783 8823
rect 14783 8789 14792 8823
rect 14740 8780 14792 8789
rect 15108 8780 15160 8832
rect 19432 8959 19484 8968
rect 19432 8925 19441 8959
rect 19441 8925 19475 8959
rect 19475 8925 19484 8959
rect 19432 8916 19484 8925
rect 22192 8916 22244 8968
rect 30748 8959 30800 8968
rect 30748 8925 30757 8959
rect 30757 8925 30791 8959
rect 30791 8925 30800 8959
rect 30748 8916 30800 8925
rect 32036 8916 32088 8968
rect 33600 8916 33652 8968
rect 33876 9027 33928 9036
rect 33876 8993 33885 9027
rect 33885 8993 33919 9027
rect 33919 8993 33928 9027
rect 33876 8984 33928 8993
rect 34428 8984 34480 9036
rect 34060 8916 34112 8968
rect 35532 8984 35584 9036
rect 16580 8891 16632 8900
rect 16580 8857 16589 8891
rect 16589 8857 16623 8891
rect 16623 8857 16632 8891
rect 16580 8848 16632 8857
rect 16672 8848 16724 8900
rect 16856 8780 16908 8832
rect 18236 8848 18288 8900
rect 18420 8848 18472 8900
rect 19708 8891 19760 8900
rect 19708 8857 19717 8891
rect 19717 8857 19751 8891
rect 19751 8857 19760 8891
rect 19708 8848 19760 8857
rect 21088 8848 21140 8900
rect 23296 8848 23348 8900
rect 25136 8848 25188 8900
rect 32864 8848 32916 8900
rect 19616 8780 19668 8832
rect 24952 8823 25004 8832
rect 24952 8789 24961 8823
rect 24961 8789 24995 8823
rect 24995 8789 25004 8823
rect 24952 8780 25004 8789
rect 27620 8823 27672 8832
rect 27620 8789 27629 8823
rect 27629 8789 27663 8823
rect 27663 8789 27672 8823
rect 28632 8823 28684 8832
rect 27620 8780 27672 8789
rect 28632 8789 28641 8823
rect 28641 8789 28675 8823
rect 28675 8789 28684 8823
rect 28632 8780 28684 8789
rect 30012 8780 30064 8832
rect 33784 8823 33836 8832
rect 33784 8789 33793 8823
rect 33793 8789 33827 8823
rect 33827 8789 33836 8823
rect 33784 8780 33836 8789
rect 34888 8823 34940 8832
rect 34888 8789 34897 8823
rect 34897 8789 34931 8823
rect 34931 8789 34940 8823
rect 34888 8780 34940 8789
rect 35256 8823 35308 8832
rect 35256 8789 35265 8823
rect 35265 8789 35299 8823
rect 35299 8789 35308 8823
rect 35256 8780 35308 8789
rect 35624 8780 35676 8832
rect 49240 8984 49292 9036
rect 43628 8916 43680 8968
rect 44180 8916 44232 8968
rect 46572 8848 46624 8900
rect 44272 8780 44324 8832
rect 7950 8678 8002 8730
rect 8014 8678 8066 8730
rect 8078 8678 8130 8730
rect 8142 8678 8194 8730
rect 8206 8678 8258 8730
rect 17950 8678 18002 8730
rect 18014 8678 18066 8730
rect 18078 8678 18130 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 27950 8678 28002 8730
rect 28014 8678 28066 8730
rect 28078 8678 28130 8730
rect 28142 8678 28194 8730
rect 28206 8678 28258 8730
rect 37950 8678 38002 8730
rect 38014 8678 38066 8730
rect 38078 8678 38130 8730
rect 38142 8678 38194 8730
rect 38206 8678 38258 8730
rect 47950 8678 48002 8730
rect 48014 8678 48066 8730
rect 48078 8678 48130 8730
rect 48142 8678 48194 8730
rect 48206 8678 48258 8730
rect 14648 8576 14700 8628
rect 1860 8483 1912 8492
rect 1860 8449 1869 8483
rect 1869 8449 1903 8483
rect 1903 8449 1912 8483
rect 1860 8440 1912 8449
rect 13820 8508 13872 8560
rect 15292 8619 15344 8628
rect 15292 8585 15301 8619
rect 15301 8585 15335 8619
rect 15335 8585 15344 8619
rect 15292 8576 15344 8585
rect 18512 8576 18564 8628
rect 18604 8619 18656 8628
rect 18604 8585 18613 8619
rect 18613 8585 18647 8619
rect 18647 8585 18656 8619
rect 18604 8576 18656 8585
rect 19984 8576 20036 8628
rect 30656 8576 30708 8628
rect 31668 8576 31720 8628
rect 16672 8440 16724 8492
rect 16856 8483 16908 8492
rect 16856 8449 16865 8483
rect 16865 8449 16899 8483
rect 16899 8449 16908 8483
rect 16856 8440 16908 8449
rect 1584 8415 1636 8424
rect 1584 8381 1593 8415
rect 1593 8381 1627 8415
rect 1627 8381 1636 8415
rect 1584 8372 1636 8381
rect 14556 8372 14608 8424
rect 16396 8372 16448 8424
rect 17868 8372 17920 8424
rect 13544 8304 13596 8356
rect 19156 8440 19208 8492
rect 19432 8440 19484 8492
rect 20260 8508 20312 8560
rect 22284 8551 22336 8560
rect 22284 8517 22293 8551
rect 22293 8517 22327 8551
rect 22327 8517 22336 8551
rect 22284 8508 22336 8517
rect 29092 8551 29144 8560
rect 29092 8517 29101 8551
rect 29101 8517 29135 8551
rect 29135 8517 29144 8551
rect 29092 8508 29144 8517
rect 29644 8508 29696 8560
rect 30748 8508 30800 8560
rect 21088 8440 21140 8492
rect 22008 8483 22060 8492
rect 22008 8449 22017 8483
rect 22017 8449 22051 8483
rect 22051 8449 22060 8483
rect 22008 8440 22060 8449
rect 23388 8440 23440 8492
rect 25044 8440 25096 8492
rect 31392 8483 31444 8492
rect 31392 8449 31401 8483
rect 31401 8449 31435 8483
rect 31435 8449 31444 8483
rect 31392 8440 31444 8449
rect 33508 8576 33560 8628
rect 34060 8619 34112 8628
rect 34060 8585 34069 8619
rect 34069 8585 34103 8619
rect 34103 8585 34112 8619
rect 34060 8576 34112 8585
rect 40224 8576 40276 8628
rect 47676 8576 47728 8628
rect 32588 8551 32640 8560
rect 32588 8517 32597 8551
rect 32597 8517 32631 8551
rect 32631 8517 32640 8551
rect 32588 8508 32640 8517
rect 34520 8508 34572 8560
rect 34888 8508 34940 8560
rect 34336 8440 34388 8492
rect 44272 8551 44324 8560
rect 44272 8517 44281 8551
rect 44281 8517 44315 8551
rect 44315 8517 44324 8551
rect 44272 8508 44324 8517
rect 49148 8551 49200 8560
rect 49148 8517 49157 8551
rect 49157 8517 49191 8551
rect 49191 8517 49200 8551
rect 49148 8508 49200 8517
rect 18420 8304 18472 8356
rect 21088 8236 21140 8288
rect 28816 8415 28868 8424
rect 28816 8381 28825 8415
rect 28825 8381 28859 8415
rect 28859 8381 28868 8415
rect 28816 8372 28868 8381
rect 29736 8372 29788 8424
rect 22652 8236 22704 8288
rect 33876 8372 33928 8424
rect 34704 8372 34756 8424
rect 35532 8372 35584 8424
rect 42708 8440 42760 8492
rect 46756 8440 46808 8492
rect 46848 8415 46900 8424
rect 46848 8381 46857 8415
rect 46857 8381 46891 8415
rect 46891 8381 46900 8415
rect 46848 8372 46900 8381
rect 40132 8304 40184 8356
rect 47860 8304 47912 8356
rect 31484 8236 31536 8288
rect 38476 8236 38528 8288
rect 2950 8134 3002 8186
rect 3014 8134 3066 8186
rect 3078 8134 3130 8186
rect 3142 8134 3194 8186
rect 3206 8134 3258 8186
rect 12950 8134 13002 8186
rect 13014 8134 13066 8186
rect 13078 8134 13130 8186
rect 13142 8134 13194 8186
rect 13206 8134 13258 8186
rect 22950 8134 23002 8186
rect 23014 8134 23066 8186
rect 23078 8134 23130 8186
rect 23142 8134 23194 8186
rect 23206 8134 23258 8186
rect 32950 8134 33002 8186
rect 33014 8134 33066 8186
rect 33078 8134 33130 8186
rect 33142 8134 33194 8186
rect 33206 8134 33258 8186
rect 42950 8134 43002 8186
rect 43014 8134 43066 8186
rect 43078 8134 43130 8186
rect 43142 8134 43194 8186
rect 43206 8134 43258 8186
rect 19708 8032 19760 8084
rect 21916 8032 21968 8084
rect 29920 8075 29972 8084
rect 29920 8041 29929 8075
rect 29929 8041 29963 8075
rect 29963 8041 29972 8075
rect 29920 8032 29972 8041
rect 35256 8032 35308 8084
rect 19248 7964 19300 8016
rect 38384 7964 38436 8016
rect 16488 7896 16540 7948
rect 18604 7896 18656 7948
rect 19432 7939 19484 7948
rect 19432 7905 19441 7939
rect 19441 7905 19475 7939
rect 19475 7905 19484 7939
rect 19432 7896 19484 7905
rect 23756 7896 23808 7948
rect 32588 7896 32640 7948
rect 35808 7896 35860 7948
rect 49240 7896 49292 7948
rect 940 7828 992 7880
rect 12808 7828 12860 7880
rect 18328 7828 18380 7880
rect 22192 7828 22244 7880
rect 30564 7828 30616 7880
rect 31760 7828 31812 7880
rect 31852 7871 31904 7880
rect 31852 7837 31861 7871
rect 31861 7837 31895 7871
rect 31895 7837 31904 7871
rect 31852 7828 31904 7837
rect 32772 7828 32824 7880
rect 38752 7871 38804 7880
rect 38752 7837 38761 7871
rect 38761 7837 38795 7871
rect 38795 7837 38804 7871
rect 38752 7828 38804 7837
rect 43720 7828 43772 7880
rect 15476 7760 15528 7812
rect 18972 7760 19024 7812
rect 19984 7760 20036 7812
rect 21088 7760 21140 7812
rect 21824 7760 21876 7812
rect 27712 7760 27764 7812
rect 40040 7760 40092 7812
rect 22744 7692 22796 7744
rect 26056 7692 26108 7744
rect 32680 7735 32732 7744
rect 32680 7701 32689 7735
rect 32689 7701 32723 7735
rect 32723 7701 32732 7735
rect 32680 7692 32732 7701
rect 32772 7735 32824 7744
rect 32772 7701 32781 7735
rect 32781 7701 32815 7735
rect 32815 7701 32824 7735
rect 32772 7692 32824 7701
rect 38660 7692 38712 7744
rect 7950 7590 8002 7642
rect 8014 7590 8066 7642
rect 8078 7590 8130 7642
rect 8142 7590 8194 7642
rect 8206 7590 8258 7642
rect 17950 7590 18002 7642
rect 18014 7590 18066 7642
rect 18078 7590 18130 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 27950 7590 28002 7642
rect 28014 7590 28066 7642
rect 28078 7590 28130 7642
rect 28142 7590 28194 7642
rect 28206 7590 28258 7642
rect 37950 7590 38002 7642
rect 38014 7590 38066 7642
rect 38078 7590 38130 7642
rect 38142 7590 38194 7642
rect 38206 7590 38258 7642
rect 47950 7590 48002 7642
rect 48014 7590 48066 7642
rect 48078 7590 48130 7642
rect 48142 7590 48194 7642
rect 48206 7590 48258 7642
rect 21180 7488 21232 7540
rect 22376 7488 22428 7540
rect 18788 7420 18840 7472
rect 940 7352 992 7404
rect 15568 7352 15620 7404
rect 16948 7284 17000 7336
rect 31484 7488 31536 7540
rect 24952 7420 25004 7472
rect 31852 7488 31904 7540
rect 38660 7488 38712 7540
rect 47584 7488 47636 7540
rect 31392 7352 31444 7404
rect 40132 7420 40184 7472
rect 49332 7420 49384 7472
rect 22652 7327 22704 7336
rect 22652 7293 22661 7327
rect 22661 7293 22695 7327
rect 22695 7293 22704 7327
rect 22652 7284 22704 7293
rect 27804 7284 27856 7336
rect 34244 7352 34296 7404
rect 42800 7352 42852 7404
rect 31760 7284 31812 7336
rect 35532 7284 35584 7336
rect 45744 7216 45796 7268
rect 20444 7148 20496 7200
rect 37924 7191 37976 7200
rect 37924 7157 37933 7191
rect 37933 7157 37967 7191
rect 37967 7157 37976 7191
rect 37924 7148 37976 7157
rect 47768 7148 47820 7200
rect 2950 7046 3002 7098
rect 3014 7046 3066 7098
rect 3078 7046 3130 7098
rect 3142 7046 3194 7098
rect 3206 7046 3258 7098
rect 12950 7046 13002 7098
rect 13014 7046 13066 7098
rect 13078 7046 13130 7098
rect 13142 7046 13194 7098
rect 13206 7046 13258 7098
rect 22950 7046 23002 7098
rect 23014 7046 23066 7098
rect 23078 7046 23130 7098
rect 23142 7046 23194 7098
rect 23206 7046 23258 7098
rect 32950 7046 33002 7098
rect 33014 7046 33066 7098
rect 33078 7046 33130 7098
rect 33142 7046 33194 7098
rect 33206 7046 33258 7098
rect 42950 7046 43002 7098
rect 43014 7046 43066 7098
rect 43078 7046 43130 7098
rect 43142 7046 43194 7098
rect 43206 7046 43258 7098
rect 37924 6876 37976 6928
rect 46940 6876 46992 6928
rect 32772 6808 32824 6860
rect 37740 6808 37792 6860
rect 49148 6851 49200 6860
rect 49148 6817 49157 6851
rect 49157 6817 49191 6851
rect 49191 6817 49200 6851
rect 49148 6808 49200 6817
rect 940 6740 992 6792
rect 1308 6672 1360 6724
rect 19248 6740 19300 6792
rect 40040 6740 40092 6792
rect 47860 6740 47912 6792
rect 27620 6672 27672 6724
rect 48872 6672 48924 6724
rect 2320 6647 2372 6656
rect 2320 6613 2329 6647
rect 2329 6613 2363 6647
rect 2363 6613 2372 6647
rect 2320 6604 2372 6613
rect 21916 6604 21968 6656
rect 7950 6502 8002 6554
rect 8014 6502 8066 6554
rect 8078 6502 8130 6554
rect 8142 6502 8194 6554
rect 8206 6502 8258 6554
rect 17950 6502 18002 6554
rect 18014 6502 18066 6554
rect 18078 6502 18130 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 27950 6502 28002 6554
rect 28014 6502 28066 6554
rect 28078 6502 28130 6554
rect 28142 6502 28194 6554
rect 28206 6502 28258 6554
rect 37950 6502 38002 6554
rect 38014 6502 38066 6554
rect 38078 6502 38130 6554
rect 38142 6502 38194 6554
rect 38206 6502 38258 6554
rect 47950 6502 48002 6554
rect 48014 6502 48066 6554
rect 48078 6502 48130 6554
rect 48142 6502 48194 6554
rect 48206 6502 48258 6554
rect 30472 6332 30524 6384
rect 40224 6332 40276 6384
rect 49240 6332 49292 6384
rect 940 6264 992 6316
rect 16396 6264 16448 6316
rect 46572 6264 46624 6316
rect 18328 6196 18380 6248
rect 1860 6128 1912 6180
rect 24952 6128 25004 6180
rect 32128 6128 32180 6180
rect 16304 6060 16356 6112
rect 19616 6060 19668 6112
rect 37648 6103 37700 6112
rect 37648 6069 37657 6103
rect 37657 6069 37691 6103
rect 37691 6069 37700 6103
rect 37648 6060 37700 6069
rect 47032 6128 47084 6180
rect 45560 6060 45612 6112
rect 2950 5958 3002 6010
rect 3014 5958 3066 6010
rect 3078 5958 3130 6010
rect 3142 5958 3194 6010
rect 3206 5958 3258 6010
rect 12950 5958 13002 6010
rect 13014 5958 13066 6010
rect 13078 5958 13130 6010
rect 13142 5958 13194 6010
rect 13206 5958 13258 6010
rect 22950 5958 23002 6010
rect 23014 5958 23066 6010
rect 23078 5958 23130 6010
rect 23142 5958 23194 6010
rect 23206 5958 23258 6010
rect 32950 5958 33002 6010
rect 33014 5958 33066 6010
rect 33078 5958 33130 6010
rect 33142 5958 33194 6010
rect 33206 5958 33258 6010
rect 42950 5958 43002 6010
rect 43014 5958 43066 6010
rect 43078 5958 43130 6010
rect 43142 5958 43194 6010
rect 43206 5958 43258 6010
rect 37648 5856 37700 5908
rect 47216 5856 47268 5908
rect 17224 5788 17276 5840
rect 49424 5720 49476 5772
rect 940 5652 992 5704
rect 2320 5695 2372 5704
rect 2320 5661 2329 5695
rect 2329 5661 2363 5695
rect 2363 5661 2372 5695
rect 2320 5652 2372 5661
rect 43720 5695 43772 5704
rect 43720 5661 43729 5695
rect 43729 5661 43763 5695
rect 43763 5661 43772 5695
rect 43720 5652 43772 5661
rect 47676 5652 47728 5704
rect 45836 5584 45888 5636
rect 18696 5516 18748 5568
rect 7950 5414 8002 5466
rect 8014 5414 8066 5466
rect 8078 5414 8130 5466
rect 8142 5414 8194 5466
rect 8206 5414 8258 5466
rect 17950 5414 18002 5466
rect 18014 5414 18066 5466
rect 18078 5414 18130 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 27950 5414 28002 5466
rect 28014 5414 28066 5466
rect 28078 5414 28130 5466
rect 28142 5414 28194 5466
rect 28206 5414 28258 5466
rect 37950 5414 38002 5466
rect 38014 5414 38066 5466
rect 38078 5414 38130 5466
rect 38142 5414 38194 5466
rect 38206 5414 38258 5466
rect 47950 5414 48002 5466
rect 48014 5414 48066 5466
rect 48078 5414 48130 5466
rect 48142 5414 48194 5466
rect 48206 5414 48258 5466
rect 37740 5287 37792 5296
rect 37740 5253 37749 5287
rect 37749 5253 37783 5287
rect 37783 5253 37792 5287
rect 37740 5244 37792 5253
rect 38476 5287 38528 5296
rect 38476 5253 38485 5287
rect 38485 5253 38519 5287
rect 38519 5253 38528 5287
rect 38476 5244 38528 5253
rect 49148 5287 49200 5296
rect 49148 5253 49157 5287
rect 49157 5253 49191 5287
rect 49191 5253 49200 5287
rect 49148 5244 49200 5253
rect 18972 5219 19024 5228
rect 18972 5185 18981 5219
rect 18981 5185 19015 5219
rect 19015 5185 19024 5219
rect 18972 5176 19024 5185
rect 940 5108 992 5160
rect 15752 5108 15804 5160
rect 19156 5151 19208 5160
rect 19156 5117 19165 5151
rect 19165 5117 19199 5151
rect 19199 5117 19208 5151
rect 24032 5176 24084 5228
rect 45744 5176 45796 5228
rect 47768 5176 47820 5228
rect 19156 5108 19208 5117
rect 48320 5108 48372 5160
rect 40040 5040 40092 5092
rect 20812 4972 20864 5024
rect 24308 4972 24360 5024
rect 26792 4972 26844 5024
rect 37280 4972 37332 5024
rect 37832 5015 37884 5024
rect 37832 4981 37841 5015
rect 37841 4981 37875 5015
rect 37875 4981 37884 5015
rect 37832 4972 37884 4981
rect 2950 4870 3002 4922
rect 3014 4870 3066 4922
rect 3078 4870 3130 4922
rect 3142 4870 3194 4922
rect 3206 4870 3258 4922
rect 12950 4870 13002 4922
rect 13014 4870 13066 4922
rect 13078 4870 13130 4922
rect 13142 4870 13194 4922
rect 13206 4870 13258 4922
rect 22950 4870 23002 4922
rect 23014 4870 23066 4922
rect 23078 4870 23130 4922
rect 23142 4870 23194 4922
rect 23206 4870 23258 4922
rect 32950 4870 33002 4922
rect 33014 4870 33066 4922
rect 33078 4870 33130 4922
rect 33142 4870 33194 4922
rect 33206 4870 33258 4922
rect 42950 4870 43002 4922
rect 43014 4870 43066 4922
rect 43078 4870 43130 4922
rect 43142 4870 43194 4922
rect 43206 4870 43258 4922
rect 37832 4768 37884 4820
rect 47124 4768 47176 4820
rect 24676 4700 24728 4752
rect 20444 4675 20496 4684
rect 20444 4641 20453 4675
rect 20453 4641 20487 4675
rect 20487 4641 20496 4675
rect 20444 4632 20496 4641
rect 21916 4675 21968 4684
rect 21916 4641 21925 4675
rect 21925 4641 21959 4675
rect 21959 4641 21968 4675
rect 21916 4632 21968 4641
rect 28724 4700 28776 4752
rect 33784 4700 33836 4752
rect 25596 4675 25648 4684
rect 25596 4641 25605 4675
rect 25605 4641 25639 4675
rect 25639 4641 25648 4675
rect 25596 4632 25648 4641
rect 36544 4632 36596 4684
rect 49424 4632 49476 4684
rect 19524 4564 19576 4616
rect 940 4496 992 4548
rect 22100 4607 22152 4616
rect 22100 4573 22109 4607
rect 22109 4573 22143 4607
rect 22143 4573 22152 4607
rect 22100 4564 22152 4573
rect 23664 4564 23716 4616
rect 27528 4564 27580 4616
rect 47584 4564 47636 4616
rect 37280 4539 37332 4548
rect 37280 4505 37289 4539
rect 37289 4505 37323 4539
rect 37323 4505 37332 4539
rect 37280 4496 37332 4505
rect 39856 4496 39908 4548
rect 21456 4428 21508 4480
rect 26148 4428 26200 4480
rect 44640 4428 44692 4480
rect 47676 4496 47728 4548
rect 49792 4428 49844 4480
rect 7950 4326 8002 4378
rect 8014 4326 8066 4378
rect 8078 4326 8130 4378
rect 8142 4326 8194 4378
rect 8206 4326 8258 4378
rect 17950 4326 18002 4378
rect 18014 4326 18066 4378
rect 18078 4326 18130 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 27950 4326 28002 4378
rect 28014 4326 28066 4378
rect 28078 4326 28130 4378
rect 28142 4326 28194 4378
rect 28206 4326 28258 4378
rect 37950 4326 38002 4378
rect 38014 4326 38066 4378
rect 38078 4326 38130 4378
rect 38142 4326 38194 4378
rect 38206 4326 38258 4378
rect 47950 4326 48002 4378
rect 48014 4326 48066 4378
rect 48078 4326 48130 4378
rect 48142 4326 48194 4378
rect 48206 4326 48258 4378
rect 20720 4224 20772 4276
rect 21640 4224 21692 4276
rect 25596 4224 25648 4276
rect 1676 4199 1728 4208
rect 1676 4165 1685 4199
rect 1685 4165 1719 4199
rect 1719 4165 1728 4199
rect 1676 4156 1728 4165
rect 940 4088 992 4140
rect 18328 4088 18380 4140
rect 22652 4131 22704 4140
rect 22652 4097 22670 4131
rect 22670 4097 22704 4131
rect 22652 4088 22704 4097
rect 1860 4063 1912 4072
rect 1860 4029 1869 4063
rect 1869 4029 1903 4063
rect 1903 4029 1912 4063
rect 1860 4020 1912 4029
rect 22100 4020 22152 4072
rect 24124 4063 24176 4072
rect 24124 4029 24133 4063
rect 24133 4029 24167 4063
rect 24167 4029 24176 4063
rect 24124 4020 24176 4029
rect 24308 4063 24360 4072
rect 24308 4029 24317 4063
rect 24317 4029 24351 4063
rect 24351 4029 24360 4063
rect 24308 4020 24360 4029
rect 24400 4020 24452 4072
rect 16948 3884 17000 3936
rect 24768 3884 24820 3936
rect 36544 4088 36596 4140
rect 46940 4088 46992 4140
rect 49332 4088 49384 4140
rect 27620 4063 27672 4072
rect 27620 4029 27629 4063
rect 27629 4029 27663 4063
rect 27663 4029 27672 4063
rect 27620 4020 27672 4029
rect 46664 4063 46716 4072
rect 46664 4029 46673 4063
rect 46673 4029 46707 4063
rect 46707 4029 46716 4063
rect 46664 4020 46716 4029
rect 34428 3884 34480 3936
rect 2950 3782 3002 3834
rect 3014 3782 3066 3834
rect 3078 3782 3130 3834
rect 3142 3782 3194 3834
rect 3206 3782 3258 3834
rect 12950 3782 13002 3834
rect 13014 3782 13066 3834
rect 13078 3782 13130 3834
rect 13142 3782 13194 3834
rect 13206 3782 13258 3834
rect 22950 3782 23002 3834
rect 23014 3782 23066 3834
rect 23078 3782 23130 3834
rect 23142 3782 23194 3834
rect 23206 3782 23258 3834
rect 32950 3782 33002 3834
rect 33014 3782 33066 3834
rect 33078 3782 33130 3834
rect 33142 3782 33194 3834
rect 33206 3782 33258 3834
rect 42950 3782 43002 3834
rect 43014 3782 43066 3834
rect 43078 3782 43130 3834
rect 43142 3782 43194 3834
rect 43206 3782 43258 3834
rect 25872 3680 25924 3732
rect 36544 3723 36596 3732
rect 36544 3689 36553 3723
rect 36553 3689 36587 3723
rect 36587 3689 36596 3723
rect 36544 3680 36596 3689
rect 45560 3723 45612 3732
rect 45560 3689 45569 3723
rect 45569 3689 45603 3723
rect 45603 3689 45612 3723
rect 45560 3680 45612 3689
rect 3332 3544 3384 3596
rect 20720 3544 20772 3596
rect 940 3476 992 3528
rect 14740 3476 14792 3528
rect 18328 3476 18380 3528
rect 18420 3476 18472 3528
rect 21916 3544 21968 3596
rect 23388 3612 23440 3664
rect 24308 3612 24360 3664
rect 20904 3519 20956 3528
rect 20904 3485 20913 3519
rect 20913 3485 20947 3519
rect 20947 3485 20956 3519
rect 20904 3476 20956 3485
rect 17868 3408 17920 3460
rect 21180 3451 21232 3460
rect 21180 3417 21189 3451
rect 21189 3417 21223 3451
rect 21223 3417 21232 3451
rect 21180 3408 21232 3417
rect 21916 3408 21968 3460
rect 12532 3340 12584 3392
rect 17224 3340 17276 3392
rect 22652 3476 22704 3528
rect 23572 3519 23624 3528
rect 23572 3485 23581 3519
rect 23581 3485 23615 3519
rect 23615 3485 23624 3519
rect 23572 3476 23624 3485
rect 24032 3587 24084 3596
rect 24032 3553 24041 3587
rect 24041 3553 24075 3587
rect 24075 3553 24084 3587
rect 24032 3544 24084 3553
rect 28908 3612 28960 3664
rect 24768 3587 24820 3596
rect 24768 3553 24777 3587
rect 24777 3553 24811 3587
rect 24811 3553 24820 3587
rect 24768 3544 24820 3553
rect 24860 3544 24912 3596
rect 25688 3544 25740 3596
rect 24492 3476 24544 3528
rect 27804 3476 27856 3528
rect 40040 3544 40092 3596
rect 45560 3476 45612 3528
rect 49148 3587 49200 3596
rect 49148 3553 49157 3587
rect 49157 3553 49191 3587
rect 49191 3553 49200 3587
rect 49148 3544 49200 3553
rect 47032 3476 47084 3528
rect 23296 3340 23348 3392
rect 23388 3340 23440 3392
rect 48688 3408 48740 3460
rect 27160 3340 27212 3392
rect 39212 3340 39264 3392
rect 7950 3238 8002 3290
rect 8014 3238 8066 3290
rect 8078 3238 8130 3290
rect 8142 3238 8194 3290
rect 8206 3238 8258 3290
rect 17950 3238 18002 3290
rect 18014 3238 18066 3290
rect 18078 3238 18130 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 27950 3238 28002 3290
rect 28014 3238 28066 3290
rect 28078 3238 28130 3290
rect 28142 3238 28194 3290
rect 28206 3238 28258 3290
rect 37950 3238 38002 3290
rect 38014 3238 38066 3290
rect 38078 3238 38130 3290
rect 38142 3238 38194 3290
rect 38206 3238 38258 3290
rect 47950 3238 48002 3290
rect 48014 3238 48066 3290
rect 48078 3238 48130 3290
rect 48142 3238 48194 3290
rect 48206 3238 48258 3290
rect 7472 3136 7524 3188
rect 17224 3136 17276 3188
rect 18420 3136 18472 3188
rect 23112 3136 23164 3188
rect 940 3000 992 3052
rect 13820 3000 13872 3052
rect 19156 3068 19208 3120
rect 22100 3068 22152 3120
rect 22652 3068 22704 3120
rect 11060 2932 11112 2984
rect 17868 2932 17920 2984
rect 14464 2864 14516 2916
rect 20812 3043 20864 3052
rect 20812 3009 20821 3043
rect 20821 3009 20855 3043
rect 20855 3009 20864 3043
rect 20812 3000 20864 3009
rect 21456 3043 21508 3052
rect 21456 3009 21465 3043
rect 21465 3009 21499 3043
rect 21499 3009 21508 3043
rect 21456 3000 21508 3009
rect 23572 3136 23624 3188
rect 23296 3068 23348 3120
rect 24492 3068 24544 3120
rect 26148 3000 26200 3052
rect 36820 3136 36872 3188
rect 27528 3068 27580 3120
rect 29644 3068 29696 3120
rect 49240 3068 49292 3120
rect 28816 3000 28868 3052
rect 39856 3000 39908 3052
rect 45836 3043 45888 3052
rect 45836 3009 45845 3043
rect 45845 3009 45879 3043
rect 45879 3009 45888 3043
rect 45836 3000 45888 3009
rect 47216 3000 47268 3052
rect 18420 2932 18472 2984
rect 20904 2932 20956 2984
rect 22008 2932 22060 2984
rect 24492 2932 24544 2984
rect 22376 2864 22428 2916
rect 22652 2907 22704 2916
rect 22652 2873 22661 2907
rect 22661 2873 22695 2907
rect 22695 2873 22704 2907
rect 22652 2864 22704 2873
rect 23112 2864 23164 2916
rect 25872 2975 25924 2984
rect 25872 2941 25881 2975
rect 25881 2941 25915 2975
rect 25915 2941 25924 2975
rect 25872 2932 25924 2941
rect 46756 2932 46808 2984
rect 46848 2975 46900 2984
rect 46848 2941 46857 2975
rect 46857 2941 46891 2975
rect 46891 2941 46900 2975
rect 46848 2932 46900 2941
rect 16396 2796 16448 2848
rect 21180 2796 21232 2848
rect 23296 2839 23348 2848
rect 23296 2805 23305 2839
rect 23305 2805 23339 2839
rect 23339 2805 23348 2839
rect 23296 2796 23348 2805
rect 23664 2839 23716 2848
rect 23664 2805 23673 2839
rect 23673 2805 23707 2839
rect 23707 2805 23716 2839
rect 23664 2796 23716 2805
rect 27528 2864 27580 2916
rect 24584 2796 24636 2848
rect 27160 2796 27212 2848
rect 27804 2796 27856 2848
rect 38108 2796 38160 2848
rect 2950 2694 3002 2746
rect 3014 2694 3066 2746
rect 3078 2694 3130 2746
rect 3142 2694 3194 2746
rect 3206 2694 3258 2746
rect 12950 2694 13002 2746
rect 13014 2694 13066 2746
rect 13078 2694 13130 2746
rect 13142 2694 13194 2746
rect 13206 2694 13258 2746
rect 22950 2694 23002 2746
rect 23014 2694 23066 2746
rect 23078 2694 23130 2746
rect 23142 2694 23194 2746
rect 23206 2694 23258 2746
rect 32950 2694 33002 2746
rect 33014 2694 33066 2746
rect 33078 2694 33130 2746
rect 33142 2694 33194 2746
rect 33206 2694 33258 2746
rect 42950 2694 43002 2746
rect 43014 2694 43066 2746
rect 43078 2694 43130 2746
rect 43142 2694 43194 2746
rect 43206 2694 43258 2746
rect 22468 2592 22520 2644
rect 28908 2592 28960 2644
rect 34428 2592 34480 2644
rect 11060 2524 11112 2576
rect 13452 2524 13504 2576
rect 940 2388 992 2440
rect 1216 2320 1268 2372
rect 1308 2252 1360 2304
rect 11704 2456 11756 2508
rect 13820 2456 13872 2508
rect 15936 2456 15988 2508
rect 9588 2388 9640 2440
rect 12532 2388 12584 2440
rect 16396 2388 16448 2440
rect 14648 2320 14700 2372
rect 19524 2388 19576 2440
rect 19616 2431 19668 2440
rect 19616 2397 19625 2431
rect 19625 2397 19659 2431
rect 19659 2397 19668 2431
rect 19616 2388 19668 2397
rect 24124 2524 24176 2576
rect 34336 2524 34388 2576
rect 20168 2456 20220 2508
rect 22284 2456 22336 2508
rect 24400 2456 24452 2508
rect 26516 2456 26568 2508
rect 36820 2456 36872 2508
rect 41328 2456 41380 2508
rect 49148 2499 49200 2508
rect 49148 2465 49157 2499
rect 49157 2465 49191 2499
rect 49191 2465 49200 2499
rect 49148 2456 49200 2465
rect 22376 2431 22428 2440
rect 22376 2397 22385 2431
rect 22385 2397 22419 2431
rect 22419 2397 22428 2431
rect 22376 2388 22428 2397
rect 24584 2431 24636 2440
rect 24584 2397 24593 2431
rect 24593 2397 24627 2431
rect 24627 2397 24636 2431
rect 24584 2388 24636 2397
rect 27160 2431 27212 2440
rect 27160 2397 27169 2431
rect 27169 2397 27203 2431
rect 27203 2397 27212 2431
rect 27160 2388 27212 2397
rect 28632 2388 28684 2440
rect 30748 2388 30800 2440
rect 32864 2388 32916 2440
rect 34980 2388 35032 2440
rect 37096 2388 37148 2440
rect 38108 2388 38160 2440
rect 43444 2388 43496 2440
rect 44640 2388 44692 2440
rect 47124 2388 47176 2440
rect 48504 2320 48556 2372
rect 28724 2252 28776 2304
rect 7950 2150 8002 2202
rect 8014 2150 8066 2202
rect 8078 2150 8130 2202
rect 8142 2150 8194 2202
rect 8206 2150 8258 2202
rect 17950 2150 18002 2202
rect 18014 2150 18066 2202
rect 18078 2150 18130 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
rect 27950 2150 28002 2202
rect 28014 2150 28066 2202
rect 28078 2150 28130 2202
rect 28142 2150 28194 2202
rect 28206 2150 28258 2202
rect 37950 2150 38002 2202
rect 38014 2150 38066 2202
rect 38078 2150 38130 2202
rect 38142 2150 38194 2202
rect 38206 2150 38258 2202
rect 47950 2150 48002 2202
rect 48014 2150 48066 2202
rect 48078 2150 48130 2202
rect 48142 2150 48194 2202
rect 48206 2150 48258 2202
<< metal2 >>
rect 1582 26200 1638 27000
rect 2226 26200 2282 27000
rect 2870 26200 2926 27000
rect 3514 26200 3570 27000
rect 4158 26200 4214 27000
rect 4802 26330 4858 27000
rect 4802 26302 5120 26330
rect 4802 26200 4858 26302
rect 1596 23254 1624 26200
rect 1584 23248 1636 23254
rect 1584 23190 1636 23196
rect 2240 22234 2268 26200
rect 2778 24440 2834 24449
rect 2778 24375 2780 24384
rect 2832 24375 2834 24384
rect 2780 24346 2832 24352
rect 2320 24200 2372 24206
rect 2320 24142 2372 24148
rect 2228 22228 2280 22234
rect 2228 22170 2280 22176
rect 1308 22092 1360 22098
rect 1308 22034 1360 22040
rect 1320 20777 1348 22034
rect 1306 20768 1362 20777
rect 1306 20703 1362 20712
rect 1768 20460 1820 20466
rect 1768 20402 1820 20408
rect 1780 18737 1808 20402
rect 2332 19174 2360 24142
rect 2884 23050 2912 26200
rect 3422 25664 3478 25673
rect 3422 25599 3478 25608
rect 3330 25256 3386 25265
rect 3436 25226 3464 25599
rect 3330 25191 3386 25200
rect 3424 25220 3476 25226
rect 3344 25090 3372 25191
rect 3424 25162 3476 25168
rect 3332 25084 3384 25090
rect 3332 25026 3384 25032
rect 3146 24848 3202 24857
rect 3146 24783 3202 24792
rect 3160 24614 3188 24783
rect 3148 24608 3200 24614
rect 3148 24550 3200 24556
rect 2950 24508 3258 24517
rect 2950 24506 2956 24508
rect 3012 24506 3036 24508
rect 3092 24506 3116 24508
rect 3172 24506 3196 24508
rect 3252 24506 3258 24508
rect 3012 24454 3014 24506
rect 3194 24454 3196 24506
rect 2950 24452 2956 24454
rect 3012 24452 3036 24454
rect 3092 24452 3116 24454
rect 3172 24452 3196 24454
rect 3252 24452 3258 24454
rect 2950 24443 3258 24452
rect 3528 24274 3556 26200
rect 3516 24268 3568 24274
rect 3516 24210 3568 24216
rect 3698 24032 3754 24041
rect 3698 23967 3754 23976
rect 3516 23724 3568 23730
rect 3516 23666 3568 23672
rect 3422 23624 3478 23633
rect 3422 23559 3424 23568
rect 3476 23559 3478 23568
rect 3424 23530 3476 23536
rect 2950 23420 3258 23429
rect 2950 23418 2956 23420
rect 3012 23418 3036 23420
rect 3092 23418 3116 23420
rect 3172 23418 3196 23420
rect 3252 23418 3258 23420
rect 3012 23366 3014 23418
rect 3194 23366 3196 23418
rect 2950 23364 2956 23366
rect 3012 23364 3036 23366
rect 3092 23364 3116 23366
rect 3172 23364 3196 23366
rect 3252 23364 3258 23366
rect 2950 23355 3258 23364
rect 3330 23216 3386 23225
rect 3330 23151 3386 23160
rect 2780 23044 2832 23050
rect 2780 22986 2832 22992
rect 2872 23044 2924 23050
rect 2872 22986 2924 22992
rect 2792 22216 2820 22986
rect 3344 22778 3372 23151
rect 3422 22808 3478 22817
rect 3332 22772 3384 22778
rect 3422 22743 3478 22752
rect 3332 22714 3384 22720
rect 2872 22704 2924 22710
rect 2872 22646 2924 22652
rect 2700 22188 2820 22216
rect 2700 21593 2728 22188
rect 2686 21584 2742 21593
rect 2686 21519 2742 21528
rect 2778 21176 2834 21185
rect 2884 21162 2912 22646
rect 2950 22332 3258 22341
rect 2950 22330 2956 22332
rect 3012 22330 3036 22332
rect 3092 22330 3116 22332
rect 3172 22330 3196 22332
rect 3252 22330 3258 22332
rect 3012 22278 3014 22330
rect 3194 22278 3196 22330
rect 2950 22276 2956 22278
rect 3012 22276 3036 22278
rect 3092 22276 3116 22278
rect 3172 22276 3196 22278
rect 3252 22276 3258 22278
rect 2950 22267 3258 22276
rect 3436 22166 3464 22743
rect 3424 22160 3476 22166
rect 3424 22102 3476 22108
rect 3332 21480 3384 21486
rect 3332 21422 3384 21428
rect 2950 21244 3258 21253
rect 2950 21242 2956 21244
rect 3012 21242 3036 21244
rect 3092 21242 3116 21244
rect 3172 21242 3196 21244
rect 3252 21242 3258 21244
rect 3012 21190 3014 21242
rect 3194 21190 3196 21242
rect 2950 21188 2956 21190
rect 3012 21188 3036 21190
rect 3092 21188 3116 21190
rect 3172 21188 3196 21190
rect 3252 21188 3258 21190
rect 2950 21179 3258 21188
rect 2834 21134 2912 21162
rect 2778 21111 2834 21120
rect 2780 20868 2832 20874
rect 2780 20810 2832 20816
rect 2792 19938 2820 20810
rect 2872 20392 2924 20398
rect 2872 20334 2924 20340
rect 2700 19910 2820 19938
rect 2700 19553 2728 19910
rect 2780 19780 2832 19786
rect 2780 19722 2832 19728
rect 2686 19544 2742 19553
rect 2686 19479 2742 19488
rect 2320 19168 2372 19174
rect 2320 19110 2372 19116
rect 2792 18873 2820 19722
rect 2884 19496 2912 20334
rect 2950 20156 3258 20165
rect 2950 20154 2956 20156
rect 3012 20154 3036 20156
rect 3092 20154 3116 20156
rect 3172 20154 3196 20156
rect 3252 20154 3258 20156
rect 3012 20102 3014 20154
rect 3194 20102 3196 20154
rect 2950 20100 2956 20102
rect 3012 20100 3036 20102
rect 3092 20100 3116 20102
rect 3172 20100 3196 20102
rect 3252 20100 3258 20102
rect 2950 20091 3258 20100
rect 3344 19961 3372 21422
rect 3330 19952 3386 19961
rect 3330 19887 3386 19896
rect 2884 19468 3004 19496
rect 2872 19372 2924 19378
rect 2872 19314 2924 19320
rect 2778 18864 2834 18873
rect 2778 18799 2834 18808
rect 1766 18728 1822 18737
rect 1766 18663 1822 18672
rect 2780 18692 2832 18698
rect 2780 18634 2832 18640
rect 2792 18306 2820 18634
rect 2884 18329 2912 19314
rect 2976 19281 3004 19468
rect 2962 19272 3018 19281
rect 2962 19207 3018 19216
rect 2950 19068 3258 19077
rect 2950 19066 2956 19068
rect 3012 19066 3036 19068
rect 3092 19066 3116 19068
rect 3172 19066 3196 19068
rect 3252 19066 3258 19068
rect 3012 19014 3014 19066
rect 3194 19014 3196 19066
rect 2950 19012 2956 19014
rect 3012 19012 3036 19014
rect 3092 19012 3116 19014
rect 3172 19012 3196 19014
rect 3252 19012 3258 19014
rect 2950 19003 3258 19012
rect 2700 18278 2820 18306
rect 2870 18320 2926 18329
rect 2700 17921 2728 18278
rect 3528 18290 3556 23666
rect 3608 22976 3660 22982
rect 3608 22918 3660 22924
rect 3620 21554 3648 22918
rect 3608 21548 3660 21554
rect 3608 21490 3660 21496
rect 3608 20460 3660 20466
rect 3608 20402 3660 20408
rect 3620 19990 3648 20402
rect 3608 19984 3660 19990
rect 3608 19926 3660 19932
rect 3712 18834 3740 23967
rect 4172 23798 4200 26200
rect 4712 24200 4764 24206
rect 4712 24142 4764 24148
rect 4620 24064 4672 24070
rect 4620 24006 4672 24012
rect 4160 23792 4212 23798
rect 4160 23734 4212 23740
rect 4632 23730 4660 24006
rect 4620 23724 4672 23730
rect 4620 23666 4672 23672
rect 4344 23248 4396 23254
rect 4344 23190 4396 23196
rect 4160 23044 4212 23050
rect 4160 22986 4212 22992
rect 3792 22092 3844 22098
rect 3792 22034 3844 22040
rect 3804 22001 3832 22034
rect 4068 22024 4120 22030
rect 3790 21992 3846 22001
rect 4068 21966 4120 21972
rect 3790 21927 3846 21936
rect 4080 21690 4108 21966
rect 4068 21684 4120 21690
rect 4068 21626 4120 21632
rect 4172 21486 4200 22986
rect 4250 22536 4306 22545
rect 4250 22471 4306 22480
rect 4160 21480 4212 21486
rect 4160 21422 4212 21428
rect 4068 21344 4120 21350
rect 4068 21286 4120 21292
rect 4080 20942 4108 21286
rect 4264 21010 4292 22471
rect 4252 21004 4304 21010
rect 4252 20946 4304 20952
rect 4068 20936 4120 20942
rect 4068 20878 4120 20884
rect 3884 20392 3936 20398
rect 3882 20360 3884 20369
rect 3936 20360 3938 20369
rect 3882 20295 3938 20304
rect 4356 19446 4384 23190
rect 4436 23112 4488 23118
rect 4436 23054 4488 23060
rect 4344 19440 4396 19446
rect 4344 19382 4396 19388
rect 3700 18828 3752 18834
rect 3700 18770 3752 18776
rect 2870 18255 2926 18264
rect 3516 18284 3568 18290
rect 3516 18226 3568 18232
rect 2780 18216 2832 18222
rect 2780 18158 2832 18164
rect 4160 18216 4212 18222
rect 4160 18158 4212 18164
rect 2686 17912 2742 17921
rect 2686 17847 2742 17856
rect 1216 17740 1268 17746
rect 1216 17682 1268 17688
rect 1228 17105 1256 17682
rect 2792 17513 2820 18158
rect 2950 17980 3258 17989
rect 2950 17978 2956 17980
rect 3012 17978 3036 17980
rect 3092 17978 3116 17980
rect 3172 17978 3196 17980
rect 3252 17978 3258 17980
rect 3012 17926 3014 17978
rect 3194 17926 3196 17978
rect 2950 17924 2956 17926
rect 3012 17924 3036 17926
rect 3092 17924 3116 17926
rect 3172 17924 3196 17926
rect 3252 17924 3258 17926
rect 2950 17915 3258 17924
rect 2778 17504 2834 17513
rect 2778 17439 2834 17448
rect 1308 17128 1360 17134
rect 1214 17096 1270 17105
rect 1308 17070 1360 17076
rect 1214 17031 1270 17040
rect 1320 16697 1348 17070
rect 2950 16892 3258 16901
rect 2950 16890 2956 16892
rect 3012 16890 3036 16892
rect 3092 16890 3116 16892
rect 3172 16890 3196 16892
rect 3252 16890 3258 16892
rect 3012 16838 3014 16890
rect 3194 16838 3196 16890
rect 2950 16836 2956 16838
rect 3012 16836 3036 16838
rect 3092 16836 3116 16838
rect 3172 16836 3196 16838
rect 3252 16836 3258 16838
rect 2950 16827 3258 16836
rect 1306 16688 1362 16697
rect 1306 16623 1362 16632
rect 1308 16516 1360 16522
rect 1308 16458 1360 16464
rect 1320 16289 1348 16458
rect 1306 16280 1362 16289
rect 1306 16215 1362 16224
rect 1768 16108 1820 16114
rect 1768 16050 1820 16056
rect 1308 16040 1360 16046
rect 1308 15982 1360 15988
rect 1320 15881 1348 15982
rect 1306 15872 1362 15881
rect 1306 15807 1362 15816
rect 1780 15706 1808 16050
rect 4172 16046 4200 18158
rect 4448 16658 4476 23054
rect 4724 21894 4752 24142
rect 4804 23520 4856 23526
rect 4804 23462 4856 23468
rect 4816 22642 4844 23462
rect 4804 22636 4856 22642
rect 4804 22578 4856 22584
rect 5092 22574 5120 26302
rect 5446 26200 5502 27000
rect 6090 26200 6146 27000
rect 6734 26200 6790 27000
rect 7378 26200 7434 27000
rect 8022 26200 8078 27000
rect 8666 26200 8722 27000
rect 9310 26200 9366 27000
rect 9954 26200 10010 27000
rect 10598 26200 10654 27000
rect 11242 26200 11298 27000
rect 11886 26200 11942 27000
rect 12530 26200 12586 27000
rect 13174 26330 13230 27000
rect 13174 26302 13400 26330
rect 13174 26200 13230 26302
rect 5460 23662 5488 26200
rect 5724 24608 5776 24614
rect 5724 24550 5776 24556
rect 5448 23656 5500 23662
rect 5448 23598 5500 23604
rect 5540 23588 5592 23594
rect 5540 23530 5592 23536
rect 5264 23112 5316 23118
rect 5316 23060 5488 23066
rect 5264 23054 5488 23060
rect 5276 23050 5488 23054
rect 5276 23044 5500 23050
rect 5276 23038 5448 23044
rect 5448 22986 5500 22992
rect 5080 22568 5132 22574
rect 5080 22510 5132 22516
rect 4896 22228 4948 22234
rect 4896 22170 4948 22176
rect 4712 21888 4764 21894
rect 4712 21830 4764 21836
rect 4908 19922 4936 22170
rect 5552 21486 5580 23530
rect 5632 21616 5684 21622
rect 5632 21558 5684 21564
rect 5540 21480 5592 21486
rect 5540 21422 5592 21428
rect 4896 19916 4948 19922
rect 4896 19858 4948 19864
rect 5356 19372 5408 19378
rect 5356 19314 5408 19320
rect 5368 17270 5396 19314
rect 5644 18426 5672 21558
rect 5736 20398 5764 24550
rect 6104 23186 6132 26200
rect 6276 24404 6328 24410
rect 6276 24346 6328 24352
rect 6092 23180 6144 23186
rect 6092 23122 6144 23128
rect 6000 22024 6052 22030
rect 6000 21966 6052 21972
rect 6012 21146 6040 21966
rect 6000 21140 6052 21146
rect 6000 21082 6052 21088
rect 5724 20392 5776 20398
rect 5724 20334 5776 20340
rect 6288 19922 6316 24346
rect 6748 24342 6776 26200
rect 6736 24336 6788 24342
rect 6736 24278 6788 24284
rect 6552 24200 6604 24206
rect 6552 24142 6604 24148
rect 6564 23866 6592 24142
rect 6552 23860 6604 23866
rect 6552 23802 6604 23808
rect 7288 23724 7340 23730
rect 7288 23666 7340 23672
rect 7104 23112 7156 23118
rect 7104 23054 7156 23060
rect 6736 22772 6788 22778
rect 6736 22714 6788 22720
rect 6460 22432 6512 22438
rect 6460 22374 6512 22380
rect 6472 20466 6500 22374
rect 6552 21548 6604 21554
rect 6552 21490 6604 21496
rect 6564 20602 6592 21490
rect 6748 21010 6776 22714
rect 7116 22234 7144 23054
rect 7104 22228 7156 22234
rect 7104 22170 7156 22176
rect 6736 21004 6788 21010
rect 6736 20946 6788 20952
rect 6552 20596 6604 20602
rect 6552 20538 6604 20544
rect 6368 20460 6420 20466
rect 6368 20402 6420 20408
rect 6460 20460 6512 20466
rect 6460 20402 6512 20408
rect 6276 19916 6328 19922
rect 6276 19858 6328 19864
rect 5632 18420 5684 18426
rect 5632 18362 5684 18368
rect 5356 17264 5408 17270
rect 5356 17206 5408 17212
rect 4436 16652 4488 16658
rect 4436 16594 4488 16600
rect 4160 16040 4212 16046
rect 4160 15982 4212 15988
rect 2950 15804 3258 15813
rect 2950 15802 2956 15804
rect 3012 15802 3036 15804
rect 3092 15802 3116 15804
rect 3172 15802 3196 15804
rect 3252 15802 3258 15804
rect 3012 15750 3014 15802
rect 3194 15750 3196 15802
rect 2950 15748 2956 15750
rect 3012 15748 3036 15750
rect 3092 15748 3116 15750
rect 3172 15748 3196 15750
rect 3252 15748 3258 15750
rect 2950 15739 3258 15748
rect 1768 15700 1820 15706
rect 1768 15642 1820 15648
rect 1308 15564 1360 15570
rect 1308 15506 1360 15512
rect 1320 15473 1348 15506
rect 1306 15464 1362 15473
rect 1306 15399 1362 15408
rect 1306 15056 1362 15065
rect 1306 14991 1362 15000
rect 1320 14958 1348 14991
rect 1308 14952 1360 14958
rect 1308 14894 1360 14900
rect 2320 14884 2372 14890
rect 2320 14826 2372 14832
rect 1306 14648 1362 14657
rect 1306 14583 1362 14592
rect 1320 14482 1348 14583
rect 1308 14476 1360 14482
rect 1308 14418 1360 14424
rect 1306 14240 1362 14249
rect 1306 14175 1362 14184
rect 1320 13870 1348 14175
rect 1308 13864 1360 13870
rect 1308 13806 1360 13812
rect 938 13016 994 13025
rect 938 12951 994 12960
rect 952 12918 980 12951
rect 940 12912 992 12918
rect 940 12854 992 12860
rect 1308 12844 1360 12850
rect 1308 12786 1360 12792
rect 1320 12617 1348 12786
rect 1306 12608 1362 12617
rect 1306 12543 1362 12552
rect 940 12232 992 12238
rect 940 12174 992 12180
rect 1030 12200 1086 12209
rect 952 11801 980 12174
rect 1030 12135 1086 12144
rect 938 11792 994 11801
rect 1044 11762 1072 12135
rect 1860 11892 1912 11898
rect 1860 11834 1912 11840
rect 938 11727 994 11736
rect 1032 11756 1084 11762
rect 1032 11698 1084 11704
rect 940 11688 992 11694
rect 940 11630 992 11636
rect 952 11393 980 11630
rect 938 11384 994 11393
rect 938 11319 994 11328
rect 1584 11144 1636 11150
rect 1584 11086 1636 11092
rect 1596 10985 1624 11086
rect 1582 10976 1638 10985
rect 1582 10911 1638 10920
rect 940 10668 992 10674
rect 940 10610 992 10616
rect 952 10577 980 10610
rect 1216 10600 1268 10606
rect 938 10568 994 10577
rect 1216 10542 1268 10548
rect 938 10503 994 10512
rect 1228 10169 1256 10542
rect 1214 10160 1270 10169
rect 1214 10095 1270 10104
rect 940 10056 992 10062
rect 940 9998 992 10004
rect 952 9761 980 9998
rect 938 9752 994 9761
rect 938 9687 994 9696
rect 940 9580 992 9586
rect 940 9522 992 9528
rect 952 9353 980 9522
rect 1766 9480 1822 9489
rect 1766 9415 1768 9424
rect 1820 9415 1822 9424
rect 1768 9386 1820 9392
rect 938 9344 994 9353
rect 938 9279 994 9288
rect 940 8968 992 8974
rect 938 8936 940 8945
rect 992 8936 994 8945
rect 938 8871 994 8880
rect 1216 8900 1268 8906
rect 1216 8842 1268 8848
rect 1228 8537 1256 8842
rect 1214 8528 1270 8537
rect 1872 8498 1900 11834
rect 1214 8463 1270 8472
rect 1860 8492 1912 8498
rect 1860 8434 1912 8440
rect 1584 8424 1636 8430
rect 1584 8366 1636 8372
rect 1596 8129 1624 8366
rect 1582 8120 1638 8129
rect 1582 8055 1638 8064
rect 940 7880 992 7886
rect 940 7822 992 7828
rect 952 7721 980 7822
rect 938 7712 994 7721
rect 938 7647 994 7656
rect 940 7404 992 7410
rect 940 7346 992 7352
rect 952 7313 980 7346
rect 938 7304 994 7313
rect 938 7239 994 7248
rect 938 6896 994 6905
rect 938 6831 994 6840
rect 952 6798 980 6831
rect 940 6792 992 6798
rect 940 6734 992 6740
rect 1308 6724 1360 6730
rect 1308 6666 1360 6672
rect 1320 6497 1348 6666
rect 2332 6662 2360 14826
rect 2950 14716 3258 14725
rect 2950 14714 2956 14716
rect 3012 14714 3036 14716
rect 3092 14714 3116 14716
rect 3172 14714 3196 14716
rect 3252 14714 3258 14716
rect 3012 14662 3014 14714
rect 3194 14662 3196 14714
rect 2950 14660 2956 14662
rect 3012 14660 3036 14662
rect 3092 14660 3116 14662
rect 3172 14660 3196 14662
rect 3252 14660 3258 14662
rect 2950 14651 3258 14660
rect 3608 14544 3660 14550
rect 3608 14486 3660 14492
rect 3620 14074 3648 14486
rect 3608 14068 3660 14074
rect 3608 14010 3660 14016
rect 3516 13932 3568 13938
rect 3516 13874 3568 13880
rect 2778 13832 2834 13841
rect 2778 13767 2834 13776
rect 2792 13326 2820 13767
rect 2950 13628 3258 13637
rect 2950 13626 2956 13628
rect 3012 13626 3036 13628
rect 3092 13626 3116 13628
rect 3172 13626 3196 13628
rect 3252 13626 3258 13628
rect 3012 13574 3014 13626
rect 3194 13574 3196 13626
rect 2950 13572 2956 13574
rect 3012 13572 3036 13574
rect 3092 13572 3116 13574
rect 3172 13572 3196 13574
rect 3252 13572 3258 13574
rect 2950 13563 3258 13572
rect 3528 13433 3556 13874
rect 3514 13424 3570 13433
rect 3514 13359 3570 13368
rect 2780 13320 2832 13326
rect 2780 13262 2832 13268
rect 2950 12540 3258 12549
rect 2950 12538 2956 12540
rect 3012 12538 3036 12540
rect 3092 12538 3116 12540
rect 3172 12538 3196 12540
rect 3252 12538 3258 12540
rect 3012 12486 3014 12538
rect 3194 12486 3196 12538
rect 2950 12484 2956 12486
rect 3012 12484 3036 12486
rect 3092 12484 3116 12486
rect 3172 12484 3196 12486
rect 3252 12484 3258 12486
rect 2950 12475 3258 12484
rect 4172 11558 4200 15982
rect 5368 12306 5396 17206
rect 5448 16652 5500 16658
rect 5448 16594 5500 16600
rect 5460 12986 5488 16594
rect 6380 16250 6408 20402
rect 7300 19786 7328 23666
rect 7392 22574 7420 26200
rect 7470 24712 7526 24721
rect 8036 24698 8064 26200
rect 7470 24647 7526 24656
rect 7852 24670 8064 24698
rect 7484 24206 7512 24647
rect 7472 24200 7524 24206
rect 7472 24142 7524 24148
rect 7472 24064 7524 24070
rect 7472 24006 7524 24012
rect 7484 22642 7512 24006
rect 7748 23248 7800 23254
rect 7748 23190 7800 23196
rect 7656 23044 7708 23050
rect 7656 22986 7708 22992
rect 7564 22704 7616 22710
rect 7564 22646 7616 22652
rect 7472 22636 7524 22642
rect 7472 22578 7524 22584
rect 7380 22568 7432 22574
rect 7380 22510 7432 22516
rect 7288 19780 7340 19786
rect 7288 19722 7340 19728
rect 7576 19378 7604 22646
rect 7668 20330 7696 22986
rect 7760 22030 7788 23190
rect 7852 23186 7880 24670
rect 8680 24274 8708 26200
rect 9220 25220 9272 25226
rect 9220 25162 9272 25168
rect 8852 25084 8904 25090
rect 8852 25026 8904 25032
rect 8668 24268 8720 24274
rect 8668 24210 8720 24216
rect 7950 23964 8258 23973
rect 7950 23962 7956 23964
rect 8012 23962 8036 23964
rect 8092 23962 8116 23964
rect 8172 23962 8196 23964
rect 8252 23962 8258 23964
rect 8012 23910 8014 23962
rect 8194 23910 8196 23962
rect 7950 23908 7956 23910
rect 8012 23908 8036 23910
rect 8092 23908 8116 23910
rect 8172 23908 8196 23910
rect 8252 23908 8258 23910
rect 7950 23899 8258 23908
rect 7840 23180 7892 23186
rect 7840 23122 7892 23128
rect 8300 23112 8352 23118
rect 8300 23054 8352 23060
rect 7950 22876 8258 22885
rect 7950 22874 7956 22876
rect 8012 22874 8036 22876
rect 8092 22874 8116 22876
rect 8172 22874 8196 22876
rect 8252 22874 8258 22876
rect 8012 22822 8014 22874
rect 8194 22822 8196 22874
rect 7950 22820 7956 22822
rect 8012 22820 8036 22822
rect 8092 22820 8116 22822
rect 8172 22820 8196 22822
rect 8252 22820 8258 22822
rect 7950 22811 8258 22820
rect 7748 22024 7800 22030
rect 7748 21966 7800 21972
rect 7950 21788 8258 21797
rect 7950 21786 7956 21788
rect 8012 21786 8036 21788
rect 8092 21786 8116 21788
rect 8172 21786 8196 21788
rect 8252 21786 8258 21788
rect 8012 21734 8014 21786
rect 8194 21734 8196 21786
rect 7950 21732 7956 21734
rect 8012 21732 8036 21734
rect 8092 21732 8116 21734
rect 8172 21732 8196 21734
rect 8252 21732 8258 21734
rect 7950 21723 8258 21732
rect 7840 20800 7892 20806
rect 7840 20742 7892 20748
rect 7656 20324 7708 20330
rect 7656 20266 7708 20272
rect 7564 19372 7616 19378
rect 7564 19314 7616 19320
rect 6828 17060 6880 17066
rect 6828 17002 6880 17008
rect 6840 16590 6868 17002
rect 7576 16590 7604 19314
rect 7852 18766 7880 20742
rect 7950 20700 8258 20709
rect 7950 20698 7956 20700
rect 8012 20698 8036 20700
rect 8092 20698 8116 20700
rect 8172 20698 8196 20700
rect 8252 20698 8258 20700
rect 8012 20646 8014 20698
rect 8194 20646 8196 20698
rect 7950 20644 7956 20646
rect 8012 20644 8036 20646
rect 8092 20644 8116 20646
rect 8172 20644 8196 20646
rect 8252 20644 8258 20646
rect 7950 20635 8258 20644
rect 8312 20602 8340 23054
rect 8864 21486 8892 25026
rect 9128 24064 9180 24070
rect 9128 24006 9180 24012
rect 9140 23118 9168 24006
rect 9128 23112 9180 23118
rect 9128 23054 9180 23060
rect 9128 22432 9180 22438
rect 9128 22374 9180 22380
rect 9140 22030 9168 22374
rect 9232 22098 9260 25162
rect 9324 23798 9352 26200
rect 9680 24200 9732 24206
rect 9680 24142 9732 24148
rect 9312 23792 9364 23798
rect 9312 23734 9364 23740
rect 9588 23656 9640 23662
rect 9588 23598 9640 23604
rect 9312 22976 9364 22982
rect 9312 22918 9364 22924
rect 9220 22092 9272 22098
rect 9220 22034 9272 22040
rect 9128 22024 9180 22030
rect 9128 21966 9180 21972
rect 8852 21480 8904 21486
rect 8852 21422 8904 21428
rect 8300 20596 8352 20602
rect 8300 20538 8352 20544
rect 9324 19922 9352 22918
rect 9600 20602 9628 23598
rect 9692 23526 9720 24142
rect 9680 23520 9732 23526
rect 9680 23462 9732 23468
rect 9968 22658 9996 26200
rect 10324 24132 10376 24138
rect 10324 24074 10376 24080
rect 9968 22630 10088 22658
rect 10060 22574 10088 22630
rect 10048 22568 10100 22574
rect 10048 22510 10100 22516
rect 10336 21690 10364 24074
rect 10612 23798 10640 26200
rect 10600 23792 10652 23798
rect 10600 23734 10652 23740
rect 11256 23186 11284 26200
rect 11900 24342 11928 26200
rect 11888 24336 11940 24342
rect 11888 24278 11940 24284
rect 12072 23656 12124 23662
rect 12072 23598 12124 23604
rect 11244 23180 11296 23186
rect 11244 23122 11296 23128
rect 10692 23112 10744 23118
rect 10692 23054 10744 23060
rect 10508 22160 10560 22166
rect 10508 22102 10560 22108
rect 9680 21684 9732 21690
rect 9680 21626 9732 21632
rect 10324 21684 10376 21690
rect 10324 21626 10376 21632
rect 9588 20596 9640 20602
rect 9588 20538 9640 20544
rect 9692 20262 9720 21626
rect 10416 21616 10468 21622
rect 10416 21558 10468 21564
rect 9864 21480 9916 21486
rect 9864 21422 9916 21428
rect 9772 20392 9824 20398
rect 9772 20334 9824 20340
rect 9680 20256 9732 20262
rect 9680 20198 9732 20204
rect 9312 19916 9364 19922
rect 9312 19858 9364 19864
rect 9496 19848 9548 19854
rect 9496 19790 9548 19796
rect 7950 19612 8258 19621
rect 7950 19610 7956 19612
rect 8012 19610 8036 19612
rect 8092 19610 8116 19612
rect 8172 19610 8196 19612
rect 8252 19610 8258 19612
rect 8012 19558 8014 19610
rect 8194 19558 8196 19610
rect 7950 19556 7956 19558
rect 8012 19556 8036 19558
rect 8092 19556 8116 19558
rect 8172 19556 8196 19558
rect 8252 19556 8258 19558
rect 7950 19547 8258 19556
rect 9312 19508 9364 19514
rect 9312 19450 9364 19456
rect 9128 19304 9180 19310
rect 9128 19246 9180 19252
rect 9140 18834 9168 19246
rect 9128 18828 9180 18834
rect 9128 18770 9180 18776
rect 7840 18760 7892 18766
rect 7840 18702 7892 18708
rect 8300 18624 8352 18630
rect 8300 18566 8352 18572
rect 7950 18524 8258 18533
rect 7950 18522 7956 18524
rect 8012 18522 8036 18524
rect 8092 18522 8116 18524
rect 8172 18522 8196 18524
rect 8252 18522 8258 18524
rect 8012 18470 8014 18522
rect 8194 18470 8196 18522
rect 7950 18468 7956 18470
rect 8012 18468 8036 18470
rect 8092 18468 8116 18470
rect 8172 18468 8196 18470
rect 8252 18468 8258 18470
rect 7950 18459 8258 18468
rect 7950 17436 8258 17445
rect 7950 17434 7956 17436
rect 8012 17434 8036 17436
rect 8092 17434 8116 17436
rect 8172 17434 8196 17436
rect 8252 17434 8258 17436
rect 8012 17382 8014 17434
rect 8194 17382 8196 17434
rect 7950 17380 7956 17382
rect 8012 17380 8036 17382
rect 8092 17380 8116 17382
rect 8172 17380 8196 17382
rect 8252 17380 8258 17382
rect 7950 17371 8258 17380
rect 8312 17202 8340 18566
rect 8300 17196 8352 17202
rect 8300 17138 8352 17144
rect 8576 16652 8628 16658
rect 8576 16594 8628 16600
rect 6828 16584 6880 16590
rect 6828 16526 6880 16532
rect 7564 16584 7616 16590
rect 7564 16526 7616 16532
rect 7950 16348 8258 16357
rect 7950 16346 7956 16348
rect 8012 16346 8036 16348
rect 8092 16346 8116 16348
rect 8172 16346 8196 16348
rect 8252 16346 8258 16348
rect 8012 16294 8014 16346
rect 8194 16294 8196 16346
rect 7950 16292 7956 16294
rect 8012 16292 8036 16294
rect 8092 16292 8116 16294
rect 8172 16292 8196 16294
rect 8252 16292 8258 16294
rect 7950 16283 8258 16292
rect 6368 16244 6420 16250
rect 6368 16186 6420 16192
rect 8588 16046 8616 16594
rect 9324 16250 9352 19450
rect 9312 16244 9364 16250
rect 9312 16186 9364 16192
rect 8576 16040 8628 16046
rect 8576 15982 8628 15988
rect 6644 15360 6696 15366
rect 6644 15302 6696 15308
rect 6656 15026 6684 15302
rect 7950 15260 8258 15269
rect 7950 15258 7956 15260
rect 8012 15258 8036 15260
rect 8092 15258 8116 15260
rect 8172 15258 8196 15260
rect 8252 15258 8258 15260
rect 8012 15206 8014 15258
rect 8194 15206 8196 15258
rect 7950 15204 7956 15206
rect 8012 15204 8036 15206
rect 8092 15204 8116 15206
rect 8172 15204 8196 15206
rect 8252 15204 8258 15206
rect 7950 15195 8258 15204
rect 6644 15020 6696 15026
rect 6644 14962 6696 14968
rect 7950 14172 8258 14181
rect 7950 14170 7956 14172
rect 8012 14170 8036 14172
rect 8092 14170 8116 14172
rect 8172 14170 8196 14172
rect 8252 14170 8258 14172
rect 8012 14118 8014 14170
rect 8194 14118 8196 14170
rect 7950 14116 7956 14118
rect 8012 14116 8036 14118
rect 8092 14116 8116 14118
rect 8172 14116 8196 14118
rect 8252 14116 8258 14118
rect 7950 14107 8258 14116
rect 8588 13258 8616 15982
rect 9508 15978 9536 19790
rect 9784 18426 9812 20334
rect 9876 18970 9904 21422
rect 10428 20602 10456 21558
rect 10416 20596 10468 20602
rect 10416 20538 10468 20544
rect 10048 20460 10100 20466
rect 10048 20402 10100 20408
rect 9864 18964 9916 18970
rect 9864 18906 9916 18912
rect 9772 18420 9824 18426
rect 9772 18362 9824 18368
rect 9864 18284 9916 18290
rect 9864 18226 9916 18232
rect 9876 16998 9904 18226
rect 10060 18154 10088 20402
rect 10416 19168 10468 19174
rect 10416 19110 10468 19116
rect 10428 18426 10456 19110
rect 10416 18420 10468 18426
rect 10416 18362 10468 18368
rect 10048 18148 10100 18154
rect 10048 18090 10100 18096
rect 10520 17762 10548 22102
rect 10704 21690 10732 23054
rect 12084 22681 12112 23598
rect 12440 23588 12492 23594
rect 12440 23530 12492 23536
rect 12070 22672 12126 22681
rect 12070 22607 12126 22616
rect 12452 22030 12480 23530
rect 12544 22574 12572 26200
rect 12950 24508 13258 24517
rect 12950 24506 12956 24508
rect 13012 24506 13036 24508
rect 13092 24506 13116 24508
rect 13172 24506 13196 24508
rect 13252 24506 13258 24508
rect 13012 24454 13014 24506
rect 13194 24454 13196 24506
rect 12950 24452 12956 24454
rect 13012 24452 13036 24454
rect 13092 24452 13116 24454
rect 13172 24452 13196 24454
rect 13252 24452 13258 24454
rect 12950 24443 13258 24452
rect 12624 24200 12676 24206
rect 12624 24142 12676 24148
rect 12532 22568 12584 22574
rect 12532 22510 12584 22516
rect 11980 22024 12032 22030
rect 12072 22024 12124 22030
rect 11980 21966 12032 21972
rect 12070 21992 12072 22001
rect 12440 22024 12492 22030
rect 12124 21992 12126 22001
rect 11428 21888 11480 21894
rect 11428 21830 11480 21836
rect 11612 21888 11664 21894
rect 11612 21830 11664 21836
rect 10692 21684 10744 21690
rect 10692 21626 10744 21632
rect 11244 21412 11296 21418
rect 11244 21354 11296 21360
rect 11150 21040 11206 21049
rect 11150 20975 11206 20984
rect 11164 20942 11192 20975
rect 10968 20936 11020 20942
rect 10968 20878 11020 20884
rect 11152 20936 11204 20942
rect 11152 20878 11204 20884
rect 10692 20596 10744 20602
rect 10692 20538 10744 20544
rect 10428 17734 10548 17762
rect 10428 17134 10456 17734
rect 10508 17672 10560 17678
rect 10508 17614 10560 17620
rect 10600 17672 10652 17678
rect 10600 17614 10652 17620
rect 10232 17128 10284 17134
rect 10232 17070 10284 17076
rect 10416 17128 10468 17134
rect 10416 17070 10468 17076
rect 9864 16992 9916 16998
rect 9864 16934 9916 16940
rect 9588 16516 9640 16522
rect 9588 16458 9640 16464
rect 9496 15972 9548 15978
rect 9496 15914 9548 15920
rect 9220 15904 9272 15910
rect 9220 15846 9272 15852
rect 9232 15162 9260 15846
rect 9220 15156 9272 15162
rect 9220 15098 9272 15104
rect 9600 15094 9628 16458
rect 9588 15088 9640 15094
rect 9588 15030 9640 15036
rect 10140 14340 10192 14346
rect 10140 14282 10192 14288
rect 10152 14249 10180 14282
rect 10138 14240 10194 14249
rect 10138 14175 10194 14184
rect 8576 13252 8628 13258
rect 8576 13194 8628 13200
rect 7950 13084 8258 13093
rect 7950 13082 7956 13084
rect 8012 13082 8036 13084
rect 8092 13082 8116 13084
rect 8172 13082 8196 13084
rect 8252 13082 8258 13084
rect 8012 13030 8014 13082
rect 8194 13030 8196 13082
rect 7950 13028 7956 13030
rect 8012 13028 8036 13030
rect 8092 13028 8116 13030
rect 8172 13028 8196 13030
rect 8252 13028 8258 13030
rect 7950 13019 8258 13028
rect 5448 12980 5500 12986
rect 5448 12922 5500 12928
rect 10244 12918 10272 17070
rect 10520 16794 10548 17614
rect 10508 16788 10560 16794
rect 10508 16730 10560 16736
rect 10612 15570 10640 17614
rect 10704 17202 10732 20538
rect 10876 19440 10928 19446
rect 10876 19382 10928 19388
rect 10888 18970 10916 19382
rect 10980 18970 11008 20878
rect 11256 20534 11284 21354
rect 11336 20596 11388 20602
rect 11336 20538 11388 20544
rect 11244 20528 11296 20534
rect 11244 20470 11296 20476
rect 11348 19854 11376 20538
rect 11440 20534 11468 21830
rect 11624 21486 11652 21830
rect 11612 21480 11664 21486
rect 11612 21422 11664 21428
rect 11520 20868 11572 20874
rect 11520 20810 11572 20816
rect 11428 20528 11480 20534
rect 11428 20470 11480 20476
rect 11060 19848 11112 19854
rect 11060 19790 11112 19796
rect 11336 19848 11388 19854
rect 11336 19790 11388 19796
rect 11072 19514 11100 19790
rect 11060 19508 11112 19514
rect 11060 19450 11112 19456
rect 11532 19174 11560 20810
rect 11702 20768 11758 20777
rect 11702 20703 11758 20712
rect 11612 19236 11664 19242
rect 11612 19178 11664 19184
rect 11336 19168 11388 19174
rect 11336 19110 11388 19116
rect 11520 19168 11572 19174
rect 11520 19110 11572 19116
rect 10876 18964 10928 18970
rect 10876 18906 10928 18912
rect 10968 18964 11020 18970
rect 10968 18906 11020 18912
rect 10692 17196 10744 17202
rect 10692 17138 10744 17144
rect 10888 16658 10916 18906
rect 11060 18828 11112 18834
rect 11060 18770 11112 18776
rect 10968 17128 11020 17134
rect 10968 17070 11020 17076
rect 10980 16726 11008 17070
rect 10968 16720 11020 16726
rect 10968 16662 11020 16668
rect 10876 16652 10928 16658
rect 10876 16594 10928 16600
rect 11072 16590 11100 18770
rect 11348 18698 11376 19110
rect 11244 18692 11296 18698
rect 11244 18634 11296 18640
rect 11336 18692 11388 18698
rect 11336 18634 11388 18640
rect 11256 18426 11284 18634
rect 11520 18624 11572 18630
rect 11520 18566 11572 18572
rect 11152 18420 11204 18426
rect 11152 18362 11204 18368
rect 11244 18420 11296 18426
rect 11244 18362 11296 18368
rect 11060 16584 11112 16590
rect 11060 16526 11112 16532
rect 11060 16448 11112 16454
rect 11060 16390 11112 16396
rect 11072 15706 11100 16390
rect 11164 16250 11192 18362
rect 11428 18148 11480 18154
rect 11428 18090 11480 18096
rect 11244 18080 11296 18086
rect 11244 18022 11296 18028
rect 11152 16244 11204 16250
rect 11152 16186 11204 16192
rect 11060 15700 11112 15706
rect 11060 15642 11112 15648
rect 10600 15564 10652 15570
rect 10600 15506 10652 15512
rect 11060 15564 11112 15570
rect 11060 15506 11112 15512
rect 10416 15496 10468 15502
rect 10416 15438 10468 15444
rect 10428 14618 10456 15438
rect 10968 15428 11020 15434
rect 10968 15370 11020 15376
rect 10980 15042 11008 15370
rect 11072 15162 11100 15506
rect 11060 15156 11112 15162
rect 11060 15098 11112 15104
rect 10980 15026 11100 15042
rect 10980 15020 11112 15026
rect 10980 15014 11060 15020
rect 11060 14962 11112 14968
rect 10784 14952 10836 14958
rect 10784 14894 10836 14900
rect 10416 14612 10468 14618
rect 10416 14554 10468 14560
rect 10324 14340 10376 14346
rect 10324 14282 10376 14288
rect 10336 13297 10364 14282
rect 10508 13320 10560 13326
rect 10322 13288 10378 13297
rect 10508 13262 10560 13268
rect 10322 13223 10378 13232
rect 10232 12912 10284 12918
rect 10232 12854 10284 12860
rect 10520 12306 10548 13262
rect 10796 13190 10824 14894
rect 10876 14816 10928 14822
rect 10876 14758 10928 14764
rect 10784 13184 10836 13190
rect 10784 13126 10836 13132
rect 10796 12306 10824 13126
rect 10888 12986 10916 14758
rect 11256 14618 11284 18022
rect 11336 16516 11388 16522
rect 11336 16458 11388 16464
rect 11348 16017 11376 16458
rect 11334 16008 11390 16017
rect 11334 15943 11390 15952
rect 11244 14612 11296 14618
rect 11244 14554 11296 14560
rect 11150 14376 11206 14385
rect 11150 14311 11152 14320
rect 11204 14311 11206 14320
rect 11152 14282 11204 14288
rect 11244 14272 11296 14278
rect 11244 14214 11296 14220
rect 11256 14006 11284 14214
rect 11244 14000 11296 14006
rect 11244 13942 11296 13948
rect 11060 13252 11112 13258
rect 11060 13194 11112 13200
rect 10876 12980 10928 12986
rect 10876 12922 10928 12928
rect 5356 12300 5408 12306
rect 5356 12242 5408 12248
rect 10508 12300 10560 12306
rect 10508 12242 10560 12248
rect 10784 12300 10836 12306
rect 10784 12242 10836 12248
rect 11072 12209 11100 13194
rect 11348 12345 11376 15943
rect 11440 15162 11468 18090
rect 11532 17202 11560 18566
rect 11624 18222 11652 19178
rect 11612 18216 11664 18222
rect 11612 18158 11664 18164
rect 11624 17746 11652 18158
rect 11612 17740 11664 17746
rect 11612 17682 11664 17688
rect 11520 17196 11572 17202
rect 11520 17138 11572 17144
rect 11520 16448 11572 16454
rect 11520 16390 11572 16396
rect 11532 16250 11560 16390
rect 11716 16266 11744 20703
rect 11888 20460 11940 20466
rect 11888 20402 11940 20408
rect 11900 16794 11928 20402
rect 11992 20262 12020 21966
rect 12440 21966 12492 21972
rect 12070 21927 12126 21936
rect 12636 21894 12664 24142
rect 12716 23860 12768 23866
rect 12716 23802 12768 23808
rect 12440 21888 12492 21894
rect 12440 21830 12492 21836
rect 12624 21888 12676 21894
rect 12624 21830 12676 21836
rect 12164 21616 12216 21622
rect 12348 21616 12400 21622
rect 12216 21564 12348 21570
rect 12164 21558 12400 21564
rect 12176 21542 12388 21558
rect 12452 20913 12480 21830
rect 12624 21548 12676 21554
rect 12624 21490 12676 21496
rect 12532 21480 12584 21486
rect 12532 21422 12584 21428
rect 12438 20904 12494 20913
rect 12438 20839 12494 20848
rect 11980 20256 12032 20262
rect 11980 20198 12032 20204
rect 11980 19848 12032 19854
rect 11980 19790 12032 19796
rect 11992 19242 12020 19790
rect 12164 19780 12216 19786
rect 12164 19722 12216 19728
rect 12256 19780 12308 19786
rect 12256 19722 12308 19728
rect 12072 19712 12124 19718
rect 12072 19654 12124 19660
rect 12084 19378 12112 19654
rect 12072 19372 12124 19378
rect 12072 19314 12124 19320
rect 11980 19236 12032 19242
rect 11980 19178 12032 19184
rect 11980 18964 12032 18970
rect 11980 18906 12032 18912
rect 11992 18748 12020 18906
rect 12176 18902 12204 19722
rect 12164 18896 12216 18902
rect 12164 18838 12216 18844
rect 11992 18720 12204 18748
rect 12176 18630 12204 18720
rect 12164 18624 12216 18630
rect 12164 18566 12216 18572
rect 11980 18420 12032 18426
rect 11980 18362 12032 18368
rect 11992 17678 12020 18362
rect 12268 18358 12296 19722
rect 12256 18352 12308 18358
rect 12256 18294 12308 18300
rect 12268 17882 12296 18294
rect 12256 17876 12308 17882
rect 12256 17818 12308 17824
rect 12070 17776 12126 17785
rect 12070 17711 12126 17720
rect 11980 17672 12032 17678
rect 11980 17614 12032 17620
rect 11888 16788 11940 16794
rect 11888 16730 11940 16736
rect 11520 16244 11572 16250
rect 11716 16238 11836 16266
rect 11520 16186 11572 16192
rect 11704 16108 11756 16114
rect 11704 16050 11756 16056
rect 11428 15156 11480 15162
rect 11428 15098 11480 15104
rect 11716 14482 11744 16050
rect 11808 15026 11836 16238
rect 11886 16144 11942 16153
rect 11886 16079 11942 16088
rect 11900 15978 11928 16079
rect 11888 15972 11940 15978
rect 11888 15914 11940 15920
rect 11992 15892 12020 17614
rect 12084 17202 12112 17711
rect 12164 17536 12216 17542
rect 12164 17478 12216 17484
rect 12072 17196 12124 17202
rect 12072 17138 12124 17144
rect 12072 16448 12124 16454
rect 12072 16390 12124 16396
rect 12084 16046 12112 16390
rect 12072 16040 12124 16046
rect 12072 15982 12124 15988
rect 11992 15864 12112 15892
rect 12084 15434 12112 15864
rect 12072 15428 12124 15434
rect 12072 15370 12124 15376
rect 11796 15020 11848 15026
rect 11796 14962 11848 14968
rect 11704 14476 11756 14482
rect 11704 14418 11756 14424
rect 11808 13870 11836 14962
rect 12084 14906 12112 15370
rect 12176 15026 12204 17478
rect 12452 17202 12480 20839
rect 12544 17814 12572 21422
rect 12636 21146 12664 21490
rect 12728 21146 12756 23802
rect 12950 23420 13258 23429
rect 12950 23418 12956 23420
rect 13012 23418 13036 23420
rect 13092 23418 13116 23420
rect 13172 23418 13196 23420
rect 13252 23418 13258 23420
rect 13012 23366 13014 23418
rect 13194 23366 13196 23418
rect 12950 23364 12956 23366
rect 13012 23364 13036 23366
rect 13092 23364 13116 23366
rect 13172 23364 13196 23366
rect 13252 23364 13258 23366
rect 12950 23355 13258 23364
rect 13372 23186 13400 26302
rect 13818 26200 13874 27000
rect 14462 26200 14518 27000
rect 15106 26330 15162 27000
rect 15028 26302 15162 26330
rect 13832 24274 13860 26200
rect 14476 24970 14504 26200
rect 14384 24942 14504 24970
rect 13820 24268 13872 24274
rect 13820 24210 13872 24216
rect 13636 24132 13688 24138
rect 13636 24074 13688 24080
rect 13728 24132 13780 24138
rect 13728 24074 13780 24080
rect 13452 24064 13504 24070
rect 13452 24006 13504 24012
rect 13464 23730 13492 24006
rect 13452 23724 13504 23730
rect 13452 23666 13504 23672
rect 13360 23180 13412 23186
rect 13360 23122 13412 23128
rect 12808 22976 12860 22982
rect 12808 22918 12860 22924
rect 12820 22642 12848 22918
rect 13360 22772 13412 22778
rect 13360 22714 13412 22720
rect 12808 22636 12860 22642
rect 12808 22578 12860 22584
rect 12950 22332 13258 22341
rect 12950 22330 12956 22332
rect 13012 22330 13036 22332
rect 13092 22330 13116 22332
rect 13172 22330 13196 22332
rect 13252 22330 13258 22332
rect 13012 22278 13014 22330
rect 13194 22278 13196 22330
rect 12950 22276 12956 22278
rect 13012 22276 13036 22278
rect 13092 22276 13116 22278
rect 13172 22276 13196 22278
rect 13252 22276 13258 22278
rect 12950 22267 13258 22276
rect 12808 21956 12860 21962
rect 12808 21898 12860 21904
rect 12624 21140 12676 21146
rect 12624 21082 12676 21088
rect 12716 21140 12768 21146
rect 12716 21082 12768 21088
rect 12716 20256 12768 20262
rect 12636 20204 12716 20210
rect 12636 20198 12768 20204
rect 12636 20182 12756 20198
rect 12636 19718 12664 20182
rect 12624 19712 12676 19718
rect 12624 19654 12676 19660
rect 12624 19508 12676 19514
rect 12624 19450 12676 19456
rect 12636 18426 12664 19450
rect 12714 19272 12770 19281
rect 12714 19207 12716 19216
rect 12768 19207 12770 19216
rect 12716 19178 12768 19184
rect 12624 18420 12676 18426
rect 12624 18362 12676 18368
rect 12716 18080 12768 18086
rect 12716 18022 12768 18028
rect 12532 17808 12584 17814
rect 12532 17750 12584 17756
rect 12728 17542 12756 18022
rect 12820 17882 12848 21898
rect 12950 21244 13258 21253
rect 12950 21242 12956 21244
rect 13012 21242 13036 21244
rect 13092 21242 13116 21244
rect 13172 21242 13196 21244
rect 13252 21242 13258 21244
rect 13012 21190 13014 21242
rect 13194 21190 13196 21242
rect 12950 21188 12956 21190
rect 13012 21188 13036 21190
rect 13092 21188 13116 21190
rect 13172 21188 13196 21190
rect 13252 21188 13258 21190
rect 12950 21179 13258 21188
rect 12950 20156 13258 20165
rect 12950 20154 12956 20156
rect 13012 20154 13036 20156
rect 13092 20154 13116 20156
rect 13172 20154 13196 20156
rect 13252 20154 13258 20156
rect 13012 20102 13014 20154
rect 13194 20102 13196 20154
rect 12950 20100 12956 20102
rect 13012 20100 13036 20102
rect 13092 20100 13116 20102
rect 13172 20100 13196 20102
rect 13252 20100 13258 20102
rect 12950 20091 13258 20100
rect 13372 19990 13400 22714
rect 13452 21616 13504 21622
rect 13452 21558 13504 21564
rect 13360 19984 13412 19990
rect 13360 19926 13412 19932
rect 13268 19712 13320 19718
rect 13268 19654 13320 19660
rect 13280 19446 13308 19654
rect 13360 19508 13412 19514
rect 13360 19450 13412 19456
rect 13268 19440 13320 19446
rect 13268 19382 13320 19388
rect 12950 19068 13258 19077
rect 12950 19066 12956 19068
rect 13012 19066 13036 19068
rect 13092 19066 13116 19068
rect 13172 19066 13196 19068
rect 13252 19066 13258 19068
rect 13012 19014 13014 19066
rect 13194 19014 13196 19066
rect 12950 19012 12956 19014
rect 13012 19012 13036 19014
rect 13092 19012 13116 19014
rect 13172 19012 13196 19014
rect 13252 19012 13258 19014
rect 12950 19003 13258 19012
rect 13372 18834 13400 19450
rect 13084 18828 13136 18834
rect 13084 18770 13136 18776
rect 13360 18828 13412 18834
rect 13360 18770 13412 18776
rect 13096 18630 13124 18770
rect 13084 18624 13136 18630
rect 13084 18566 13136 18572
rect 13372 18222 13400 18770
rect 13464 18222 13492 21558
rect 13544 21344 13596 21350
rect 13544 21286 13596 21292
rect 13556 20874 13584 21286
rect 13648 21146 13676 24074
rect 13740 22166 13768 24074
rect 14384 23798 14412 24942
rect 14464 24200 14516 24206
rect 14464 24142 14516 24148
rect 14372 23792 14424 23798
rect 14372 23734 14424 23740
rect 13820 23248 13872 23254
rect 13820 23190 13872 23196
rect 13728 22160 13780 22166
rect 13728 22102 13780 22108
rect 13832 22098 13860 23190
rect 14372 23112 14424 23118
rect 14372 23054 14424 23060
rect 13820 22092 13872 22098
rect 13820 22034 13872 22040
rect 14004 22024 14056 22030
rect 14004 21966 14056 21972
rect 13728 21684 13780 21690
rect 13780 21644 13952 21672
rect 13728 21626 13780 21632
rect 13728 21480 13780 21486
rect 13728 21422 13780 21428
rect 13636 21140 13688 21146
rect 13636 21082 13688 21088
rect 13636 21004 13688 21010
rect 13636 20946 13688 20952
rect 13544 20868 13596 20874
rect 13544 20810 13596 20816
rect 13648 20602 13676 20946
rect 13636 20596 13688 20602
rect 13636 20538 13688 20544
rect 13634 20496 13690 20505
rect 13634 20431 13636 20440
rect 13688 20431 13690 20440
rect 13636 20402 13688 20408
rect 13544 19984 13596 19990
rect 13544 19926 13596 19932
rect 13360 18216 13412 18222
rect 13360 18158 13412 18164
rect 13452 18216 13504 18222
rect 13452 18158 13504 18164
rect 12950 17980 13258 17989
rect 12950 17978 12956 17980
rect 13012 17978 13036 17980
rect 13092 17978 13116 17980
rect 13172 17978 13196 17980
rect 13252 17978 13258 17980
rect 13012 17926 13014 17978
rect 13194 17926 13196 17978
rect 12950 17924 12956 17926
rect 13012 17924 13036 17926
rect 13092 17924 13116 17926
rect 13172 17924 13196 17926
rect 13252 17924 13258 17926
rect 12950 17915 13258 17924
rect 12808 17876 12860 17882
rect 12808 17818 12860 17824
rect 12716 17536 12768 17542
rect 12716 17478 12768 17484
rect 12624 17332 12676 17338
rect 12624 17274 12676 17280
rect 13360 17332 13412 17338
rect 13360 17274 13412 17280
rect 12440 17196 12492 17202
rect 12440 17138 12492 17144
rect 12256 17128 12308 17134
rect 12256 17070 12308 17076
rect 12268 16726 12296 17070
rect 12256 16720 12308 16726
rect 12256 16662 12308 16668
rect 12532 16720 12584 16726
rect 12532 16662 12584 16668
rect 12636 16674 12664 17274
rect 12950 16892 13258 16901
rect 12950 16890 12956 16892
rect 13012 16890 13036 16892
rect 13092 16890 13116 16892
rect 13172 16890 13196 16892
rect 13252 16890 13258 16892
rect 13012 16838 13014 16890
rect 13194 16838 13196 16890
rect 12950 16836 12956 16838
rect 13012 16836 13036 16838
rect 13092 16836 13116 16838
rect 13172 16836 13196 16838
rect 13252 16836 13258 16838
rect 12950 16827 13258 16836
rect 12440 16584 12492 16590
rect 12440 16526 12492 16532
rect 12348 16176 12400 16182
rect 12348 16118 12400 16124
rect 12256 16040 12308 16046
rect 12256 15982 12308 15988
rect 12268 15706 12296 15982
rect 12256 15700 12308 15706
rect 12256 15642 12308 15648
rect 12360 15502 12388 16118
rect 12452 16046 12480 16526
rect 12440 16040 12492 16046
rect 12440 15982 12492 15988
rect 12348 15496 12400 15502
rect 12348 15438 12400 15444
rect 12452 15366 12480 15982
rect 12440 15360 12492 15366
rect 12440 15302 12492 15308
rect 12256 15156 12308 15162
rect 12256 15098 12308 15104
rect 12164 15020 12216 15026
rect 12164 14962 12216 14968
rect 12084 14878 12204 14906
rect 12268 14890 12296 15098
rect 11980 14068 12032 14074
rect 11980 14010 12032 14016
rect 11796 13864 11848 13870
rect 11796 13806 11848 13812
rect 11334 12336 11390 12345
rect 11334 12271 11390 12280
rect 11058 12200 11114 12209
rect 11058 12135 11114 12144
rect 7950 11996 8258 12005
rect 7950 11994 7956 11996
rect 8012 11994 8036 11996
rect 8092 11994 8116 11996
rect 8172 11994 8196 11996
rect 8252 11994 8258 11996
rect 8012 11942 8014 11994
rect 8194 11942 8196 11994
rect 7950 11940 7956 11942
rect 8012 11940 8036 11942
rect 8092 11940 8116 11942
rect 8172 11940 8196 11942
rect 8252 11940 8258 11942
rect 7950 11931 8258 11940
rect 4160 11552 4212 11558
rect 4160 11494 4212 11500
rect 2950 11452 3258 11461
rect 2950 11450 2956 11452
rect 3012 11450 3036 11452
rect 3092 11450 3116 11452
rect 3172 11450 3196 11452
rect 3252 11450 3258 11452
rect 3012 11398 3014 11450
rect 3194 11398 3196 11450
rect 2950 11396 2956 11398
rect 3012 11396 3036 11398
rect 3092 11396 3116 11398
rect 3172 11396 3196 11398
rect 3252 11396 3258 11398
rect 2950 11387 3258 11396
rect 7950 10908 8258 10917
rect 7950 10906 7956 10908
rect 8012 10906 8036 10908
rect 8092 10906 8116 10908
rect 8172 10906 8196 10908
rect 8252 10906 8258 10908
rect 8012 10854 8014 10906
rect 8194 10854 8196 10906
rect 7950 10852 7956 10854
rect 8012 10852 8036 10854
rect 8092 10852 8116 10854
rect 8172 10852 8196 10854
rect 8252 10852 8258 10854
rect 7950 10843 8258 10852
rect 11888 10464 11940 10470
rect 11888 10406 11940 10412
rect 2950 10364 3258 10373
rect 2950 10362 2956 10364
rect 3012 10362 3036 10364
rect 3092 10362 3116 10364
rect 3172 10362 3196 10364
rect 3252 10362 3258 10364
rect 3012 10310 3014 10362
rect 3194 10310 3196 10362
rect 2950 10308 2956 10310
rect 3012 10308 3036 10310
rect 3092 10308 3116 10310
rect 3172 10308 3196 10310
rect 3252 10308 3258 10310
rect 2950 10299 3258 10308
rect 11900 10130 11928 10406
rect 11888 10124 11940 10130
rect 11888 10066 11940 10072
rect 11992 10062 12020 14010
rect 12176 13326 12204 14878
rect 12256 14884 12308 14890
rect 12256 14826 12308 14832
rect 12256 14612 12308 14618
rect 12256 14554 12308 14560
rect 12164 13320 12216 13326
rect 12164 13262 12216 13268
rect 12176 12866 12204 13262
rect 12268 12986 12296 14554
rect 12544 14550 12572 16662
rect 12636 16646 12756 16674
rect 12624 16516 12676 16522
rect 12624 16458 12676 16464
rect 12636 14550 12664 16458
rect 12728 16182 12756 16646
rect 13268 16448 13320 16454
rect 13268 16390 13320 16396
rect 12716 16176 12768 16182
rect 12716 16118 12768 16124
rect 12808 16040 12860 16046
rect 12808 15982 12860 15988
rect 12716 15904 12768 15910
rect 12716 15846 12768 15852
rect 12532 14544 12584 14550
rect 12532 14486 12584 14492
rect 12624 14544 12676 14550
rect 12624 14486 12676 14492
rect 12624 14340 12676 14346
rect 12624 14282 12676 14288
rect 12532 14272 12584 14278
rect 12532 14214 12584 14220
rect 12440 13796 12492 13802
rect 12440 13738 12492 13744
rect 12452 13190 12480 13738
rect 12440 13184 12492 13190
rect 12440 13126 12492 13132
rect 12256 12980 12308 12986
rect 12256 12922 12308 12928
rect 12176 12838 12296 12866
rect 12164 12776 12216 12782
rect 12164 12718 12216 12724
rect 12176 12102 12204 12718
rect 12268 12238 12296 12838
rect 12440 12776 12492 12782
rect 12440 12718 12492 12724
rect 12452 12458 12480 12718
rect 12360 12430 12480 12458
rect 12256 12232 12308 12238
rect 12256 12174 12308 12180
rect 12164 12096 12216 12102
rect 12164 12038 12216 12044
rect 12176 11014 12204 12038
rect 12268 11082 12296 12174
rect 12360 11830 12388 12430
rect 12348 11824 12400 11830
rect 12348 11766 12400 11772
rect 12256 11076 12308 11082
rect 12256 11018 12308 11024
rect 12164 11008 12216 11014
rect 12164 10950 12216 10956
rect 12072 10532 12124 10538
rect 12072 10474 12124 10480
rect 12084 10130 12112 10474
rect 12176 10130 12204 10950
rect 12544 10266 12572 14214
rect 12636 13530 12664 14282
rect 12624 13524 12676 13530
rect 12624 13466 12676 13472
rect 12624 12640 12676 12646
rect 12624 12582 12676 12588
rect 12532 10260 12584 10266
rect 12532 10202 12584 10208
rect 12440 10192 12492 10198
rect 12440 10134 12492 10140
rect 12072 10124 12124 10130
rect 12072 10066 12124 10072
rect 12164 10124 12216 10130
rect 12164 10066 12216 10072
rect 11980 10056 12032 10062
rect 11980 9998 12032 10004
rect 7950 9820 8258 9829
rect 7950 9818 7956 9820
rect 8012 9818 8036 9820
rect 8092 9818 8116 9820
rect 8172 9818 8196 9820
rect 8252 9818 8258 9820
rect 8012 9766 8014 9818
rect 8194 9766 8196 9818
rect 7950 9764 7956 9766
rect 8012 9764 8036 9766
rect 8092 9764 8116 9766
rect 8172 9764 8196 9766
rect 8252 9764 8258 9766
rect 7950 9755 8258 9764
rect 12452 9654 12480 10134
rect 12636 9654 12664 12582
rect 12728 12306 12756 15846
rect 12820 13954 12848 15982
rect 13280 15892 13308 16390
rect 13372 16250 13400 17274
rect 13556 16522 13584 19926
rect 13740 19281 13768 21422
rect 13924 21078 13952 21644
rect 13912 21072 13964 21078
rect 13912 21014 13964 21020
rect 14016 20942 14044 21966
rect 14188 21072 14240 21078
rect 14188 21014 14240 21020
rect 14004 20936 14056 20942
rect 14004 20878 14056 20884
rect 13912 20868 13964 20874
rect 13912 20810 13964 20816
rect 13820 19712 13872 19718
rect 13924 19700 13952 20810
rect 13872 19672 13952 19700
rect 13820 19654 13872 19660
rect 13726 19272 13782 19281
rect 13726 19207 13782 19216
rect 13740 18834 13768 19207
rect 13728 18828 13780 18834
rect 13728 18770 13780 18776
rect 13832 18358 13860 19654
rect 14016 19174 14044 20878
rect 14004 19168 14056 19174
rect 14004 19110 14056 19116
rect 13820 18352 13872 18358
rect 13820 18294 13872 18300
rect 14016 17746 14044 19110
rect 14200 18057 14228 21014
rect 14384 20602 14412 23054
rect 14372 20596 14424 20602
rect 14372 20538 14424 20544
rect 14280 19848 14332 19854
rect 14280 19790 14332 19796
rect 14292 19446 14320 19790
rect 14280 19440 14332 19446
rect 14280 19382 14332 19388
rect 14186 18048 14242 18057
rect 14186 17983 14242 17992
rect 13820 17740 13872 17746
rect 13820 17682 13872 17688
rect 14004 17740 14056 17746
rect 14004 17682 14056 17688
rect 13636 17672 13688 17678
rect 13636 17614 13688 17620
rect 13544 16516 13596 16522
rect 13544 16458 13596 16464
rect 13360 16244 13412 16250
rect 13360 16186 13412 16192
rect 13280 15864 13400 15892
rect 12950 15804 13258 15813
rect 12950 15802 12956 15804
rect 13012 15802 13036 15804
rect 13092 15802 13116 15804
rect 13172 15802 13196 15804
rect 13252 15802 13258 15804
rect 13012 15750 13014 15802
rect 13194 15750 13196 15802
rect 12950 15748 12956 15750
rect 13012 15748 13036 15750
rect 13092 15748 13116 15750
rect 13172 15748 13196 15750
rect 13252 15748 13258 15750
rect 12950 15739 13258 15748
rect 13268 15700 13320 15706
rect 13268 15642 13320 15648
rect 13280 15434 13308 15642
rect 13372 15570 13400 15864
rect 13452 15632 13504 15638
rect 13452 15574 13504 15580
rect 13360 15564 13412 15570
rect 13360 15506 13412 15512
rect 13268 15428 13320 15434
rect 13268 15370 13320 15376
rect 13174 15056 13230 15065
rect 13174 14991 13176 15000
rect 13228 14991 13230 15000
rect 13176 14962 13228 14968
rect 13188 14890 13216 14962
rect 13176 14884 13228 14890
rect 13176 14826 13228 14832
rect 12950 14716 13258 14725
rect 12950 14714 12956 14716
rect 13012 14714 13036 14716
rect 13092 14714 13116 14716
rect 13172 14714 13196 14716
rect 13252 14714 13258 14716
rect 13012 14662 13014 14714
rect 13194 14662 13196 14714
rect 12950 14660 12956 14662
rect 13012 14660 13036 14662
rect 13092 14660 13116 14662
rect 13172 14660 13196 14662
rect 13252 14660 13258 14662
rect 12950 14651 13258 14660
rect 13176 14476 13228 14482
rect 13176 14418 13228 14424
rect 12820 13926 12940 13954
rect 12808 13864 12860 13870
rect 12808 13806 12860 13812
rect 12820 13394 12848 13806
rect 12912 13734 12940 13926
rect 13188 13870 13216 14418
rect 13176 13864 13228 13870
rect 13176 13806 13228 13812
rect 12900 13728 12952 13734
rect 12900 13670 12952 13676
rect 12950 13628 13258 13637
rect 12950 13626 12956 13628
rect 13012 13626 13036 13628
rect 13092 13626 13116 13628
rect 13172 13626 13196 13628
rect 13252 13626 13258 13628
rect 13012 13574 13014 13626
rect 13194 13574 13196 13626
rect 12950 13572 12956 13574
rect 13012 13572 13036 13574
rect 13092 13572 13116 13574
rect 13172 13572 13196 13574
rect 13252 13572 13258 13574
rect 12950 13563 13258 13572
rect 12808 13388 12860 13394
rect 12808 13330 12860 13336
rect 12820 12782 12848 13330
rect 12900 13320 12952 13326
rect 12900 13262 12952 13268
rect 12808 12776 12860 12782
rect 12808 12718 12860 12724
rect 12912 12628 12940 13262
rect 13360 12776 13412 12782
rect 13360 12718 13412 12724
rect 12820 12600 12940 12628
rect 12716 12300 12768 12306
rect 12716 12242 12768 12248
rect 12716 11688 12768 11694
rect 12716 11630 12768 11636
rect 12728 11286 12756 11630
rect 12716 11280 12768 11286
rect 12716 11222 12768 11228
rect 12440 9648 12492 9654
rect 12440 9590 12492 9596
rect 12624 9648 12676 9654
rect 12624 9590 12676 9596
rect 12728 9518 12756 11222
rect 12820 10606 12848 12600
rect 12950 12540 13258 12549
rect 12950 12538 12956 12540
rect 13012 12538 13036 12540
rect 13092 12538 13116 12540
rect 13172 12538 13196 12540
rect 13252 12538 13258 12540
rect 13012 12486 13014 12538
rect 13194 12486 13196 12538
rect 12950 12484 12956 12486
rect 13012 12484 13036 12486
rect 13092 12484 13116 12486
rect 13172 12484 13196 12486
rect 13252 12484 13258 12486
rect 12950 12475 13258 12484
rect 13372 12238 13400 12718
rect 13464 12434 13492 15574
rect 13544 15360 13596 15366
rect 13544 15302 13596 15308
rect 13556 14482 13584 15302
rect 13544 14476 13596 14482
rect 13544 14418 13596 14424
rect 13648 13954 13676 17614
rect 13728 16108 13780 16114
rect 13728 16050 13780 16056
rect 13740 15162 13768 16050
rect 13728 15156 13780 15162
rect 13728 15098 13780 15104
rect 13832 15094 13860 17682
rect 14476 17270 14504 24142
rect 15028 22574 15056 26302
rect 15106 26200 15162 26302
rect 15750 26200 15806 27000
rect 16394 26330 16450 27000
rect 16132 26302 16450 26330
rect 15764 23186 15792 26200
rect 16028 24336 16080 24342
rect 16028 24278 16080 24284
rect 15752 23180 15804 23186
rect 15752 23122 15804 23128
rect 15108 23112 15160 23118
rect 15108 23054 15160 23060
rect 15016 22568 15068 22574
rect 15016 22510 15068 22516
rect 14740 22500 14792 22506
rect 14740 22442 14792 22448
rect 14556 21480 14608 21486
rect 14556 21422 14608 21428
rect 14568 21010 14596 21422
rect 14556 21004 14608 21010
rect 14556 20946 14608 20952
rect 14648 20800 14700 20806
rect 14648 20742 14700 20748
rect 14660 19961 14688 20742
rect 14752 20058 14780 22442
rect 14924 21956 14976 21962
rect 14924 21898 14976 21904
rect 14832 21616 14884 21622
rect 14832 21558 14884 21564
rect 14844 20806 14872 21558
rect 14832 20800 14884 20806
rect 14832 20742 14884 20748
rect 14844 20398 14872 20742
rect 14832 20392 14884 20398
rect 14832 20334 14884 20340
rect 14740 20052 14792 20058
rect 14740 19994 14792 20000
rect 14646 19952 14702 19961
rect 14646 19887 14702 19896
rect 14648 19848 14700 19854
rect 14648 19790 14700 19796
rect 14556 17604 14608 17610
rect 14556 17546 14608 17552
rect 14188 17264 14240 17270
rect 14186 17232 14188 17241
rect 14464 17264 14516 17270
rect 14240 17232 14242 17241
rect 14464 17206 14516 17212
rect 14186 17167 14242 17176
rect 13912 16652 13964 16658
rect 13912 16594 13964 16600
rect 13924 16096 13952 16594
rect 14464 16448 14516 16454
rect 14464 16390 14516 16396
rect 14372 16176 14424 16182
rect 14370 16144 14372 16153
rect 14424 16144 14426 16153
rect 14004 16108 14056 16114
rect 13924 16068 14004 16096
rect 13820 15088 13872 15094
rect 13820 15030 13872 15036
rect 13728 14816 13780 14822
rect 13924 14770 13952 16068
rect 14370 16079 14426 16088
rect 14004 16050 14056 16056
rect 14096 16040 14148 16046
rect 14096 15982 14148 15988
rect 14002 14920 14058 14929
rect 14002 14855 14058 14864
rect 13780 14764 13952 14770
rect 13728 14758 13952 14764
rect 13740 14742 13952 14758
rect 13728 14272 13780 14278
rect 13728 14214 13780 14220
rect 13556 13926 13676 13954
rect 13556 12617 13584 13926
rect 13636 13864 13688 13870
rect 13636 13806 13688 13812
rect 13648 12782 13676 13806
rect 13636 12776 13688 12782
rect 13636 12718 13688 12724
rect 13542 12608 13598 12617
rect 13542 12543 13598 12552
rect 13464 12406 13584 12434
rect 13360 12232 13412 12238
rect 13360 12174 13412 12180
rect 12950 11452 13258 11461
rect 12950 11450 12956 11452
rect 13012 11450 13036 11452
rect 13092 11450 13116 11452
rect 13172 11450 13196 11452
rect 13252 11450 13258 11452
rect 13012 11398 13014 11450
rect 13194 11398 13196 11450
rect 12950 11396 12956 11398
rect 13012 11396 13036 11398
rect 13092 11396 13116 11398
rect 13172 11396 13196 11398
rect 13252 11396 13258 11398
rect 12950 11387 13258 11396
rect 12808 10600 12860 10606
rect 12808 10542 12860 10548
rect 12950 10364 13258 10373
rect 12950 10362 12956 10364
rect 13012 10362 13036 10364
rect 13092 10362 13116 10364
rect 13172 10362 13196 10364
rect 13252 10362 13258 10364
rect 13012 10310 13014 10362
rect 13194 10310 13196 10362
rect 12950 10308 12956 10310
rect 13012 10308 13036 10310
rect 13092 10308 13116 10310
rect 13172 10308 13196 10310
rect 13252 10308 13258 10310
rect 12950 10299 13258 10308
rect 13372 10130 13400 12174
rect 13452 12164 13504 12170
rect 13452 12106 13504 12112
rect 13464 11762 13492 12106
rect 13452 11756 13504 11762
rect 13452 11698 13504 11704
rect 13452 11008 13504 11014
rect 13452 10950 13504 10956
rect 13464 10674 13492 10950
rect 13452 10668 13504 10674
rect 13452 10610 13504 10616
rect 13360 10124 13412 10130
rect 13360 10066 13412 10072
rect 13268 10056 13320 10062
rect 13266 10024 13268 10033
rect 13320 10024 13322 10033
rect 13266 9959 13322 9968
rect 13452 9988 13504 9994
rect 13452 9930 13504 9936
rect 12716 9512 12768 9518
rect 12716 9454 12768 9460
rect 12808 9444 12860 9450
rect 12808 9386 12860 9392
rect 12164 9376 12216 9382
rect 12164 9318 12216 9324
rect 2950 9276 3258 9285
rect 2950 9274 2956 9276
rect 3012 9274 3036 9276
rect 3092 9274 3116 9276
rect 3172 9274 3196 9276
rect 3252 9274 3258 9276
rect 3012 9222 3014 9274
rect 3194 9222 3196 9274
rect 2950 9220 2956 9222
rect 3012 9220 3036 9222
rect 3092 9220 3116 9222
rect 3172 9220 3196 9222
rect 3252 9220 3258 9222
rect 2950 9211 3258 9220
rect 12176 9178 12204 9318
rect 12164 9172 12216 9178
rect 12164 9114 12216 9120
rect 7950 8732 8258 8741
rect 7950 8730 7956 8732
rect 8012 8730 8036 8732
rect 8092 8730 8116 8732
rect 8172 8730 8196 8732
rect 8252 8730 8258 8732
rect 8012 8678 8014 8730
rect 8194 8678 8196 8730
rect 7950 8676 7956 8678
rect 8012 8676 8036 8678
rect 8092 8676 8116 8678
rect 8172 8676 8196 8678
rect 8252 8676 8258 8678
rect 7950 8667 8258 8676
rect 2950 8188 3258 8197
rect 2950 8186 2956 8188
rect 3012 8186 3036 8188
rect 3092 8186 3116 8188
rect 3172 8186 3196 8188
rect 3252 8186 3258 8188
rect 3012 8134 3014 8186
rect 3194 8134 3196 8186
rect 2950 8132 2956 8134
rect 3012 8132 3036 8134
rect 3092 8132 3116 8134
rect 3172 8132 3196 8134
rect 3252 8132 3258 8134
rect 2950 8123 3258 8132
rect 12820 7886 12848 9386
rect 12950 9276 13258 9285
rect 12950 9274 12956 9276
rect 13012 9274 13036 9276
rect 13092 9274 13116 9276
rect 13172 9274 13196 9276
rect 13252 9274 13258 9276
rect 13012 9222 13014 9274
rect 13194 9222 13196 9274
rect 12950 9220 12956 9222
rect 13012 9220 13036 9222
rect 13092 9220 13116 9222
rect 13172 9220 13196 9222
rect 13252 9220 13258 9222
rect 12950 9211 13258 9220
rect 12950 8188 13258 8197
rect 12950 8186 12956 8188
rect 13012 8186 13036 8188
rect 13092 8186 13116 8188
rect 13172 8186 13196 8188
rect 13252 8186 13258 8188
rect 13012 8134 13014 8186
rect 13194 8134 13196 8186
rect 12950 8132 12956 8134
rect 13012 8132 13036 8134
rect 13092 8132 13116 8134
rect 13172 8132 13196 8134
rect 13252 8132 13258 8134
rect 12950 8123 13258 8132
rect 12808 7880 12860 7886
rect 12808 7822 12860 7828
rect 7950 7644 8258 7653
rect 7950 7642 7956 7644
rect 8012 7642 8036 7644
rect 8092 7642 8116 7644
rect 8172 7642 8196 7644
rect 8252 7642 8258 7644
rect 8012 7590 8014 7642
rect 8194 7590 8196 7642
rect 7950 7588 7956 7590
rect 8012 7588 8036 7590
rect 8092 7588 8116 7590
rect 8172 7588 8196 7590
rect 8252 7588 8258 7590
rect 7950 7579 8258 7588
rect 2950 7100 3258 7109
rect 2950 7098 2956 7100
rect 3012 7098 3036 7100
rect 3092 7098 3116 7100
rect 3172 7098 3196 7100
rect 3252 7098 3258 7100
rect 3012 7046 3014 7098
rect 3194 7046 3196 7098
rect 2950 7044 2956 7046
rect 3012 7044 3036 7046
rect 3092 7044 3116 7046
rect 3172 7044 3196 7046
rect 3252 7044 3258 7046
rect 2950 7035 3258 7044
rect 12950 7100 13258 7109
rect 12950 7098 12956 7100
rect 13012 7098 13036 7100
rect 13092 7098 13116 7100
rect 13172 7098 13196 7100
rect 13252 7098 13258 7100
rect 13012 7046 13014 7098
rect 13194 7046 13196 7098
rect 12950 7044 12956 7046
rect 13012 7044 13036 7046
rect 13092 7044 13116 7046
rect 13172 7044 13196 7046
rect 13252 7044 13258 7046
rect 12950 7035 13258 7044
rect 2320 6656 2372 6662
rect 2320 6598 2372 6604
rect 7950 6556 8258 6565
rect 7950 6554 7956 6556
rect 8012 6554 8036 6556
rect 8092 6554 8116 6556
rect 8172 6554 8196 6556
rect 8252 6554 8258 6556
rect 8012 6502 8014 6554
rect 8194 6502 8196 6554
rect 7950 6500 7956 6502
rect 8012 6500 8036 6502
rect 8092 6500 8116 6502
rect 8172 6500 8196 6502
rect 8252 6500 8258 6502
rect 1306 6488 1362 6497
rect 7950 6491 8258 6500
rect 1306 6423 1362 6432
rect 940 6316 992 6322
rect 940 6258 992 6264
rect 952 6089 980 6258
rect 1860 6180 1912 6186
rect 1860 6122 1912 6128
rect 938 6080 994 6089
rect 938 6015 994 6024
rect 940 5704 992 5710
rect 938 5672 940 5681
rect 992 5672 994 5681
rect 938 5607 994 5616
rect 940 5160 992 5166
rect 940 5102 992 5108
rect 952 4865 980 5102
rect 938 4856 994 4865
rect 938 4791 994 4800
rect 940 4548 992 4554
rect 940 4490 992 4496
rect 952 4457 980 4490
rect 938 4448 994 4457
rect 938 4383 994 4392
rect 1676 4208 1728 4214
rect 1676 4150 1728 4156
rect 940 4140 992 4146
rect 940 4082 992 4088
rect 952 3641 980 4082
rect 1688 4049 1716 4150
rect 1872 4078 1900 6122
rect 2950 6012 3258 6021
rect 2950 6010 2956 6012
rect 3012 6010 3036 6012
rect 3092 6010 3116 6012
rect 3172 6010 3196 6012
rect 3252 6010 3258 6012
rect 3012 5958 3014 6010
rect 3194 5958 3196 6010
rect 2950 5956 2956 5958
rect 3012 5956 3036 5958
rect 3092 5956 3116 5958
rect 3172 5956 3196 5958
rect 3252 5956 3258 5958
rect 2950 5947 3258 5956
rect 12950 6012 13258 6021
rect 12950 6010 12956 6012
rect 13012 6010 13036 6012
rect 13092 6010 13116 6012
rect 13172 6010 13196 6012
rect 13252 6010 13258 6012
rect 13012 5958 13014 6010
rect 13194 5958 13196 6010
rect 12950 5956 12956 5958
rect 13012 5956 13036 5958
rect 13092 5956 13116 5958
rect 13172 5956 13196 5958
rect 13252 5956 13258 5958
rect 12950 5947 13258 5956
rect 2320 5704 2372 5710
rect 2320 5646 2372 5652
rect 2332 5273 2360 5646
rect 7950 5468 8258 5477
rect 7950 5466 7956 5468
rect 8012 5466 8036 5468
rect 8092 5466 8116 5468
rect 8172 5466 8196 5468
rect 8252 5466 8258 5468
rect 8012 5414 8014 5466
rect 8194 5414 8196 5466
rect 7950 5412 7956 5414
rect 8012 5412 8036 5414
rect 8092 5412 8116 5414
rect 8172 5412 8196 5414
rect 8252 5412 8258 5414
rect 7950 5403 8258 5412
rect 2318 5264 2374 5273
rect 2318 5199 2374 5208
rect 2950 4924 3258 4933
rect 2950 4922 2956 4924
rect 3012 4922 3036 4924
rect 3092 4922 3116 4924
rect 3172 4922 3196 4924
rect 3252 4922 3258 4924
rect 3012 4870 3014 4922
rect 3194 4870 3196 4922
rect 2950 4868 2956 4870
rect 3012 4868 3036 4870
rect 3092 4868 3116 4870
rect 3172 4868 3196 4870
rect 3252 4868 3258 4870
rect 2950 4859 3258 4868
rect 12950 4924 13258 4933
rect 12950 4922 12956 4924
rect 13012 4922 13036 4924
rect 13092 4922 13116 4924
rect 13172 4922 13196 4924
rect 13252 4922 13258 4924
rect 13012 4870 13014 4922
rect 13194 4870 13196 4922
rect 12950 4868 12956 4870
rect 13012 4868 13036 4870
rect 13092 4868 13116 4870
rect 13172 4868 13196 4870
rect 13252 4868 13258 4870
rect 12950 4859 13258 4868
rect 7950 4380 8258 4389
rect 7950 4378 7956 4380
rect 8012 4378 8036 4380
rect 8092 4378 8116 4380
rect 8172 4378 8196 4380
rect 8252 4378 8258 4380
rect 8012 4326 8014 4378
rect 8194 4326 8196 4378
rect 7950 4324 7956 4326
rect 8012 4324 8036 4326
rect 8092 4324 8116 4326
rect 8172 4324 8196 4326
rect 8252 4324 8258 4326
rect 7950 4315 8258 4324
rect 1860 4072 1912 4078
rect 1674 4040 1730 4049
rect 1860 4014 1912 4020
rect 1674 3975 1730 3984
rect 2950 3836 3258 3845
rect 2950 3834 2956 3836
rect 3012 3834 3036 3836
rect 3092 3834 3116 3836
rect 3172 3834 3196 3836
rect 3252 3834 3258 3836
rect 3012 3782 3014 3834
rect 3194 3782 3196 3834
rect 2950 3780 2956 3782
rect 3012 3780 3036 3782
rect 3092 3780 3116 3782
rect 3172 3780 3196 3782
rect 3252 3780 3258 3782
rect 2950 3771 3258 3780
rect 12950 3836 13258 3845
rect 12950 3834 12956 3836
rect 13012 3834 13036 3836
rect 13092 3834 13116 3836
rect 13172 3834 13196 3836
rect 13252 3834 13258 3836
rect 13012 3782 13014 3834
rect 13194 3782 13196 3834
rect 12950 3780 12956 3782
rect 13012 3780 13036 3782
rect 13092 3780 13116 3782
rect 13172 3780 13196 3782
rect 13252 3780 13258 3782
rect 12950 3771 13258 3780
rect 938 3632 994 3641
rect 5354 3632 5410 3641
rect 938 3567 994 3576
rect 3332 3596 3384 3602
rect 5354 3567 5410 3576
rect 3332 3538 3384 3544
rect 940 3528 992 3534
rect 940 3470 992 3476
rect 1122 3496 1178 3505
rect 952 3233 980 3470
rect 1122 3431 1178 3440
rect 938 3224 994 3233
rect 938 3159 994 3168
rect 940 3052 992 3058
rect 940 2994 992 3000
rect 952 2825 980 2994
rect 938 2816 994 2825
rect 938 2751 994 2760
rect 940 2440 992 2446
rect 938 2408 940 2417
rect 992 2408 994 2417
rect 938 2343 994 2352
rect 1136 800 1164 3431
rect 2950 2748 3258 2757
rect 2950 2746 2956 2748
rect 3012 2746 3036 2748
rect 3092 2746 3116 2748
rect 3172 2746 3196 2748
rect 3252 2746 3258 2748
rect 3012 2694 3014 2746
rect 3194 2694 3196 2746
rect 2950 2692 2956 2694
rect 3012 2692 3036 2694
rect 3092 2692 3116 2694
rect 3172 2692 3196 2694
rect 3252 2692 3258 2694
rect 2950 2683 3258 2692
rect 1216 2372 1268 2378
rect 1216 2314 1268 2320
rect 1228 2009 1256 2314
rect 1308 2304 1360 2310
rect 1308 2246 1360 2252
rect 1214 2000 1270 2009
rect 1214 1935 1270 1944
rect 1320 1601 1348 2246
rect 3344 1850 3372 3538
rect 3252 1822 3372 1850
rect 1306 1592 1362 1601
rect 1306 1527 1362 1536
rect 3252 800 3280 1822
rect 5368 800 5396 3567
rect 12532 3392 12584 3398
rect 12532 3334 12584 3340
rect 7950 3292 8258 3301
rect 7950 3290 7956 3292
rect 8012 3290 8036 3292
rect 8092 3290 8116 3292
rect 8172 3290 8196 3292
rect 8252 3290 8258 3292
rect 8012 3238 8014 3290
rect 8194 3238 8196 3290
rect 7950 3236 7956 3238
rect 8012 3236 8036 3238
rect 8092 3236 8116 3238
rect 8172 3236 8196 3238
rect 8252 3236 8258 3238
rect 7950 3227 8258 3236
rect 7472 3188 7524 3194
rect 7472 3130 7524 3136
rect 7484 800 7512 3130
rect 11060 2984 11112 2990
rect 11060 2926 11112 2932
rect 11072 2582 11100 2926
rect 11060 2576 11112 2582
rect 11060 2518 11112 2524
rect 11704 2508 11756 2514
rect 11704 2450 11756 2456
rect 9588 2440 9640 2446
rect 9588 2382 9640 2388
rect 7950 2204 8258 2213
rect 7950 2202 7956 2204
rect 8012 2202 8036 2204
rect 8092 2202 8116 2204
rect 8172 2202 8196 2204
rect 8252 2202 8258 2204
rect 8012 2150 8014 2202
rect 8194 2150 8196 2202
rect 7950 2148 7956 2150
rect 8012 2148 8036 2150
rect 8092 2148 8116 2150
rect 8172 2148 8196 2150
rect 8252 2148 8258 2150
rect 7950 2139 8258 2148
rect 9600 800 9628 2382
rect 11716 800 11744 2450
rect 12544 2446 12572 3334
rect 12950 2748 13258 2757
rect 12950 2746 12956 2748
rect 13012 2746 13036 2748
rect 13092 2746 13116 2748
rect 13172 2746 13196 2748
rect 13252 2746 13258 2748
rect 13012 2694 13014 2746
rect 13194 2694 13196 2746
rect 12950 2692 12956 2694
rect 13012 2692 13036 2694
rect 13092 2692 13116 2694
rect 13172 2692 13196 2694
rect 13252 2692 13258 2694
rect 12950 2683 13258 2692
rect 13464 2582 13492 9930
rect 13556 8974 13584 12406
rect 13636 12300 13688 12306
rect 13636 12242 13688 12248
rect 13648 10690 13676 12242
rect 13740 11354 13768 14214
rect 13832 11762 13860 14742
rect 14016 14464 14044 14855
rect 13924 14436 14044 14464
rect 13820 11756 13872 11762
rect 13820 11698 13872 11704
rect 13728 11348 13780 11354
rect 13728 11290 13780 11296
rect 13924 11286 13952 14436
rect 14108 11558 14136 15982
rect 14476 15978 14504 16390
rect 14464 15972 14516 15978
rect 14464 15914 14516 15920
rect 14372 15904 14424 15910
rect 14372 15846 14424 15852
rect 14384 15502 14412 15846
rect 14568 15638 14596 17546
rect 14556 15632 14608 15638
rect 14556 15574 14608 15580
rect 14372 15496 14424 15502
rect 14372 15438 14424 15444
rect 14188 15088 14240 15094
rect 14188 15030 14240 15036
rect 14200 14006 14228 15030
rect 14568 14074 14596 15574
rect 14556 14068 14608 14074
rect 14556 14010 14608 14016
rect 14188 14000 14240 14006
rect 14188 13942 14240 13948
rect 14200 12986 14228 13942
rect 14556 13320 14608 13326
rect 14556 13262 14608 13268
rect 14188 12980 14240 12986
rect 14188 12922 14240 12928
rect 14280 12640 14332 12646
rect 14280 12582 14332 12588
rect 14292 12306 14320 12582
rect 14568 12306 14596 13262
rect 14660 12918 14688 19790
rect 14740 19780 14792 19786
rect 14740 19722 14792 19728
rect 14752 15910 14780 19722
rect 14832 18692 14884 18698
rect 14832 18634 14884 18640
rect 14844 18426 14872 18634
rect 14832 18420 14884 18426
rect 14832 18362 14884 18368
rect 14830 18184 14886 18193
rect 14830 18119 14886 18128
rect 14844 16658 14872 18119
rect 14832 16652 14884 16658
rect 14832 16594 14884 16600
rect 14936 16425 14964 21898
rect 15120 17882 15148 23054
rect 15660 22432 15712 22438
rect 15660 22374 15712 22380
rect 15476 21344 15528 21350
rect 15476 21286 15528 21292
rect 15292 21140 15344 21146
rect 15292 21082 15344 21088
rect 15304 19514 15332 21082
rect 15384 20460 15436 20466
rect 15384 20402 15436 20408
rect 15396 20369 15424 20402
rect 15382 20360 15438 20369
rect 15382 20295 15438 20304
rect 15292 19508 15344 19514
rect 15292 19450 15344 19456
rect 15200 18828 15252 18834
rect 15200 18770 15252 18776
rect 15292 18828 15344 18834
rect 15292 18770 15344 18776
rect 15212 18222 15240 18770
rect 15200 18216 15252 18222
rect 15200 18158 15252 18164
rect 15108 17876 15160 17882
rect 15108 17818 15160 17824
rect 15304 17610 15332 18770
rect 15488 18426 15516 21286
rect 15672 20534 15700 22374
rect 15844 20868 15896 20874
rect 15844 20810 15896 20816
rect 15660 20528 15712 20534
rect 15660 20470 15712 20476
rect 15856 19530 15884 20810
rect 15764 19502 15884 19530
rect 15764 19446 15792 19502
rect 15752 19440 15804 19446
rect 15752 19382 15804 19388
rect 15658 18864 15714 18873
rect 15764 18834 15792 19382
rect 15844 19372 15896 19378
rect 15844 19314 15896 19320
rect 15658 18799 15714 18808
rect 15752 18828 15804 18834
rect 15568 18624 15620 18630
rect 15568 18566 15620 18572
rect 15384 18420 15436 18426
rect 15384 18362 15436 18368
rect 15476 18420 15528 18426
rect 15476 18362 15528 18368
rect 15292 17604 15344 17610
rect 15292 17546 15344 17552
rect 15016 17128 15068 17134
rect 15016 17070 15068 17076
rect 14922 16416 14978 16425
rect 14922 16351 14978 16360
rect 14832 16040 14884 16046
rect 14832 15982 14884 15988
rect 14740 15904 14792 15910
rect 14740 15846 14792 15852
rect 14844 15366 14872 15982
rect 15028 15688 15056 17070
rect 15292 17060 15344 17066
rect 15292 17002 15344 17008
rect 15108 16652 15160 16658
rect 15108 16594 15160 16600
rect 15120 16046 15148 16594
rect 15304 16182 15332 17002
rect 15396 16250 15424 18362
rect 15580 17338 15608 18566
rect 15568 17332 15620 17338
rect 15568 17274 15620 17280
rect 15672 17202 15700 18799
rect 15752 18770 15804 18776
rect 15660 17196 15712 17202
rect 15660 17138 15712 17144
rect 15752 17196 15804 17202
rect 15752 17138 15804 17144
rect 15476 16992 15528 16998
rect 15476 16934 15528 16940
rect 15384 16244 15436 16250
rect 15384 16186 15436 16192
rect 15292 16176 15344 16182
rect 15292 16118 15344 16124
rect 15108 16040 15160 16046
rect 15108 15982 15160 15988
rect 15028 15660 15148 15688
rect 15016 15564 15068 15570
rect 15016 15506 15068 15512
rect 14832 15360 14884 15366
rect 14832 15302 14884 15308
rect 14738 15192 14794 15201
rect 14738 15127 14794 15136
rect 14648 12912 14700 12918
rect 14648 12854 14700 12860
rect 14752 12434 14780 15127
rect 15028 14958 15056 15506
rect 15120 15201 15148 15660
rect 15304 15502 15332 16118
rect 15384 15972 15436 15978
rect 15384 15914 15436 15920
rect 15292 15496 15344 15502
rect 15292 15438 15344 15444
rect 15106 15192 15162 15201
rect 15106 15127 15162 15136
rect 15016 14952 15068 14958
rect 15016 14894 15068 14900
rect 14924 14476 14976 14482
rect 14924 14418 14976 14424
rect 14936 13190 14964 14418
rect 14924 13184 14976 13190
rect 14924 13126 14976 13132
rect 14660 12406 14780 12434
rect 14280 12300 14332 12306
rect 14280 12242 14332 12248
rect 14556 12300 14608 12306
rect 14556 12242 14608 12248
rect 14660 12170 14688 12406
rect 14464 12164 14516 12170
rect 14464 12106 14516 12112
rect 14648 12164 14700 12170
rect 14648 12106 14700 12112
rect 14476 11880 14504 12106
rect 14556 11892 14608 11898
rect 14476 11852 14556 11880
rect 14556 11834 14608 11840
rect 14096 11552 14148 11558
rect 14096 11494 14148 11500
rect 14832 11552 14884 11558
rect 14832 11494 14884 11500
rect 13912 11280 13964 11286
rect 13912 11222 13964 11228
rect 14844 11218 14872 11494
rect 13820 11212 13872 11218
rect 13820 11154 13872 11160
rect 14832 11212 14884 11218
rect 14832 11154 14884 11160
rect 13648 10662 13768 10690
rect 13648 10266 13676 10662
rect 13740 10606 13768 10662
rect 13728 10600 13780 10606
rect 13728 10542 13780 10548
rect 13636 10260 13688 10266
rect 13636 10202 13688 10208
rect 13544 8968 13596 8974
rect 13544 8910 13596 8916
rect 13648 8378 13676 10202
rect 13832 10062 13860 11154
rect 14740 11144 14792 11150
rect 14740 11086 14792 11092
rect 14462 10704 14518 10713
rect 14372 10668 14424 10674
rect 14462 10639 14464 10648
rect 14372 10610 14424 10616
rect 14516 10639 14518 10648
rect 14464 10610 14516 10616
rect 13820 10056 13872 10062
rect 13820 9998 13872 10004
rect 13832 9654 13860 9998
rect 13820 9648 13872 9654
rect 13820 9590 13872 9596
rect 13832 8974 13860 9590
rect 14384 9178 14412 10610
rect 14372 9172 14424 9178
rect 14372 9114 14424 9120
rect 13820 8968 13872 8974
rect 13820 8910 13872 8916
rect 13832 8566 13860 8910
rect 13820 8560 13872 8566
rect 13820 8502 13872 8508
rect 13556 8362 13676 8378
rect 13544 8356 13676 8362
rect 13596 8350 13676 8356
rect 13544 8298 13596 8304
rect 13832 3058 13860 8502
rect 13820 3052 13872 3058
rect 13820 2994 13872 3000
rect 14476 2922 14504 10610
rect 14556 9988 14608 9994
rect 14556 9930 14608 9936
rect 14568 9110 14596 9930
rect 14556 9104 14608 9110
rect 14556 9046 14608 9052
rect 14752 8922 14780 11086
rect 14936 10606 14964 13126
rect 15028 12434 15056 14894
rect 15292 14068 15344 14074
rect 15292 14010 15344 14016
rect 15106 13696 15162 13705
rect 15106 13631 15162 13640
rect 15120 13394 15148 13631
rect 15108 13388 15160 13394
rect 15108 13330 15160 13336
rect 15200 13184 15252 13190
rect 15200 13126 15252 13132
rect 15028 12406 15148 12434
rect 15014 12200 15070 12209
rect 15014 12135 15070 12144
rect 14924 10600 14976 10606
rect 14924 10542 14976 10548
rect 15028 9654 15056 12135
rect 15120 11218 15148 12406
rect 15212 11218 15240 13126
rect 15304 12102 15332 14010
rect 15396 13394 15424 15914
rect 15488 14414 15516 16934
rect 15660 16584 15712 16590
rect 15660 16526 15712 16532
rect 15568 15700 15620 15706
rect 15568 15642 15620 15648
rect 15476 14408 15528 14414
rect 15476 14350 15528 14356
rect 15384 13388 15436 13394
rect 15384 13330 15436 13336
rect 15580 13258 15608 15642
rect 15672 15162 15700 16526
rect 15660 15156 15712 15162
rect 15660 15098 15712 15104
rect 15660 14272 15712 14278
rect 15660 14214 15712 14220
rect 15672 13841 15700 14214
rect 15658 13832 15714 13841
rect 15658 13767 15714 13776
rect 15568 13252 15620 13258
rect 15568 13194 15620 13200
rect 15660 13252 15712 13258
rect 15660 13194 15712 13200
rect 15384 12844 15436 12850
rect 15384 12786 15436 12792
rect 15396 12102 15424 12786
rect 15566 12608 15622 12617
rect 15566 12543 15622 12552
rect 15580 12374 15608 12543
rect 15568 12368 15620 12374
rect 15474 12336 15530 12345
rect 15568 12310 15620 12316
rect 15474 12271 15530 12280
rect 15292 12096 15344 12102
rect 15292 12038 15344 12044
rect 15384 12096 15436 12102
rect 15384 12038 15436 12044
rect 15396 11778 15424 12038
rect 15304 11750 15424 11778
rect 15488 11762 15516 12271
rect 15476 11756 15528 11762
rect 15304 11626 15332 11750
rect 15476 11698 15528 11704
rect 15292 11620 15344 11626
rect 15292 11562 15344 11568
rect 15108 11212 15160 11218
rect 15108 11154 15160 11160
rect 15200 11212 15252 11218
rect 15200 11154 15252 11160
rect 15292 10600 15344 10606
rect 15292 10542 15344 10548
rect 15016 9648 15068 9654
rect 15016 9590 15068 9596
rect 15200 9512 15252 9518
rect 15304 9466 15332 10542
rect 15672 10538 15700 13194
rect 15764 11778 15792 17138
rect 15856 16776 15884 19314
rect 15936 19304 15988 19310
rect 15936 19246 15988 19252
rect 15948 18970 15976 19246
rect 15936 18964 15988 18970
rect 15936 18906 15988 18912
rect 15948 17066 15976 18906
rect 16040 18766 16068 24278
rect 16132 23798 16160 26302
rect 16394 26200 16450 26302
rect 17038 26330 17094 27000
rect 17038 26302 17264 26330
rect 17038 26200 17094 26302
rect 16580 24200 16632 24206
rect 16580 24142 16632 24148
rect 16120 23792 16172 23798
rect 16120 23734 16172 23740
rect 16592 23633 16620 24142
rect 16578 23624 16634 23633
rect 16578 23559 16634 23568
rect 16580 23520 16632 23526
rect 16580 23462 16632 23468
rect 16304 21888 16356 21894
rect 16304 21830 16356 21836
rect 16488 21888 16540 21894
rect 16488 21830 16540 21836
rect 16120 21616 16172 21622
rect 16120 21558 16172 21564
rect 16132 20874 16160 21558
rect 16316 21350 16344 21830
rect 16500 21622 16528 21830
rect 16488 21616 16540 21622
rect 16488 21558 16540 21564
rect 16396 21480 16448 21486
rect 16396 21422 16448 21428
rect 16304 21344 16356 21350
rect 16304 21286 16356 21292
rect 16120 20868 16172 20874
rect 16120 20810 16172 20816
rect 16120 20460 16172 20466
rect 16120 20402 16172 20408
rect 16028 18760 16080 18766
rect 16028 18702 16080 18708
rect 16132 18426 16160 20402
rect 16316 19922 16344 21286
rect 16408 20058 16436 21422
rect 16488 20800 16540 20806
rect 16486 20768 16488 20777
rect 16540 20768 16542 20777
rect 16486 20703 16542 20712
rect 16396 20052 16448 20058
rect 16396 19994 16448 20000
rect 16304 19916 16356 19922
rect 16304 19858 16356 19864
rect 16488 19372 16540 19378
rect 16488 19314 16540 19320
rect 16212 19168 16264 19174
rect 16212 19110 16264 19116
rect 16224 18737 16252 19110
rect 16210 18728 16266 18737
rect 16210 18663 16266 18672
rect 16120 18420 16172 18426
rect 16120 18362 16172 18368
rect 16500 18329 16528 19314
rect 16592 18970 16620 23462
rect 17040 23112 17092 23118
rect 17040 23054 17092 23060
rect 17052 22710 17080 23054
rect 17040 22704 17092 22710
rect 17040 22646 17092 22652
rect 17052 21418 17080 22646
rect 17132 22568 17184 22574
rect 17132 22510 17184 22516
rect 17144 22234 17172 22510
rect 17132 22228 17184 22234
rect 17132 22170 17184 22176
rect 17144 21690 17172 22170
rect 17236 22166 17264 26302
rect 17682 26200 17738 27000
rect 18326 26200 18382 27000
rect 18970 26200 19026 27000
rect 19614 26200 19670 27000
rect 20258 26330 20314 27000
rect 20258 26302 20576 26330
rect 20258 26200 20314 26302
rect 17592 24676 17644 24682
rect 17592 24618 17644 24624
rect 17604 24206 17632 24618
rect 17696 24274 17724 26200
rect 17776 24608 17828 24614
rect 17776 24550 17828 24556
rect 17684 24268 17736 24274
rect 17684 24210 17736 24216
rect 17592 24200 17644 24206
rect 17592 24142 17644 24148
rect 17592 23316 17644 23322
rect 17592 23258 17644 23264
rect 17316 23044 17368 23050
rect 17316 22986 17368 22992
rect 17500 23044 17552 23050
rect 17500 22986 17552 22992
rect 17224 22160 17276 22166
rect 17224 22102 17276 22108
rect 17132 21684 17184 21690
rect 17132 21626 17184 21632
rect 17040 21412 17092 21418
rect 17040 21354 17092 21360
rect 17052 21010 17080 21354
rect 17040 21004 17092 21010
rect 17040 20946 17092 20952
rect 17052 20466 17080 20946
rect 17040 20460 17092 20466
rect 17040 20402 17092 20408
rect 16764 20392 16816 20398
rect 16764 20334 16816 20340
rect 16670 19816 16726 19825
rect 16670 19751 16672 19760
rect 16724 19751 16726 19760
rect 16672 19722 16724 19728
rect 16580 18964 16632 18970
rect 16580 18906 16632 18912
rect 16776 18426 16804 20334
rect 16856 20324 16908 20330
rect 16856 20266 16908 20272
rect 16868 19514 16896 20266
rect 16948 19780 17000 19786
rect 16948 19722 17000 19728
rect 16856 19508 16908 19514
rect 16856 19450 16908 19456
rect 16764 18420 16816 18426
rect 16764 18362 16816 18368
rect 16486 18320 16542 18329
rect 16486 18255 16542 18264
rect 16028 18216 16080 18222
rect 16028 18158 16080 18164
rect 16396 18216 16448 18222
rect 16396 18158 16448 18164
rect 16488 18216 16540 18222
rect 16488 18158 16540 18164
rect 16040 17882 16068 18158
rect 16028 17876 16080 17882
rect 16028 17818 16080 17824
rect 15936 17060 15988 17066
rect 15936 17002 15988 17008
rect 16028 16788 16080 16794
rect 15856 16748 15976 16776
rect 15844 16652 15896 16658
rect 15844 16594 15896 16600
rect 15856 13258 15884 16594
rect 15948 14906 15976 16748
rect 16028 16730 16080 16736
rect 16120 16788 16172 16794
rect 16120 16730 16172 16736
rect 16040 16590 16068 16730
rect 16028 16584 16080 16590
rect 16026 16552 16028 16561
rect 16080 16552 16082 16561
rect 16026 16487 16082 16496
rect 16132 16454 16160 16730
rect 16304 16652 16356 16658
rect 16304 16594 16356 16600
rect 16120 16448 16172 16454
rect 16120 16390 16172 16396
rect 16316 16114 16344 16594
rect 16304 16108 16356 16114
rect 16304 16050 16356 16056
rect 16120 16040 16172 16046
rect 16120 15982 16172 15988
rect 16132 15570 16160 15982
rect 16120 15564 16172 15570
rect 16120 15506 16172 15512
rect 16304 15564 16356 15570
rect 16304 15506 16356 15512
rect 16316 15473 16344 15506
rect 16302 15464 16358 15473
rect 16120 15428 16172 15434
rect 16302 15399 16358 15408
rect 16120 15370 16172 15376
rect 15948 14878 16068 14906
rect 15936 14816 15988 14822
rect 15936 14758 15988 14764
rect 15948 14074 15976 14758
rect 15936 14068 15988 14074
rect 15936 14010 15988 14016
rect 15936 13728 15988 13734
rect 15936 13670 15988 13676
rect 15844 13252 15896 13258
rect 15844 13194 15896 13200
rect 15842 12880 15898 12889
rect 15842 12815 15844 12824
rect 15896 12815 15898 12824
rect 15844 12786 15896 12792
rect 15948 12102 15976 13670
rect 16040 12764 16068 14878
rect 16132 12986 16160 15370
rect 16210 14512 16266 14521
rect 16210 14447 16212 14456
rect 16264 14447 16266 14456
rect 16212 14418 16264 14424
rect 16316 13258 16344 15399
rect 16408 13308 16436 18158
rect 16500 16538 16528 18158
rect 16764 18148 16816 18154
rect 16764 18090 16816 18096
rect 16672 17536 16724 17542
rect 16672 17478 16724 17484
rect 16580 17196 16632 17202
rect 16580 17138 16632 17144
rect 16592 17105 16620 17138
rect 16578 17096 16634 17105
rect 16578 17031 16634 17040
rect 16500 16510 16620 16538
rect 16486 16416 16542 16425
rect 16486 16351 16542 16360
rect 16500 16250 16528 16351
rect 16488 16244 16540 16250
rect 16488 16186 16540 16192
rect 16592 16130 16620 16510
rect 16500 16102 16620 16130
rect 16500 13734 16528 16102
rect 16580 13864 16632 13870
rect 16580 13806 16632 13812
rect 16488 13728 16540 13734
rect 16488 13670 16540 13676
rect 16408 13280 16528 13308
rect 16304 13252 16356 13258
rect 16304 13194 16356 13200
rect 16316 13025 16344 13194
rect 16500 13138 16528 13280
rect 16408 13110 16528 13138
rect 16302 13016 16358 13025
rect 16120 12980 16172 12986
rect 16302 12951 16358 12960
rect 16120 12922 16172 12928
rect 16302 12880 16358 12889
rect 16302 12815 16358 12824
rect 16212 12776 16264 12782
rect 16040 12736 16212 12764
rect 16212 12718 16264 12724
rect 16120 12640 16172 12646
rect 16120 12582 16172 12588
rect 16028 12436 16080 12442
rect 16028 12378 16080 12384
rect 15936 12096 15988 12102
rect 15936 12038 15988 12044
rect 15764 11762 15884 11778
rect 15764 11756 15896 11762
rect 15764 11750 15844 11756
rect 15660 10532 15712 10538
rect 15660 10474 15712 10480
rect 15568 10464 15620 10470
rect 15568 10406 15620 10412
rect 15474 9616 15530 9625
rect 15474 9551 15530 9560
rect 15252 9460 15332 9466
rect 15200 9454 15332 9460
rect 15212 9438 15332 9454
rect 15108 9172 15160 9178
rect 15108 9114 15160 9120
rect 14830 9072 14886 9081
rect 14830 9007 14832 9016
rect 14884 9007 14886 9016
rect 14832 8978 14884 8984
rect 14660 8894 14780 8922
rect 14556 8832 14608 8838
rect 14556 8774 14608 8780
rect 14568 8430 14596 8774
rect 14660 8634 14688 8894
rect 15120 8838 15148 9114
rect 14740 8832 14792 8838
rect 14740 8774 14792 8780
rect 15108 8832 15160 8838
rect 15108 8774 15160 8780
rect 14648 8628 14700 8634
rect 14648 8570 14700 8576
rect 14556 8424 14608 8430
rect 14556 8366 14608 8372
rect 14464 2916 14516 2922
rect 14464 2858 14516 2864
rect 13452 2576 13504 2582
rect 13452 2518 13504 2524
rect 13820 2508 13872 2514
rect 13820 2450 13872 2456
rect 12532 2440 12584 2446
rect 12532 2382 12584 2388
rect 13832 800 13860 2450
rect 14660 2378 14688 8570
rect 14752 3534 14780 8774
rect 15304 8634 15332 9438
rect 15292 8628 15344 8634
rect 15292 8570 15344 8576
rect 15488 7818 15516 9551
rect 15476 7812 15528 7818
rect 15476 7754 15528 7760
rect 15580 7410 15608 10406
rect 15568 7404 15620 7410
rect 15568 7346 15620 7352
rect 15764 5166 15792 11750
rect 15844 11698 15896 11704
rect 15948 10538 15976 12038
rect 16040 10810 16068 12378
rect 16028 10804 16080 10810
rect 16028 10746 16080 10752
rect 15936 10532 15988 10538
rect 15936 10474 15988 10480
rect 15948 9926 15976 10474
rect 16132 10130 16160 12582
rect 16212 12096 16264 12102
rect 16212 12038 16264 12044
rect 16224 10674 16252 12038
rect 16212 10668 16264 10674
rect 16212 10610 16264 10616
rect 16120 10124 16172 10130
rect 16120 10066 16172 10072
rect 16120 9988 16172 9994
rect 16120 9930 16172 9936
rect 16212 9988 16264 9994
rect 16212 9930 16264 9936
rect 15936 9920 15988 9926
rect 15936 9862 15988 9868
rect 16132 9722 16160 9930
rect 16120 9716 16172 9722
rect 16120 9658 16172 9664
rect 16224 8906 16252 9930
rect 16212 8900 16264 8906
rect 16212 8842 16264 8848
rect 16316 6118 16344 12815
rect 16408 12442 16436 13110
rect 16486 13016 16542 13025
rect 16486 12951 16542 12960
rect 16500 12850 16528 12951
rect 16488 12844 16540 12850
rect 16488 12786 16540 12792
rect 16396 12436 16448 12442
rect 16396 12378 16448 12384
rect 16396 12164 16448 12170
rect 16396 12106 16448 12112
rect 16408 11762 16436 12106
rect 16592 11830 16620 13806
rect 16580 11824 16632 11830
rect 16580 11766 16632 11772
rect 16396 11756 16448 11762
rect 16396 11698 16448 11704
rect 16408 10062 16436 11698
rect 16684 11354 16712 17478
rect 16776 15706 16804 18090
rect 16960 16726 16988 19722
rect 17052 19446 17080 20402
rect 17328 19990 17356 22986
rect 17408 22772 17460 22778
rect 17408 22714 17460 22720
rect 17420 22234 17448 22714
rect 17512 22438 17540 22986
rect 17500 22432 17552 22438
rect 17500 22374 17552 22380
rect 17408 22228 17460 22234
rect 17408 22170 17460 22176
rect 17604 22094 17632 23258
rect 17420 22066 17632 22094
rect 17420 21690 17448 22066
rect 17788 21690 17816 24550
rect 17950 23964 18258 23973
rect 17950 23962 17956 23964
rect 18012 23962 18036 23964
rect 18092 23962 18116 23964
rect 18172 23962 18196 23964
rect 18252 23962 18258 23964
rect 18012 23910 18014 23962
rect 18194 23910 18196 23962
rect 17950 23908 17956 23910
rect 18012 23908 18036 23910
rect 18092 23908 18116 23910
rect 18172 23908 18196 23910
rect 18252 23908 18258 23910
rect 17950 23899 18258 23908
rect 18340 23798 18368 26200
rect 18328 23792 18380 23798
rect 18328 23734 18380 23740
rect 18788 23724 18840 23730
rect 18788 23666 18840 23672
rect 17960 23656 18012 23662
rect 17960 23598 18012 23604
rect 17972 23322 18000 23598
rect 18800 23526 18828 23666
rect 18788 23520 18840 23526
rect 18788 23462 18840 23468
rect 17960 23316 18012 23322
rect 17960 23258 18012 23264
rect 18696 23044 18748 23050
rect 18696 22986 18748 22992
rect 17950 22876 18258 22885
rect 17950 22874 17956 22876
rect 18012 22874 18036 22876
rect 18092 22874 18116 22876
rect 18172 22874 18196 22876
rect 18252 22874 18258 22876
rect 18012 22822 18014 22874
rect 18194 22822 18196 22874
rect 17950 22820 17956 22822
rect 18012 22820 18036 22822
rect 18092 22820 18116 22822
rect 18172 22820 18196 22822
rect 18252 22820 18258 22822
rect 17950 22811 18258 22820
rect 18708 22710 18736 22986
rect 18696 22704 18748 22710
rect 18696 22646 18748 22652
rect 18880 22704 18932 22710
rect 18880 22646 18932 22652
rect 18604 22568 18656 22574
rect 18604 22510 18656 22516
rect 17950 21788 18258 21797
rect 17950 21786 17956 21788
rect 18012 21786 18036 21788
rect 18092 21786 18116 21788
rect 18172 21786 18196 21788
rect 18252 21786 18258 21788
rect 18012 21734 18014 21786
rect 18194 21734 18196 21786
rect 17950 21732 17956 21734
rect 18012 21732 18036 21734
rect 18092 21732 18116 21734
rect 18172 21732 18196 21734
rect 18252 21732 18258 21734
rect 17950 21723 18258 21732
rect 17408 21684 17460 21690
rect 17408 21626 17460 21632
rect 17776 21684 17828 21690
rect 17776 21626 17828 21632
rect 17776 21548 17828 21554
rect 17776 21490 17828 21496
rect 17788 21146 17816 21490
rect 18616 21486 18644 22510
rect 18708 21894 18736 22646
rect 18696 21888 18748 21894
rect 18696 21830 18748 21836
rect 18604 21480 18656 21486
rect 18604 21422 18656 21428
rect 17776 21140 17828 21146
rect 17776 21082 17828 21088
rect 18708 20874 18736 21830
rect 18788 21616 18840 21622
rect 18788 21558 18840 21564
rect 18696 20868 18748 20874
rect 18696 20810 18748 20816
rect 17950 20700 18258 20709
rect 17950 20698 17956 20700
rect 18012 20698 18036 20700
rect 18092 20698 18116 20700
rect 18172 20698 18196 20700
rect 18252 20698 18258 20700
rect 18012 20646 18014 20698
rect 18194 20646 18196 20698
rect 17950 20644 17956 20646
rect 18012 20644 18036 20646
rect 18092 20644 18116 20646
rect 18172 20644 18196 20646
rect 18252 20644 18258 20646
rect 17950 20635 18258 20644
rect 18708 20534 18736 20810
rect 18696 20528 18748 20534
rect 18696 20470 18748 20476
rect 18800 20262 18828 21558
rect 18892 21146 18920 22646
rect 18984 22166 19012 26200
rect 19064 24744 19116 24750
rect 19064 24686 19116 24692
rect 19076 23798 19104 24686
rect 19432 24336 19484 24342
rect 19628 24290 19656 26200
rect 20076 24608 20128 24614
rect 20076 24550 20128 24556
rect 19432 24278 19484 24284
rect 19064 23792 19116 23798
rect 19064 23734 19116 23740
rect 19064 22976 19116 22982
rect 19064 22918 19116 22924
rect 18972 22160 19024 22166
rect 18972 22102 19024 22108
rect 19076 21350 19104 22918
rect 19444 22094 19472 24278
rect 19536 24274 19656 24290
rect 19524 24268 19656 24274
rect 19576 24262 19656 24268
rect 19524 24210 19576 24216
rect 20088 23594 20116 24550
rect 20548 24342 20576 26302
rect 20902 26200 20958 27000
rect 21546 26330 21602 27000
rect 22190 26330 22246 27000
rect 21546 26302 21956 26330
rect 21546 26200 21602 26302
rect 20536 24336 20588 24342
rect 20536 24278 20588 24284
rect 20916 24274 20944 26200
rect 21456 24608 21508 24614
rect 21456 24550 21508 24556
rect 20904 24268 20956 24274
rect 20904 24210 20956 24216
rect 20444 23860 20496 23866
rect 20444 23802 20496 23808
rect 20456 23746 20484 23802
rect 20168 23724 20220 23730
rect 20168 23666 20220 23672
rect 20272 23718 20484 23746
rect 20536 23792 20588 23798
rect 20536 23734 20588 23740
rect 20076 23588 20128 23594
rect 20076 23530 20128 23536
rect 20180 22710 20208 23666
rect 20272 23662 20300 23718
rect 20260 23656 20312 23662
rect 20548 23610 20576 23734
rect 21468 23730 21496 24550
rect 21456 23724 21508 23730
rect 21456 23666 21508 23672
rect 20260 23598 20312 23604
rect 20456 23582 20576 23610
rect 20352 23520 20404 23526
rect 20352 23462 20404 23468
rect 20364 23186 20392 23462
rect 20352 23180 20404 23186
rect 20352 23122 20404 23128
rect 20168 22704 20220 22710
rect 20456 22658 20484 23582
rect 20536 23520 20588 23526
rect 20536 23462 20588 23468
rect 21272 23520 21324 23526
rect 21272 23462 21324 23468
rect 20548 22817 20576 23462
rect 20720 23180 20772 23186
rect 20720 23122 20772 23128
rect 20628 23044 20680 23050
rect 20628 22986 20680 22992
rect 20534 22808 20590 22817
rect 20640 22778 20668 22986
rect 20534 22743 20590 22752
rect 20628 22772 20680 22778
rect 20168 22646 20220 22652
rect 20180 22094 20208 22646
rect 20364 22630 20484 22658
rect 20364 22386 20392 22630
rect 20364 22358 20484 22386
rect 19444 22066 19564 22094
rect 20180 22066 20392 22094
rect 19248 21888 19300 21894
rect 19248 21830 19300 21836
rect 19064 21344 19116 21350
rect 19064 21286 19116 21292
rect 18880 21140 18932 21146
rect 18880 21082 18932 21088
rect 18420 20256 18472 20262
rect 18420 20198 18472 20204
rect 18788 20256 18840 20262
rect 18788 20198 18840 20204
rect 17316 19984 17368 19990
rect 17316 19926 17368 19932
rect 17224 19712 17276 19718
rect 17408 19712 17460 19718
rect 17276 19672 17356 19700
rect 17224 19654 17276 19660
rect 17040 19440 17092 19446
rect 17040 19382 17092 19388
rect 17224 19372 17276 19378
rect 17224 19314 17276 19320
rect 17236 18970 17264 19314
rect 17224 18964 17276 18970
rect 17224 18906 17276 18912
rect 17328 18850 17356 19672
rect 17408 19654 17460 19660
rect 18328 19712 18380 19718
rect 18432 19689 18460 20198
rect 18512 19712 18564 19718
rect 18328 19654 18380 19660
rect 18418 19680 18474 19689
rect 17420 19417 17448 19654
rect 17950 19612 18258 19621
rect 17950 19610 17956 19612
rect 18012 19610 18036 19612
rect 18092 19610 18116 19612
rect 18172 19610 18196 19612
rect 18252 19610 18258 19612
rect 18012 19558 18014 19610
rect 18194 19558 18196 19610
rect 17950 19556 17956 19558
rect 18012 19556 18036 19558
rect 18092 19556 18116 19558
rect 18172 19556 18196 19558
rect 18252 19556 18258 19558
rect 17950 19547 18258 19556
rect 17406 19408 17462 19417
rect 17406 19343 17462 19352
rect 17328 18834 17448 18850
rect 17328 18828 17460 18834
rect 17328 18822 17408 18828
rect 17408 18770 17460 18776
rect 18340 18714 18368 19654
rect 18512 19654 18564 19660
rect 18418 19615 18474 19624
rect 18524 18970 18552 19654
rect 18604 19440 18656 19446
rect 18604 19382 18656 19388
rect 18512 18964 18564 18970
rect 18512 18906 18564 18912
rect 18156 18698 18368 18714
rect 18144 18692 18368 18698
rect 18196 18686 18368 18692
rect 18418 18728 18474 18737
rect 18418 18663 18474 18672
rect 18144 18634 18196 18640
rect 18328 18624 18380 18630
rect 18328 18566 18380 18572
rect 17950 18524 18258 18533
rect 17950 18522 17956 18524
rect 18012 18522 18036 18524
rect 18092 18522 18116 18524
rect 18172 18522 18196 18524
rect 18252 18522 18258 18524
rect 18012 18470 18014 18522
rect 18194 18470 18196 18522
rect 17950 18468 17956 18470
rect 18012 18468 18036 18470
rect 18092 18468 18116 18470
rect 18172 18468 18196 18470
rect 18252 18468 18258 18470
rect 17950 18459 18258 18468
rect 17316 18420 17368 18426
rect 17316 18362 17368 18368
rect 17132 17740 17184 17746
rect 17132 17682 17184 17688
rect 16948 16720 17000 16726
rect 16948 16662 17000 16668
rect 17144 16658 17172 17682
rect 17224 17536 17276 17542
rect 17224 17478 17276 17484
rect 17236 16794 17264 17478
rect 17224 16788 17276 16794
rect 17224 16730 17276 16736
rect 17132 16652 17184 16658
rect 17132 16594 17184 16600
rect 16856 16176 16908 16182
rect 16856 16118 16908 16124
rect 16764 15700 16816 15706
rect 16764 15642 16816 15648
rect 16868 14929 16896 16118
rect 16948 15700 17000 15706
rect 16948 15642 17000 15648
rect 16960 15366 16988 15642
rect 16948 15360 17000 15366
rect 16948 15302 17000 15308
rect 17040 15360 17092 15366
rect 17040 15302 17092 15308
rect 16854 14920 16910 14929
rect 16854 14855 16910 14864
rect 16948 14884 17000 14890
rect 16948 14826 17000 14832
rect 16856 14612 16908 14618
rect 16856 14554 16908 14560
rect 16764 14272 16816 14278
rect 16762 14240 16764 14249
rect 16816 14240 16818 14249
rect 16762 14175 16818 14184
rect 16764 14068 16816 14074
rect 16764 14010 16816 14016
rect 16672 11348 16724 11354
rect 16672 11290 16724 11296
rect 16488 11280 16540 11286
rect 16488 11222 16540 11228
rect 16396 10056 16448 10062
rect 16396 9998 16448 10004
rect 16396 8424 16448 8430
rect 16396 8366 16448 8372
rect 16408 6322 16436 8366
rect 16500 7954 16528 11222
rect 16776 11150 16804 14010
rect 16868 12782 16896 14554
rect 16960 14482 16988 14826
rect 16948 14476 17000 14482
rect 16948 14418 17000 14424
rect 16856 12776 16908 12782
rect 16856 12718 16908 12724
rect 16868 12306 16896 12718
rect 16856 12300 16908 12306
rect 16856 12242 16908 12248
rect 16856 12164 16908 12170
rect 16856 12106 16908 12112
rect 16868 11694 16896 12106
rect 16856 11688 16908 11694
rect 16856 11630 16908 11636
rect 16764 11144 16816 11150
rect 16764 11086 16816 11092
rect 16580 10056 16632 10062
rect 16580 9998 16632 10004
rect 16592 8906 16620 9998
rect 16672 9648 16724 9654
rect 16672 9590 16724 9596
rect 16684 8906 16712 9590
rect 16868 9518 16896 11630
rect 16948 11144 17000 11150
rect 16948 11086 17000 11092
rect 16960 10674 16988 11086
rect 16948 10668 17000 10674
rect 16948 10610 17000 10616
rect 16948 9920 17000 9926
rect 16948 9862 17000 9868
rect 16856 9512 16908 9518
rect 16856 9454 16908 9460
rect 16868 9382 16896 9454
rect 16856 9376 16908 9382
rect 16856 9318 16908 9324
rect 16580 8900 16632 8906
rect 16580 8842 16632 8848
rect 16672 8900 16724 8906
rect 16672 8842 16724 8848
rect 16684 8498 16712 8842
rect 16868 8838 16896 9318
rect 16856 8832 16908 8838
rect 16856 8774 16908 8780
rect 16868 8498 16896 8774
rect 16672 8492 16724 8498
rect 16672 8434 16724 8440
rect 16856 8492 16908 8498
rect 16856 8434 16908 8440
rect 16488 7948 16540 7954
rect 16488 7890 16540 7896
rect 16960 7342 16988 9862
rect 17052 9178 17080 15302
rect 17328 14958 17356 18362
rect 18236 18080 18288 18086
rect 18236 18022 18288 18028
rect 17776 17604 17828 17610
rect 17776 17546 17828 17552
rect 17788 17202 17816 17546
rect 18248 17524 18276 18022
rect 18340 17882 18368 18566
rect 18328 17876 18380 17882
rect 18328 17818 18380 17824
rect 18248 17496 18368 17524
rect 17950 17436 18258 17445
rect 17950 17434 17956 17436
rect 18012 17434 18036 17436
rect 18092 17434 18116 17436
rect 18172 17434 18196 17436
rect 18252 17434 18258 17436
rect 18012 17382 18014 17434
rect 18194 17382 18196 17434
rect 17950 17380 17956 17382
rect 18012 17380 18036 17382
rect 18092 17380 18116 17382
rect 18172 17380 18196 17382
rect 18252 17380 18258 17382
rect 17950 17371 18258 17380
rect 17776 17196 17828 17202
rect 17776 17138 17828 17144
rect 17684 16516 17736 16522
rect 17684 16458 17736 16464
rect 17592 15972 17644 15978
rect 17592 15914 17644 15920
rect 17406 15192 17462 15201
rect 17406 15127 17462 15136
rect 17420 14958 17448 15127
rect 17316 14952 17368 14958
rect 17316 14894 17368 14900
rect 17408 14952 17460 14958
rect 17408 14894 17460 14900
rect 17224 14884 17276 14890
rect 17224 14826 17276 14832
rect 17236 14618 17264 14826
rect 17224 14612 17276 14618
rect 17224 14554 17276 14560
rect 17222 14512 17278 14521
rect 17222 14447 17278 14456
rect 17236 12306 17264 14447
rect 17328 13870 17356 14894
rect 17500 14884 17552 14890
rect 17500 14826 17552 14832
rect 17408 14272 17460 14278
rect 17408 14214 17460 14220
rect 17316 13864 17368 13870
rect 17316 13806 17368 13812
rect 17420 13190 17448 14214
rect 17512 14074 17540 14826
rect 17604 14074 17632 15914
rect 17696 15910 17724 16458
rect 17684 15904 17736 15910
rect 17684 15846 17736 15852
rect 17500 14068 17552 14074
rect 17500 14010 17552 14016
rect 17592 14068 17644 14074
rect 17592 14010 17644 14016
rect 17696 13954 17724 15846
rect 17604 13926 17724 13954
rect 17604 13190 17632 13926
rect 17684 13796 17736 13802
rect 17684 13738 17736 13744
rect 17696 13530 17724 13738
rect 17684 13524 17736 13530
rect 17684 13466 17736 13472
rect 17408 13184 17460 13190
rect 17408 13126 17460 13132
rect 17592 13184 17644 13190
rect 17592 13126 17644 13132
rect 17224 12300 17276 12306
rect 17224 12242 17276 12248
rect 17236 12209 17264 12242
rect 17222 12200 17278 12209
rect 17222 12135 17278 12144
rect 17224 12096 17276 12102
rect 17224 12038 17276 12044
rect 17236 11257 17264 12038
rect 17604 11830 17632 13126
rect 17592 11824 17644 11830
rect 17592 11766 17644 11772
rect 17222 11248 17278 11257
rect 17222 11183 17278 11192
rect 17040 9172 17092 9178
rect 17040 9114 17092 9120
rect 16948 7336 17000 7342
rect 16948 7278 17000 7284
rect 16396 6316 16448 6322
rect 16396 6258 16448 6264
rect 16304 6112 16356 6118
rect 16304 6054 16356 6060
rect 15752 5160 15804 5166
rect 15752 5102 15804 5108
rect 16960 3942 16988 7278
rect 17236 5846 17264 11183
rect 17696 10470 17724 13466
rect 17788 12850 17816 17138
rect 18340 16454 18368 17496
rect 18328 16448 18380 16454
rect 18328 16390 18380 16396
rect 17950 16348 18258 16357
rect 17950 16346 17956 16348
rect 18012 16346 18036 16348
rect 18092 16346 18116 16348
rect 18172 16346 18196 16348
rect 18252 16346 18258 16348
rect 18012 16294 18014 16346
rect 18194 16294 18196 16346
rect 17950 16292 17956 16294
rect 18012 16292 18036 16294
rect 18092 16292 18116 16294
rect 18172 16292 18196 16294
rect 18252 16292 18258 16294
rect 17950 16283 18258 16292
rect 17868 16176 17920 16182
rect 17868 16118 17920 16124
rect 17880 14074 17908 16118
rect 18432 15706 18460 18663
rect 18616 18426 18644 19382
rect 18800 19174 18828 20198
rect 18892 19922 18920 21082
rect 18972 20256 19024 20262
rect 18972 20198 19024 20204
rect 18880 19916 18932 19922
rect 18880 19858 18932 19864
rect 18878 19680 18934 19689
rect 18878 19615 18934 19624
rect 18788 19168 18840 19174
rect 18788 19110 18840 19116
rect 18604 18420 18656 18426
rect 18604 18362 18656 18368
rect 18786 18048 18842 18057
rect 18786 17983 18842 17992
rect 18696 17604 18748 17610
rect 18696 17546 18748 17552
rect 18708 17134 18736 17546
rect 18800 17338 18828 17983
rect 18788 17332 18840 17338
rect 18788 17274 18840 17280
rect 18696 17128 18748 17134
rect 18696 17070 18748 17076
rect 18512 16788 18564 16794
rect 18512 16730 18564 16736
rect 18420 15700 18472 15706
rect 18420 15642 18472 15648
rect 18328 15564 18380 15570
rect 18328 15506 18380 15512
rect 17950 15260 18258 15269
rect 17950 15258 17956 15260
rect 18012 15258 18036 15260
rect 18092 15258 18116 15260
rect 18172 15258 18196 15260
rect 18252 15258 18258 15260
rect 18012 15206 18014 15258
rect 18194 15206 18196 15258
rect 17950 15204 17956 15206
rect 18012 15204 18036 15206
rect 18092 15204 18116 15206
rect 18172 15204 18196 15206
rect 18252 15204 18258 15206
rect 17950 15195 18258 15204
rect 18340 15144 18368 15506
rect 18432 15502 18460 15642
rect 18420 15496 18472 15502
rect 18420 15438 18472 15444
rect 18248 15116 18368 15144
rect 18052 15088 18104 15094
rect 18052 15030 18104 15036
rect 18064 14822 18092 15030
rect 18248 15026 18276 15116
rect 18236 15020 18288 15026
rect 18236 14962 18288 14968
rect 18328 15020 18380 15026
rect 18328 14962 18380 14968
rect 18052 14816 18104 14822
rect 18052 14758 18104 14764
rect 17958 14512 18014 14521
rect 17958 14447 18014 14456
rect 17972 14414 18000 14447
rect 17960 14408 18012 14414
rect 17960 14350 18012 14356
rect 17950 14172 18258 14181
rect 17950 14170 17956 14172
rect 18012 14170 18036 14172
rect 18092 14170 18116 14172
rect 18172 14170 18196 14172
rect 18252 14170 18258 14172
rect 18012 14118 18014 14170
rect 18194 14118 18196 14170
rect 17950 14116 17956 14118
rect 18012 14116 18036 14118
rect 18092 14116 18116 14118
rect 18172 14116 18196 14118
rect 18252 14116 18258 14118
rect 17950 14107 18258 14116
rect 17868 14068 17920 14074
rect 17868 14010 17920 14016
rect 17958 13288 18014 13297
rect 17958 13223 18014 13232
rect 17972 13190 18000 13223
rect 17960 13184 18012 13190
rect 17960 13126 18012 13132
rect 17950 13084 18258 13093
rect 17950 13082 17956 13084
rect 18012 13082 18036 13084
rect 18092 13082 18116 13084
rect 18172 13082 18196 13084
rect 18252 13082 18258 13084
rect 18012 13030 18014 13082
rect 18194 13030 18196 13082
rect 17950 13028 17956 13030
rect 18012 13028 18036 13030
rect 18092 13028 18116 13030
rect 18172 13028 18196 13030
rect 18252 13028 18258 13030
rect 17950 13019 18258 13028
rect 17776 12844 17828 12850
rect 17776 12786 17828 12792
rect 17788 12238 17816 12786
rect 18236 12640 18288 12646
rect 18236 12582 18288 12588
rect 18248 12238 18276 12582
rect 17776 12232 17828 12238
rect 17774 12200 17776 12209
rect 18236 12232 18288 12238
rect 17828 12200 17830 12209
rect 18236 12174 18288 12180
rect 17774 12135 17830 12144
rect 17950 11996 18258 12005
rect 17950 11994 17956 11996
rect 18012 11994 18036 11996
rect 18092 11994 18116 11996
rect 18172 11994 18196 11996
rect 18252 11994 18258 11996
rect 18012 11942 18014 11994
rect 18194 11942 18196 11994
rect 17950 11940 17956 11942
rect 18012 11940 18036 11942
rect 18092 11940 18116 11942
rect 18172 11940 18196 11942
rect 18252 11940 18258 11942
rect 17950 11931 18258 11940
rect 18144 11620 18196 11626
rect 18144 11562 18196 11568
rect 17868 11144 17920 11150
rect 17868 11086 17920 11092
rect 17684 10464 17736 10470
rect 17684 10406 17736 10412
rect 17696 10130 17724 10406
rect 17880 10282 17908 11086
rect 18156 11014 18184 11562
rect 18340 11558 18368 14962
rect 18420 14952 18472 14958
rect 18420 14894 18472 14900
rect 18432 14822 18460 14894
rect 18420 14816 18472 14822
rect 18420 14758 18472 14764
rect 18432 13682 18460 14758
rect 18524 13802 18552 16730
rect 18708 16658 18736 17070
rect 18696 16652 18748 16658
rect 18696 16594 18748 16600
rect 18800 16538 18828 17274
rect 18892 16572 18920 19615
rect 18984 18834 19012 20198
rect 18972 18828 19024 18834
rect 18972 18770 19024 18776
rect 19076 18698 19104 21286
rect 19154 20632 19210 20641
rect 19154 20567 19156 20576
rect 19208 20567 19210 20576
rect 19156 20538 19208 20544
rect 19064 18692 19116 18698
rect 19064 18634 19116 18640
rect 18972 18352 19024 18358
rect 18972 18294 19024 18300
rect 18984 17746 19012 18294
rect 18972 17740 19024 17746
rect 18972 17682 19024 17688
rect 19168 17354 19196 20538
rect 19260 19514 19288 21830
rect 19536 20942 19564 22066
rect 20364 21622 20392 22066
rect 20456 21962 20484 22358
rect 20444 21956 20496 21962
rect 20444 21898 20496 21904
rect 20548 21690 20576 22743
rect 20628 22714 20680 22720
rect 20536 21684 20588 21690
rect 20536 21626 20588 21632
rect 20352 21616 20404 21622
rect 20352 21558 20404 21564
rect 20732 21486 20760 23122
rect 20996 22228 21048 22234
rect 20996 22170 21048 22176
rect 21008 21690 21036 22170
rect 21284 22030 21312 23462
rect 21928 23118 21956 26302
rect 22190 26302 22324 26330
rect 22190 26200 22246 26302
rect 22100 24744 22152 24750
rect 22100 24686 22152 24692
rect 22008 23316 22060 23322
rect 22008 23258 22060 23264
rect 21916 23112 21968 23118
rect 21916 23054 21968 23060
rect 22020 23050 22048 23258
rect 22112 23254 22140 24686
rect 22192 24200 22244 24206
rect 22192 24142 22244 24148
rect 22204 23322 22232 24142
rect 22192 23316 22244 23322
rect 22192 23258 22244 23264
rect 22100 23248 22152 23254
rect 22100 23190 22152 23196
rect 22008 23044 22060 23050
rect 22008 22986 22060 22992
rect 22112 22982 22140 23190
rect 22296 23050 22324 26302
rect 22834 26200 22890 27000
rect 23478 26200 23534 27000
rect 24122 26200 24178 27000
rect 24766 26200 24822 27000
rect 25410 26200 25466 27000
rect 26054 26330 26110 27000
rect 26054 26302 26188 26330
rect 26054 26200 26110 26302
rect 22848 23322 22876 26200
rect 22950 24508 23258 24517
rect 22950 24506 22956 24508
rect 23012 24506 23036 24508
rect 23092 24506 23116 24508
rect 23172 24506 23196 24508
rect 23252 24506 23258 24508
rect 23012 24454 23014 24506
rect 23194 24454 23196 24506
rect 22950 24452 22956 24454
rect 23012 24452 23036 24454
rect 23092 24452 23116 24454
rect 23172 24452 23196 24454
rect 23252 24452 23258 24454
rect 22950 24443 23258 24452
rect 23492 23866 23520 26200
rect 24032 24812 24084 24818
rect 24032 24754 24084 24760
rect 24044 24410 24072 24754
rect 24136 24410 24164 26200
rect 24780 24614 24808 26200
rect 24768 24608 24820 24614
rect 24768 24550 24820 24556
rect 24032 24404 24084 24410
rect 24032 24346 24084 24352
rect 24124 24404 24176 24410
rect 24124 24346 24176 24352
rect 23572 24336 23624 24342
rect 23572 24278 23624 24284
rect 24952 24336 25004 24342
rect 24952 24278 25004 24284
rect 23480 23860 23532 23866
rect 23480 23802 23532 23808
rect 23480 23724 23532 23730
rect 23480 23666 23532 23672
rect 23296 23656 23348 23662
rect 23296 23598 23348 23604
rect 22950 23420 23258 23429
rect 22950 23418 22956 23420
rect 23012 23418 23036 23420
rect 23092 23418 23116 23420
rect 23172 23418 23196 23420
rect 23252 23418 23258 23420
rect 23012 23366 23014 23418
rect 23194 23366 23196 23418
rect 22950 23364 22956 23366
rect 23012 23364 23036 23366
rect 23092 23364 23116 23366
rect 23172 23364 23196 23366
rect 23252 23364 23258 23366
rect 22950 23355 23258 23364
rect 22836 23316 22888 23322
rect 22836 23258 22888 23264
rect 23308 23254 23336 23598
rect 23388 23316 23440 23322
rect 23388 23258 23440 23264
rect 23296 23248 23348 23254
rect 23296 23190 23348 23196
rect 22744 23180 22796 23186
rect 22744 23122 22796 23128
rect 22284 23044 22336 23050
rect 22284 22986 22336 22992
rect 21916 22976 21968 22982
rect 21916 22918 21968 22924
rect 22100 22976 22152 22982
rect 22100 22918 22152 22924
rect 22192 22976 22244 22982
rect 22192 22918 22244 22924
rect 21732 22160 21784 22166
rect 21732 22102 21784 22108
rect 21272 22024 21324 22030
rect 21272 21966 21324 21972
rect 21548 21888 21600 21894
rect 21548 21830 21600 21836
rect 20996 21684 21048 21690
rect 20996 21626 21048 21632
rect 20720 21480 20772 21486
rect 20720 21422 20772 21428
rect 20260 21344 20312 21350
rect 20260 21286 20312 21292
rect 19524 20936 19576 20942
rect 19524 20878 19576 20884
rect 19432 20528 19484 20534
rect 19432 20470 19484 20476
rect 19338 19952 19394 19961
rect 19338 19887 19394 19896
rect 19248 19508 19300 19514
rect 19248 19450 19300 19456
rect 19248 18624 19300 18630
rect 19352 18601 19380 19887
rect 19444 19378 19472 20470
rect 19616 20392 19668 20398
rect 19616 20334 19668 20340
rect 19628 19446 19656 20334
rect 19616 19440 19668 19446
rect 19616 19382 19668 19388
rect 19432 19372 19484 19378
rect 19432 19314 19484 19320
rect 19248 18566 19300 18572
rect 19338 18592 19394 18601
rect 19260 18465 19288 18566
rect 19338 18527 19394 18536
rect 19246 18456 19302 18465
rect 19246 18391 19302 18400
rect 19524 18284 19576 18290
rect 19524 18226 19576 18232
rect 19246 17776 19302 17785
rect 19246 17711 19302 17720
rect 19076 17326 19196 17354
rect 18892 16544 19012 16572
rect 18616 16510 18828 16538
rect 18616 14600 18644 16510
rect 18696 16448 18748 16454
rect 18696 16390 18748 16396
rect 18788 16448 18840 16454
rect 18788 16390 18840 16396
rect 18880 16448 18932 16454
rect 18880 16390 18932 16396
rect 18708 16046 18736 16390
rect 18800 16182 18828 16390
rect 18892 16182 18920 16390
rect 18788 16176 18840 16182
rect 18788 16118 18840 16124
rect 18880 16176 18932 16182
rect 18880 16118 18932 16124
rect 18696 16040 18748 16046
rect 18696 15982 18748 15988
rect 18984 15892 19012 16544
rect 18708 15864 19012 15892
rect 18708 15094 18736 15864
rect 19076 15570 19104 17326
rect 19156 17264 19208 17270
rect 19156 17206 19208 17212
rect 19168 15706 19196 17206
rect 19156 15700 19208 15706
rect 19156 15642 19208 15648
rect 19260 15586 19288 17711
rect 19064 15564 19116 15570
rect 19064 15506 19116 15512
rect 19168 15558 19288 15586
rect 18878 15464 18934 15473
rect 18878 15399 18934 15408
rect 18892 15162 18920 15399
rect 18880 15156 18932 15162
rect 18880 15098 18932 15104
rect 18696 15088 18748 15094
rect 18696 15030 18748 15036
rect 18788 15020 18840 15026
rect 18788 14962 18840 14968
rect 18616 14572 18736 14600
rect 18602 14512 18658 14521
rect 18602 14447 18658 14456
rect 18616 14346 18644 14447
rect 18604 14340 18656 14346
rect 18604 14282 18656 14288
rect 18708 14278 18736 14572
rect 18696 14272 18748 14278
rect 18696 14214 18748 14220
rect 18512 13796 18564 13802
rect 18512 13738 18564 13744
rect 18432 13654 18552 13682
rect 18328 11552 18380 11558
rect 18328 11494 18380 11500
rect 18420 11280 18472 11286
rect 18420 11222 18472 11228
rect 18144 11008 18196 11014
rect 18144 10950 18196 10956
rect 17950 10908 18258 10917
rect 17950 10906 17956 10908
rect 18012 10906 18036 10908
rect 18092 10906 18116 10908
rect 18172 10906 18196 10908
rect 18252 10906 18258 10908
rect 18012 10854 18014 10906
rect 18194 10854 18196 10906
rect 17950 10852 17956 10854
rect 18012 10852 18036 10854
rect 18092 10852 18116 10854
rect 18172 10852 18196 10854
rect 18252 10852 18258 10854
rect 17950 10843 18258 10852
rect 17880 10266 18000 10282
rect 17880 10260 18012 10266
rect 17880 10254 17960 10260
rect 17684 10124 17736 10130
rect 17684 10066 17736 10072
rect 17880 9178 17908 10254
rect 17960 10202 18012 10208
rect 17972 9982 18368 10010
rect 17972 9926 18000 9982
rect 17960 9920 18012 9926
rect 17960 9862 18012 9868
rect 17950 9820 18258 9829
rect 17950 9818 17956 9820
rect 18012 9818 18036 9820
rect 18092 9818 18116 9820
rect 18172 9818 18196 9820
rect 18252 9818 18258 9820
rect 18012 9766 18014 9818
rect 18194 9766 18196 9818
rect 17950 9764 17956 9766
rect 18012 9764 18036 9766
rect 18092 9764 18116 9766
rect 18172 9764 18196 9766
rect 18252 9764 18258 9766
rect 17950 9755 18258 9764
rect 18236 9580 18288 9586
rect 18236 9522 18288 9528
rect 17868 9172 17920 9178
rect 17868 9114 17920 9120
rect 17880 8430 17908 9114
rect 18248 8906 18276 9522
rect 18236 8900 18288 8906
rect 18236 8842 18288 8848
rect 17950 8732 18258 8741
rect 17950 8730 17956 8732
rect 18012 8730 18036 8732
rect 18092 8730 18116 8732
rect 18172 8730 18196 8732
rect 18252 8730 18258 8732
rect 18012 8678 18014 8730
rect 18194 8678 18196 8730
rect 17950 8676 17956 8678
rect 18012 8676 18036 8678
rect 18092 8676 18116 8678
rect 18172 8676 18196 8678
rect 18252 8676 18258 8678
rect 17950 8667 18258 8676
rect 17868 8424 17920 8430
rect 17868 8366 17920 8372
rect 18340 7886 18368 9982
rect 18432 9081 18460 11222
rect 18524 11218 18552 13654
rect 18800 13297 18828 14962
rect 18972 13864 19024 13870
rect 18972 13806 19024 13812
rect 18984 13394 19012 13806
rect 18972 13388 19024 13394
rect 18972 13330 19024 13336
rect 18786 13288 18842 13297
rect 18786 13223 18842 13232
rect 18604 13184 18656 13190
rect 18604 13126 18656 13132
rect 18512 11212 18564 11218
rect 18512 11154 18564 11160
rect 18616 10810 18644 13126
rect 18696 12300 18748 12306
rect 18696 12242 18748 12248
rect 18708 11014 18736 12242
rect 18696 11008 18748 11014
rect 18696 10950 18748 10956
rect 18604 10804 18656 10810
rect 18604 10746 18656 10752
rect 18604 9512 18656 9518
rect 18604 9454 18656 9460
rect 18418 9072 18474 9081
rect 18418 9007 18474 9016
rect 18512 9036 18564 9042
rect 18512 8978 18564 8984
rect 18420 8900 18472 8906
rect 18420 8842 18472 8848
rect 18432 8362 18460 8842
rect 18524 8634 18552 8978
rect 18616 8634 18644 9454
rect 18512 8628 18564 8634
rect 18512 8570 18564 8576
rect 18604 8628 18656 8634
rect 18604 8570 18656 8576
rect 18420 8356 18472 8362
rect 18420 8298 18472 8304
rect 18616 7954 18644 8570
rect 18604 7948 18656 7954
rect 18604 7890 18656 7896
rect 18328 7880 18380 7886
rect 18328 7822 18380 7828
rect 17950 7644 18258 7653
rect 17950 7642 17956 7644
rect 18012 7642 18036 7644
rect 18092 7642 18116 7644
rect 18172 7642 18196 7644
rect 18252 7642 18258 7644
rect 18012 7590 18014 7642
rect 18194 7590 18196 7642
rect 17950 7588 17956 7590
rect 18012 7588 18036 7590
rect 18092 7588 18116 7590
rect 18172 7588 18196 7590
rect 18252 7588 18258 7590
rect 17950 7579 18258 7588
rect 17950 6556 18258 6565
rect 17950 6554 17956 6556
rect 18012 6554 18036 6556
rect 18092 6554 18116 6556
rect 18172 6554 18196 6556
rect 18252 6554 18258 6556
rect 18012 6502 18014 6554
rect 18194 6502 18196 6554
rect 17950 6500 17956 6502
rect 18012 6500 18036 6502
rect 18092 6500 18116 6502
rect 18172 6500 18196 6502
rect 18252 6500 18258 6502
rect 17950 6491 18258 6500
rect 18328 6248 18380 6254
rect 18328 6190 18380 6196
rect 17224 5840 17276 5846
rect 17224 5782 17276 5788
rect 17950 5468 18258 5477
rect 17950 5466 17956 5468
rect 18012 5466 18036 5468
rect 18092 5466 18116 5468
rect 18172 5466 18196 5468
rect 18252 5466 18258 5468
rect 18012 5414 18014 5466
rect 18194 5414 18196 5466
rect 17950 5412 17956 5414
rect 18012 5412 18036 5414
rect 18092 5412 18116 5414
rect 18172 5412 18196 5414
rect 18252 5412 18258 5414
rect 17950 5403 18258 5412
rect 17950 4380 18258 4389
rect 17950 4378 17956 4380
rect 18012 4378 18036 4380
rect 18092 4378 18116 4380
rect 18172 4378 18196 4380
rect 18252 4378 18258 4380
rect 18012 4326 18014 4378
rect 18194 4326 18196 4378
rect 17950 4324 17956 4326
rect 18012 4324 18036 4326
rect 18092 4324 18116 4326
rect 18172 4324 18196 4326
rect 18252 4324 18258 4326
rect 17950 4315 18258 4324
rect 18340 4146 18368 6190
rect 18708 5574 18736 10950
rect 18800 7478 18828 13223
rect 18984 12918 19012 13330
rect 18972 12912 19024 12918
rect 18972 12854 19024 12860
rect 18880 11212 18932 11218
rect 18880 11154 18932 11160
rect 18892 9654 18920 11154
rect 19168 11150 19196 15558
rect 19536 15162 19564 18226
rect 19628 17270 19656 19382
rect 19892 19372 19944 19378
rect 19892 19314 19944 19320
rect 19706 18592 19762 18601
rect 19706 18527 19762 18536
rect 19616 17264 19668 17270
rect 19616 17206 19668 17212
rect 19616 16652 19668 16658
rect 19616 16594 19668 16600
rect 19524 15156 19576 15162
rect 19524 15098 19576 15104
rect 19248 14816 19300 14822
rect 19248 14758 19300 14764
rect 19260 14482 19288 14758
rect 19432 14544 19484 14550
rect 19432 14486 19484 14492
rect 19248 14476 19300 14482
rect 19248 14418 19300 14424
rect 19340 14340 19392 14346
rect 19340 14282 19392 14288
rect 19352 13938 19380 14282
rect 19340 13932 19392 13938
rect 19340 13874 19392 13880
rect 19248 12844 19300 12850
rect 19248 12786 19300 12792
rect 19156 11144 19208 11150
rect 19156 11086 19208 11092
rect 18972 11076 19024 11082
rect 18972 11018 19024 11024
rect 18984 10810 19012 11018
rect 18972 10804 19024 10810
rect 18972 10746 19024 10752
rect 19156 10668 19208 10674
rect 19156 10610 19208 10616
rect 18972 10600 19024 10606
rect 18972 10542 19024 10548
rect 18880 9648 18932 9654
rect 18880 9590 18932 9596
rect 18984 9178 19012 10542
rect 19064 10464 19116 10470
rect 19064 10406 19116 10412
rect 19076 10062 19104 10406
rect 19064 10056 19116 10062
rect 19064 9998 19116 10004
rect 18972 9172 19024 9178
rect 18972 9114 19024 9120
rect 19168 8498 19196 10610
rect 19260 10266 19288 12786
rect 19444 10810 19472 14486
rect 19524 14272 19576 14278
rect 19524 14214 19576 14220
rect 19536 14006 19564 14214
rect 19628 14074 19656 16594
rect 19720 14278 19748 18527
rect 19904 17252 19932 19314
rect 20272 17610 20300 21286
rect 20732 20942 20760 21422
rect 20996 21072 21048 21078
rect 20996 21014 21048 21020
rect 20720 20936 20772 20942
rect 20640 20884 20720 20890
rect 20640 20878 20772 20884
rect 20640 20862 20760 20878
rect 20812 20868 20864 20874
rect 20640 20602 20668 20862
rect 20812 20810 20864 20816
rect 20628 20596 20680 20602
rect 20628 20538 20680 20544
rect 20536 19848 20588 19854
rect 20536 19790 20588 19796
rect 20352 19372 20404 19378
rect 20352 19314 20404 19320
rect 20260 17604 20312 17610
rect 20260 17546 20312 17552
rect 19982 17368 20038 17377
rect 19982 17303 20038 17312
rect 19996 17270 20024 17303
rect 19984 17264 20036 17270
rect 19904 17224 19984 17252
rect 19800 16448 19852 16454
rect 19800 16390 19852 16396
rect 19812 16250 19840 16390
rect 19800 16244 19852 16250
rect 19800 16186 19852 16192
rect 19904 16182 19932 17224
rect 19984 17206 20036 17212
rect 20076 17128 20128 17134
rect 20076 17070 20128 17076
rect 20088 16402 20116 17070
rect 20260 16584 20312 16590
rect 20260 16526 20312 16532
rect 20168 16448 20220 16454
rect 20088 16396 20168 16402
rect 20088 16390 20220 16396
rect 20088 16374 20208 16390
rect 19892 16176 19944 16182
rect 19892 16118 19944 16124
rect 19904 15910 19932 16118
rect 19892 15904 19944 15910
rect 19892 15846 19944 15852
rect 19984 15360 20036 15366
rect 19984 15302 20036 15308
rect 19892 14408 19944 14414
rect 19892 14350 19944 14356
rect 19800 14340 19852 14346
rect 19800 14282 19852 14288
rect 19708 14272 19760 14278
rect 19708 14214 19760 14220
rect 19616 14068 19668 14074
rect 19616 14010 19668 14016
rect 19524 14000 19576 14006
rect 19524 13942 19576 13948
rect 19524 12776 19576 12782
rect 19524 12718 19576 12724
rect 19432 10804 19484 10810
rect 19432 10746 19484 10752
rect 19536 10742 19564 12718
rect 19812 11898 19840 14282
rect 19800 11892 19852 11898
rect 19800 11834 19852 11840
rect 19800 11688 19852 11694
rect 19800 11630 19852 11636
rect 19616 11348 19668 11354
rect 19616 11290 19668 11296
rect 19524 10736 19576 10742
rect 19338 10704 19394 10713
rect 19524 10678 19576 10684
rect 19338 10639 19340 10648
rect 19392 10639 19394 10648
rect 19340 10610 19392 10616
rect 19248 10260 19300 10266
rect 19248 10202 19300 10208
rect 19628 9654 19656 11290
rect 19812 11286 19840 11630
rect 19904 11626 19932 14350
rect 19996 12986 20024 15302
rect 20088 14958 20116 16374
rect 20272 16250 20300 16526
rect 20260 16244 20312 16250
rect 20260 16186 20312 16192
rect 20364 15162 20392 19314
rect 20548 19009 20576 19790
rect 20824 19514 20852 20810
rect 21008 20602 21036 21014
rect 20996 20596 21048 20602
rect 20996 20538 21048 20544
rect 20812 19508 20864 19514
rect 20812 19450 20864 19456
rect 20534 19000 20590 19009
rect 20534 18935 20590 18944
rect 20444 18624 20496 18630
rect 20444 18566 20496 18572
rect 20456 15706 20484 18566
rect 20548 17746 20576 18935
rect 21008 18834 21036 20538
rect 21272 20528 21324 20534
rect 21178 20496 21234 20505
rect 21272 20470 21324 20476
rect 21178 20431 21234 20440
rect 21088 19168 21140 19174
rect 21088 19110 21140 19116
rect 21100 18902 21128 19110
rect 21088 18896 21140 18902
rect 21088 18838 21140 18844
rect 20996 18828 21048 18834
rect 20996 18770 21048 18776
rect 20720 18624 20772 18630
rect 21192 18578 21220 20431
rect 21284 19786 21312 20470
rect 21364 20392 21416 20398
rect 21364 20334 21416 20340
rect 21272 19780 21324 19786
rect 21272 19722 21324 19728
rect 21284 18698 21312 19722
rect 21376 19156 21404 20334
rect 21456 19712 21508 19718
rect 21456 19654 21508 19660
rect 21468 19281 21496 19654
rect 21560 19378 21588 21830
rect 21640 21548 21692 21554
rect 21640 21490 21692 21496
rect 21548 19372 21600 19378
rect 21548 19314 21600 19320
rect 21454 19272 21510 19281
rect 21454 19207 21510 19216
rect 21376 19128 21496 19156
rect 21272 18692 21324 18698
rect 21272 18634 21324 18640
rect 20720 18566 20772 18572
rect 20536 17740 20588 17746
rect 20536 17682 20588 17688
rect 20548 16658 20576 17682
rect 20628 17604 20680 17610
rect 20628 17546 20680 17552
rect 20640 17513 20668 17546
rect 20626 17504 20682 17513
rect 20626 17439 20682 17448
rect 20536 16652 20588 16658
rect 20536 16594 20588 16600
rect 20732 16522 20760 18566
rect 21100 18550 21220 18578
rect 21284 18578 21312 18634
rect 21284 18550 21404 18578
rect 20996 18284 21048 18290
rect 20996 18226 21048 18232
rect 20904 18216 20956 18222
rect 20904 18158 20956 18164
rect 20916 17338 20944 18158
rect 21008 17610 21036 18226
rect 20996 17604 21048 17610
rect 20996 17546 21048 17552
rect 21008 17377 21036 17546
rect 20994 17368 21050 17377
rect 20904 17332 20956 17338
rect 20994 17303 21050 17312
rect 20904 17274 20956 17280
rect 21008 16522 21036 17303
rect 20720 16516 20772 16522
rect 20720 16458 20772 16464
rect 20996 16516 21048 16522
rect 20996 16458 21048 16464
rect 20720 16040 20772 16046
rect 20720 15982 20772 15988
rect 20444 15700 20496 15706
rect 20444 15642 20496 15648
rect 20352 15156 20404 15162
rect 20352 15098 20404 15104
rect 20444 15156 20496 15162
rect 20444 15098 20496 15104
rect 20364 14958 20392 15098
rect 20076 14952 20128 14958
rect 20076 14894 20128 14900
rect 20352 14952 20404 14958
rect 20352 14894 20404 14900
rect 20456 14550 20484 15098
rect 20628 14816 20680 14822
rect 20628 14758 20680 14764
rect 20536 14612 20588 14618
rect 20536 14554 20588 14560
rect 20444 14544 20496 14550
rect 20444 14486 20496 14492
rect 20074 14104 20130 14113
rect 20074 14039 20130 14048
rect 20088 14006 20116 14039
rect 20076 14000 20128 14006
rect 20128 13960 20300 13988
rect 20076 13942 20128 13948
rect 20076 13320 20128 13326
rect 20076 13262 20128 13268
rect 20088 12986 20116 13262
rect 19984 12980 20036 12986
rect 19984 12922 20036 12928
rect 20076 12980 20128 12986
rect 20076 12922 20128 12928
rect 20272 12782 20300 13960
rect 20168 12776 20220 12782
rect 20168 12718 20220 12724
rect 20260 12776 20312 12782
rect 20260 12718 20312 12724
rect 20180 12434 20208 12718
rect 20088 12406 20208 12434
rect 19984 12300 20036 12306
rect 19984 12242 20036 12248
rect 19892 11620 19944 11626
rect 19892 11562 19944 11568
rect 19800 11280 19852 11286
rect 19800 11222 19852 11228
rect 19708 10600 19760 10606
rect 19708 10542 19760 10548
rect 19616 9648 19668 9654
rect 19616 9590 19668 9596
rect 19432 8968 19484 8974
rect 19432 8910 19484 8916
rect 19444 8498 19472 8910
rect 19628 8838 19656 9590
rect 19720 8906 19748 10542
rect 19708 8900 19760 8906
rect 19708 8842 19760 8848
rect 19616 8832 19668 8838
rect 19616 8774 19668 8780
rect 19156 8492 19208 8498
rect 19156 8434 19208 8440
rect 19432 8492 19484 8498
rect 19432 8434 19484 8440
rect 19248 8016 19300 8022
rect 19248 7958 19300 7964
rect 18972 7812 19024 7818
rect 18972 7754 19024 7760
rect 18788 7472 18840 7478
rect 18788 7414 18840 7420
rect 18696 5568 18748 5574
rect 18696 5510 18748 5516
rect 18984 5234 19012 7754
rect 19260 6798 19288 7958
rect 19444 7954 19472 8434
rect 19720 8090 19748 8842
rect 19996 8634 20024 12242
rect 20088 11558 20116 12406
rect 20168 11756 20220 11762
rect 20168 11698 20220 11704
rect 20076 11552 20128 11558
rect 20076 11494 20128 11500
rect 20180 11354 20208 11698
rect 20168 11348 20220 11354
rect 20168 11290 20220 11296
rect 20548 10810 20576 14554
rect 20640 14414 20668 14758
rect 20732 14482 20760 15982
rect 20904 15904 20956 15910
rect 20904 15846 20956 15852
rect 20916 15609 20944 15846
rect 20902 15600 20958 15609
rect 20902 15535 20958 15544
rect 21100 15094 21128 18550
rect 21270 18456 21326 18465
rect 21270 18391 21326 18400
rect 21180 18080 21232 18086
rect 21180 18022 21232 18028
rect 21192 16289 21220 18022
rect 21178 16280 21234 16289
rect 21178 16215 21234 16224
rect 20812 15088 20864 15094
rect 20812 15030 20864 15036
rect 21088 15088 21140 15094
rect 21088 15030 21140 15036
rect 21180 15088 21232 15094
rect 21180 15030 21232 15036
rect 20720 14476 20772 14482
rect 20720 14418 20772 14424
rect 20628 14408 20680 14414
rect 20628 14350 20680 14356
rect 20720 12844 20772 12850
rect 20720 12786 20772 12792
rect 20628 12436 20680 12442
rect 20628 12378 20680 12384
rect 20640 11558 20668 12378
rect 20628 11552 20680 11558
rect 20628 11494 20680 11500
rect 20732 10962 20760 12786
rect 20824 12442 20852 15030
rect 20904 15020 20956 15026
rect 20904 14962 20956 14968
rect 20916 13530 20944 14962
rect 20996 14952 21048 14958
rect 20996 14894 21048 14900
rect 20904 13524 20956 13530
rect 20904 13466 20956 13472
rect 20812 12436 20864 12442
rect 20812 12378 20864 12384
rect 21008 11801 21036 14894
rect 21192 13705 21220 15030
rect 21178 13696 21234 13705
rect 21178 13631 21234 13640
rect 21284 13326 21312 18391
rect 21376 18290 21404 18550
rect 21364 18284 21416 18290
rect 21364 18226 21416 18232
rect 21468 18086 21496 19128
rect 21548 18624 21600 18630
rect 21548 18566 21600 18572
rect 21560 18222 21588 18566
rect 21548 18216 21600 18222
rect 21548 18158 21600 18164
rect 21456 18080 21508 18086
rect 21456 18022 21508 18028
rect 21468 15570 21496 18022
rect 21652 17814 21680 21490
rect 21744 20262 21772 22102
rect 21928 21350 21956 22918
rect 22008 22568 22060 22574
rect 22008 22510 22060 22516
rect 22020 21486 22048 22510
rect 22008 21480 22060 21486
rect 22008 21422 22060 21428
rect 21916 21344 21968 21350
rect 21916 21286 21968 21292
rect 22112 21010 22140 22918
rect 22204 21049 22232 22918
rect 22282 22808 22338 22817
rect 22282 22743 22338 22752
rect 22652 22772 22704 22778
rect 22296 22710 22324 22743
rect 22652 22714 22704 22720
rect 22284 22704 22336 22710
rect 22284 22646 22336 22652
rect 22376 22228 22428 22234
rect 22376 22170 22428 22176
rect 22284 21956 22336 21962
rect 22284 21898 22336 21904
rect 22296 21865 22324 21898
rect 22282 21856 22338 21865
rect 22282 21791 22338 21800
rect 22284 21616 22336 21622
rect 22284 21558 22336 21564
rect 22190 21040 22246 21049
rect 22100 21004 22152 21010
rect 22190 20975 22246 20984
rect 22100 20946 22152 20952
rect 22296 20890 22324 21558
rect 22388 21146 22416 22170
rect 22560 21684 22612 21690
rect 22560 21626 22612 21632
rect 22376 21140 22428 21146
rect 22376 21082 22428 21088
rect 22468 21072 22520 21078
rect 22468 21014 22520 21020
rect 22376 21004 22428 21010
rect 22376 20946 22428 20952
rect 21836 20874 22324 20890
rect 21824 20868 22324 20874
rect 21876 20862 22324 20868
rect 21824 20810 21876 20816
rect 21836 20534 21864 20810
rect 22008 20800 22060 20806
rect 22008 20742 22060 20748
rect 22100 20800 22152 20806
rect 22100 20742 22152 20748
rect 21824 20528 21876 20534
rect 21824 20470 21876 20476
rect 21732 20256 21784 20262
rect 21732 20198 21784 20204
rect 21916 20256 21968 20262
rect 21916 20198 21968 20204
rect 21744 20074 21772 20198
rect 21744 20046 21864 20074
rect 21836 19990 21864 20046
rect 21824 19984 21876 19990
rect 21824 19926 21876 19932
rect 21824 18896 21876 18902
rect 21824 18838 21876 18844
rect 21640 17808 21692 17814
rect 21640 17750 21692 17756
rect 21836 17524 21864 18838
rect 21928 17882 21956 20198
rect 22020 18086 22048 20742
rect 22112 20602 22140 20742
rect 22100 20596 22152 20602
rect 22100 20538 22152 20544
rect 22388 20482 22416 20946
rect 22112 20454 22416 20482
rect 22112 18170 22140 20454
rect 22376 20324 22428 20330
rect 22376 20266 22428 20272
rect 22388 19334 22416 20266
rect 22204 19306 22416 19334
rect 22204 18834 22232 19306
rect 22480 19242 22508 21014
rect 22572 21010 22600 21626
rect 22560 21004 22612 21010
rect 22560 20946 22612 20952
rect 22560 20528 22612 20534
rect 22560 20470 22612 20476
rect 22468 19236 22520 19242
rect 22468 19178 22520 19184
rect 22282 19000 22338 19009
rect 22282 18935 22338 18944
rect 22192 18828 22244 18834
rect 22192 18770 22244 18776
rect 22296 18766 22324 18935
rect 22284 18760 22336 18766
rect 22284 18702 22336 18708
rect 22296 18358 22324 18702
rect 22374 18456 22430 18465
rect 22374 18391 22430 18400
rect 22284 18352 22336 18358
rect 22284 18294 22336 18300
rect 22388 18290 22416 18391
rect 22376 18284 22428 18290
rect 22376 18226 22428 18232
rect 22468 18216 22520 18222
rect 22112 18142 22232 18170
rect 22468 18158 22520 18164
rect 22008 18080 22060 18086
rect 22008 18022 22060 18028
rect 21916 17876 21968 17882
rect 21916 17818 21968 17824
rect 22204 17785 22232 18142
rect 22190 17776 22246 17785
rect 22190 17711 22246 17720
rect 22480 17626 22508 18158
rect 22192 17604 22244 17610
rect 22192 17546 22244 17552
rect 22388 17598 22508 17626
rect 21916 17536 21968 17542
rect 21836 17496 21916 17524
rect 21916 17478 21968 17484
rect 21928 16794 21956 17478
rect 22008 16992 22060 16998
rect 22008 16934 22060 16940
rect 22020 16794 22048 16934
rect 21916 16788 21968 16794
rect 21916 16730 21968 16736
rect 22008 16788 22060 16794
rect 22008 16730 22060 16736
rect 21640 15632 21692 15638
rect 21640 15574 21692 15580
rect 21364 15564 21416 15570
rect 21364 15506 21416 15512
rect 21456 15564 21508 15570
rect 21456 15506 21508 15512
rect 21376 14482 21404 15506
rect 21548 15360 21600 15366
rect 21548 15302 21600 15308
rect 21364 14476 21416 14482
rect 21364 14418 21416 14424
rect 21456 14476 21508 14482
rect 21456 14418 21508 14424
rect 21376 14074 21404 14418
rect 21468 14346 21496 14418
rect 21456 14340 21508 14346
rect 21456 14282 21508 14288
rect 21364 14068 21416 14074
rect 21364 14010 21416 14016
rect 21456 13388 21508 13394
rect 21456 13330 21508 13336
rect 21272 13320 21324 13326
rect 21272 13262 21324 13268
rect 21272 12776 21324 12782
rect 21272 12718 21324 12724
rect 21180 12096 21232 12102
rect 21180 12038 21232 12044
rect 20994 11792 21050 11801
rect 20994 11727 21050 11736
rect 20732 10934 20944 10962
rect 20536 10804 20588 10810
rect 20536 10746 20588 10752
rect 20720 10804 20772 10810
rect 20720 10746 20772 10752
rect 20626 10704 20682 10713
rect 20732 10690 20760 10746
rect 20682 10662 20760 10690
rect 20626 10639 20682 10648
rect 20260 10124 20312 10130
rect 20260 10066 20312 10072
rect 19984 8628 20036 8634
rect 19984 8570 20036 8576
rect 19708 8084 19760 8090
rect 19708 8026 19760 8032
rect 19432 7948 19484 7954
rect 19432 7890 19484 7896
rect 19996 7818 20024 8570
rect 20272 8566 20300 10066
rect 20812 9988 20864 9994
rect 20812 9930 20864 9936
rect 20824 9518 20852 9930
rect 20812 9512 20864 9518
rect 20812 9454 20864 9460
rect 20916 9382 20944 10934
rect 21008 10266 21036 11727
rect 20996 10260 21048 10266
rect 20996 10202 21048 10208
rect 21088 9648 21140 9654
rect 21088 9590 21140 9596
rect 20996 9580 21048 9586
rect 20996 9522 21048 9528
rect 20904 9376 20956 9382
rect 20904 9318 20956 9324
rect 21008 9042 21036 9522
rect 20996 9036 21048 9042
rect 20996 8978 21048 8984
rect 21100 8906 21128 9590
rect 21088 8900 21140 8906
rect 21088 8842 21140 8848
rect 20260 8560 20312 8566
rect 20260 8502 20312 8508
rect 21100 8498 21128 8842
rect 21088 8492 21140 8498
rect 21088 8434 21140 8440
rect 21100 8294 21128 8434
rect 21088 8288 21140 8294
rect 21088 8230 21140 8236
rect 21100 7818 21128 8230
rect 19984 7812 20036 7818
rect 19984 7754 20036 7760
rect 21088 7812 21140 7818
rect 21088 7754 21140 7760
rect 21192 7546 21220 12038
rect 21284 11354 21312 12718
rect 21468 12306 21496 13330
rect 21456 12300 21508 12306
rect 21456 12242 21508 12248
rect 21456 11688 21508 11694
rect 21456 11630 21508 11636
rect 21272 11348 21324 11354
rect 21272 11290 21324 11296
rect 21468 11218 21496 11630
rect 21560 11558 21588 15302
rect 21652 14074 21680 15574
rect 21732 15360 21784 15366
rect 21732 15302 21784 15308
rect 21744 15201 21772 15302
rect 21730 15192 21786 15201
rect 21730 15127 21732 15136
rect 21784 15127 21786 15136
rect 21732 15098 21784 15104
rect 22100 15020 22152 15026
rect 22100 14962 22152 14968
rect 21640 14068 21692 14074
rect 21640 14010 21692 14016
rect 22008 13864 22060 13870
rect 22008 13806 22060 13812
rect 21640 13320 21692 13326
rect 21640 13262 21692 13268
rect 21548 11552 21600 11558
rect 21548 11494 21600 11500
rect 21456 11212 21508 11218
rect 21456 11154 21508 11160
rect 21180 7540 21232 7546
rect 21180 7482 21232 7488
rect 20444 7200 20496 7206
rect 20444 7142 20496 7148
rect 19248 6792 19300 6798
rect 19248 6734 19300 6740
rect 19616 6112 19668 6118
rect 19616 6054 19668 6060
rect 18972 5228 19024 5234
rect 18972 5170 19024 5176
rect 19156 5160 19208 5166
rect 19156 5102 19208 5108
rect 18328 4140 18380 4146
rect 18328 4082 18380 4088
rect 16948 3936 17000 3942
rect 16948 3878 17000 3884
rect 18340 3534 18368 4082
rect 14740 3528 14792 3534
rect 14740 3470 14792 3476
rect 18328 3528 18380 3534
rect 18328 3470 18380 3476
rect 18420 3528 18472 3534
rect 18420 3470 18472 3476
rect 17868 3460 17920 3466
rect 17868 3402 17920 3408
rect 17224 3392 17276 3398
rect 17224 3334 17276 3340
rect 17236 3194 17264 3334
rect 17224 3188 17276 3194
rect 17224 3130 17276 3136
rect 17880 2990 17908 3402
rect 17950 3292 18258 3301
rect 17950 3290 17956 3292
rect 18012 3290 18036 3292
rect 18092 3290 18116 3292
rect 18172 3290 18196 3292
rect 18252 3290 18258 3292
rect 18012 3238 18014 3290
rect 18194 3238 18196 3290
rect 17950 3236 17956 3238
rect 18012 3236 18036 3238
rect 18092 3236 18116 3238
rect 18172 3236 18196 3238
rect 18252 3236 18258 3238
rect 17950 3227 18258 3236
rect 18432 3194 18460 3470
rect 18420 3188 18472 3194
rect 18420 3130 18472 3136
rect 19168 3126 19196 5102
rect 19524 4616 19576 4622
rect 19524 4558 19576 4564
rect 19156 3120 19208 3126
rect 19156 3062 19208 3068
rect 17868 2984 17920 2990
rect 17868 2926 17920 2932
rect 18420 2984 18472 2990
rect 18420 2926 18472 2932
rect 16396 2848 16448 2854
rect 16396 2790 16448 2796
rect 15936 2508 15988 2514
rect 15936 2450 15988 2456
rect 14648 2372 14700 2378
rect 14648 2314 14700 2320
rect 15948 800 15976 2450
rect 16408 2446 16436 2790
rect 16396 2440 16448 2446
rect 16396 2382 16448 2388
rect 17950 2204 18258 2213
rect 17950 2202 17956 2204
rect 18012 2202 18036 2204
rect 18092 2202 18116 2204
rect 18172 2202 18196 2204
rect 18252 2202 18258 2204
rect 18012 2150 18014 2202
rect 18194 2150 18196 2202
rect 17950 2148 17956 2150
rect 18012 2148 18036 2150
rect 18092 2148 18116 2150
rect 18172 2148 18196 2150
rect 18252 2148 18258 2150
rect 17950 2139 18258 2148
rect 18064 870 18184 898
rect 18064 800 18092 870
rect 1122 0 1178 800
rect 3238 0 3294 800
rect 5354 0 5410 800
rect 7470 0 7526 800
rect 9586 0 9642 800
rect 11702 0 11758 800
rect 13818 0 13874 800
rect 15934 0 15990 800
rect 18050 0 18106 800
rect 18156 762 18184 870
rect 18432 762 18460 2926
rect 19536 2446 19564 4558
rect 19628 2446 19656 6054
rect 20456 4690 20484 7142
rect 20812 5024 20864 5030
rect 20812 4966 20864 4972
rect 20444 4684 20496 4690
rect 20444 4626 20496 4632
rect 20720 4276 20772 4282
rect 20720 4218 20772 4224
rect 20732 3602 20760 4218
rect 20720 3596 20772 3602
rect 20720 3538 20772 3544
rect 20824 3058 20852 4966
rect 21456 4480 21508 4486
rect 21456 4422 21508 4428
rect 20904 3528 20956 3534
rect 20904 3470 20956 3476
rect 20812 3052 20864 3058
rect 20812 2994 20864 3000
rect 20916 2990 20944 3470
rect 21180 3460 21232 3466
rect 21180 3402 21232 3408
rect 20904 2984 20956 2990
rect 20904 2926 20956 2932
rect 21192 2854 21220 3402
rect 21468 3058 21496 4422
rect 21652 4282 21680 13262
rect 21916 12844 21968 12850
rect 21916 12786 21968 12792
rect 21824 11144 21876 11150
rect 21824 11086 21876 11092
rect 21732 10736 21784 10742
rect 21732 10678 21784 10684
rect 21744 10266 21772 10678
rect 21732 10260 21784 10266
rect 21732 10202 21784 10208
rect 21836 9994 21864 11086
rect 21824 9988 21876 9994
rect 21824 9930 21876 9936
rect 21928 8090 21956 12786
rect 22020 11694 22048 13806
rect 22112 12442 22140 14962
rect 22204 13530 22232 17546
rect 22282 15600 22338 15609
rect 22282 15535 22338 15544
rect 22296 13870 22324 15535
rect 22388 14385 22416 17598
rect 22468 17536 22520 17542
rect 22468 17478 22520 17484
rect 22480 16794 22508 17478
rect 22468 16788 22520 16794
rect 22468 16730 22520 16736
rect 22468 16652 22520 16658
rect 22468 16594 22520 16600
rect 22480 14550 22508 16594
rect 22572 15162 22600 20470
rect 22664 18222 22692 22714
rect 22756 22710 22784 23122
rect 22744 22704 22796 22710
rect 22744 22646 22796 22652
rect 22756 21622 22784 22646
rect 22950 22332 23258 22341
rect 22950 22330 22956 22332
rect 23012 22330 23036 22332
rect 23092 22330 23116 22332
rect 23172 22330 23196 22332
rect 23252 22330 23258 22332
rect 23012 22278 23014 22330
rect 23194 22278 23196 22330
rect 22950 22276 22956 22278
rect 23012 22276 23036 22278
rect 23092 22276 23116 22278
rect 23172 22276 23196 22278
rect 23252 22276 23258 22278
rect 22950 22267 23258 22276
rect 23204 22228 23256 22234
rect 23204 22170 23256 22176
rect 23216 22098 23244 22170
rect 23400 22166 23428 23258
rect 23388 22160 23440 22166
rect 23388 22102 23440 22108
rect 23204 22092 23256 22098
rect 23204 22034 23256 22040
rect 23386 21992 23442 22001
rect 23386 21927 23442 21936
rect 22836 21888 22888 21894
rect 22836 21830 22888 21836
rect 23112 21888 23164 21894
rect 23112 21830 23164 21836
rect 22744 21616 22796 21622
rect 22744 21558 22796 21564
rect 22848 19990 22876 21830
rect 23124 21690 23152 21830
rect 23112 21684 23164 21690
rect 23112 21626 23164 21632
rect 23400 21486 23428 21927
rect 23492 21894 23520 23666
rect 23480 21888 23532 21894
rect 23480 21830 23532 21836
rect 23388 21480 23440 21486
rect 23388 21422 23440 21428
rect 22950 21244 23258 21253
rect 22950 21242 22956 21244
rect 23012 21242 23036 21244
rect 23092 21242 23116 21244
rect 23172 21242 23196 21244
rect 23252 21242 23258 21244
rect 23012 21190 23014 21242
rect 23194 21190 23196 21242
rect 22950 21188 22956 21190
rect 23012 21188 23036 21190
rect 23092 21188 23116 21190
rect 23172 21188 23196 21190
rect 23252 21188 23258 21190
rect 22950 21179 23258 21188
rect 23296 20800 23348 20806
rect 23296 20742 23348 20748
rect 22950 20156 23258 20165
rect 22950 20154 22956 20156
rect 23012 20154 23036 20156
rect 23092 20154 23116 20156
rect 23172 20154 23196 20156
rect 23252 20154 23258 20156
rect 23012 20102 23014 20154
rect 23194 20102 23196 20154
rect 22950 20100 22956 20102
rect 23012 20100 23036 20102
rect 23092 20100 23116 20102
rect 23172 20100 23196 20102
rect 23252 20100 23258 20102
rect 22950 20091 23258 20100
rect 23308 20058 23336 20742
rect 23388 20392 23440 20398
rect 23388 20334 23440 20340
rect 23296 20052 23348 20058
rect 23296 19994 23348 20000
rect 22836 19984 22888 19990
rect 22836 19926 22888 19932
rect 22744 19712 22796 19718
rect 22744 19654 22796 19660
rect 22836 19712 22888 19718
rect 22836 19654 22888 19660
rect 22756 18873 22784 19654
rect 22742 18864 22798 18873
rect 22742 18799 22798 18808
rect 22744 18352 22796 18358
rect 22744 18294 22796 18300
rect 22652 18216 22704 18222
rect 22652 18158 22704 18164
rect 22652 17672 22704 17678
rect 22652 17614 22704 17620
rect 22664 17338 22692 17614
rect 22652 17332 22704 17338
rect 22652 17274 22704 17280
rect 22756 17202 22784 18294
rect 22848 17882 22876 19654
rect 23400 19378 23428 20334
rect 23388 19372 23440 19378
rect 23584 19334 23612 24278
rect 24964 24177 24992 24278
rect 25136 24268 25188 24274
rect 25136 24210 25188 24216
rect 24950 24168 25006 24177
rect 24950 24103 25006 24112
rect 24860 23656 24912 23662
rect 25148 23610 25176 24210
rect 25424 24206 25452 26200
rect 26054 24848 26110 24857
rect 26054 24783 26110 24792
rect 26068 24206 26096 24783
rect 26160 24342 26188 26302
rect 26698 26200 26754 27000
rect 27342 26200 27398 27000
rect 27986 26200 28042 27000
rect 28630 26330 28686 27000
rect 28630 26302 28948 26330
rect 28630 26200 28686 26302
rect 26330 24712 26386 24721
rect 26330 24647 26386 24656
rect 26148 24336 26200 24342
rect 26148 24278 26200 24284
rect 26344 24274 26372 24647
rect 26332 24268 26384 24274
rect 26332 24210 26384 24216
rect 26712 24206 26740 26200
rect 25412 24200 25464 24206
rect 25412 24142 25464 24148
rect 26056 24200 26108 24206
rect 26056 24142 26108 24148
rect 26700 24200 26752 24206
rect 26700 24142 26752 24148
rect 26424 24132 26476 24138
rect 26424 24074 26476 24080
rect 27252 24132 27304 24138
rect 27252 24074 27304 24080
rect 26240 24064 26292 24070
rect 26240 24006 26292 24012
rect 25228 23792 25280 23798
rect 25228 23734 25280 23740
rect 24860 23598 24912 23604
rect 24768 23588 24820 23594
rect 24768 23530 24820 23536
rect 24780 23361 24808 23530
rect 24766 23352 24822 23361
rect 24766 23287 24822 23296
rect 24676 23044 24728 23050
rect 24676 22986 24728 22992
rect 23664 22976 23716 22982
rect 23664 22918 23716 22924
rect 23676 22574 23704 22918
rect 23664 22568 23716 22574
rect 23664 22510 23716 22516
rect 23664 22432 23716 22438
rect 24688 22409 24716 22986
rect 24872 22778 24900 23598
rect 25056 23582 25176 23610
rect 24950 23216 25006 23225
rect 24950 23151 25006 23160
rect 24964 23118 24992 23151
rect 24952 23112 25004 23118
rect 24952 23054 25004 23060
rect 24768 22772 24820 22778
rect 24768 22714 24820 22720
rect 24860 22772 24912 22778
rect 24860 22714 24912 22720
rect 23664 22374 23716 22380
rect 24674 22400 24730 22409
rect 23676 20534 23704 22374
rect 24674 22335 24730 22344
rect 24780 22098 24808 22714
rect 24872 22642 24900 22714
rect 25056 22710 25084 23582
rect 25240 23526 25268 23734
rect 26252 23633 26280 24006
rect 26436 23882 26464 24074
rect 26344 23854 26464 23882
rect 26238 23624 26294 23633
rect 26238 23559 26294 23568
rect 25136 23520 25188 23526
rect 25136 23462 25188 23468
rect 25228 23520 25280 23526
rect 25228 23462 25280 23468
rect 25148 23254 25176 23462
rect 25136 23248 25188 23254
rect 25136 23190 25188 23196
rect 25688 23112 25740 23118
rect 25688 23054 25740 23060
rect 25320 23044 25372 23050
rect 25320 22986 25372 22992
rect 25136 22976 25188 22982
rect 25136 22918 25188 22924
rect 25148 22710 25176 22918
rect 25044 22704 25096 22710
rect 25044 22646 25096 22652
rect 25136 22704 25188 22710
rect 25136 22646 25188 22652
rect 24860 22636 24912 22642
rect 24860 22578 24912 22584
rect 24584 22092 24636 22098
rect 24584 22034 24636 22040
rect 24768 22092 24820 22098
rect 24768 22034 24820 22040
rect 23940 22024 23992 22030
rect 23940 21966 23992 21972
rect 23756 21412 23808 21418
rect 23756 21354 23808 21360
rect 23768 20874 23796 21354
rect 23756 20868 23808 20874
rect 23756 20810 23808 20816
rect 23664 20528 23716 20534
rect 23664 20470 23716 20476
rect 23756 20460 23808 20466
rect 23756 20402 23808 20408
rect 23664 20256 23716 20262
rect 23664 20198 23716 20204
rect 23388 19314 23440 19320
rect 23296 19304 23348 19310
rect 23296 19246 23348 19252
rect 23492 19306 23612 19334
rect 23676 19310 23704 20198
rect 22950 19068 23258 19077
rect 22950 19066 22956 19068
rect 23012 19066 23036 19068
rect 23092 19066 23116 19068
rect 23172 19066 23196 19068
rect 23252 19066 23258 19068
rect 23012 19014 23014 19066
rect 23194 19014 23196 19066
rect 22950 19012 22956 19014
rect 23012 19012 23036 19014
rect 23092 19012 23116 19014
rect 23172 19012 23196 19014
rect 23252 19012 23258 19014
rect 22950 19003 23258 19012
rect 23020 18692 23072 18698
rect 23020 18634 23072 18640
rect 23032 18154 23060 18634
rect 23308 18290 23336 19246
rect 23492 19174 23520 19306
rect 23664 19304 23716 19310
rect 23664 19246 23716 19252
rect 23480 19168 23532 19174
rect 23480 19110 23532 19116
rect 23296 18284 23348 18290
rect 23296 18226 23348 18232
rect 23020 18148 23072 18154
rect 23020 18090 23072 18096
rect 22950 17980 23258 17989
rect 22950 17978 22956 17980
rect 23012 17978 23036 17980
rect 23092 17978 23116 17980
rect 23172 17978 23196 17980
rect 23252 17978 23258 17980
rect 23012 17926 23014 17978
rect 23194 17926 23196 17978
rect 22950 17924 22956 17926
rect 23012 17924 23036 17926
rect 23092 17924 23116 17926
rect 23172 17924 23196 17926
rect 23252 17924 23258 17926
rect 22950 17915 23258 17924
rect 22836 17876 22888 17882
rect 22836 17818 22888 17824
rect 23112 17604 23164 17610
rect 23112 17546 23164 17552
rect 23124 17270 23152 17546
rect 23112 17264 23164 17270
rect 23112 17206 23164 17212
rect 22744 17196 22796 17202
rect 22744 17138 22796 17144
rect 22744 16992 22796 16998
rect 22744 16934 22796 16940
rect 22560 15156 22612 15162
rect 22560 15098 22612 15104
rect 22652 14952 22704 14958
rect 22652 14894 22704 14900
rect 22468 14544 22520 14550
rect 22468 14486 22520 14492
rect 22374 14376 22430 14385
rect 22374 14311 22430 14320
rect 22284 13864 22336 13870
rect 22284 13806 22336 13812
rect 22192 13524 22244 13530
rect 22192 13466 22244 13472
rect 22192 12640 22244 12646
rect 22192 12582 22244 12588
rect 22100 12436 22152 12442
rect 22100 12378 22152 12384
rect 22204 12238 22232 12582
rect 22192 12232 22244 12238
rect 22192 12174 22244 12180
rect 22296 11830 22324 13806
rect 22480 13394 22508 14486
rect 22558 14376 22614 14385
rect 22558 14311 22614 14320
rect 22468 13388 22520 13394
rect 22468 13330 22520 13336
rect 22572 13274 22600 14311
rect 22480 13246 22600 13274
rect 22376 13184 22428 13190
rect 22376 13126 22428 13132
rect 22388 12753 22416 13126
rect 22374 12744 22430 12753
rect 22374 12679 22430 12688
rect 22284 11824 22336 11830
rect 22284 11766 22336 11772
rect 22008 11688 22060 11694
rect 22008 11630 22060 11636
rect 22284 11620 22336 11626
rect 22284 11562 22336 11568
rect 22100 11552 22152 11558
rect 22100 11494 22152 11500
rect 22008 10600 22060 10606
rect 22008 10542 22060 10548
rect 22020 10130 22048 10542
rect 22008 10124 22060 10130
rect 22008 10066 22060 10072
rect 22020 9042 22048 10066
rect 22008 9036 22060 9042
rect 22008 8978 22060 8984
rect 22020 8498 22048 8978
rect 22008 8492 22060 8498
rect 22008 8434 22060 8440
rect 21916 8084 21968 8090
rect 21916 8026 21968 8032
rect 21824 7812 21876 7818
rect 21824 7754 21876 7760
rect 21836 4434 21864 7754
rect 21916 6656 21968 6662
rect 21916 6598 21968 6604
rect 21928 4690 21956 6598
rect 21916 4684 21968 4690
rect 21916 4626 21968 4632
rect 21836 4406 21956 4434
rect 21640 4276 21692 4282
rect 21640 4218 21692 4224
rect 21928 3602 21956 4406
rect 21916 3596 21968 3602
rect 21916 3538 21968 3544
rect 21928 3466 21956 3538
rect 21916 3460 21968 3466
rect 21916 3402 21968 3408
rect 21456 3052 21508 3058
rect 21456 2994 21508 3000
rect 22020 2990 22048 8434
rect 22112 7698 22140 11494
rect 22296 9178 22324 11562
rect 22284 9172 22336 9178
rect 22284 9114 22336 9120
rect 22192 8968 22244 8974
rect 22192 8910 22244 8916
rect 22204 7886 22232 8910
rect 22296 8566 22324 9114
rect 22284 8560 22336 8566
rect 22284 8502 22336 8508
rect 22192 7880 22244 7886
rect 22192 7822 22244 7828
rect 22112 7670 22232 7698
rect 22100 4616 22152 4622
rect 22100 4558 22152 4564
rect 22112 4078 22140 4558
rect 22100 4072 22152 4078
rect 22100 4014 22152 4020
rect 22112 3126 22140 4014
rect 22204 3505 22232 7670
rect 22388 7546 22416 12679
rect 22480 12186 22508 13246
rect 22560 12776 22612 12782
rect 22560 12718 22612 12724
rect 22572 12306 22600 12718
rect 22664 12646 22692 14894
rect 22756 14890 22784 16934
rect 22950 16892 23258 16901
rect 22950 16890 22956 16892
rect 23012 16890 23036 16892
rect 23092 16890 23116 16892
rect 23172 16890 23196 16892
rect 23252 16890 23258 16892
rect 23012 16838 23014 16890
rect 23194 16838 23196 16890
rect 22950 16836 22956 16838
rect 23012 16836 23036 16838
rect 23092 16836 23116 16838
rect 23172 16836 23196 16838
rect 23252 16836 23258 16838
rect 22950 16827 23258 16836
rect 22836 16448 22888 16454
rect 22836 16390 22888 16396
rect 22848 15502 22876 16390
rect 22950 15804 23258 15813
rect 22950 15802 22956 15804
rect 23012 15802 23036 15804
rect 23092 15802 23116 15804
rect 23172 15802 23196 15804
rect 23252 15802 23258 15804
rect 23012 15750 23014 15802
rect 23194 15750 23196 15802
rect 22950 15748 22956 15750
rect 23012 15748 23036 15750
rect 23092 15748 23116 15750
rect 23172 15748 23196 15750
rect 23252 15748 23258 15750
rect 22950 15739 23258 15748
rect 22836 15496 22888 15502
rect 22836 15438 22888 15444
rect 22744 14884 22796 14890
rect 22744 14826 22796 14832
rect 22950 14716 23258 14725
rect 22950 14714 22956 14716
rect 23012 14714 23036 14716
rect 23092 14714 23116 14716
rect 23172 14714 23196 14716
rect 23252 14714 23258 14716
rect 23012 14662 23014 14714
rect 23194 14662 23196 14714
rect 22950 14660 22956 14662
rect 23012 14660 23036 14662
rect 23092 14660 23116 14662
rect 23172 14660 23196 14662
rect 23252 14660 23258 14662
rect 22950 14651 23258 14660
rect 22744 14340 22796 14346
rect 22744 14282 22796 14288
rect 22756 14006 22784 14282
rect 22744 14000 22796 14006
rect 22744 13942 22796 13948
rect 22836 13728 22888 13734
rect 22836 13670 22888 13676
rect 22848 13530 22876 13670
rect 22950 13628 23258 13637
rect 22950 13626 22956 13628
rect 23012 13626 23036 13628
rect 23092 13626 23116 13628
rect 23172 13626 23196 13628
rect 23252 13626 23258 13628
rect 23012 13574 23014 13626
rect 23194 13574 23196 13626
rect 22950 13572 22956 13574
rect 23012 13572 23036 13574
rect 23092 13572 23116 13574
rect 23172 13572 23196 13574
rect 23252 13572 23258 13574
rect 22950 13563 23258 13572
rect 22836 13524 22888 13530
rect 22836 13466 22888 13472
rect 23204 13320 23256 13326
rect 23204 13262 23256 13268
rect 22836 12844 22888 12850
rect 22836 12786 22888 12792
rect 22652 12640 22704 12646
rect 22652 12582 22704 12588
rect 22560 12300 22612 12306
rect 22560 12242 22612 12248
rect 22480 12158 22600 12186
rect 22466 12064 22522 12073
rect 22466 11999 22522 12008
rect 22480 11830 22508 11999
rect 22468 11824 22520 11830
rect 22468 11766 22520 11772
rect 22480 10062 22508 11766
rect 22468 10056 22520 10062
rect 22468 9998 22520 10004
rect 22572 9654 22600 12158
rect 22848 11558 22876 12786
rect 23216 12782 23244 13262
rect 23204 12776 23256 12782
rect 23204 12718 23256 12724
rect 22950 12540 23258 12549
rect 22950 12538 22956 12540
rect 23012 12538 23036 12540
rect 23092 12538 23116 12540
rect 23172 12538 23196 12540
rect 23252 12538 23258 12540
rect 23012 12486 23014 12538
rect 23194 12486 23196 12538
rect 22950 12484 22956 12486
rect 23012 12484 23036 12486
rect 23092 12484 23116 12486
rect 23172 12484 23196 12486
rect 23252 12484 23258 12486
rect 22950 12475 23258 12484
rect 23204 12436 23256 12442
rect 23204 12378 23256 12384
rect 23216 12102 23244 12378
rect 23308 12374 23336 18226
rect 23480 18148 23532 18154
rect 23480 18090 23532 18096
rect 23492 17270 23520 18090
rect 23676 17746 23704 19246
rect 23768 18154 23796 20402
rect 23848 19848 23900 19854
rect 23848 19790 23900 19796
rect 23860 18630 23888 19790
rect 23952 19514 23980 21966
rect 24216 21480 24268 21486
rect 24216 21422 24268 21428
rect 24228 20777 24256 21422
rect 24214 20768 24270 20777
rect 24214 20703 24270 20712
rect 24124 20528 24176 20534
rect 24124 20470 24176 20476
rect 24136 20398 24164 20470
rect 24124 20392 24176 20398
rect 24124 20334 24176 20340
rect 24136 20058 24164 20334
rect 24124 20052 24176 20058
rect 24124 19994 24176 20000
rect 23940 19508 23992 19514
rect 23940 19450 23992 19456
rect 23848 18624 23900 18630
rect 23848 18566 23900 18572
rect 23756 18148 23808 18154
rect 23756 18090 23808 18096
rect 23848 18080 23900 18086
rect 23848 18022 23900 18028
rect 23940 18080 23992 18086
rect 23940 18022 23992 18028
rect 23860 17882 23888 18022
rect 23848 17876 23900 17882
rect 23848 17818 23900 17824
rect 23664 17740 23716 17746
rect 23664 17682 23716 17688
rect 23664 17536 23716 17542
rect 23664 17478 23716 17484
rect 23756 17536 23808 17542
rect 23756 17478 23808 17484
rect 23480 17264 23532 17270
rect 23480 17206 23532 17212
rect 23388 16992 23440 16998
rect 23388 16934 23440 16940
rect 23572 16992 23624 16998
rect 23572 16934 23624 16940
rect 23400 16454 23428 16934
rect 23584 16658 23612 16934
rect 23676 16794 23704 17478
rect 23664 16788 23716 16794
rect 23664 16730 23716 16736
rect 23572 16652 23624 16658
rect 23572 16594 23624 16600
rect 23388 16448 23440 16454
rect 23388 16390 23440 16396
rect 23388 16108 23440 16114
rect 23388 16050 23440 16056
rect 23296 12368 23348 12374
rect 23296 12310 23348 12316
rect 23204 12096 23256 12102
rect 23204 12038 23256 12044
rect 23308 11830 23336 12310
rect 23400 12102 23428 16050
rect 23480 16040 23532 16046
rect 23480 15982 23532 15988
rect 23492 15706 23520 15982
rect 23480 15700 23532 15706
rect 23480 15642 23532 15648
rect 23664 15564 23716 15570
rect 23664 15506 23716 15512
rect 23572 14340 23624 14346
rect 23572 14282 23624 14288
rect 23584 14006 23612 14282
rect 23676 14113 23704 15506
rect 23768 15162 23796 17478
rect 23952 16726 23980 18022
rect 23940 16720 23992 16726
rect 23940 16662 23992 16668
rect 23848 15904 23900 15910
rect 23848 15846 23900 15852
rect 23756 15156 23808 15162
rect 23756 15098 23808 15104
rect 23662 14104 23718 14113
rect 23718 14062 23796 14090
rect 23662 14039 23718 14048
rect 23572 14000 23624 14006
rect 23572 13942 23624 13948
rect 23664 13864 23716 13870
rect 23664 13806 23716 13812
rect 23572 13388 23624 13394
rect 23572 13330 23624 13336
rect 23480 13184 23532 13190
rect 23480 13126 23532 13132
rect 23388 12096 23440 12102
rect 23388 12038 23440 12044
rect 23296 11824 23348 11830
rect 23296 11766 23348 11772
rect 23388 11824 23440 11830
rect 23388 11766 23440 11772
rect 22836 11552 22888 11558
rect 22836 11494 22888 11500
rect 23296 11552 23348 11558
rect 23296 11494 23348 11500
rect 22950 11452 23258 11461
rect 22950 11450 22956 11452
rect 23012 11450 23036 11452
rect 23092 11450 23116 11452
rect 23172 11450 23196 11452
rect 23252 11450 23258 11452
rect 23012 11398 23014 11450
rect 23194 11398 23196 11450
rect 22950 11396 22956 11398
rect 23012 11396 23036 11398
rect 23092 11396 23116 11398
rect 23172 11396 23196 11398
rect 23252 11396 23258 11398
rect 22950 11387 23258 11396
rect 23308 11257 23336 11494
rect 23294 11248 23350 11257
rect 23400 11218 23428 11766
rect 23492 11354 23520 13126
rect 23480 11348 23532 11354
rect 23480 11290 23532 11296
rect 23294 11183 23296 11192
rect 23348 11183 23350 11192
rect 23388 11212 23440 11218
rect 23296 11154 23348 11160
rect 23388 11154 23440 11160
rect 23296 11076 23348 11082
rect 23296 11018 23348 11024
rect 22950 10364 23258 10373
rect 22950 10362 22956 10364
rect 23012 10362 23036 10364
rect 23092 10362 23116 10364
rect 23172 10362 23196 10364
rect 23252 10362 23258 10364
rect 23012 10310 23014 10362
rect 23194 10310 23196 10362
rect 22950 10308 22956 10310
rect 23012 10308 23036 10310
rect 23092 10308 23116 10310
rect 23172 10308 23196 10310
rect 23252 10308 23258 10310
rect 22950 10299 23258 10308
rect 23308 10266 23336 11018
rect 23388 10668 23440 10674
rect 23388 10610 23440 10616
rect 23296 10260 23348 10266
rect 23296 10202 23348 10208
rect 23400 9994 23428 10610
rect 23388 9988 23440 9994
rect 23388 9930 23440 9936
rect 23400 9674 23428 9930
rect 23584 9926 23612 13330
rect 23676 12238 23704 13806
rect 23768 13802 23796 14062
rect 23756 13796 23808 13802
rect 23756 13738 23808 13744
rect 23860 13394 23888 15846
rect 24136 14958 24164 19994
rect 24596 18970 24624 22034
rect 25228 21956 25280 21962
rect 25228 21898 25280 21904
rect 24952 21888 25004 21894
rect 25136 21888 25188 21894
rect 25004 21836 25136 21842
rect 24952 21830 25188 21836
rect 24964 21814 25176 21830
rect 24768 21684 24820 21690
rect 24768 21626 24820 21632
rect 24780 20942 24808 21626
rect 25136 21548 25188 21554
rect 25136 21490 25188 21496
rect 25148 21457 25176 21490
rect 25134 21448 25190 21457
rect 25134 21383 25190 21392
rect 24768 20936 24820 20942
rect 25044 20936 25096 20942
rect 24768 20878 24820 20884
rect 25042 20904 25044 20913
rect 25096 20904 25098 20913
rect 25042 20839 25098 20848
rect 24952 20800 25004 20806
rect 24952 20742 25004 20748
rect 24674 19272 24730 19281
rect 24674 19207 24730 19216
rect 24688 18970 24716 19207
rect 24584 18964 24636 18970
rect 24584 18906 24636 18912
rect 24676 18964 24728 18970
rect 24676 18906 24728 18912
rect 24492 18828 24544 18834
rect 24492 18770 24544 18776
rect 24306 17776 24362 17785
rect 24306 17711 24362 17720
rect 24320 17270 24348 17711
rect 24308 17264 24360 17270
rect 24308 17206 24360 17212
rect 24504 17134 24532 18770
rect 24860 18624 24912 18630
rect 24860 18566 24912 18572
rect 24674 18048 24730 18057
rect 24674 17983 24730 17992
rect 24492 17128 24544 17134
rect 24492 17070 24544 17076
rect 24492 16176 24544 16182
rect 24490 16144 24492 16153
rect 24544 16144 24546 16153
rect 24490 16079 24546 16088
rect 24688 15502 24716 17983
rect 24872 16017 24900 18566
rect 24964 18193 24992 20742
rect 25148 20505 25176 21383
rect 25134 20496 25190 20505
rect 25134 20431 25190 20440
rect 25240 20330 25268 21898
rect 25332 20942 25360 22986
rect 25594 22672 25650 22681
rect 25594 22607 25650 22616
rect 25504 22160 25556 22166
rect 25504 22102 25556 22108
rect 25412 21480 25464 21486
rect 25412 21422 25464 21428
rect 25320 20936 25372 20942
rect 25320 20878 25372 20884
rect 25320 20800 25372 20806
rect 25320 20742 25372 20748
rect 25228 20324 25280 20330
rect 25228 20266 25280 20272
rect 25136 19916 25188 19922
rect 25136 19858 25188 19864
rect 25148 19514 25176 19858
rect 25136 19508 25188 19514
rect 25136 19450 25188 19456
rect 25042 19136 25098 19145
rect 25042 19071 25098 19080
rect 25056 18834 25084 19071
rect 25044 18828 25096 18834
rect 25044 18770 25096 18776
rect 25056 18601 25084 18770
rect 25148 18698 25176 19450
rect 25332 18902 25360 20742
rect 25424 20602 25452 21422
rect 25412 20596 25464 20602
rect 25412 20538 25464 20544
rect 25516 20466 25544 22102
rect 25504 20460 25556 20466
rect 25504 20402 25556 20408
rect 25608 20398 25636 22607
rect 25596 20392 25648 20398
rect 25596 20334 25648 20340
rect 25596 20256 25648 20262
rect 25596 20198 25648 20204
rect 25608 19922 25636 20198
rect 25596 19916 25648 19922
rect 25596 19858 25648 19864
rect 25320 18896 25372 18902
rect 25320 18838 25372 18844
rect 25700 18834 25728 23054
rect 26148 22500 26200 22506
rect 26148 22442 26200 22448
rect 26160 22098 26188 22442
rect 26148 22092 26200 22098
rect 26344 22094 26372 23854
rect 26424 23792 26476 23798
rect 26424 23734 26476 23740
rect 26436 23050 26464 23734
rect 27160 23724 27212 23730
rect 27160 23666 27212 23672
rect 26608 23520 26660 23526
rect 26608 23462 26660 23468
rect 26620 23186 26648 23462
rect 26608 23180 26660 23186
rect 26608 23122 26660 23128
rect 26976 23180 27028 23186
rect 26976 23122 27028 23128
rect 26698 23080 26754 23089
rect 26424 23044 26476 23050
rect 26698 23015 26754 23024
rect 26424 22986 26476 22992
rect 26436 22710 26464 22986
rect 26424 22704 26476 22710
rect 26424 22646 26476 22652
rect 26608 22432 26660 22438
rect 26608 22374 26660 22380
rect 26422 22264 26478 22273
rect 26422 22199 26478 22208
rect 26436 22098 26464 22199
rect 26620 22166 26648 22374
rect 26608 22160 26660 22166
rect 26608 22102 26660 22108
rect 26148 22034 26200 22040
rect 26252 22066 26372 22094
rect 26424 22092 26476 22098
rect 26252 21894 26280 22066
rect 26424 22034 26476 22040
rect 25872 21888 25924 21894
rect 25872 21830 25924 21836
rect 26240 21888 26292 21894
rect 26240 21830 26292 21836
rect 26516 21888 26568 21894
rect 26608 21888 26660 21894
rect 26516 21830 26568 21836
rect 26606 21856 26608 21865
rect 26660 21856 26662 21865
rect 25884 20505 25912 21830
rect 26148 21344 26200 21350
rect 26148 21286 26200 21292
rect 26240 21344 26292 21350
rect 26240 21286 26292 21292
rect 26160 21078 26188 21286
rect 26148 21072 26200 21078
rect 26148 21014 26200 21020
rect 26252 20806 26280 21286
rect 26422 21040 26478 21049
rect 26332 21004 26384 21010
rect 26422 20975 26478 20984
rect 26332 20946 26384 20952
rect 26240 20800 26292 20806
rect 26240 20742 26292 20748
rect 25870 20496 25926 20505
rect 25870 20431 25926 20440
rect 26146 20360 26202 20369
rect 26056 20324 26108 20330
rect 26146 20295 26202 20304
rect 26056 20266 26108 20272
rect 25962 20224 26018 20233
rect 25962 20159 26018 20168
rect 25976 19417 26004 20159
rect 25962 19408 26018 19417
rect 25872 19372 25924 19378
rect 25962 19343 26018 19352
rect 25872 19314 25924 19320
rect 25780 19168 25832 19174
rect 25780 19110 25832 19116
rect 25688 18828 25740 18834
rect 25688 18770 25740 18776
rect 25136 18692 25188 18698
rect 25136 18634 25188 18640
rect 25042 18592 25098 18601
rect 25042 18527 25098 18536
rect 25700 18358 25728 18770
rect 25792 18426 25820 19110
rect 25780 18420 25832 18426
rect 25780 18362 25832 18368
rect 25688 18352 25740 18358
rect 25688 18294 25740 18300
rect 25504 18216 25556 18222
rect 24950 18184 25006 18193
rect 25504 18158 25556 18164
rect 24950 18119 25006 18128
rect 25412 17672 25464 17678
rect 25412 17614 25464 17620
rect 25320 17196 25372 17202
rect 25320 17138 25372 17144
rect 25228 17128 25280 17134
rect 25228 17070 25280 17076
rect 25136 16516 25188 16522
rect 25136 16458 25188 16464
rect 25044 16040 25096 16046
rect 24858 16008 24914 16017
rect 25044 15982 25096 15988
rect 24858 15943 24914 15952
rect 24858 15600 24914 15609
rect 24858 15535 24860 15544
rect 24912 15535 24914 15544
rect 24860 15506 24912 15512
rect 24676 15496 24728 15502
rect 24676 15438 24728 15444
rect 24860 15088 24912 15094
rect 24860 15030 24912 15036
rect 24400 15020 24452 15026
rect 24400 14962 24452 14968
rect 24124 14952 24176 14958
rect 24124 14894 24176 14900
rect 24412 14482 24440 14962
rect 24768 14884 24820 14890
rect 24768 14826 24820 14832
rect 24400 14476 24452 14482
rect 24400 14418 24452 14424
rect 23940 13728 23992 13734
rect 23940 13670 23992 13676
rect 23848 13388 23900 13394
rect 23848 13330 23900 13336
rect 23952 12986 23980 13670
rect 24216 13252 24268 13258
rect 24216 13194 24268 13200
rect 23940 12980 23992 12986
rect 23940 12922 23992 12928
rect 23940 12776 23992 12782
rect 23940 12718 23992 12724
rect 23756 12300 23808 12306
rect 23756 12242 23808 12248
rect 23664 12232 23716 12238
rect 23664 12174 23716 12180
rect 23768 12102 23796 12242
rect 23756 12096 23808 12102
rect 23754 12064 23756 12073
rect 23808 12064 23810 12073
rect 23754 11999 23810 12008
rect 23848 11756 23900 11762
rect 23848 11698 23900 11704
rect 23664 11688 23716 11694
rect 23664 11630 23716 11636
rect 23676 11218 23704 11630
rect 23664 11212 23716 11218
rect 23664 11154 23716 11160
rect 23572 9920 23624 9926
rect 23572 9862 23624 9868
rect 22560 9648 22612 9654
rect 22560 9590 22612 9596
rect 23308 9646 23428 9674
rect 23584 9654 23612 9862
rect 23572 9648 23624 9654
rect 22950 9276 23258 9285
rect 22950 9274 22956 9276
rect 23012 9274 23036 9276
rect 23092 9274 23116 9276
rect 23172 9274 23196 9276
rect 23252 9274 23258 9276
rect 23012 9222 23014 9274
rect 23194 9222 23196 9274
rect 22950 9220 22956 9222
rect 23012 9220 23036 9222
rect 23092 9220 23116 9222
rect 23172 9220 23196 9222
rect 23252 9220 23258 9222
rect 22950 9211 23258 9220
rect 23308 8906 23336 9646
rect 23572 9590 23624 9596
rect 23676 9586 23704 11154
rect 23756 11144 23808 11150
rect 23756 11086 23808 11092
rect 23768 10538 23796 11086
rect 23756 10532 23808 10538
rect 23756 10474 23808 10480
rect 23664 9580 23716 9586
rect 23664 9522 23716 9528
rect 23296 8900 23348 8906
rect 23296 8842 23348 8848
rect 23308 8480 23336 8842
rect 23388 8492 23440 8498
rect 23308 8452 23388 8480
rect 23388 8434 23440 8440
rect 22652 8288 22704 8294
rect 22652 8230 22704 8236
rect 22376 7540 22428 7546
rect 22376 7482 22428 7488
rect 22664 7342 22692 8230
rect 22950 8188 23258 8197
rect 22950 8186 22956 8188
rect 23012 8186 23036 8188
rect 23092 8186 23116 8188
rect 23172 8186 23196 8188
rect 23252 8186 23258 8188
rect 23012 8134 23014 8186
rect 23194 8134 23196 8186
rect 22950 8132 22956 8134
rect 23012 8132 23036 8134
rect 23092 8132 23116 8134
rect 23172 8132 23196 8134
rect 23252 8132 23258 8134
rect 22950 8123 23258 8132
rect 22744 7744 22796 7750
rect 22744 7686 22796 7692
rect 22652 7336 22704 7342
rect 22652 7278 22704 7284
rect 22652 4140 22704 4146
rect 22652 4082 22704 4088
rect 22664 3534 22692 4082
rect 22652 3528 22704 3534
rect 22190 3496 22246 3505
rect 22652 3470 22704 3476
rect 22756 3482 22784 7686
rect 22950 7100 23258 7109
rect 22950 7098 22956 7100
rect 23012 7098 23036 7100
rect 23092 7098 23116 7100
rect 23172 7098 23196 7100
rect 23252 7098 23258 7100
rect 23012 7046 23014 7098
rect 23194 7046 23196 7098
rect 22950 7044 22956 7046
rect 23012 7044 23036 7046
rect 23092 7044 23116 7046
rect 23172 7044 23196 7046
rect 23252 7044 23258 7046
rect 22950 7035 23258 7044
rect 22950 6012 23258 6021
rect 22950 6010 22956 6012
rect 23012 6010 23036 6012
rect 23092 6010 23116 6012
rect 23172 6010 23196 6012
rect 23252 6010 23258 6012
rect 23012 5958 23014 6010
rect 23194 5958 23196 6010
rect 22950 5956 22956 5958
rect 23012 5956 23036 5958
rect 23092 5956 23116 5958
rect 23172 5956 23196 5958
rect 23252 5956 23258 5958
rect 22950 5947 23258 5956
rect 22950 4924 23258 4933
rect 22950 4922 22956 4924
rect 23012 4922 23036 4924
rect 23092 4922 23116 4924
rect 23172 4922 23196 4924
rect 23252 4922 23258 4924
rect 23012 4870 23014 4922
rect 23194 4870 23196 4922
rect 22950 4868 22956 4870
rect 23012 4868 23036 4870
rect 23092 4868 23116 4870
rect 23172 4868 23196 4870
rect 23252 4868 23258 4870
rect 22950 4859 23258 4868
rect 22950 3836 23258 3845
rect 22950 3834 22956 3836
rect 23012 3834 23036 3836
rect 23092 3834 23116 3836
rect 23172 3834 23196 3836
rect 23252 3834 23258 3836
rect 23012 3782 23014 3834
rect 23194 3782 23196 3834
rect 22950 3780 22956 3782
rect 23012 3780 23036 3782
rect 23092 3780 23116 3782
rect 23172 3780 23196 3782
rect 23252 3780 23258 3782
rect 22950 3771 23258 3780
rect 23400 3670 23428 8434
rect 23768 7954 23796 10474
rect 23860 9110 23888 11698
rect 23952 11694 23980 12718
rect 23940 11688 23992 11694
rect 23940 11630 23992 11636
rect 24228 10810 24256 13194
rect 24308 12776 24360 12782
rect 24308 12718 24360 12724
rect 24320 12238 24348 12718
rect 24308 12232 24360 12238
rect 24308 12174 24360 12180
rect 24216 10804 24268 10810
rect 24216 10746 24268 10752
rect 23848 9104 23900 9110
rect 23848 9046 23900 9052
rect 23756 7948 23808 7954
rect 23756 7890 23808 7896
rect 24032 5228 24084 5234
rect 24032 5170 24084 5176
rect 23664 4616 23716 4622
rect 23664 4558 23716 4564
rect 23388 3664 23440 3670
rect 23388 3606 23440 3612
rect 23572 3528 23624 3534
rect 22190 3431 22246 3440
rect 22756 3454 23428 3482
rect 23572 3470 23624 3476
rect 22100 3120 22152 3126
rect 22100 3062 22152 3068
rect 22652 3120 22704 3126
rect 22652 3062 22704 3068
rect 22008 2984 22060 2990
rect 22008 2926 22060 2932
rect 22664 2922 22692 3062
rect 22376 2916 22428 2922
rect 22376 2858 22428 2864
rect 22652 2916 22704 2922
rect 22652 2858 22704 2864
rect 21180 2848 21232 2854
rect 21180 2790 21232 2796
rect 20168 2508 20220 2514
rect 20168 2450 20220 2456
rect 22284 2508 22336 2514
rect 22284 2450 22336 2456
rect 19524 2440 19576 2446
rect 19524 2382 19576 2388
rect 19616 2440 19668 2446
rect 19616 2382 19668 2388
rect 20180 800 20208 2450
rect 22296 800 22324 2450
rect 22388 2446 22416 2858
rect 22756 2774 22784 3454
rect 23400 3398 23428 3454
rect 23296 3392 23348 3398
rect 23296 3334 23348 3340
rect 23388 3392 23440 3398
rect 23388 3334 23440 3340
rect 23112 3188 23164 3194
rect 23112 3130 23164 3136
rect 23124 2922 23152 3130
rect 23308 3126 23336 3334
rect 23584 3194 23612 3470
rect 23572 3188 23624 3194
rect 23572 3130 23624 3136
rect 23296 3120 23348 3126
rect 23296 3062 23348 3068
rect 23112 2916 23164 2922
rect 23112 2858 23164 2864
rect 23308 2854 23336 3062
rect 23676 2854 23704 4558
rect 24044 3602 24072 5170
rect 24308 5024 24360 5030
rect 24308 4966 24360 4972
rect 24320 4078 24348 4966
rect 24412 4078 24440 14418
rect 24676 14000 24728 14006
rect 24674 13968 24676 13977
rect 24728 13968 24730 13977
rect 24674 13903 24730 13912
rect 24584 12232 24636 12238
rect 24584 12174 24636 12180
rect 24596 11218 24624 12174
rect 24584 11212 24636 11218
rect 24584 11154 24636 11160
rect 24676 10600 24728 10606
rect 24676 10542 24728 10548
rect 24688 10266 24716 10542
rect 24780 10538 24808 14826
rect 24872 14822 24900 15030
rect 24860 14816 24912 14822
rect 24860 14758 24912 14764
rect 24952 14816 25004 14822
rect 24952 14758 25004 14764
rect 24964 14550 24992 14758
rect 24952 14544 25004 14550
rect 24952 14486 25004 14492
rect 24952 14408 25004 14414
rect 24952 14350 25004 14356
rect 24860 14340 24912 14346
rect 24860 14282 24912 14288
rect 24872 13938 24900 14282
rect 24860 13932 24912 13938
rect 24860 13874 24912 13880
rect 24860 13388 24912 13394
rect 24860 13330 24912 13336
rect 24872 11694 24900 13330
rect 24964 13326 24992 14350
rect 24952 13320 25004 13326
rect 24952 13262 25004 13268
rect 25056 12986 25084 15982
rect 25148 15162 25176 16458
rect 25136 15156 25188 15162
rect 25136 15098 25188 15104
rect 25136 14816 25188 14822
rect 25136 14758 25188 14764
rect 25044 12980 25096 12986
rect 25044 12922 25096 12928
rect 25056 12434 25084 12922
rect 24964 12406 25084 12434
rect 24964 12170 24992 12406
rect 24952 12164 25004 12170
rect 24952 12106 25004 12112
rect 24860 11688 24912 11694
rect 24860 11630 24912 11636
rect 24872 11218 24900 11630
rect 24860 11212 24912 11218
rect 24860 11154 24912 11160
rect 24860 10600 24912 10606
rect 24860 10542 24912 10548
rect 24768 10532 24820 10538
rect 24768 10474 24820 10480
rect 24676 10260 24728 10266
rect 24676 10202 24728 10208
rect 24688 4758 24716 10202
rect 24872 9994 24900 10542
rect 24860 9988 24912 9994
rect 24860 9930 24912 9936
rect 25044 9580 25096 9586
rect 25044 9522 25096 9528
rect 24952 8832 25004 8838
rect 24952 8774 25004 8780
rect 24964 7478 24992 8774
rect 25056 8498 25084 9522
rect 25148 8906 25176 14758
rect 25240 14006 25268 17070
rect 25228 14000 25280 14006
rect 25228 13942 25280 13948
rect 25332 13530 25360 17138
rect 25424 16658 25452 17614
rect 25412 16652 25464 16658
rect 25412 16594 25464 16600
rect 25424 16250 25452 16594
rect 25516 16590 25544 18158
rect 25686 17640 25742 17649
rect 25884 17626 25912 19314
rect 26068 19292 26096 20266
rect 26160 19446 26188 20295
rect 26148 19440 26200 19446
rect 26146 19408 26148 19417
rect 26240 19440 26292 19446
rect 26200 19408 26202 19417
rect 26240 19382 26292 19388
rect 26146 19343 26202 19352
rect 26068 19264 26188 19292
rect 25964 18216 26016 18222
rect 25964 18158 26016 18164
rect 25686 17575 25688 17584
rect 25740 17575 25742 17584
rect 25792 17598 25912 17626
rect 25688 17546 25740 17552
rect 25596 17536 25648 17542
rect 25596 17478 25648 17484
rect 25608 17241 25636 17478
rect 25594 17232 25650 17241
rect 25594 17167 25650 17176
rect 25608 16998 25636 17167
rect 25792 17066 25820 17598
rect 25872 17536 25924 17542
rect 25872 17478 25924 17484
rect 25780 17060 25832 17066
rect 25780 17002 25832 17008
rect 25596 16992 25648 16998
rect 25596 16934 25648 16940
rect 25884 16658 25912 17478
rect 25872 16652 25924 16658
rect 25872 16594 25924 16600
rect 25504 16584 25556 16590
rect 25504 16526 25556 16532
rect 25412 16244 25464 16250
rect 25412 16186 25464 16192
rect 25780 16176 25832 16182
rect 25780 16118 25832 16124
rect 25410 15464 25466 15473
rect 25410 15399 25412 15408
rect 25464 15399 25466 15408
rect 25412 15370 25464 15376
rect 25424 14822 25452 15370
rect 25688 15088 25740 15094
rect 25688 15030 25740 15036
rect 25504 15020 25556 15026
rect 25504 14962 25556 14968
rect 25412 14816 25464 14822
rect 25412 14758 25464 14764
rect 25516 14618 25544 14962
rect 25504 14612 25556 14618
rect 25504 14554 25556 14560
rect 25412 14476 25464 14482
rect 25412 14418 25464 14424
rect 25424 14006 25452 14418
rect 25596 14340 25648 14346
rect 25516 14300 25596 14328
rect 25412 14000 25464 14006
rect 25412 13942 25464 13948
rect 25516 13870 25544 14300
rect 25596 14282 25648 14288
rect 25504 13864 25556 13870
rect 25504 13806 25556 13812
rect 25320 13524 25372 13530
rect 25320 13466 25372 13472
rect 25516 13394 25544 13806
rect 25504 13388 25556 13394
rect 25504 13330 25556 13336
rect 25596 13320 25648 13326
rect 25596 13262 25648 13268
rect 25320 13184 25372 13190
rect 25320 13126 25372 13132
rect 25332 12889 25360 13126
rect 25318 12880 25374 12889
rect 25318 12815 25374 12824
rect 25412 12844 25464 12850
rect 25412 12786 25464 12792
rect 25424 12170 25452 12786
rect 25412 12164 25464 12170
rect 25412 12106 25464 12112
rect 25320 11756 25372 11762
rect 25424 11744 25452 12106
rect 25608 12102 25636 13262
rect 25700 12424 25728 15030
rect 25792 14346 25820 16118
rect 25884 14958 25912 16594
rect 25976 16454 26004 18158
rect 26056 18080 26108 18086
rect 26054 18048 26056 18057
rect 26108 18048 26110 18057
rect 26054 17983 26110 17992
rect 26160 17270 26188 19264
rect 26252 18290 26280 19382
rect 26240 18284 26292 18290
rect 26240 18226 26292 18232
rect 26344 17746 26372 20946
rect 26436 20806 26464 20975
rect 26424 20800 26476 20806
rect 26424 20742 26476 20748
rect 26528 19174 26556 21830
rect 26606 21791 26662 21800
rect 26608 20596 26660 20602
rect 26608 20538 26660 20544
rect 26620 19514 26648 20538
rect 26608 19508 26660 19514
rect 26608 19450 26660 19456
rect 26516 19168 26568 19174
rect 26516 19110 26568 19116
rect 26620 18698 26648 19450
rect 26608 18692 26660 18698
rect 26608 18634 26660 18640
rect 26516 18216 26568 18222
rect 26516 18158 26568 18164
rect 26332 17740 26384 17746
rect 26332 17682 26384 17688
rect 26344 17513 26372 17682
rect 26330 17504 26386 17513
rect 26330 17439 26386 17448
rect 26148 17264 26200 17270
rect 26148 17206 26200 17212
rect 26240 16652 26292 16658
rect 26240 16594 26292 16600
rect 26054 16552 26110 16561
rect 26252 16538 26280 16594
rect 26110 16510 26280 16538
rect 26054 16487 26110 16496
rect 25964 16448 26016 16454
rect 25964 16390 26016 16396
rect 25976 16250 26004 16390
rect 25964 16244 26016 16250
rect 25964 16186 26016 16192
rect 26068 15502 26096 16487
rect 26330 16280 26386 16289
rect 26330 16215 26332 16224
rect 26384 16215 26386 16224
rect 26332 16186 26384 16192
rect 26148 16108 26200 16114
rect 26148 16050 26200 16056
rect 26160 16017 26188 16050
rect 26146 16008 26202 16017
rect 26146 15943 26202 15952
rect 26528 15706 26556 18158
rect 26620 17513 26648 18634
rect 26606 17504 26662 17513
rect 26606 17439 26662 17448
rect 26620 16522 26648 17439
rect 26608 16516 26660 16522
rect 26608 16458 26660 16464
rect 26620 16182 26648 16458
rect 26608 16176 26660 16182
rect 26608 16118 26660 16124
rect 26516 15700 26568 15706
rect 26516 15642 26568 15648
rect 26238 15600 26294 15609
rect 26238 15535 26294 15544
rect 26424 15564 26476 15570
rect 26252 15502 26280 15535
rect 26424 15506 26476 15512
rect 26516 15564 26568 15570
rect 26516 15506 26568 15512
rect 26056 15496 26108 15502
rect 26056 15438 26108 15444
rect 26240 15496 26292 15502
rect 26240 15438 26292 15444
rect 26148 15428 26200 15434
rect 26148 15370 26200 15376
rect 26160 15065 26188 15370
rect 26146 15056 26202 15065
rect 26146 14991 26202 15000
rect 25872 14952 25924 14958
rect 26148 14952 26200 14958
rect 25872 14894 25924 14900
rect 26146 14920 26148 14929
rect 26200 14920 26202 14929
rect 26146 14855 26202 14864
rect 26056 14612 26108 14618
rect 26056 14554 26108 14560
rect 25780 14340 25832 14346
rect 25780 14282 25832 14288
rect 25792 14006 25820 14282
rect 26068 14074 26096 14554
rect 26056 14068 26108 14074
rect 26056 14010 26108 14016
rect 25780 14000 25832 14006
rect 25778 13968 25780 13977
rect 25832 13968 25834 13977
rect 25778 13903 25834 13912
rect 25792 12850 25820 13903
rect 26252 13734 26280 15438
rect 26332 14816 26384 14822
rect 26332 14758 26384 14764
rect 26240 13728 26292 13734
rect 26240 13670 26292 13676
rect 26238 12880 26294 12889
rect 25780 12844 25832 12850
rect 26238 12815 26294 12824
rect 25780 12786 25832 12792
rect 25872 12436 25924 12442
rect 25700 12396 25872 12424
rect 25596 12096 25648 12102
rect 25596 12038 25648 12044
rect 25372 11716 25452 11744
rect 25320 11698 25372 11704
rect 25332 11082 25360 11698
rect 25320 11076 25372 11082
rect 25320 11018 25372 11024
rect 25332 9994 25360 11018
rect 25596 10532 25648 10538
rect 25596 10474 25648 10480
rect 25320 9988 25372 9994
rect 25320 9930 25372 9936
rect 25332 9586 25360 9930
rect 25608 9722 25636 10474
rect 25596 9716 25648 9722
rect 25596 9658 25648 9664
rect 25320 9580 25372 9586
rect 25320 9522 25372 9528
rect 25412 9376 25464 9382
rect 25412 9318 25464 9324
rect 25424 9042 25452 9318
rect 25412 9036 25464 9042
rect 25412 8978 25464 8984
rect 25136 8900 25188 8906
rect 25136 8842 25188 8848
rect 25044 8492 25096 8498
rect 25044 8434 25096 8440
rect 24952 7472 25004 7478
rect 24952 7414 25004 7420
rect 24964 6186 24992 7414
rect 24952 6180 25004 6186
rect 24952 6122 25004 6128
rect 24676 4752 24728 4758
rect 24676 4694 24728 4700
rect 25596 4684 25648 4690
rect 25596 4626 25648 4632
rect 25608 4282 25636 4626
rect 25596 4276 25648 4282
rect 25596 4218 25648 4224
rect 24124 4072 24176 4078
rect 24124 4014 24176 4020
rect 24308 4072 24360 4078
rect 24308 4014 24360 4020
rect 24400 4072 24452 4078
rect 24400 4014 24452 4020
rect 24032 3596 24084 3602
rect 24032 3538 24084 3544
rect 23296 2848 23348 2854
rect 23296 2790 23348 2796
rect 23664 2848 23716 2854
rect 23664 2790 23716 2796
rect 22480 2746 22784 2774
rect 22950 2748 23258 2757
rect 22950 2746 22956 2748
rect 23012 2746 23036 2748
rect 23092 2746 23116 2748
rect 23172 2746 23196 2748
rect 23252 2746 23258 2748
rect 22480 2650 22508 2746
rect 23012 2694 23014 2746
rect 23194 2694 23196 2746
rect 22950 2692 22956 2694
rect 23012 2692 23036 2694
rect 23092 2692 23116 2694
rect 23172 2692 23196 2694
rect 23252 2692 23258 2694
rect 22950 2683 23258 2692
rect 22468 2644 22520 2650
rect 22468 2586 22520 2592
rect 24136 2582 24164 4014
rect 24308 3664 24360 3670
rect 24412 3641 24440 4014
rect 24768 3936 24820 3942
rect 24768 3878 24820 3884
rect 24308 3606 24360 3612
rect 24398 3632 24454 3641
rect 24320 3210 24348 3606
rect 24780 3602 24808 3878
rect 25700 3602 25728 12396
rect 25872 12378 25924 12384
rect 26252 12170 26280 12815
rect 26344 12646 26372 14758
rect 26436 14074 26464 15506
rect 26424 14068 26476 14074
rect 26424 14010 26476 14016
rect 26436 12782 26464 14010
rect 26424 12776 26476 12782
rect 26424 12718 26476 12724
rect 26332 12640 26384 12646
rect 26332 12582 26384 12588
rect 26332 12436 26384 12442
rect 26332 12378 26384 12384
rect 26240 12164 26292 12170
rect 26240 12106 26292 12112
rect 26344 11898 26372 12378
rect 26332 11892 26384 11898
rect 26332 11834 26384 11840
rect 26528 11354 26556 15506
rect 26608 15360 26660 15366
rect 26608 15302 26660 15308
rect 26620 13462 26648 15302
rect 26712 15162 26740 23015
rect 26988 22506 27016 23122
rect 27172 22506 27200 23666
rect 26976 22500 27028 22506
rect 26976 22442 27028 22448
rect 27160 22500 27212 22506
rect 27160 22442 27212 22448
rect 27068 22092 27120 22098
rect 27068 22034 27120 22040
rect 26884 20800 26936 20806
rect 26884 20742 26936 20748
rect 26790 19816 26846 19825
rect 26790 19751 26792 19760
rect 26844 19751 26846 19760
rect 26792 19722 26844 19728
rect 26896 19242 26924 20742
rect 26976 20392 27028 20398
rect 26976 20334 27028 20340
rect 26988 19718 27016 20334
rect 26976 19712 27028 19718
rect 26976 19654 27028 19660
rect 26884 19236 26936 19242
rect 26884 19178 26936 19184
rect 26792 18284 26844 18290
rect 26792 18226 26844 18232
rect 26804 17610 26832 18226
rect 26792 17604 26844 17610
rect 26792 17546 26844 17552
rect 26792 15972 26844 15978
rect 26792 15914 26844 15920
rect 26700 15156 26752 15162
rect 26700 15098 26752 15104
rect 26700 14272 26752 14278
rect 26700 14214 26752 14220
rect 26712 14006 26740 14214
rect 26700 14000 26752 14006
rect 26700 13942 26752 13948
rect 26608 13456 26660 13462
rect 26608 13398 26660 13404
rect 26712 13394 26740 13942
rect 26700 13388 26752 13394
rect 26700 13330 26752 13336
rect 26712 12850 26740 13330
rect 26700 12844 26752 12850
rect 26700 12786 26752 12792
rect 26804 12442 26832 15914
rect 26896 14550 26924 19178
rect 26988 17202 27016 19654
rect 27080 18834 27108 22034
rect 27160 21888 27212 21894
rect 27160 21830 27212 21836
rect 27172 20602 27200 21830
rect 27264 21690 27292 24074
rect 27356 23798 27384 26200
rect 27804 24812 27856 24818
rect 27804 24754 27856 24760
rect 27436 24744 27488 24750
rect 27436 24686 27488 24692
rect 27344 23792 27396 23798
rect 27344 23734 27396 23740
rect 27448 23730 27476 24686
rect 27712 24064 27764 24070
rect 27712 24006 27764 24012
rect 27436 23724 27488 23730
rect 27436 23666 27488 23672
rect 27620 23656 27672 23662
rect 27620 23598 27672 23604
rect 27632 22710 27660 23598
rect 27436 22704 27488 22710
rect 27436 22646 27488 22652
rect 27620 22704 27672 22710
rect 27620 22646 27672 22652
rect 27344 22636 27396 22642
rect 27344 22578 27396 22584
rect 27252 21684 27304 21690
rect 27252 21626 27304 21632
rect 27356 21185 27384 22578
rect 27448 21894 27476 22646
rect 27620 22568 27672 22574
rect 27620 22510 27672 22516
rect 27632 22137 27660 22510
rect 27618 22128 27674 22137
rect 27618 22063 27674 22072
rect 27724 22030 27752 24006
rect 27816 23866 27844 24754
rect 28000 24274 28028 26200
rect 28816 24880 28868 24886
rect 28816 24822 28868 24828
rect 28724 24336 28776 24342
rect 28724 24278 28776 24284
rect 27988 24268 28040 24274
rect 27988 24210 28040 24216
rect 28736 24206 28764 24278
rect 28724 24200 28776 24206
rect 28724 24142 28776 24148
rect 28448 24064 28500 24070
rect 28448 24006 28500 24012
rect 27950 23964 28258 23973
rect 27950 23962 27956 23964
rect 28012 23962 28036 23964
rect 28092 23962 28116 23964
rect 28172 23962 28196 23964
rect 28252 23962 28258 23964
rect 28012 23910 28014 23962
rect 28194 23910 28196 23962
rect 27950 23908 27956 23910
rect 28012 23908 28036 23910
rect 28092 23908 28116 23910
rect 28172 23908 28196 23910
rect 28252 23908 28258 23910
rect 27950 23899 28258 23908
rect 27804 23860 27856 23866
rect 27804 23802 27856 23808
rect 27894 23352 27950 23361
rect 27804 23316 27856 23322
rect 27894 23287 27896 23296
rect 27804 23258 27856 23264
rect 27948 23287 27950 23296
rect 27896 23258 27948 23264
rect 27816 22234 27844 23258
rect 28356 22976 28408 22982
rect 28356 22918 28408 22924
rect 27950 22876 28258 22885
rect 27950 22874 27956 22876
rect 28012 22874 28036 22876
rect 28092 22874 28116 22876
rect 28172 22874 28196 22876
rect 28252 22874 28258 22876
rect 28012 22822 28014 22874
rect 28194 22822 28196 22874
rect 27950 22820 27956 22822
rect 28012 22820 28036 22822
rect 28092 22820 28116 22822
rect 28172 22820 28196 22822
rect 28252 22820 28258 22822
rect 27950 22811 28258 22820
rect 27896 22704 27948 22710
rect 27896 22646 27948 22652
rect 27804 22228 27856 22234
rect 27804 22170 27856 22176
rect 27802 22128 27858 22137
rect 27908 22098 27936 22646
rect 27802 22063 27858 22072
rect 27896 22092 27948 22098
rect 27712 22024 27764 22030
rect 27712 21966 27764 21972
rect 27436 21888 27488 21894
rect 27436 21830 27488 21836
rect 27816 21690 27844 22063
rect 27896 22034 27948 22040
rect 27950 21788 28258 21797
rect 27950 21786 27956 21788
rect 28012 21786 28036 21788
rect 28092 21786 28116 21788
rect 28172 21786 28196 21788
rect 28252 21786 28258 21788
rect 28012 21734 28014 21786
rect 28194 21734 28196 21786
rect 27950 21732 27956 21734
rect 28012 21732 28036 21734
rect 28092 21732 28116 21734
rect 28172 21732 28196 21734
rect 28252 21732 28258 21734
rect 27950 21723 28258 21732
rect 27712 21684 27764 21690
rect 27712 21626 27764 21632
rect 27804 21684 27856 21690
rect 27804 21626 27856 21632
rect 27436 21616 27488 21622
rect 27724 21593 27752 21626
rect 27710 21584 27766 21593
rect 27488 21564 27568 21570
rect 27436 21558 27568 21564
rect 27448 21542 27568 21558
rect 27342 21176 27398 21185
rect 27342 21111 27398 21120
rect 27160 20596 27212 20602
rect 27160 20538 27212 20544
rect 27436 20528 27488 20534
rect 27356 20488 27436 20516
rect 27160 19984 27212 19990
rect 27160 19926 27212 19932
rect 27172 19446 27200 19926
rect 27252 19712 27304 19718
rect 27252 19654 27304 19660
rect 27160 19440 27212 19446
rect 27160 19382 27212 19388
rect 27160 18896 27212 18902
rect 27160 18838 27212 18844
rect 27068 18828 27120 18834
rect 27068 18770 27120 18776
rect 26976 17196 27028 17202
rect 26976 17138 27028 17144
rect 27172 16250 27200 18838
rect 27264 18426 27292 19654
rect 27252 18420 27304 18426
rect 27252 18362 27304 18368
rect 27356 16794 27384 20488
rect 27436 20470 27488 20476
rect 27540 20346 27568 21542
rect 27710 21519 27766 21528
rect 27896 21548 27948 21554
rect 27896 21490 27948 21496
rect 27908 21146 27936 21490
rect 28264 21480 28316 21486
rect 28264 21422 28316 21428
rect 27804 21140 27856 21146
rect 27804 21082 27856 21088
rect 27896 21140 27948 21146
rect 27896 21082 27948 21088
rect 27816 21010 27844 21082
rect 27804 21004 27856 21010
rect 27804 20946 27856 20952
rect 27618 20904 27674 20913
rect 27618 20839 27674 20848
rect 27632 20806 27660 20839
rect 27620 20800 27672 20806
rect 27620 20742 27672 20748
rect 27710 20768 27766 20777
rect 27448 20318 27568 20346
rect 27448 18170 27476 20318
rect 27528 19916 27580 19922
rect 27528 19858 27580 19864
rect 27540 19514 27568 19858
rect 27632 19786 27660 20742
rect 27710 20703 27766 20712
rect 27724 20602 27752 20703
rect 27712 20596 27764 20602
rect 27712 20538 27764 20544
rect 27620 19780 27672 19786
rect 27620 19722 27672 19728
rect 27528 19508 27580 19514
rect 27528 19450 27580 19456
rect 27712 19440 27764 19446
rect 27712 19382 27764 19388
rect 27528 19236 27580 19242
rect 27528 19178 27580 19184
rect 27540 18902 27568 19178
rect 27528 18896 27580 18902
rect 27528 18838 27580 18844
rect 27540 18290 27568 18838
rect 27620 18624 27672 18630
rect 27620 18566 27672 18572
rect 27632 18426 27660 18566
rect 27620 18420 27672 18426
rect 27620 18362 27672 18368
rect 27528 18284 27580 18290
rect 27528 18226 27580 18232
rect 27448 18142 27568 18170
rect 27436 17332 27488 17338
rect 27436 17274 27488 17280
rect 27448 17202 27476 17274
rect 27436 17196 27488 17202
rect 27436 17138 27488 17144
rect 27540 17082 27568 18142
rect 27620 18080 27672 18086
rect 27620 18022 27672 18028
rect 27448 17054 27568 17082
rect 27344 16788 27396 16794
rect 27344 16730 27396 16736
rect 27160 16244 27212 16250
rect 27160 16186 27212 16192
rect 27448 14822 27476 17054
rect 27632 16946 27660 18022
rect 27724 17320 27752 19382
rect 27816 19310 27844 20946
rect 28276 20788 28304 21422
rect 28368 20913 28396 22918
rect 28460 21865 28488 24006
rect 28632 23520 28684 23526
rect 28632 23462 28684 23468
rect 28540 21888 28592 21894
rect 28446 21856 28502 21865
rect 28540 21830 28592 21836
rect 28446 21791 28502 21800
rect 28448 21684 28500 21690
rect 28448 21626 28500 21632
rect 28460 21010 28488 21626
rect 28552 21321 28580 21830
rect 28644 21350 28672 23462
rect 28828 22094 28856 24822
rect 28920 24342 28948 26302
rect 29274 26200 29330 27000
rect 29918 26200 29974 27000
rect 30562 26200 30618 27000
rect 31206 26200 31262 27000
rect 31850 26330 31906 27000
rect 31850 26302 32168 26330
rect 31850 26200 31906 26302
rect 29288 24682 29316 26200
rect 29092 24676 29144 24682
rect 29092 24618 29144 24624
rect 29276 24676 29328 24682
rect 29276 24618 29328 24624
rect 28908 24336 28960 24342
rect 28908 24278 28960 24284
rect 29104 24138 29132 24618
rect 29092 24132 29144 24138
rect 29092 24074 29144 24080
rect 29184 24064 29236 24070
rect 29184 24006 29236 24012
rect 29000 23520 29052 23526
rect 29000 23462 29052 23468
rect 29012 23225 29040 23462
rect 28998 23216 29054 23225
rect 28998 23151 29054 23160
rect 29000 22568 29052 22574
rect 29000 22510 29052 22516
rect 29090 22536 29146 22545
rect 28908 22432 28960 22438
rect 28908 22374 28960 22380
rect 28920 22098 28948 22374
rect 28736 22066 28856 22094
rect 28908 22092 28960 22098
rect 28632 21344 28684 21350
rect 28538 21312 28594 21321
rect 28632 21286 28684 21292
rect 28538 21247 28594 21256
rect 28448 21004 28500 21010
rect 28448 20946 28500 20952
rect 28354 20904 28410 20913
rect 28736 20890 28764 22066
rect 28908 22034 28960 22040
rect 28814 21856 28870 21865
rect 28814 21791 28870 21800
rect 28354 20839 28410 20848
rect 28644 20862 28764 20890
rect 28644 20806 28672 20862
rect 28632 20800 28684 20806
rect 28276 20760 28396 20788
rect 27950 20700 28258 20709
rect 27950 20698 27956 20700
rect 28012 20698 28036 20700
rect 28092 20698 28116 20700
rect 28172 20698 28196 20700
rect 28252 20698 28258 20700
rect 28012 20646 28014 20698
rect 28194 20646 28196 20698
rect 27950 20644 27956 20646
rect 28012 20644 28036 20646
rect 28092 20644 28116 20646
rect 28172 20644 28196 20646
rect 28252 20644 28258 20646
rect 27950 20635 28258 20644
rect 27896 20392 27948 20398
rect 27896 20334 27948 20340
rect 27908 19922 27936 20334
rect 28262 19952 28318 19961
rect 27896 19916 27948 19922
rect 28368 19938 28396 20760
rect 28632 20742 28684 20748
rect 28724 20800 28776 20806
rect 28724 20742 28776 20748
rect 28540 20596 28592 20602
rect 28540 20538 28592 20544
rect 28552 20369 28580 20538
rect 28538 20360 28594 20369
rect 28538 20295 28594 20304
rect 28446 20224 28502 20233
rect 28446 20159 28502 20168
rect 28318 19910 28396 19938
rect 28262 19887 28318 19896
rect 27896 19858 27948 19864
rect 28276 19700 28304 19887
rect 28276 19672 28396 19700
rect 27950 19612 28258 19621
rect 27950 19610 27956 19612
rect 28012 19610 28036 19612
rect 28092 19610 28116 19612
rect 28172 19610 28196 19612
rect 28252 19610 28258 19612
rect 28012 19558 28014 19610
rect 28194 19558 28196 19610
rect 27950 19556 27956 19558
rect 28012 19556 28036 19558
rect 28092 19556 28116 19558
rect 28172 19556 28196 19558
rect 28252 19556 28258 19558
rect 27950 19547 28258 19556
rect 27988 19508 28040 19514
rect 27988 19450 28040 19456
rect 28000 19334 28028 19450
rect 27804 19304 27856 19310
rect 27804 19246 27856 19252
rect 27908 19306 28028 19334
rect 27908 18612 27936 19306
rect 28368 19009 28396 19672
rect 28354 19000 28410 19009
rect 28354 18935 28410 18944
rect 27816 18584 27936 18612
rect 27816 18086 27844 18584
rect 27950 18524 28258 18533
rect 27950 18522 27956 18524
rect 28012 18522 28036 18524
rect 28092 18522 28116 18524
rect 28172 18522 28196 18524
rect 28252 18522 28258 18524
rect 28012 18470 28014 18522
rect 28194 18470 28196 18522
rect 27950 18468 27956 18470
rect 28012 18468 28036 18470
rect 28092 18468 28116 18470
rect 28172 18468 28196 18470
rect 28252 18468 28258 18470
rect 27950 18459 28258 18468
rect 27804 18080 27856 18086
rect 27804 18022 27856 18028
rect 28356 17808 28408 17814
rect 28356 17750 28408 17756
rect 27804 17604 27856 17610
rect 27804 17546 27856 17552
rect 27816 17513 27844 17546
rect 27802 17504 27858 17513
rect 27802 17439 27858 17448
rect 27950 17436 28258 17445
rect 27950 17434 27956 17436
rect 28012 17434 28036 17436
rect 28092 17434 28116 17436
rect 28172 17434 28196 17436
rect 28252 17434 28258 17436
rect 28012 17382 28014 17434
rect 28194 17382 28196 17434
rect 27950 17380 27956 17382
rect 28012 17380 28036 17382
rect 28092 17380 28116 17382
rect 28172 17380 28196 17382
rect 28252 17380 28258 17382
rect 27950 17371 28258 17380
rect 27724 17292 27936 17320
rect 27710 17232 27766 17241
rect 27710 17167 27712 17176
rect 27764 17167 27766 17176
rect 27712 17138 27764 17144
rect 27804 17128 27856 17134
rect 27802 17096 27804 17105
rect 27856 17096 27858 17105
rect 27802 17031 27858 17040
rect 27632 16918 27752 16946
rect 27620 16788 27672 16794
rect 27620 16730 27672 16736
rect 27526 15056 27582 15065
rect 27526 14991 27528 15000
rect 27580 14991 27582 15000
rect 27528 14962 27580 14968
rect 27436 14816 27488 14822
rect 27436 14758 27488 14764
rect 26884 14544 26936 14550
rect 26884 14486 26936 14492
rect 27632 14074 27660 16730
rect 27724 16153 27752 16918
rect 27908 16504 27936 17292
rect 27988 17128 28040 17134
rect 27988 17070 28040 17076
rect 28000 16794 28028 17070
rect 28368 16998 28396 17750
rect 28356 16992 28408 16998
rect 28356 16934 28408 16940
rect 27988 16788 28040 16794
rect 27988 16730 28040 16736
rect 27816 16476 27936 16504
rect 27710 16144 27766 16153
rect 27710 16079 27766 16088
rect 27724 14498 27752 16079
rect 27816 14618 27844 16476
rect 27950 16348 28258 16357
rect 27950 16346 27956 16348
rect 28012 16346 28036 16348
rect 28092 16346 28116 16348
rect 28172 16346 28196 16348
rect 28252 16346 28258 16348
rect 28012 16294 28014 16346
rect 28194 16294 28196 16346
rect 27950 16292 27956 16294
rect 28012 16292 28036 16294
rect 28092 16292 28116 16294
rect 28172 16292 28196 16294
rect 28252 16292 28258 16294
rect 27950 16283 28258 16292
rect 28368 15502 28396 16934
rect 28356 15496 28408 15502
rect 28356 15438 28408 15444
rect 28460 15434 28488 20159
rect 28538 20088 28594 20097
rect 28538 20023 28594 20032
rect 28552 19922 28580 20023
rect 28540 19916 28592 19922
rect 28540 19858 28592 19864
rect 28632 19916 28684 19922
rect 28632 19858 28684 19864
rect 28538 19680 28594 19689
rect 28538 19615 28594 19624
rect 28552 17864 28580 19615
rect 28644 19378 28672 19858
rect 28736 19514 28764 20742
rect 28828 20346 28856 21791
rect 28920 21486 28948 22034
rect 28908 21480 28960 21486
rect 28908 21422 28960 21428
rect 28908 21344 28960 21350
rect 28908 21286 28960 21292
rect 28920 20482 28948 21286
rect 29012 20602 29040 22510
rect 29090 22471 29146 22480
rect 29104 21622 29132 22471
rect 29092 21616 29144 21622
rect 29092 21558 29144 21564
rect 29104 21350 29132 21558
rect 29092 21344 29144 21350
rect 29092 21286 29144 21292
rect 29000 20596 29052 20602
rect 29000 20538 29052 20544
rect 28920 20454 29040 20482
rect 29012 20346 29040 20454
rect 28828 20318 28948 20346
rect 29012 20318 29132 20346
rect 28816 19848 28868 19854
rect 28816 19790 28868 19796
rect 28828 19514 28856 19790
rect 28920 19718 28948 20318
rect 29000 19984 29052 19990
rect 29000 19926 29052 19932
rect 28908 19712 28960 19718
rect 28908 19654 28960 19660
rect 28724 19508 28776 19514
rect 28724 19450 28776 19456
rect 28816 19508 28868 19514
rect 28816 19450 28868 19456
rect 28632 19372 28684 19378
rect 28632 19314 28684 19320
rect 28816 18216 28868 18222
rect 28816 18158 28868 18164
rect 28552 17836 28764 17864
rect 28540 17740 28592 17746
rect 28540 17682 28592 17688
rect 28552 16114 28580 17682
rect 28632 17604 28684 17610
rect 28632 17546 28684 17552
rect 28644 17202 28672 17546
rect 28632 17196 28684 17202
rect 28632 17138 28684 17144
rect 28736 17116 28764 17836
rect 28828 17542 28856 18158
rect 28920 18154 28948 19654
rect 29012 18358 29040 19926
rect 29000 18352 29052 18358
rect 29000 18294 29052 18300
rect 28908 18148 28960 18154
rect 28908 18090 28960 18096
rect 28816 17536 28868 17542
rect 28816 17478 28868 17484
rect 28908 17536 28960 17542
rect 28908 17478 28960 17484
rect 28920 17338 28948 17478
rect 29104 17338 29132 20318
rect 29196 18630 29224 24006
rect 29736 23656 29788 23662
rect 29736 23598 29788 23604
rect 29276 23588 29328 23594
rect 29276 23530 29328 23536
rect 29368 23588 29420 23594
rect 29368 23530 29420 23536
rect 29288 22234 29316 23530
rect 29276 22228 29328 22234
rect 29276 22170 29328 22176
rect 29276 21344 29328 21350
rect 29276 21286 29328 21292
rect 29288 18698 29316 21286
rect 29380 21010 29408 23530
rect 29748 23322 29776 23598
rect 29736 23316 29788 23322
rect 29736 23258 29788 23264
rect 29552 22092 29604 22098
rect 29552 22034 29604 22040
rect 29564 21894 29592 22034
rect 29828 22024 29880 22030
rect 29932 22001 29960 26200
rect 30472 24064 30524 24070
rect 30472 24006 30524 24012
rect 30012 23656 30064 23662
rect 30012 23598 30064 23604
rect 30024 23118 30052 23598
rect 30288 23520 30340 23526
rect 30288 23462 30340 23468
rect 30300 23186 30328 23462
rect 30288 23180 30340 23186
rect 30288 23122 30340 23128
rect 30012 23112 30064 23118
rect 30012 23054 30064 23060
rect 30024 22778 30052 23054
rect 30104 22976 30156 22982
rect 30104 22918 30156 22924
rect 30012 22772 30064 22778
rect 30012 22714 30064 22720
rect 29828 21966 29880 21972
rect 29918 21992 29974 22001
rect 29552 21888 29604 21894
rect 29552 21830 29604 21836
rect 29736 21412 29788 21418
rect 29736 21354 29788 21360
rect 29552 21344 29604 21350
rect 29552 21286 29604 21292
rect 29458 21040 29514 21049
rect 29368 21004 29420 21010
rect 29458 20975 29514 20984
rect 29368 20946 29420 20952
rect 29368 20868 29420 20874
rect 29368 20810 29420 20816
rect 29380 20398 29408 20810
rect 29472 20777 29500 20975
rect 29458 20768 29514 20777
rect 29458 20703 29514 20712
rect 29368 20392 29420 20398
rect 29368 20334 29420 20340
rect 29276 18692 29328 18698
rect 29276 18634 29328 18640
rect 29184 18624 29236 18630
rect 29184 18566 29236 18572
rect 28908 17332 28960 17338
rect 28908 17274 28960 17280
rect 29092 17332 29144 17338
rect 29092 17274 29144 17280
rect 28736 17088 28856 17116
rect 28724 16992 28776 16998
rect 28724 16934 28776 16940
rect 28540 16108 28592 16114
rect 28540 16050 28592 16056
rect 28552 15570 28580 16050
rect 28540 15564 28592 15570
rect 28540 15506 28592 15512
rect 28448 15428 28500 15434
rect 28448 15370 28500 15376
rect 27950 15260 28258 15269
rect 27950 15258 27956 15260
rect 28012 15258 28036 15260
rect 28092 15258 28116 15260
rect 28172 15258 28196 15260
rect 28252 15258 28258 15260
rect 28012 15206 28014 15258
rect 28194 15206 28196 15258
rect 27950 15204 27956 15206
rect 28012 15204 28036 15206
rect 28092 15204 28116 15206
rect 28172 15204 28196 15206
rect 28252 15204 28258 15206
rect 27950 15195 28258 15204
rect 28356 15020 28408 15026
rect 28356 14962 28408 14968
rect 27804 14612 27856 14618
rect 27804 14554 27856 14560
rect 28264 14612 28316 14618
rect 28264 14554 28316 14560
rect 27724 14470 27844 14498
rect 28276 14482 28304 14554
rect 27712 14408 27764 14414
rect 27712 14350 27764 14356
rect 27620 14068 27672 14074
rect 27620 14010 27672 14016
rect 27160 13932 27212 13938
rect 27160 13874 27212 13880
rect 26792 12436 26844 12442
rect 26792 12378 26844 12384
rect 27068 12164 27120 12170
rect 27068 12106 27120 12112
rect 26792 11824 26844 11830
rect 26792 11766 26844 11772
rect 26516 11348 26568 11354
rect 26516 11290 26568 11296
rect 26528 10606 26556 11290
rect 26516 10600 26568 10606
rect 26516 10542 26568 10548
rect 26146 9616 26202 9625
rect 26056 9580 26108 9586
rect 26146 9551 26148 9560
rect 26056 9522 26108 9528
rect 26200 9551 26202 9560
rect 26148 9522 26200 9528
rect 26068 7750 26096 9522
rect 26160 9110 26188 9522
rect 26804 9450 26832 11766
rect 26884 11144 26936 11150
rect 26936 11104 27016 11132
rect 26884 11086 26936 11092
rect 26988 10062 27016 11104
rect 26976 10056 27028 10062
rect 26976 9998 27028 10004
rect 26884 9988 26936 9994
rect 26884 9930 26936 9936
rect 26896 9518 26924 9930
rect 26988 9518 27016 9998
rect 26884 9512 26936 9518
rect 26884 9454 26936 9460
rect 26976 9512 27028 9518
rect 26976 9454 27028 9460
rect 26792 9444 26844 9450
rect 26792 9386 26844 9392
rect 26148 9104 26200 9110
rect 26148 9046 26200 9052
rect 26056 7744 26108 7750
rect 26056 7686 26108 7692
rect 26804 5030 26832 9386
rect 27080 9178 27108 12106
rect 27068 9172 27120 9178
rect 27068 9114 27120 9120
rect 26792 5024 26844 5030
rect 26792 4966 26844 4972
rect 26148 4480 26200 4486
rect 26148 4422 26200 4428
rect 25872 3732 25924 3738
rect 25872 3674 25924 3680
rect 24398 3567 24454 3576
rect 24768 3596 24820 3602
rect 24768 3538 24820 3544
rect 24860 3596 24912 3602
rect 24860 3538 24912 3544
rect 25688 3596 25740 3602
rect 25688 3538 25740 3544
rect 24492 3528 24544 3534
rect 24872 3482 24900 3538
rect 24544 3476 24900 3482
rect 24492 3470 24900 3476
rect 24504 3454 24900 3470
rect 24320 3182 24532 3210
rect 24504 3126 24532 3182
rect 24492 3120 24544 3126
rect 24492 3062 24544 3068
rect 24504 2990 24532 3062
rect 25884 2990 25912 3674
rect 26160 3058 26188 4422
rect 27172 3398 27200 13874
rect 27632 13870 27660 14010
rect 27620 13864 27672 13870
rect 27620 13806 27672 13812
rect 27620 12980 27672 12986
rect 27620 12922 27672 12928
rect 27528 12300 27580 12306
rect 27528 12242 27580 12248
rect 27252 12096 27304 12102
rect 27252 12038 27304 12044
rect 27344 12096 27396 12102
rect 27344 12038 27396 12044
rect 27264 11218 27292 12038
rect 27356 11762 27384 12038
rect 27434 11792 27490 11801
rect 27344 11756 27396 11762
rect 27434 11727 27490 11736
rect 27344 11698 27396 11704
rect 27448 11694 27476 11727
rect 27436 11688 27488 11694
rect 27436 11630 27488 11636
rect 27344 11552 27396 11558
rect 27344 11494 27396 11500
rect 27252 11212 27304 11218
rect 27252 11154 27304 11160
rect 27356 9994 27384 11494
rect 27540 11354 27568 12242
rect 27632 11898 27660 12922
rect 27724 12073 27752 14350
rect 27816 13530 27844 14470
rect 28264 14476 28316 14482
rect 28264 14418 28316 14424
rect 27950 14172 28258 14181
rect 27950 14170 27956 14172
rect 28012 14170 28036 14172
rect 28092 14170 28116 14172
rect 28172 14170 28196 14172
rect 28252 14170 28258 14172
rect 28012 14118 28014 14170
rect 28194 14118 28196 14170
rect 27950 14116 27956 14118
rect 28012 14116 28036 14118
rect 28092 14116 28116 14118
rect 28172 14116 28196 14118
rect 28252 14116 28258 14118
rect 27950 14107 28258 14116
rect 27804 13524 27856 13530
rect 27804 13466 27856 13472
rect 27816 13190 27844 13466
rect 27804 13184 27856 13190
rect 27804 13126 27856 13132
rect 27950 13084 28258 13093
rect 27950 13082 27956 13084
rect 28012 13082 28036 13084
rect 28092 13082 28116 13084
rect 28172 13082 28196 13084
rect 28252 13082 28258 13084
rect 28012 13030 28014 13082
rect 28194 13030 28196 13082
rect 27950 13028 27956 13030
rect 28012 13028 28036 13030
rect 28092 13028 28116 13030
rect 28172 13028 28196 13030
rect 28252 13028 28258 13030
rect 27950 13019 28258 13028
rect 27988 12844 28040 12850
rect 27988 12786 28040 12792
rect 27804 12776 27856 12782
rect 27804 12718 27856 12724
rect 27710 12064 27766 12073
rect 27710 11999 27766 12008
rect 27620 11892 27672 11898
rect 27620 11834 27672 11840
rect 27528 11348 27580 11354
rect 27528 11290 27580 11296
rect 27724 11098 27752 11999
rect 27816 11694 27844 12718
rect 28000 12102 28028 12786
rect 27988 12096 28040 12102
rect 27988 12038 28040 12044
rect 27950 11996 28258 12005
rect 27950 11994 27956 11996
rect 28012 11994 28036 11996
rect 28092 11994 28116 11996
rect 28172 11994 28196 11996
rect 28252 11994 28258 11996
rect 28012 11942 28014 11994
rect 28194 11942 28196 11994
rect 27950 11940 27956 11942
rect 28012 11940 28036 11942
rect 28092 11940 28116 11942
rect 28172 11940 28196 11942
rect 28252 11940 28258 11942
rect 27950 11931 28258 11940
rect 27804 11688 27856 11694
rect 27804 11630 27856 11636
rect 28368 11626 28396 14962
rect 28448 14612 28500 14618
rect 28448 14554 28500 14560
rect 28460 13326 28488 14554
rect 28632 13388 28684 13394
rect 28632 13330 28684 13336
rect 28448 13320 28500 13326
rect 28448 13262 28500 13268
rect 28448 12096 28500 12102
rect 28448 12038 28500 12044
rect 28460 11762 28488 12038
rect 28448 11756 28500 11762
rect 28448 11698 28500 11704
rect 28356 11620 28408 11626
rect 28356 11562 28408 11568
rect 27724 11070 27844 11098
rect 27528 10668 27580 10674
rect 27528 10610 27580 10616
rect 27344 9988 27396 9994
rect 27344 9930 27396 9936
rect 27540 4622 27568 10610
rect 27712 9172 27764 9178
rect 27712 9114 27764 9120
rect 27620 8832 27672 8838
rect 27620 8774 27672 8780
rect 27632 6730 27660 8774
rect 27724 7818 27752 9114
rect 27712 7812 27764 7818
rect 27712 7754 27764 7760
rect 27816 7342 27844 11070
rect 27950 10908 28258 10917
rect 27950 10906 27956 10908
rect 28012 10906 28036 10908
rect 28092 10906 28116 10908
rect 28172 10906 28196 10908
rect 28252 10906 28258 10908
rect 28012 10854 28014 10906
rect 28194 10854 28196 10906
rect 27950 10852 27956 10854
rect 28012 10852 28036 10854
rect 28092 10852 28116 10854
rect 28172 10852 28196 10854
rect 28252 10852 28258 10854
rect 27950 10843 28258 10852
rect 28368 10452 28396 11562
rect 28644 11218 28672 13330
rect 28736 11218 28764 16934
rect 28828 16182 28856 17088
rect 29092 17060 29144 17066
rect 29092 17002 29144 17008
rect 28816 16176 28868 16182
rect 28816 16118 28868 16124
rect 28828 14482 28856 16118
rect 28816 14476 28868 14482
rect 28816 14418 28868 14424
rect 28828 13433 28856 14418
rect 28908 13864 28960 13870
rect 28908 13806 28960 13812
rect 28814 13424 28870 13433
rect 28814 13359 28870 13368
rect 28816 12436 28868 12442
rect 28816 12378 28868 12384
rect 28828 11830 28856 12378
rect 28920 12170 28948 13806
rect 29000 13456 29052 13462
rect 29000 13398 29052 13404
rect 29012 12782 29040 13398
rect 29000 12776 29052 12782
rect 29000 12718 29052 12724
rect 28908 12164 28960 12170
rect 28908 12106 28960 12112
rect 28920 11898 28948 12106
rect 28908 11892 28960 11898
rect 28908 11834 28960 11840
rect 28816 11824 28868 11830
rect 28816 11766 28868 11772
rect 28632 11212 28684 11218
rect 28632 11154 28684 11160
rect 28724 11212 28776 11218
rect 28724 11154 28776 11160
rect 28632 11008 28684 11014
rect 28828 10996 28856 11766
rect 28684 10968 28856 10996
rect 28632 10950 28684 10956
rect 28540 10532 28592 10538
rect 28540 10474 28592 10480
rect 28448 10464 28500 10470
rect 28368 10424 28448 10452
rect 28448 10406 28500 10412
rect 28552 9926 28580 10474
rect 28644 9994 28672 10950
rect 28920 10742 28948 11834
rect 29104 11354 29132 17002
rect 29196 16522 29224 18566
rect 29472 17338 29500 20703
rect 29564 19922 29592 21286
rect 29644 20460 29696 20466
rect 29644 20402 29696 20408
rect 29656 20369 29684 20402
rect 29642 20360 29698 20369
rect 29642 20295 29698 20304
rect 29552 19916 29604 19922
rect 29552 19858 29604 19864
rect 29644 19508 29696 19514
rect 29644 19450 29696 19456
rect 29656 18426 29684 19450
rect 29748 18970 29776 21354
rect 29840 20466 29868 21966
rect 29918 21927 29974 21936
rect 30012 21480 30064 21486
rect 30012 21422 30064 21428
rect 29918 21312 29974 21321
rect 29918 21247 29974 21256
rect 29932 21049 29960 21247
rect 29918 21040 29974 21049
rect 29918 20975 29974 20984
rect 29828 20460 29880 20466
rect 29828 20402 29880 20408
rect 29932 20398 29960 20975
rect 29920 20392 29972 20398
rect 29920 20334 29972 20340
rect 30024 20058 30052 21422
rect 30116 21146 30144 22918
rect 30380 22500 30432 22506
rect 30380 22442 30432 22448
rect 30288 22432 30340 22438
rect 30288 22374 30340 22380
rect 30300 22273 30328 22374
rect 30286 22264 30342 22273
rect 30286 22199 30342 22208
rect 30392 21962 30420 22442
rect 30484 22098 30512 24006
rect 30576 23322 30604 26200
rect 31220 24698 31248 26200
rect 32140 24954 32168 26302
rect 32494 26200 32550 27000
rect 33138 26200 33194 27000
rect 33782 26200 33838 27000
rect 34426 26330 34482 27000
rect 34518 26344 34574 26353
rect 34426 26302 34518 26330
rect 34426 26200 34482 26302
rect 34518 26279 34574 26288
rect 35070 26200 35126 27000
rect 35714 26200 35770 27000
rect 36358 26330 36414 27000
rect 36358 26302 36676 26330
rect 36358 26200 36414 26302
rect 32128 24948 32180 24954
rect 32128 24890 32180 24896
rect 31220 24670 31340 24698
rect 31208 24608 31260 24614
rect 31208 24550 31260 24556
rect 31220 24206 31248 24550
rect 31208 24200 31260 24206
rect 31208 24142 31260 24148
rect 30748 23792 30800 23798
rect 30748 23734 30800 23740
rect 30564 23316 30616 23322
rect 30564 23258 30616 23264
rect 30656 23248 30708 23254
rect 30656 23190 30708 23196
rect 30472 22092 30524 22098
rect 30472 22034 30524 22040
rect 30380 21956 30432 21962
rect 30380 21898 30432 21904
rect 30484 21554 30512 22034
rect 30472 21548 30524 21554
rect 30472 21490 30524 21496
rect 30380 21344 30432 21350
rect 30668 21332 30696 23190
rect 30760 22982 30788 23734
rect 30840 23044 30892 23050
rect 30840 22986 30892 22992
rect 30748 22976 30800 22982
rect 30748 22918 30800 22924
rect 30760 22710 30788 22918
rect 30748 22704 30800 22710
rect 30748 22646 30800 22652
rect 30852 22574 30880 22986
rect 31208 22976 31260 22982
rect 31208 22918 31260 22924
rect 31114 22672 31170 22681
rect 31114 22607 31170 22616
rect 30748 22568 30800 22574
rect 30748 22510 30800 22516
rect 30840 22568 30892 22574
rect 30840 22510 30892 22516
rect 30760 22137 30788 22510
rect 30746 22128 30802 22137
rect 30746 22063 30802 22072
rect 31128 21962 31156 22607
rect 31220 21962 31248 22918
rect 31312 22234 31340 24670
rect 31484 24404 31536 24410
rect 31484 24346 31536 24352
rect 31496 23526 31524 24346
rect 31852 24336 31904 24342
rect 31852 24278 31904 24284
rect 32310 24304 32366 24313
rect 31484 23520 31536 23526
rect 31484 23462 31536 23468
rect 31668 23520 31720 23526
rect 31668 23462 31720 23468
rect 31680 23186 31708 23462
rect 31668 23180 31720 23186
rect 31668 23122 31720 23128
rect 31576 23044 31628 23050
rect 31576 22986 31628 22992
rect 31484 22432 31536 22438
rect 31482 22400 31484 22409
rect 31536 22400 31538 22409
rect 31482 22335 31538 22344
rect 31300 22228 31352 22234
rect 31300 22170 31352 22176
rect 31588 22098 31616 22986
rect 31760 22976 31812 22982
rect 31760 22918 31812 22924
rect 31666 22808 31722 22817
rect 31666 22743 31722 22752
rect 31680 22642 31708 22743
rect 31668 22636 31720 22642
rect 31668 22578 31720 22584
rect 31576 22092 31628 22098
rect 31576 22034 31628 22040
rect 31116 21956 31168 21962
rect 31116 21898 31168 21904
rect 31208 21956 31260 21962
rect 31208 21898 31260 21904
rect 31128 21690 31156 21898
rect 31300 21888 31352 21894
rect 31300 21830 31352 21836
rect 31392 21888 31444 21894
rect 31392 21830 31444 21836
rect 31116 21684 31168 21690
rect 31116 21626 31168 21632
rect 31024 21548 31076 21554
rect 31024 21490 31076 21496
rect 30840 21344 30892 21350
rect 30668 21304 30840 21332
rect 30380 21286 30432 21292
rect 30840 21286 30892 21292
rect 30286 21176 30342 21185
rect 30104 21140 30156 21146
rect 30286 21111 30288 21120
rect 30104 21082 30156 21088
rect 30340 21111 30342 21120
rect 30288 21082 30340 21088
rect 30288 20936 30340 20942
rect 30288 20878 30340 20884
rect 30104 20392 30156 20398
rect 30102 20360 30104 20369
rect 30196 20392 30248 20398
rect 30156 20360 30158 20369
rect 30196 20334 30248 20340
rect 30102 20295 30158 20304
rect 30012 20052 30064 20058
rect 30012 19994 30064 20000
rect 30010 19680 30066 19689
rect 30010 19615 30066 19624
rect 29920 19440 29972 19446
rect 29920 19382 29972 19388
rect 29736 18964 29788 18970
rect 29736 18906 29788 18912
rect 29828 18624 29880 18630
rect 29828 18566 29880 18572
rect 29644 18420 29696 18426
rect 29644 18362 29696 18368
rect 29734 17776 29790 17785
rect 29734 17711 29790 17720
rect 29460 17332 29512 17338
rect 29460 17274 29512 17280
rect 29552 17196 29604 17202
rect 29552 17138 29604 17144
rect 29276 16788 29328 16794
rect 29276 16730 29328 16736
rect 29184 16516 29236 16522
rect 29184 16458 29236 16464
rect 29288 14958 29316 16730
rect 29564 14958 29592 17138
rect 29748 15638 29776 17711
rect 29736 15632 29788 15638
rect 29736 15574 29788 15580
rect 29644 15360 29696 15366
rect 29644 15302 29696 15308
rect 29276 14952 29328 14958
rect 29276 14894 29328 14900
rect 29552 14952 29604 14958
rect 29552 14894 29604 14900
rect 29460 14884 29512 14890
rect 29460 14826 29512 14832
rect 29472 14793 29500 14826
rect 29458 14784 29514 14793
rect 29458 14719 29514 14728
rect 29564 14249 29592 14894
rect 29550 14240 29606 14249
rect 29550 14175 29606 14184
rect 29552 13252 29604 13258
rect 29552 13194 29604 13200
rect 29564 12918 29592 13194
rect 29552 12912 29604 12918
rect 29552 12854 29604 12860
rect 29564 12442 29592 12854
rect 29552 12436 29604 12442
rect 29656 12434 29684 15302
rect 29736 15020 29788 15026
rect 29736 14962 29788 14968
rect 29748 13326 29776 14962
rect 29840 13394 29868 18566
rect 29932 17134 29960 19382
rect 30024 19378 30052 19615
rect 30208 19446 30236 20334
rect 30300 19854 30328 20878
rect 30288 19848 30340 19854
rect 30288 19790 30340 19796
rect 30196 19440 30248 19446
rect 30196 19382 30248 19388
rect 30012 19372 30064 19378
rect 30012 19314 30064 19320
rect 30024 18329 30052 19314
rect 30194 19272 30250 19281
rect 30194 19207 30250 19216
rect 30208 18834 30236 19207
rect 30196 18828 30248 18834
rect 30196 18770 30248 18776
rect 30288 18828 30340 18834
rect 30288 18770 30340 18776
rect 30010 18320 30066 18329
rect 30010 18255 30066 18264
rect 30194 18320 30250 18329
rect 30194 18255 30250 18264
rect 30208 18086 30236 18255
rect 30196 18080 30248 18086
rect 30196 18022 30248 18028
rect 30104 17876 30156 17882
rect 30104 17818 30156 17824
rect 29920 17128 29972 17134
rect 29920 17070 29972 17076
rect 29932 15978 29960 17070
rect 30012 16652 30064 16658
rect 30012 16594 30064 16600
rect 29920 15972 29972 15978
rect 29920 15914 29972 15920
rect 30024 15586 30052 16594
rect 29932 15558 30052 15586
rect 29828 13388 29880 13394
rect 29828 13330 29880 13336
rect 29736 13320 29788 13326
rect 29736 13262 29788 13268
rect 29656 12406 29776 12434
rect 29552 12378 29604 12384
rect 29748 11558 29776 12406
rect 29736 11552 29788 11558
rect 29736 11494 29788 11500
rect 29092 11348 29144 11354
rect 29092 11290 29144 11296
rect 29276 11348 29328 11354
rect 29276 11290 29328 11296
rect 28908 10736 28960 10742
rect 28908 10678 28960 10684
rect 29092 10260 29144 10266
rect 29092 10202 29144 10208
rect 28632 9988 28684 9994
rect 28632 9930 28684 9936
rect 28908 9988 28960 9994
rect 28908 9930 28960 9936
rect 28540 9920 28592 9926
rect 28540 9862 28592 9868
rect 27950 9820 28258 9829
rect 27950 9818 27956 9820
rect 28012 9818 28036 9820
rect 28092 9818 28116 9820
rect 28172 9818 28196 9820
rect 28252 9818 28258 9820
rect 28012 9766 28014 9818
rect 28194 9766 28196 9818
rect 27950 9764 27956 9766
rect 28012 9764 28036 9766
rect 28092 9764 28116 9766
rect 28172 9764 28196 9766
rect 28252 9764 28258 9766
rect 27950 9755 28258 9764
rect 28920 9586 28948 9930
rect 28908 9580 28960 9586
rect 28908 9522 28960 9528
rect 28630 8936 28686 8945
rect 28630 8871 28686 8880
rect 28644 8838 28672 8871
rect 28632 8832 28684 8838
rect 28632 8774 28684 8780
rect 27950 8732 28258 8741
rect 27950 8730 27956 8732
rect 28012 8730 28036 8732
rect 28092 8730 28116 8732
rect 28172 8730 28196 8732
rect 28252 8730 28258 8732
rect 28012 8678 28014 8730
rect 28194 8678 28196 8730
rect 27950 8676 27956 8678
rect 28012 8676 28036 8678
rect 28092 8676 28116 8678
rect 28172 8676 28196 8678
rect 28252 8676 28258 8678
rect 27950 8667 28258 8676
rect 29104 8566 29132 10202
rect 29288 9722 29316 11290
rect 29736 11144 29788 11150
rect 29736 11086 29788 11092
rect 29748 10606 29776 11086
rect 29932 10792 29960 15558
rect 30012 15496 30064 15502
rect 30012 15438 30064 15444
rect 30024 14414 30052 15438
rect 30116 14822 30144 17818
rect 30208 16522 30236 18022
rect 30196 16516 30248 16522
rect 30196 16458 30248 16464
rect 30196 15972 30248 15978
rect 30196 15914 30248 15920
rect 30104 14816 30156 14822
rect 30104 14758 30156 14764
rect 30012 14408 30064 14414
rect 30012 14350 30064 14356
rect 30208 13954 30236 15914
rect 30300 15586 30328 18770
rect 30392 18290 30420 21286
rect 30852 20602 30880 21286
rect 30840 20596 30892 20602
rect 30840 20538 30892 20544
rect 30564 20256 30616 20262
rect 30564 20198 30616 20204
rect 30472 18760 30524 18766
rect 30472 18702 30524 18708
rect 30380 18284 30432 18290
rect 30380 18226 30432 18232
rect 30484 18086 30512 18702
rect 30472 18080 30524 18086
rect 30472 18022 30524 18028
rect 30380 17876 30432 17882
rect 30380 17818 30432 17824
rect 30392 17542 30420 17818
rect 30380 17536 30432 17542
rect 30380 17478 30432 17484
rect 30576 17134 30604 20198
rect 30838 19952 30894 19961
rect 30838 19887 30894 19896
rect 30852 19718 30880 19887
rect 30932 19780 30984 19786
rect 30932 19722 30984 19728
rect 30656 19712 30708 19718
rect 30840 19712 30892 19718
rect 30656 19654 30708 19660
rect 30760 19672 30840 19700
rect 30668 19446 30696 19654
rect 30656 19440 30708 19446
rect 30656 19382 30708 19388
rect 30760 19145 30788 19672
rect 30840 19654 30892 19660
rect 30944 19378 30972 19722
rect 30840 19372 30892 19378
rect 30840 19314 30892 19320
rect 30932 19372 30984 19378
rect 30932 19314 30984 19320
rect 30746 19136 30802 19145
rect 30746 19071 30802 19080
rect 30654 18592 30710 18601
rect 30654 18527 30710 18536
rect 30564 17128 30616 17134
rect 30564 17070 30616 17076
rect 30472 17060 30524 17066
rect 30472 17002 30524 17008
rect 30484 16250 30512 17002
rect 30668 16726 30696 18527
rect 30748 18352 30800 18358
rect 30748 18294 30800 18300
rect 30656 16720 30708 16726
rect 30656 16662 30708 16668
rect 30472 16244 30524 16250
rect 30472 16186 30524 16192
rect 30300 15558 30420 15586
rect 30288 15428 30340 15434
rect 30288 15370 30340 15376
rect 30300 14482 30328 15370
rect 30392 15366 30420 15558
rect 30484 15434 30512 16186
rect 30656 16176 30708 16182
rect 30656 16118 30708 16124
rect 30472 15428 30524 15434
rect 30472 15370 30524 15376
rect 30380 15360 30432 15366
rect 30380 15302 30432 15308
rect 30392 14958 30420 15302
rect 30380 14952 30432 14958
rect 30380 14894 30432 14900
rect 30380 14544 30432 14550
rect 30380 14486 30432 14492
rect 30288 14476 30340 14482
rect 30288 14418 30340 14424
rect 30116 13926 30236 13954
rect 30116 13462 30144 13926
rect 30104 13456 30156 13462
rect 30104 13398 30156 13404
rect 30116 12850 30144 13398
rect 30288 13388 30340 13394
rect 30288 13330 30340 13336
rect 30196 13252 30248 13258
rect 30196 13194 30248 13200
rect 30208 12918 30236 13194
rect 30196 12912 30248 12918
rect 30196 12854 30248 12860
rect 30104 12844 30156 12850
rect 30104 12786 30156 12792
rect 30012 12640 30064 12646
rect 30012 12582 30064 12588
rect 30024 12306 30052 12582
rect 30012 12300 30064 12306
rect 30012 12242 30064 12248
rect 30300 11098 30328 13330
rect 30392 12714 30420 14486
rect 30668 14006 30696 16118
rect 30760 15094 30788 18294
rect 30852 17678 30880 19314
rect 30932 17740 30984 17746
rect 30932 17682 30984 17688
rect 30840 17672 30892 17678
rect 30840 17614 30892 17620
rect 30944 17270 30972 17682
rect 30932 17264 30984 17270
rect 30932 17206 30984 17212
rect 31036 17116 31064 21490
rect 31208 21480 31260 21486
rect 31208 21422 31260 21428
rect 31220 21146 31248 21422
rect 31208 21140 31260 21146
rect 31208 21082 31260 21088
rect 31114 20904 31170 20913
rect 31114 20839 31170 20848
rect 31128 20641 31156 20839
rect 31208 20800 31260 20806
rect 31208 20742 31260 20748
rect 31114 20632 31170 20641
rect 31114 20567 31116 20576
rect 31168 20567 31170 20576
rect 31116 20538 31168 20544
rect 31116 20256 31168 20262
rect 31116 20198 31168 20204
rect 30852 17088 31064 17116
rect 30748 15088 30800 15094
rect 30748 15030 30800 15036
rect 30656 14000 30708 14006
rect 30656 13942 30708 13948
rect 30668 13258 30696 13942
rect 30656 13252 30708 13258
rect 30656 13194 30708 13200
rect 30668 12850 30696 13194
rect 30656 12844 30708 12850
rect 30656 12786 30708 12792
rect 30380 12708 30432 12714
rect 30380 12650 30432 12656
rect 30760 12306 30788 15030
rect 30852 13870 30880 17088
rect 30932 16992 30984 16998
rect 30932 16934 30984 16940
rect 31024 16992 31076 16998
rect 31024 16934 31076 16940
rect 30944 16250 30972 16934
rect 31036 16794 31064 16934
rect 31024 16788 31076 16794
rect 31024 16730 31076 16736
rect 31128 16250 31156 20198
rect 31220 18426 31248 20742
rect 31312 20262 31340 21830
rect 31300 20256 31352 20262
rect 31300 20198 31352 20204
rect 31404 20058 31432 21830
rect 31588 21486 31616 22034
rect 31484 21480 31536 21486
rect 31484 21422 31536 21428
rect 31576 21480 31628 21486
rect 31576 21422 31628 21428
rect 31496 20874 31524 21422
rect 31484 20868 31536 20874
rect 31484 20810 31536 20816
rect 31588 20398 31616 21422
rect 31576 20392 31628 20398
rect 31576 20334 31628 20340
rect 31392 20052 31444 20058
rect 31392 19994 31444 20000
rect 31588 19446 31616 20334
rect 31772 19922 31800 22918
rect 31760 19916 31812 19922
rect 31760 19858 31812 19864
rect 31864 19802 31892 24278
rect 32310 24239 32366 24248
rect 31944 24064 31996 24070
rect 31944 24006 31996 24012
rect 31726 19774 31892 19802
rect 31726 19666 31754 19774
rect 31726 19638 31800 19666
rect 31772 19514 31800 19638
rect 31760 19508 31812 19514
rect 31760 19450 31812 19456
rect 31300 19440 31352 19446
rect 31300 19382 31352 19388
rect 31576 19440 31628 19446
rect 31576 19382 31628 19388
rect 31208 18420 31260 18426
rect 31208 18362 31260 18368
rect 31312 17202 31340 19382
rect 31576 18352 31628 18358
rect 31576 18294 31628 18300
rect 31484 17536 31536 17542
rect 31484 17478 31536 17484
rect 31300 17196 31352 17202
rect 31300 17138 31352 17144
rect 31392 16652 31444 16658
rect 31392 16594 31444 16600
rect 31300 16448 31352 16454
rect 31300 16390 31352 16396
rect 30932 16244 30984 16250
rect 30932 16186 30984 16192
rect 31116 16244 31168 16250
rect 31116 16186 31168 16192
rect 31208 16040 31260 16046
rect 31208 15982 31260 15988
rect 31116 15360 31168 15366
rect 31116 15302 31168 15308
rect 31128 15162 31156 15302
rect 31116 15156 31168 15162
rect 31116 15098 31168 15104
rect 31116 14952 31168 14958
rect 31116 14894 31168 14900
rect 31128 14414 31156 14894
rect 30932 14408 30984 14414
rect 30932 14350 30984 14356
rect 31116 14408 31168 14414
rect 31116 14350 31168 14356
rect 30840 13864 30892 13870
rect 30840 13806 30892 13812
rect 30944 13734 30972 14350
rect 31024 14272 31076 14278
rect 31024 14214 31076 14220
rect 30932 13728 30984 13734
rect 30932 13670 30984 13676
rect 30748 12300 30800 12306
rect 30748 12242 30800 12248
rect 30472 11756 30524 11762
rect 30472 11698 30524 11704
rect 30208 11070 30420 11098
rect 29932 10764 30052 10792
rect 29920 10668 29972 10674
rect 29920 10610 29972 10616
rect 29736 10600 29788 10606
rect 29736 10542 29788 10548
rect 29276 9716 29328 9722
rect 29276 9658 29328 9664
rect 29644 9580 29696 9586
rect 29644 9522 29696 9528
rect 29656 8566 29684 9522
rect 29748 9518 29776 10542
rect 29736 9512 29788 9518
rect 29736 9454 29788 9460
rect 29748 9382 29776 9454
rect 29736 9376 29788 9382
rect 29736 9318 29788 9324
rect 29092 8560 29144 8566
rect 29092 8502 29144 8508
rect 29644 8560 29696 8566
rect 29644 8502 29696 8508
rect 28816 8424 28868 8430
rect 28816 8366 28868 8372
rect 27950 7644 28258 7653
rect 27950 7642 27956 7644
rect 28012 7642 28036 7644
rect 28092 7642 28116 7644
rect 28172 7642 28196 7644
rect 28252 7642 28258 7644
rect 28012 7590 28014 7642
rect 28194 7590 28196 7642
rect 27950 7588 27956 7590
rect 28012 7588 28036 7590
rect 28092 7588 28116 7590
rect 28172 7588 28196 7590
rect 28252 7588 28258 7590
rect 27950 7579 28258 7588
rect 27804 7336 27856 7342
rect 27804 7278 27856 7284
rect 27620 6724 27672 6730
rect 27620 6666 27672 6672
rect 27950 6556 28258 6565
rect 27950 6554 27956 6556
rect 28012 6554 28036 6556
rect 28092 6554 28116 6556
rect 28172 6554 28196 6556
rect 28252 6554 28258 6556
rect 28012 6502 28014 6554
rect 28194 6502 28196 6554
rect 27950 6500 27956 6502
rect 28012 6500 28036 6502
rect 28092 6500 28116 6502
rect 28172 6500 28196 6502
rect 28252 6500 28258 6502
rect 27950 6491 28258 6500
rect 27950 5468 28258 5477
rect 27950 5466 27956 5468
rect 28012 5466 28036 5468
rect 28092 5466 28116 5468
rect 28172 5466 28196 5468
rect 28252 5466 28258 5468
rect 28012 5414 28014 5466
rect 28194 5414 28196 5466
rect 27950 5412 27956 5414
rect 28012 5412 28036 5414
rect 28092 5412 28116 5414
rect 28172 5412 28196 5414
rect 28252 5412 28258 5414
rect 27950 5403 28258 5412
rect 28724 4752 28776 4758
rect 28724 4694 28776 4700
rect 27528 4616 27580 4622
rect 27528 4558 27580 4564
rect 27950 4380 28258 4389
rect 27950 4378 27956 4380
rect 28012 4378 28036 4380
rect 28092 4378 28116 4380
rect 28172 4378 28196 4380
rect 28252 4378 28258 4380
rect 28012 4326 28014 4378
rect 28194 4326 28196 4378
rect 27950 4324 27956 4326
rect 28012 4324 28036 4326
rect 28092 4324 28116 4326
rect 28172 4324 28196 4326
rect 28252 4324 28258 4326
rect 27950 4315 28258 4324
rect 27620 4072 27672 4078
rect 27620 4014 27672 4020
rect 27632 3505 27660 4014
rect 27804 3528 27856 3534
rect 27618 3496 27674 3505
rect 27804 3470 27856 3476
rect 27618 3431 27674 3440
rect 27160 3392 27212 3398
rect 27160 3334 27212 3340
rect 27528 3120 27580 3126
rect 27528 3062 27580 3068
rect 26148 3052 26200 3058
rect 26148 2994 26200 3000
rect 24492 2984 24544 2990
rect 24492 2926 24544 2932
rect 25872 2984 25924 2990
rect 25872 2926 25924 2932
rect 27540 2922 27568 3062
rect 27528 2916 27580 2922
rect 27528 2858 27580 2864
rect 27816 2854 27844 3470
rect 27950 3292 28258 3301
rect 27950 3290 27956 3292
rect 28012 3290 28036 3292
rect 28092 3290 28116 3292
rect 28172 3290 28196 3292
rect 28252 3290 28258 3292
rect 28012 3238 28014 3290
rect 28194 3238 28196 3290
rect 27950 3236 27956 3238
rect 28012 3236 28036 3238
rect 28092 3236 28116 3238
rect 28172 3236 28196 3238
rect 28252 3236 28258 3238
rect 27950 3227 28258 3236
rect 24584 2848 24636 2854
rect 24584 2790 24636 2796
rect 27160 2848 27212 2854
rect 27160 2790 27212 2796
rect 27804 2848 27856 2854
rect 27804 2790 27856 2796
rect 24124 2576 24176 2582
rect 24124 2518 24176 2524
rect 24400 2508 24452 2514
rect 24400 2450 24452 2456
rect 22376 2440 22428 2446
rect 22376 2382 22428 2388
rect 24412 800 24440 2450
rect 24596 2446 24624 2790
rect 26516 2508 26568 2514
rect 26516 2450 26568 2456
rect 24584 2440 24636 2446
rect 24584 2382 24636 2388
rect 26528 800 26556 2450
rect 27172 2446 27200 2790
rect 27160 2440 27212 2446
rect 27160 2382 27212 2388
rect 28632 2440 28684 2446
rect 28632 2382 28684 2388
rect 27950 2204 28258 2213
rect 27950 2202 27956 2204
rect 28012 2202 28036 2204
rect 28092 2202 28116 2204
rect 28172 2202 28196 2204
rect 28252 2202 28258 2204
rect 28012 2150 28014 2202
rect 28194 2150 28196 2202
rect 27950 2148 27956 2150
rect 28012 2148 28036 2150
rect 28092 2148 28116 2150
rect 28172 2148 28196 2150
rect 28252 2148 28258 2150
rect 27950 2139 28258 2148
rect 28644 800 28672 2382
rect 28736 2310 28764 4694
rect 28828 3058 28856 8366
rect 28908 3664 28960 3670
rect 28908 3606 28960 3612
rect 28816 3052 28868 3058
rect 28816 2994 28868 3000
rect 28920 2650 28948 3606
rect 29656 3126 29684 8502
rect 29748 8430 29776 9318
rect 29736 8424 29788 8430
rect 29736 8366 29788 8372
rect 29932 8090 29960 10610
rect 30024 9518 30052 10764
rect 30208 10266 30236 11070
rect 30288 11008 30340 11014
rect 30288 10950 30340 10956
rect 30300 10742 30328 10950
rect 30392 10742 30420 11070
rect 30288 10736 30340 10742
rect 30288 10678 30340 10684
rect 30380 10736 30432 10742
rect 30380 10678 30432 10684
rect 30380 10600 30432 10606
rect 30380 10542 30432 10548
rect 30196 10260 30248 10266
rect 30196 10202 30248 10208
rect 30392 9722 30420 10542
rect 30484 10266 30512 11698
rect 31036 11218 31064 14214
rect 31116 13728 31168 13734
rect 31116 13670 31168 13676
rect 31128 13190 31156 13670
rect 31116 13184 31168 13190
rect 31116 13126 31168 13132
rect 31116 12844 31168 12850
rect 31116 12786 31168 12792
rect 31128 12238 31156 12786
rect 31220 12782 31248 15982
rect 31312 15706 31340 16390
rect 31300 15700 31352 15706
rect 31300 15642 31352 15648
rect 31300 14816 31352 14822
rect 31300 14758 31352 14764
rect 31312 14482 31340 14758
rect 31300 14476 31352 14482
rect 31300 14418 31352 14424
rect 31312 14074 31340 14418
rect 31300 14068 31352 14074
rect 31300 14010 31352 14016
rect 31208 12776 31260 12782
rect 31208 12718 31260 12724
rect 31404 12434 31432 16594
rect 31312 12406 31432 12434
rect 31208 12300 31260 12306
rect 31208 12242 31260 12248
rect 31116 12232 31168 12238
rect 31116 12174 31168 12180
rect 31024 11212 31076 11218
rect 31024 11154 31076 11160
rect 31128 10742 31156 12174
rect 31220 11762 31248 12242
rect 31208 11756 31260 11762
rect 31208 11698 31260 11704
rect 31116 10736 31168 10742
rect 31116 10678 31168 10684
rect 31208 10532 31260 10538
rect 31208 10474 31260 10480
rect 30472 10260 30524 10266
rect 30472 10202 30524 10208
rect 30380 9716 30432 9722
rect 30380 9658 30432 9664
rect 30012 9512 30064 9518
rect 30012 9454 30064 9460
rect 30104 9512 30156 9518
rect 30104 9454 30156 9460
rect 30024 9042 30052 9454
rect 30116 9110 30144 9454
rect 30104 9104 30156 9110
rect 30104 9046 30156 9052
rect 30012 9036 30064 9042
rect 30012 8978 30064 8984
rect 30024 8838 30052 8978
rect 30012 8832 30064 8838
rect 30012 8774 30064 8780
rect 29920 8084 29972 8090
rect 29920 8026 29972 8032
rect 30484 6390 30512 10202
rect 31220 10130 31248 10474
rect 31312 10146 31340 12406
rect 31392 12096 31444 12102
rect 31392 12038 31444 12044
rect 31404 11694 31432 12038
rect 31392 11688 31444 11694
rect 31392 11630 31444 11636
rect 31392 11076 31444 11082
rect 31392 11018 31444 11024
rect 31404 10266 31432 11018
rect 31496 10985 31524 17478
rect 31588 16658 31616 18294
rect 31668 17740 31720 17746
rect 31668 17682 31720 17688
rect 31576 16652 31628 16658
rect 31576 16594 31628 16600
rect 31680 14822 31708 17682
rect 31772 16250 31800 19450
rect 31956 19378 31984 24006
rect 32126 23080 32182 23089
rect 32126 23015 32128 23024
rect 32180 23015 32182 23024
rect 32128 22986 32180 22992
rect 32220 22228 32272 22234
rect 32220 22170 32272 22176
rect 32232 20942 32260 22170
rect 32220 20936 32272 20942
rect 32220 20878 32272 20884
rect 32036 20800 32088 20806
rect 32036 20742 32088 20748
rect 32048 19854 32076 20742
rect 32218 20088 32274 20097
rect 32324 20074 32352 24239
rect 32404 23656 32456 23662
rect 32404 23598 32456 23604
rect 32416 22098 32444 23598
rect 32508 22778 32536 26200
rect 32864 24812 32916 24818
rect 32864 24754 32916 24760
rect 32680 23724 32732 23730
rect 32680 23666 32732 23672
rect 32586 22944 32642 22953
rect 32586 22879 32642 22888
rect 32496 22772 32548 22778
rect 32496 22714 32548 22720
rect 32600 22710 32628 22879
rect 32588 22704 32640 22710
rect 32588 22646 32640 22652
rect 32404 22092 32456 22098
rect 32404 22034 32456 22040
rect 32692 21894 32720 23666
rect 32876 23662 32904 24754
rect 33152 24721 33180 26200
rect 33138 24712 33194 24721
rect 33138 24647 33194 24656
rect 32950 24508 33258 24517
rect 32950 24506 32956 24508
rect 33012 24506 33036 24508
rect 33092 24506 33116 24508
rect 33172 24506 33196 24508
rect 33252 24506 33258 24508
rect 33012 24454 33014 24506
rect 33194 24454 33196 24506
rect 32950 24452 32956 24454
rect 33012 24452 33036 24454
rect 33092 24452 33116 24454
rect 33172 24452 33196 24454
rect 33252 24452 33258 24454
rect 32950 24443 33258 24452
rect 32864 23656 32916 23662
rect 32770 23624 32826 23633
rect 32864 23598 32916 23604
rect 33324 23656 33376 23662
rect 33324 23598 33376 23604
rect 32770 23559 32826 23568
rect 32680 21888 32732 21894
rect 32494 21856 32550 21865
rect 32680 21830 32732 21836
rect 32494 21791 32550 21800
rect 32508 21622 32536 21791
rect 32496 21616 32548 21622
rect 32496 21558 32548 21564
rect 32508 20806 32536 21558
rect 32680 21412 32732 21418
rect 32680 21354 32732 21360
rect 32496 20800 32548 20806
rect 32496 20742 32548 20748
rect 32496 20528 32548 20534
rect 32496 20470 32548 20476
rect 32274 20046 32352 20074
rect 32218 20023 32274 20032
rect 32128 19916 32180 19922
rect 32128 19858 32180 19864
rect 32036 19848 32088 19854
rect 32036 19790 32088 19796
rect 31944 19372 31996 19378
rect 31944 19314 31996 19320
rect 31852 18624 31904 18630
rect 31852 18566 31904 18572
rect 31864 16522 31892 18566
rect 31956 17610 31984 19314
rect 32140 19310 32168 19858
rect 32128 19304 32180 19310
rect 32128 19246 32180 19252
rect 32036 18284 32088 18290
rect 32036 18226 32088 18232
rect 31944 17604 31996 17610
rect 31944 17546 31996 17552
rect 32048 17338 32076 18226
rect 32232 17610 32260 20023
rect 32508 19938 32536 20470
rect 32588 20392 32640 20398
rect 32588 20334 32640 20340
rect 32600 20233 32628 20334
rect 32586 20224 32642 20233
rect 32586 20159 32642 20168
rect 32416 19910 32536 19938
rect 32416 19378 32444 19910
rect 32692 19514 32720 21354
rect 32588 19508 32640 19514
rect 32588 19450 32640 19456
rect 32680 19508 32732 19514
rect 32680 19450 32732 19456
rect 32404 19372 32456 19378
rect 32404 19314 32456 19320
rect 32416 18222 32444 19314
rect 32496 18964 32548 18970
rect 32496 18906 32548 18912
rect 32508 18766 32536 18906
rect 32496 18760 32548 18766
rect 32496 18702 32548 18708
rect 32496 18624 32548 18630
rect 32496 18566 32548 18572
rect 32404 18216 32456 18222
rect 32404 18158 32456 18164
rect 32220 17604 32272 17610
rect 32220 17546 32272 17552
rect 32036 17332 32088 17338
rect 32036 17274 32088 17280
rect 31852 16516 31904 16522
rect 31852 16458 31904 16464
rect 31760 16244 31812 16250
rect 31760 16186 31812 16192
rect 31944 16040 31996 16046
rect 31944 15982 31996 15988
rect 31760 15360 31812 15366
rect 31760 15302 31812 15308
rect 31772 15026 31800 15302
rect 31760 15020 31812 15026
rect 31760 14962 31812 14968
rect 31668 14816 31720 14822
rect 31668 14758 31720 14764
rect 31668 14544 31720 14550
rect 31668 14486 31720 14492
rect 31680 14346 31708 14486
rect 31668 14340 31720 14346
rect 31668 14282 31720 14288
rect 31668 14068 31720 14074
rect 31668 14010 31720 14016
rect 31576 12844 31628 12850
rect 31576 12786 31628 12792
rect 31588 12238 31616 12786
rect 31576 12232 31628 12238
rect 31576 12174 31628 12180
rect 31680 11082 31708 14010
rect 31760 13796 31812 13802
rect 31760 13738 31812 13744
rect 31772 13394 31800 13738
rect 31760 13388 31812 13394
rect 31760 13330 31812 13336
rect 31852 13388 31904 13394
rect 31852 13330 31904 13336
rect 31772 12850 31800 13330
rect 31864 12918 31892 13330
rect 31956 12986 31984 15982
rect 32048 15366 32076 17274
rect 32312 17196 32364 17202
rect 32312 17138 32364 17144
rect 32220 17128 32272 17134
rect 32220 17070 32272 17076
rect 32232 15978 32260 17070
rect 32324 16658 32352 17138
rect 32312 16652 32364 16658
rect 32312 16594 32364 16600
rect 32404 16244 32456 16250
rect 32404 16186 32456 16192
rect 32220 15972 32272 15978
rect 32220 15914 32272 15920
rect 32128 15904 32180 15910
rect 32128 15846 32180 15852
rect 32036 15360 32088 15366
rect 32036 15302 32088 15308
rect 32036 15156 32088 15162
rect 32036 15098 32088 15104
rect 32048 14396 32076 15098
rect 32140 14498 32168 15846
rect 32232 15706 32260 15914
rect 32312 15904 32364 15910
rect 32312 15846 32364 15852
rect 32220 15700 32272 15706
rect 32220 15642 32272 15648
rect 32324 15162 32352 15846
rect 32416 15570 32444 16186
rect 32404 15564 32456 15570
rect 32404 15506 32456 15512
rect 32404 15360 32456 15366
rect 32404 15302 32456 15308
rect 32312 15156 32364 15162
rect 32312 15098 32364 15104
rect 32220 14884 32272 14890
rect 32220 14826 32272 14832
rect 32232 14793 32260 14826
rect 32218 14784 32274 14793
rect 32218 14719 32274 14728
rect 32140 14482 32352 14498
rect 32140 14476 32364 14482
rect 32140 14470 32312 14476
rect 32312 14418 32364 14424
rect 32220 14408 32272 14414
rect 32048 14368 32168 14396
rect 32036 14272 32088 14278
rect 32036 14214 32088 14220
rect 32048 14006 32076 14214
rect 32036 14000 32088 14006
rect 32036 13942 32088 13948
rect 32036 13524 32088 13530
rect 32036 13466 32088 13472
rect 31944 12980 31996 12986
rect 31944 12922 31996 12928
rect 31852 12912 31904 12918
rect 31852 12854 31904 12860
rect 31760 12844 31812 12850
rect 31760 12786 31812 12792
rect 31956 12594 31984 12922
rect 31864 12566 31984 12594
rect 31760 12436 31812 12442
rect 31760 12378 31812 12384
rect 31772 11830 31800 12378
rect 31760 11824 31812 11830
rect 31760 11766 31812 11772
rect 31864 11234 31892 12566
rect 31942 12472 31998 12481
rect 31942 12407 31998 12416
rect 31956 11778 31984 12407
rect 32048 11937 32076 13466
rect 32140 12730 32168 14368
rect 32416 14362 32444 15302
rect 32508 14521 32536 18566
rect 32600 15094 32628 19450
rect 32784 18970 32812 23559
rect 32950 23420 33258 23429
rect 32950 23418 32956 23420
rect 33012 23418 33036 23420
rect 33092 23418 33116 23420
rect 33172 23418 33196 23420
rect 33252 23418 33258 23420
rect 33012 23366 33014 23418
rect 33194 23366 33196 23418
rect 32950 23364 32956 23366
rect 33012 23364 33036 23366
rect 33092 23364 33116 23366
rect 33172 23364 33196 23366
rect 33252 23364 33258 23366
rect 32950 23355 33258 23364
rect 33048 23316 33100 23322
rect 33048 23258 33100 23264
rect 32956 23248 33008 23254
rect 32876 23208 32956 23236
rect 32876 21418 32904 23208
rect 32956 23190 33008 23196
rect 33060 22982 33088 23258
rect 33336 23186 33364 23598
rect 33324 23180 33376 23186
rect 33324 23122 33376 23128
rect 33336 23066 33364 23122
rect 33152 23038 33364 23066
rect 33690 23080 33746 23089
rect 33048 22976 33100 22982
rect 33048 22918 33100 22924
rect 33060 22574 33088 22918
rect 33152 22642 33180 23038
rect 33690 23015 33746 23024
rect 33324 22976 33376 22982
rect 33324 22918 33376 22924
rect 33336 22710 33364 22918
rect 33704 22710 33732 23015
rect 33324 22704 33376 22710
rect 33324 22646 33376 22652
rect 33692 22704 33744 22710
rect 33692 22646 33744 22652
rect 33140 22636 33192 22642
rect 33140 22578 33192 22584
rect 33048 22568 33100 22574
rect 33048 22510 33100 22516
rect 32950 22332 33258 22341
rect 32950 22330 32956 22332
rect 33012 22330 33036 22332
rect 33092 22330 33116 22332
rect 33172 22330 33196 22332
rect 33252 22330 33258 22332
rect 33012 22278 33014 22330
rect 33194 22278 33196 22330
rect 32950 22276 32956 22278
rect 33012 22276 33036 22278
rect 33092 22276 33116 22278
rect 33172 22276 33196 22278
rect 33252 22276 33258 22278
rect 32950 22267 33258 22276
rect 33416 21888 33468 21894
rect 33416 21830 33468 21836
rect 33428 21622 33456 21830
rect 33704 21622 33732 22646
rect 33416 21616 33468 21622
rect 33416 21558 33468 21564
rect 33692 21616 33744 21622
rect 33692 21558 33744 21564
rect 33416 21480 33468 21486
rect 33796 21457 33824 26200
rect 35084 24834 35112 26200
rect 35084 24806 35204 24834
rect 35072 24676 35124 24682
rect 35072 24618 35124 24624
rect 34980 24608 35032 24614
rect 34980 24550 35032 24556
rect 33968 24064 34020 24070
rect 33968 24006 34020 24012
rect 34888 24064 34940 24070
rect 34888 24006 34940 24012
rect 33980 23866 34008 24006
rect 33968 23860 34020 23866
rect 33968 23802 34020 23808
rect 34152 23792 34204 23798
rect 34152 23734 34204 23740
rect 34336 23792 34388 23798
rect 34900 23746 34928 24006
rect 34992 23882 35020 24550
rect 35084 24206 35112 24618
rect 35072 24200 35124 24206
rect 35072 24142 35124 24148
rect 34992 23854 35112 23882
rect 34336 23734 34388 23740
rect 33876 23656 33928 23662
rect 34164 23644 34192 23734
rect 34244 23656 34296 23662
rect 34164 23616 34244 23644
rect 33876 23598 33928 23604
rect 34244 23598 34296 23604
rect 33888 22574 33916 23598
rect 34348 23089 34376 23734
rect 34808 23718 34928 23746
rect 34702 23352 34758 23361
rect 34702 23287 34704 23296
rect 34756 23287 34758 23296
rect 34704 23258 34756 23264
rect 34612 23180 34664 23186
rect 34612 23122 34664 23128
rect 34334 23080 34390 23089
rect 34334 23015 34390 23024
rect 33876 22568 33928 22574
rect 33876 22510 33928 22516
rect 33888 22166 33916 22510
rect 33876 22160 33928 22166
rect 33876 22102 33928 22108
rect 34152 22024 34204 22030
rect 34150 21992 34152 22001
rect 34204 21992 34206 22001
rect 34150 21927 34206 21936
rect 33876 21616 33928 21622
rect 33876 21558 33928 21564
rect 33416 21422 33468 21428
rect 33782 21448 33838 21457
rect 32864 21412 32916 21418
rect 32864 21354 32916 21360
rect 32950 21244 33258 21253
rect 32950 21242 32956 21244
rect 33012 21242 33036 21244
rect 33092 21242 33116 21244
rect 33172 21242 33196 21244
rect 33252 21242 33258 21244
rect 33012 21190 33014 21242
rect 33194 21190 33196 21242
rect 32950 21188 32956 21190
rect 33012 21188 33036 21190
rect 33092 21188 33116 21190
rect 33172 21188 33196 21190
rect 33252 21188 33258 21190
rect 32950 21179 33258 21188
rect 33140 21140 33192 21146
rect 33140 21082 33192 21088
rect 33152 20874 33180 21082
rect 33428 21010 33456 21422
rect 33782 21383 33838 21392
rect 33416 21004 33468 21010
rect 33416 20946 33468 20952
rect 33692 21004 33744 21010
rect 33692 20946 33744 20952
rect 33140 20868 33192 20874
rect 33140 20810 33192 20816
rect 32864 20800 32916 20806
rect 32864 20742 32916 20748
rect 32876 19514 32904 20742
rect 33428 20602 33456 20946
rect 33416 20596 33468 20602
rect 33416 20538 33468 20544
rect 33600 20392 33652 20398
rect 33600 20334 33652 20340
rect 33612 20233 33640 20334
rect 33598 20224 33654 20233
rect 32950 20156 33258 20165
rect 33598 20159 33654 20168
rect 32950 20154 32956 20156
rect 33012 20154 33036 20156
rect 33092 20154 33116 20156
rect 33172 20154 33196 20156
rect 33252 20154 33258 20156
rect 33012 20102 33014 20154
rect 33194 20102 33196 20154
rect 32950 20100 32956 20102
rect 33012 20100 33036 20102
rect 33092 20100 33116 20102
rect 33172 20100 33196 20102
rect 33252 20100 33258 20102
rect 32950 20091 33258 20100
rect 33508 19984 33560 19990
rect 33508 19926 33560 19932
rect 33416 19916 33468 19922
rect 33416 19858 33468 19864
rect 32864 19508 32916 19514
rect 32864 19450 32916 19456
rect 33428 19334 33456 19858
rect 33520 19514 33548 19926
rect 33508 19508 33560 19514
rect 33508 19450 33560 19456
rect 32864 19304 32916 19310
rect 33428 19306 33548 19334
rect 32864 19246 32916 19252
rect 32772 18964 32824 18970
rect 32772 18906 32824 18912
rect 32772 17876 32824 17882
rect 32772 17818 32824 17824
rect 32680 17808 32732 17814
rect 32680 17750 32732 17756
rect 32692 17134 32720 17750
rect 32680 17128 32732 17134
rect 32680 17070 32732 17076
rect 32784 16250 32812 17818
rect 32772 16244 32824 16250
rect 32772 16186 32824 16192
rect 32876 16046 32904 19246
rect 33324 19168 33376 19174
rect 33324 19110 33376 19116
rect 32950 19068 33258 19077
rect 32950 19066 32956 19068
rect 33012 19066 33036 19068
rect 33092 19066 33116 19068
rect 33172 19066 33196 19068
rect 33252 19066 33258 19068
rect 33012 19014 33014 19066
rect 33194 19014 33196 19066
rect 32950 19012 32956 19014
rect 33012 19012 33036 19014
rect 33092 19012 33116 19014
rect 33172 19012 33196 19014
rect 33252 19012 33258 19014
rect 32950 19003 33258 19012
rect 32956 18964 33008 18970
rect 32956 18906 33008 18912
rect 32968 18834 32996 18906
rect 33046 18864 33102 18873
rect 32956 18828 33008 18834
rect 33046 18799 33048 18808
rect 32956 18770 33008 18776
rect 33100 18799 33102 18808
rect 33048 18770 33100 18776
rect 33060 18601 33088 18770
rect 33046 18592 33102 18601
rect 33046 18527 33102 18536
rect 32950 17980 33258 17989
rect 32950 17978 32956 17980
rect 33012 17978 33036 17980
rect 33092 17978 33116 17980
rect 33172 17978 33196 17980
rect 33252 17978 33258 17980
rect 33012 17926 33014 17978
rect 33194 17926 33196 17978
rect 32950 17924 32956 17926
rect 33012 17924 33036 17926
rect 33092 17924 33116 17926
rect 33172 17924 33196 17926
rect 33252 17924 33258 17926
rect 32950 17915 33258 17924
rect 33232 17740 33284 17746
rect 33336 17728 33364 19110
rect 33416 18624 33468 18630
rect 33416 18566 33468 18572
rect 33428 18222 33456 18566
rect 33416 18216 33468 18222
rect 33416 18158 33468 18164
rect 33284 17700 33364 17728
rect 33232 17682 33284 17688
rect 32950 16892 33258 16901
rect 32950 16890 32956 16892
rect 33012 16890 33036 16892
rect 33092 16890 33116 16892
rect 33172 16890 33196 16892
rect 33252 16890 33258 16892
rect 33012 16838 33014 16890
rect 33194 16838 33196 16890
rect 32950 16836 32956 16838
rect 33012 16836 33036 16838
rect 33092 16836 33116 16838
rect 33172 16836 33196 16838
rect 33252 16836 33258 16838
rect 32950 16827 33258 16836
rect 33324 16652 33376 16658
rect 33428 16640 33456 18158
rect 33376 16612 33456 16640
rect 33324 16594 33376 16600
rect 33324 16108 33376 16114
rect 33324 16050 33376 16056
rect 32864 16040 32916 16046
rect 32864 15982 32916 15988
rect 32950 15804 33258 15813
rect 32950 15802 32956 15804
rect 33012 15802 33036 15804
rect 33092 15802 33116 15804
rect 33172 15802 33196 15804
rect 33252 15802 33258 15804
rect 33012 15750 33014 15802
rect 33194 15750 33196 15802
rect 32950 15748 32956 15750
rect 33012 15748 33036 15750
rect 33092 15748 33116 15750
rect 33172 15748 33196 15750
rect 33252 15748 33258 15750
rect 32950 15739 33258 15748
rect 32588 15088 32640 15094
rect 32588 15030 32640 15036
rect 32680 14952 32732 14958
rect 32680 14894 32732 14900
rect 32772 14952 32824 14958
rect 32772 14894 32824 14900
rect 32494 14512 32550 14521
rect 32494 14447 32550 14456
rect 32220 14350 32272 14356
rect 32232 13870 32260 14350
rect 32324 14334 32444 14362
rect 32220 13864 32272 13870
rect 32220 13806 32272 13812
rect 32140 12702 32260 12730
rect 32128 12640 32180 12646
rect 32128 12582 32180 12588
rect 32034 11928 32090 11937
rect 32034 11863 32090 11872
rect 32140 11830 32168 12582
rect 32128 11824 32180 11830
rect 31956 11750 32076 11778
rect 32128 11766 32180 11772
rect 31944 11688 31996 11694
rect 32048 11676 32076 11750
rect 32048 11648 32168 11676
rect 31944 11630 31996 11636
rect 31772 11206 31892 11234
rect 31668 11076 31720 11082
rect 31668 11018 31720 11024
rect 31772 11014 31800 11206
rect 31760 11008 31812 11014
rect 31482 10976 31538 10985
rect 31956 10962 31984 11630
rect 31760 10950 31812 10956
rect 31482 10911 31538 10920
rect 31864 10934 31984 10962
rect 31760 10804 31812 10810
rect 31760 10746 31812 10752
rect 31772 10606 31800 10746
rect 31760 10600 31812 10606
rect 31760 10542 31812 10548
rect 31392 10260 31444 10266
rect 31392 10202 31444 10208
rect 31668 10192 31720 10198
rect 30748 10124 30800 10130
rect 30748 10066 30800 10072
rect 31208 10124 31260 10130
rect 31312 10118 31432 10146
rect 31668 10134 31720 10140
rect 31208 10066 31260 10072
rect 30564 9988 30616 9994
rect 30564 9930 30616 9936
rect 30656 9988 30708 9994
rect 30656 9930 30708 9936
rect 30576 7886 30604 9930
rect 30668 9722 30696 9930
rect 30656 9716 30708 9722
rect 30656 9658 30708 9664
rect 30668 8634 30696 9658
rect 30760 8974 30788 10066
rect 31404 9926 31432 10118
rect 31392 9920 31444 9926
rect 31392 9862 31444 9868
rect 31404 9722 31432 9862
rect 31300 9716 31352 9722
rect 31300 9658 31352 9664
rect 31392 9716 31444 9722
rect 31392 9658 31444 9664
rect 31312 9586 31340 9658
rect 31300 9580 31352 9586
rect 31300 9522 31352 9528
rect 30748 8968 30800 8974
rect 30748 8910 30800 8916
rect 30656 8628 30708 8634
rect 30656 8570 30708 8576
rect 30760 8566 30788 8910
rect 31680 8634 31708 10134
rect 31864 8945 31892 10934
rect 31944 10804 31996 10810
rect 31944 10746 31996 10752
rect 31956 10538 31984 10746
rect 32036 10736 32088 10742
rect 32036 10678 32088 10684
rect 31944 10532 31996 10538
rect 31944 10474 31996 10480
rect 32048 9994 32076 10678
rect 32036 9988 32088 9994
rect 32036 9930 32088 9936
rect 32048 9654 32076 9930
rect 32036 9648 32088 9654
rect 32036 9590 32088 9596
rect 32048 8974 32076 9590
rect 32036 8968 32088 8974
rect 31850 8936 31906 8945
rect 32036 8910 32088 8916
rect 31850 8871 31906 8880
rect 31668 8628 31720 8634
rect 31668 8570 31720 8576
rect 30748 8560 30800 8566
rect 30748 8502 30800 8508
rect 31392 8492 31444 8498
rect 31392 8434 31444 8440
rect 30564 7880 30616 7886
rect 30564 7822 30616 7828
rect 31404 7410 31432 8434
rect 31484 8288 31536 8294
rect 31484 8230 31536 8236
rect 31496 7546 31524 8230
rect 31760 7880 31812 7886
rect 31760 7822 31812 7828
rect 31852 7880 31904 7886
rect 31852 7822 31904 7828
rect 31484 7540 31536 7546
rect 31484 7482 31536 7488
rect 31392 7404 31444 7410
rect 31392 7346 31444 7352
rect 31772 7342 31800 7822
rect 31864 7546 31892 7822
rect 31852 7540 31904 7546
rect 31852 7482 31904 7488
rect 31760 7336 31812 7342
rect 31760 7278 31812 7284
rect 30472 6384 30524 6390
rect 30472 6326 30524 6332
rect 32140 6186 32168 11648
rect 32232 11626 32260 12702
rect 32324 12481 32352 14334
rect 32692 14278 32720 14894
rect 32496 14272 32548 14278
rect 32496 14214 32548 14220
rect 32680 14272 32732 14278
rect 32680 14214 32732 14220
rect 32310 12472 32366 12481
rect 32310 12407 32366 12416
rect 32508 12345 32536 14214
rect 32680 14000 32732 14006
rect 32586 13968 32642 13977
rect 32680 13942 32732 13948
rect 32586 13903 32642 13912
rect 32600 13870 32628 13903
rect 32692 13870 32720 13942
rect 32588 13864 32640 13870
rect 32588 13806 32640 13812
rect 32680 13864 32732 13870
rect 32680 13806 32732 13812
rect 32494 12336 32550 12345
rect 32494 12271 32550 12280
rect 32494 12200 32550 12209
rect 32494 12135 32496 12144
rect 32548 12135 32550 12144
rect 32496 12106 32548 12112
rect 32310 11928 32366 11937
rect 32310 11863 32366 11872
rect 32220 11620 32272 11626
rect 32220 11562 32272 11568
rect 32324 10282 32352 11863
rect 32600 11626 32628 13806
rect 32784 12986 32812 14894
rect 32950 14716 33258 14725
rect 32950 14714 32956 14716
rect 33012 14714 33036 14716
rect 33092 14714 33116 14716
rect 33172 14714 33196 14716
rect 33252 14714 33258 14716
rect 33012 14662 33014 14714
rect 33194 14662 33196 14714
rect 32950 14660 32956 14662
rect 33012 14660 33036 14662
rect 33092 14660 33116 14662
rect 33172 14660 33196 14662
rect 33252 14660 33258 14662
rect 32950 14651 33258 14660
rect 33336 14618 33364 16050
rect 33520 15570 33548 19306
rect 33704 18630 33732 20946
rect 33888 20534 33916 21558
rect 34624 21010 34652 23122
rect 34808 22545 34836 23718
rect 34888 23588 34940 23594
rect 34888 23530 34940 23536
rect 34794 22536 34850 22545
rect 34794 22471 34850 22480
rect 34900 22094 34928 23530
rect 35084 22982 35112 23854
rect 35176 23322 35204 24806
rect 35728 24682 35756 26200
rect 36544 24812 36596 24818
rect 36544 24754 36596 24760
rect 36268 24744 36320 24750
rect 36268 24686 36320 24692
rect 35716 24676 35768 24682
rect 35716 24618 35768 24624
rect 35624 24064 35676 24070
rect 35624 24006 35676 24012
rect 35256 23792 35308 23798
rect 35256 23734 35308 23740
rect 35164 23316 35216 23322
rect 35164 23258 35216 23264
rect 35072 22976 35124 22982
rect 35072 22918 35124 22924
rect 35164 22976 35216 22982
rect 35164 22918 35216 22924
rect 34900 22066 35020 22094
rect 34796 21888 34848 21894
rect 34796 21830 34848 21836
rect 34704 21548 34756 21554
rect 34704 21490 34756 21496
rect 34612 21004 34664 21010
rect 34612 20946 34664 20952
rect 34716 20942 34744 21490
rect 34808 21078 34836 21830
rect 34888 21684 34940 21690
rect 34888 21626 34940 21632
rect 34796 21072 34848 21078
rect 34796 21014 34848 21020
rect 34704 20936 34756 20942
rect 34704 20878 34756 20884
rect 34428 20868 34480 20874
rect 34428 20810 34480 20816
rect 34440 20534 34468 20810
rect 34518 20632 34574 20641
rect 34518 20567 34574 20576
rect 33876 20528 33928 20534
rect 33876 20470 33928 20476
rect 34428 20528 34480 20534
rect 34428 20470 34480 20476
rect 34060 20256 34112 20262
rect 34060 20198 34112 20204
rect 34072 19854 34100 20198
rect 34060 19848 34112 19854
rect 34060 19790 34112 19796
rect 34072 19718 34100 19790
rect 34060 19712 34112 19718
rect 34060 19654 34112 19660
rect 34336 19508 34388 19514
rect 34336 19450 34388 19456
rect 33966 19408 34022 19417
rect 33966 19343 34022 19352
rect 33980 19310 34008 19343
rect 33968 19304 34020 19310
rect 33968 19246 34020 19252
rect 33692 18624 33744 18630
rect 33692 18566 33744 18572
rect 33600 18216 33652 18222
rect 33600 18158 33652 18164
rect 33612 17338 33640 18158
rect 34244 17536 34296 17542
rect 34244 17478 34296 17484
rect 33600 17332 33652 17338
rect 33600 17274 33652 17280
rect 33876 16992 33928 16998
rect 33876 16934 33928 16940
rect 34060 16992 34112 16998
rect 34060 16934 34112 16940
rect 33600 16448 33652 16454
rect 33600 16390 33652 16396
rect 33508 15564 33560 15570
rect 33508 15506 33560 15512
rect 33416 15020 33468 15026
rect 33416 14962 33468 14968
rect 33428 14618 33456 14962
rect 33324 14612 33376 14618
rect 33324 14554 33376 14560
rect 33416 14612 33468 14618
rect 33416 14554 33468 14560
rect 32864 14476 32916 14482
rect 32864 14418 32916 14424
rect 33416 14476 33468 14482
rect 33416 14418 33468 14424
rect 32772 12980 32824 12986
rect 32772 12922 32824 12928
rect 32784 12209 32812 12922
rect 32876 12442 32904 14418
rect 32950 13628 33258 13637
rect 32950 13626 32956 13628
rect 33012 13626 33036 13628
rect 33092 13626 33116 13628
rect 33172 13626 33196 13628
rect 33252 13626 33258 13628
rect 33012 13574 33014 13626
rect 33194 13574 33196 13626
rect 32950 13572 32956 13574
rect 33012 13572 33036 13574
rect 33092 13572 33116 13574
rect 33172 13572 33196 13574
rect 33252 13572 33258 13574
rect 32950 13563 33258 13572
rect 32950 12540 33258 12549
rect 32950 12538 32956 12540
rect 33012 12538 33036 12540
rect 33092 12538 33116 12540
rect 33172 12538 33196 12540
rect 33252 12538 33258 12540
rect 33012 12486 33014 12538
rect 33194 12486 33196 12538
rect 32950 12484 32956 12486
rect 33012 12484 33036 12486
rect 33092 12484 33116 12486
rect 33172 12484 33196 12486
rect 33252 12484 33258 12486
rect 32950 12475 33258 12484
rect 32864 12436 32916 12442
rect 32864 12378 32916 12384
rect 32954 12336 33010 12345
rect 32954 12271 33010 12280
rect 32770 12200 32826 12209
rect 32826 12158 32904 12186
rect 32770 12135 32826 12144
rect 32588 11620 32640 11626
rect 32588 11562 32640 11568
rect 32772 11348 32824 11354
rect 32876 11336 32904 12158
rect 32968 11626 32996 12271
rect 33322 12200 33378 12209
rect 33322 12135 33378 12144
rect 32956 11620 33008 11626
rect 32956 11562 33008 11568
rect 32950 11452 33258 11461
rect 32950 11450 32956 11452
rect 33012 11450 33036 11452
rect 33092 11450 33116 11452
rect 33172 11450 33196 11452
rect 33252 11450 33258 11452
rect 33012 11398 33014 11450
rect 33194 11398 33196 11450
rect 32950 11396 32956 11398
rect 33012 11396 33036 11398
rect 33092 11396 33116 11398
rect 33172 11396 33196 11398
rect 33252 11396 33258 11398
rect 32950 11387 33258 11396
rect 32876 11308 32996 11336
rect 32772 11290 32824 11296
rect 32588 11280 32640 11286
rect 32588 11222 32640 11228
rect 32784 11234 32812 11290
rect 32324 10254 32536 10282
rect 32220 10124 32272 10130
rect 32220 10066 32272 10072
rect 32404 10124 32456 10130
rect 32404 10066 32456 10072
rect 32232 9654 32260 10066
rect 32220 9648 32272 9654
rect 32220 9590 32272 9596
rect 32312 9512 32364 9518
rect 32312 9454 32364 9460
rect 32324 9110 32352 9454
rect 32416 9382 32444 10066
rect 32508 9586 32536 10254
rect 32496 9580 32548 9586
rect 32496 9522 32548 9528
rect 32404 9376 32456 9382
rect 32404 9318 32456 9324
rect 32312 9104 32364 9110
rect 32312 9046 32364 9052
rect 32600 8566 32628 11222
rect 32784 11206 32904 11234
rect 32772 11076 32824 11082
rect 32772 11018 32824 11024
rect 32784 10742 32812 11018
rect 32772 10736 32824 10742
rect 32772 10678 32824 10684
rect 32680 10464 32732 10470
rect 32680 10406 32732 10412
rect 32692 10198 32720 10406
rect 32680 10192 32732 10198
rect 32680 10134 32732 10140
rect 32772 10192 32824 10198
rect 32772 10134 32824 10140
rect 32680 9920 32732 9926
rect 32680 9862 32732 9868
rect 32692 9178 32720 9862
rect 32680 9172 32732 9178
rect 32680 9114 32732 9120
rect 32784 8922 32812 10134
rect 32692 8894 32812 8922
rect 32876 8906 32904 11206
rect 32968 10606 32996 11308
rect 33336 11082 33364 12135
rect 33324 11076 33376 11082
rect 33324 11018 33376 11024
rect 32956 10600 33008 10606
rect 32956 10542 33008 10548
rect 32950 10364 33258 10373
rect 32950 10362 32956 10364
rect 33012 10362 33036 10364
rect 33092 10362 33116 10364
rect 33172 10362 33196 10364
rect 33252 10362 33258 10364
rect 33012 10310 33014 10362
rect 33194 10310 33196 10362
rect 32950 10308 32956 10310
rect 33012 10308 33036 10310
rect 33092 10308 33116 10310
rect 33172 10308 33196 10310
rect 33252 10308 33258 10310
rect 32950 10299 33258 10308
rect 33428 10062 33456 14418
rect 33520 11914 33548 15506
rect 33612 14482 33640 16390
rect 33784 16040 33836 16046
rect 33784 15982 33836 15988
rect 33692 15360 33744 15366
rect 33692 15302 33744 15308
rect 33704 15162 33732 15302
rect 33692 15156 33744 15162
rect 33692 15098 33744 15104
rect 33600 14476 33652 14482
rect 33600 14418 33652 14424
rect 33796 14346 33824 15982
rect 33784 14340 33836 14346
rect 33784 14282 33836 14288
rect 33692 13932 33744 13938
rect 33692 13874 33744 13880
rect 33600 13864 33652 13870
rect 33600 13806 33652 13812
rect 33612 13326 33640 13806
rect 33704 13462 33732 13874
rect 33692 13456 33744 13462
rect 33692 13398 33744 13404
rect 33600 13320 33652 13326
rect 33600 13262 33652 13268
rect 33612 12050 33640 13262
rect 33704 12850 33732 13398
rect 33796 13394 33824 14282
rect 33888 13530 33916 16934
rect 33968 16788 34020 16794
rect 33968 16730 34020 16736
rect 33980 16250 34008 16730
rect 34072 16658 34100 16934
rect 34060 16652 34112 16658
rect 34060 16594 34112 16600
rect 34060 16448 34112 16454
rect 34060 16390 34112 16396
rect 33968 16244 34020 16250
rect 33968 16186 34020 16192
rect 34072 15706 34100 16390
rect 34060 15700 34112 15706
rect 34112 15660 34192 15688
rect 34060 15642 34112 15648
rect 34060 15496 34112 15502
rect 34060 15438 34112 15444
rect 34072 15162 34100 15438
rect 34060 15156 34112 15162
rect 34060 15098 34112 15104
rect 34164 14958 34192 15660
rect 34152 14952 34204 14958
rect 34152 14894 34204 14900
rect 34060 14544 34112 14550
rect 34060 14486 34112 14492
rect 34072 14074 34100 14486
rect 34256 14278 34284 17478
rect 34244 14272 34296 14278
rect 34244 14214 34296 14220
rect 34060 14068 34112 14074
rect 34060 14010 34112 14016
rect 33876 13524 33928 13530
rect 33876 13466 33928 13472
rect 33874 13424 33930 13433
rect 33784 13388 33836 13394
rect 33874 13359 33876 13368
rect 33784 13330 33836 13336
rect 33928 13359 33930 13368
rect 34060 13388 34112 13394
rect 33876 13330 33928 13336
rect 34060 13330 34112 13336
rect 33876 13252 33928 13258
rect 33876 13194 33928 13200
rect 33692 12844 33744 12850
rect 33692 12786 33744 12792
rect 33704 12209 33732 12786
rect 33888 12442 33916 13194
rect 33876 12436 33928 12442
rect 33876 12378 33928 12384
rect 33690 12200 33746 12209
rect 33690 12135 33692 12144
rect 33744 12135 33746 12144
rect 33692 12106 33744 12112
rect 33612 12022 33916 12050
rect 33520 11886 33732 11914
rect 33508 11688 33560 11694
rect 33508 11630 33560 11636
rect 33520 10606 33548 11630
rect 33508 10600 33560 10606
rect 33508 10542 33560 10548
rect 33520 10130 33548 10542
rect 33598 10160 33654 10169
rect 33508 10124 33560 10130
rect 33598 10095 33654 10104
rect 33508 10066 33560 10072
rect 33416 10056 33468 10062
rect 33416 9998 33468 10004
rect 33520 9586 33548 10066
rect 33508 9580 33560 9586
rect 33508 9522 33560 9528
rect 32950 9276 33258 9285
rect 32950 9274 32956 9276
rect 33012 9274 33036 9276
rect 33092 9274 33116 9276
rect 33172 9274 33196 9276
rect 33252 9274 33258 9276
rect 33012 9222 33014 9274
rect 33194 9222 33196 9274
rect 32950 9220 32956 9222
rect 33012 9220 33036 9222
rect 33092 9220 33116 9222
rect 33172 9220 33196 9222
rect 33252 9220 33258 9222
rect 32950 9211 33258 9220
rect 32864 8900 32916 8906
rect 32588 8560 32640 8566
rect 32588 8502 32640 8508
rect 32600 7954 32628 8502
rect 32588 7948 32640 7954
rect 32588 7890 32640 7896
rect 32692 7750 32720 8894
rect 32864 8842 32916 8848
rect 33520 8634 33548 9522
rect 33612 9489 33640 10095
rect 33704 9518 33732 11886
rect 33784 11076 33836 11082
rect 33784 11018 33836 11024
rect 33796 10985 33824 11018
rect 33782 10976 33838 10985
rect 33782 10911 33838 10920
rect 33888 9908 33916 12022
rect 33968 11620 34020 11626
rect 33968 11562 34020 11568
rect 33980 11354 34008 11562
rect 33968 11348 34020 11354
rect 33968 11290 34020 11296
rect 34072 10690 34100 13330
rect 34152 13320 34204 13326
rect 34152 13262 34204 13268
rect 33980 10662 34100 10690
rect 33980 10033 34008 10662
rect 33966 10024 34022 10033
rect 33966 9959 34022 9968
rect 33796 9880 33916 9908
rect 33692 9512 33744 9518
rect 33598 9480 33654 9489
rect 33692 9454 33744 9460
rect 33598 9415 33654 9424
rect 33612 8974 33640 9415
rect 33600 8968 33652 8974
rect 33600 8910 33652 8916
rect 33796 8838 33824 9880
rect 33876 9444 33928 9450
rect 33876 9386 33928 9392
rect 33888 9042 33916 9386
rect 33876 9036 33928 9042
rect 33876 8978 33928 8984
rect 33784 8832 33836 8838
rect 33784 8774 33836 8780
rect 33508 8628 33560 8634
rect 33508 8570 33560 8576
rect 32950 8188 33258 8197
rect 32950 8186 32956 8188
rect 33012 8186 33036 8188
rect 33092 8186 33116 8188
rect 33172 8186 33196 8188
rect 33252 8186 33258 8188
rect 33012 8134 33014 8186
rect 33194 8134 33196 8186
rect 32950 8132 32956 8134
rect 33012 8132 33036 8134
rect 33092 8132 33116 8134
rect 33172 8132 33196 8134
rect 33252 8132 33258 8134
rect 32950 8123 33258 8132
rect 32772 7880 32824 7886
rect 32772 7822 32824 7828
rect 32784 7750 32812 7822
rect 32680 7744 32732 7750
rect 32680 7686 32732 7692
rect 32772 7744 32824 7750
rect 32772 7686 32824 7692
rect 32784 6866 32812 7686
rect 32950 7100 33258 7109
rect 32950 7098 32956 7100
rect 33012 7098 33036 7100
rect 33092 7098 33116 7100
rect 33172 7098 33196 7100
rect 33252 7098 33258 7100
rect 33012 7046 33014 7098
rect 33194 7046 33196 7098
rect 32950 7044 32956 7046
rect 33012 7044 33036 7046
rect 33092 7044 33116 7046
rect 33172 7044 33196 7046
rect 33252 7044 33258 7046
rect 32950 7035 33258 7044
rect 32772 6860 32824 6866
rect 32772 6802 32824 6808
rect 32128 6180 32180 6186
rect 32128 6122 32180 6128
rect 32950 6012 33258 6021
rect 32950 6010 32956 6012
rect 33012 6010 33036 6012
rect 33092 6010 33116 6012
rect 33172 6010 33196 6012
rect 33252 6010 33258 6012
rect 33012 5958 33014 6010
rect 33194 5958 33196 6010
rect 32950 5956 32956 5958
rect 33012 5956 33036 5958
rect 33092 5956 33116 5958
rect 33172 5956 33196 5958
rect 33252 5956 33258 5958
rect 32950 5947 33258 5956
rect 32950 4924 33258 4933
rect 32950 4922 32956 4924
rect 33012 4922 33036 4924
rect 33092 4922 33116 4924
rect 33172 4922 33196 4924
rect 33252 4922 33258 4924
rect 33012 4870 33014 4922
rect 33194 4870 33196 4922
rect 32950 4868 32956 4870
rect 33012 4868 33036 4870
rect 33092 4868 33116 4870
rect 33172 4868 33196 4870
rect 33252 4868 33258 4870
rect 32950 4859 33258 4868
rect 33796 4758 33824 8774
rect 33888 8430 33916 8978
rect 34060 8968 34112 8974
rect 34060 8910 34112 8916
rect 34072 8634 34100 8910
rect 34060 8628 34112 8634
rect 34060 8570 34112 8576
rect 33876 8424 33928 8430
rect 33876 8366 33928 8372
rect 33784 4752 33836 4758
rect 33784 4694 33836 4700
rect 32950 3836 33258 3845
rect 32950 3834 32956 3836
rect 33012 3834 33036 3836
rect 33092 3834 33116 3836
rect 33172 3834 33196 3836
rect 33252 3834 33258 3836
rect 33012 3782 33014 3834
rect 33194 3782 33196 3834
rect 32950 3780 32956 3782
rect 33012 3780 33036 3782
rect 33092 3780 33116 3782
rect 33172 3780 33196 3782
rect 33252 3780 33258 3782
rect 32950 3771 33258 3780
rect 29644 3120 29696 3126
rect 29644 3062 29696 3068
rect 34164 2774 34192 13262
rect 34256 10985 34284 14214
rect 34242 10976 34298 10985
rect 34242 10911 34298 10920
rect 34244 10804 34296 10810
rect 34244 10746 34296 10752
rect 34256 7410 34284 10746
rect 34348 10169 34376 19450
rect 34440 18465 34468 20470
rect 34532 20466 34560 20567
rect 34612 20528 34664 20534
rect 34612 20470 34664 20476
rect 34520 20460 34572 20466
rect 34520 20402 34572 20408
rect 34532 19310 34560 20402
rect 34624 19378 34652 20470
rect 34704 20052 34756 20058
rect 34704 19994 34756 20000
rect 34612 19372 34664 19378
rect 34612 19314 34664 19320
rect 34520 19304 34572 19310
rect 34520 19246 34572 19252
rect 34426 18456 34482 18465
rect 34426 18391 34482 18400
rect 34440 17270 34468 18391
rect 34612 17876 34664 17882
rect 34612 17818 34664 17824
rect 34520 17536 34572 17542
rect 34520 17478 34572 17484
rect 34428 17264 34480 17270
rect 34428 17206 34480 17212
rect 34440 16522 34468 17206
rect 34428 16516 34480 16522
rect 34428 16458 34480 16464
rect 34440 15434 34468 16458
rect 34428 15428 34480 15434
rect 34428 15370 34480 15376
rect 34440 13938 34468 15370
rect 34532 15366 34560 17478
rect 34624 17270 34652 17818
rect 34612 17264 34664 17270
rect 34612 17206 34664 17212
rect 34624 16590 34652 17206
rect 34612 16584 34664 16590
rect 34612 16526 34664 16532
rect 34520 15360 34572 15366
rect 34520 15302 34572 15308
rect 34520 14340 34572 14346
rect 34520 14282 34572 14288
rect 34428 13932 34480 13938
rect 34428 13874 34480 13880
rect 34532 12102 34560 14282
rect 34624 12918 34652 16526
rect 34716 13870 34744 19994
rect 34900 18834 34928 21626
rect 34888 18828 34940 18834
rect 34888 18770 34940 18776
rect 34992 18306 35020 22066
rect 35084 19786 35112 22918
rect 35176 21010 35204 22918
rect 35268 22574 35296 23734
rect 35636 23594 35664 24006
rect 35624 23588 35676 23594
rect 35624 23530 35676 23536
rect 35348 23520 35400 23526
rect 35348 23462 35400 23468
rect 35440 23520 35492 23526
rect 35440 23462 35492 23468
rect 35360 23050 35388 23462
rect 35348 23044 35400 23050
rect 35348 22986 35400 22992
rect 35452 22817 35480 23462
rect 36174 23216 36230 23225
rect 36174 23151 36230 23160
rect 35806 23080 35862 23089
rect 35806 23015 35808 23024
rect 35860 23015 35862 23024
rect 35808 22986 35860 22992
rect 35438 22808 35494 22817
rect 35438 22743 35494 22752
rect 35256 22568 35308 22574
rect 35256 22510 35308 22516
rect 35256 22432 35308 22438
rect 35254 22400 35256 22409
rect 35308 22400 35310 22409
rect 35254 22335 35310 22344
rect 35164 21004 35216 21010
rect 35164 20946 35216 20952
rect 35176 20398 35204 20946
rect 35164 20392 35216 20398
rect 35164 20334 35216 20340
rect 35268 19922 35296 22335
rect 35820 22234 35848 22986
rect 36084 22636 36136 22642
rect 36084 22578 36136 22584
rect 35808 22228 35860 22234
rect 35808 22170 35860 22176
rect 35900 22092 35952 22098
rect 35900 22034 35952 22040
rect 35808 21888 35860 21894
rect 35808 21830 35860 21836
rect 35624 21344 35676 21350
rect 35624 21286 35676 21292
rect 35348 20460 35400 20466
rect 35348 20402 35400 20408
rect 35256 19916 35308 19922
rect 35256 19858 35308 19864
rect 35360 19802 35388 20402
rect 35440 19916 35492 19922
rect 35440 19858 35492 19864
rect 35072 19780 35124 19786
rect 35072 19722 35124 19728
rect 35176 19774 35388 19802
rect 35176 19378 35204 19774
rect 35256 19440 35308 19446
rect 35256 19382 35308 19388
rect 35072 19372 35124 19378
rect 35072 19314 35124 19320
rect 35164 19372 35216 19378
rect 35164 19314 35216 19320
rect 34900 18278 35020 18306
rect 34900 17814 34928 18278
rect 34888 17808 34940 17814
rect 35084 17785 35112 19314
rect 34888 17750 34940 17756
rect 35070 17776 35126 17785
rect 35070 17711 35126 17720
rect 35072 17672 35124 17678
rect 35072 17614 35124 17620
rect 35084 17338 35112 17614
rect 35072 17332 35124 17338
rect 35072 17274 35124 17280
rect 35176 17218 35204 19314
rect 35268 18834 35296 19382
rect 35256 18828 35308 18834
rect 35256 18770 35308 18776
rect 35348 18624 35400 18630
rect 35348 18566 35400 18572
rect 35254 18456 35310 18465
rect 35254 18391 35310 18400
rect 35268 18358 35296 18391
rect 35256 18352 35308 18358
rect 35256 18294 35308 18300
rect 35360 18222 35388 18566
rect 35348 18216 35400 18222
rect 35348 18158 35400 18164
rect 35084 17190 35204 17218
rect 34796 17128 34848 17134
rect 34796 17070 34848 17076
rect 34888 17128 34940 17134
rect 34888 17070 34940 17076
rect 34808 16794 34836 17070
rect 34796 16788 34848 16794
rect 34796 16730 34848 16736
rect 34900 16046 34928 17070
rect 34888 16040 34940 16046
rect 34888 15982 34940 15988
rect 34796 15632 34848 15638
rect 34796 15574 34848 15580
rect 34808 14074 34836 15574
rect 34900 15502 34928 15982
rect 34888 15496 34940 15502
rect 34888 15438 34940 15444
rect 34900 14482 34928 15438
rect 35084 15042 35112 17190
rect 35164 15564 35216 15570
rect 35164 15506 35216 15512
rect 35176 15162 35204 15506
rect 35256 15360 35308 15366
rect 35256 15302 35308 15308
rect 35164 15156 35216 15162
rect 35164 15098 35216 15104
rect 35084 15014 35204 15042
rect 34980 14952 35032 14958
rect 34980 14894 35032 14900
rect 34888 14476 34940 14482
rect 34888 14418 34940 14424
rect 34886 14240 34942 14249
rect 34886 14175 34942 14184
rect 34796 14068 34848 14074
rect 34796 14010 34848 14016
rect 34704 13864 34756 13870
rect 34704 13806 34756 13812
rect 34796 13728 34848 13734
rect 34796 13670 34848 13676
rect 34702 13288 34758 13297
rect 34702 13223 34704 13232
rect 34756 13223 34758 13232
rect 34704 13194 34756 13200
rect 34612 12912 34664 12918
rect 34612 12854 34664 12860
rect 34520 12096 34572 12102
rect 34520 12038 34572 12044
rect 34624 11830 34652 12854
rect 34612 11824 34664 11830
rect 34612 11766 34664 11772
rect 34428 11144 34480 11150
rect 34428 11086 34480 11092
rect 34334 10160 34390 10169
rect 34334 10095 34390 10104
rect 34336 9988 34388 9994
rect 34336 9930 34388 9936
rect 34348 8498 34376 9930
rect 34440 9042 34468 11086
rect 34520 9920 34572 9926
rect 34520 9862 34572 9868
rect 34428 9036 34480 9042
rect 34428 8978 34480 8984
rect 34532 8566 34560 9862
rect 34520 8560 34572 8566
rect 34520 8502 34572 8508
rect 34336 8492 34388 8498
rect 34336 8434 34388 8440
rect 34716 8430 34744 13194
rect 34808 12646 34836 13670
rect 34900 12918 34928 14175
rect 34888 12912 34940 12918
rect 34888 12854 34940 12860
rect 34888 12776 34940 12782
rect 34888 12718 34940 12724
rect 34796 12640 34848 12646
rect 34796 12582 34848 12588
rect 34900 12306 34928 12718
rect 34888 12300 34940 12306
rect 34888 12242 34940 12248
rect 34900 11762 34928 12242
rect 34888 11756 34940 11762
rect 34888 11698 34940 11704
rect 34796 11688 34848 11694
rect 34796 11630 34848 11636
rect 34808 11150 34836 11630
rect 34796 11144 34848 11150
rect 34796 11086 34848 11092
rect 34888 10804 34940 10810
rect 34888 10746 34940 10752
rect 34900 10266 34928 10746
rect 34888 10260 34940 10266
rect 34888 10202 34940 10208
rect 34992 9110 35020 14894
rect 35072 13728 35124 13734
rect 35072 13670 35124 13676
rect 35084 10810 35112 13670
rect 35176 13394 35204 15014
rect 35268 14346 35296 15302
rect 35452 14770 35480 19858
rect 35636 16726 35664 21286
rect 35820 20602 35848 21830
rect 35912 21010 35940 22034
rect 36096 21865 36124 22578
rect 36188 22574 36216 23151
rect 36280 22953 36308 24686
rect 36556 24274 36584 24754
rect 36544 24268 36596 24274
rect 36544 24210 36596 24216
rect 36360 24200 36412 24206
rect 36360 24142 36412 24148
rect 36266 22944 36322 22953
rect 36266 22879 36322 22888
rect 36176 22568 36228 22574
rect 36174 22536 36176 22545
rect 36228 22536 36230 22545
rect 36174 22471 36230 22480
rect 36174 22264 36230 22273
rect 36174 22199 36230 22208
rect 36082 21856 36138 21865
rect 36082 21791 36138 21800
rect 36188 21486 36216 22199
rect 36280 21622 36308 22879
rect 36372 22778 36400 24142
rect 36544 23656 36596 23662
rect 36542 23624 36544 23633
rect 36596 23624 36598 23633
rect 36542 23559 36598 23568
rect 36648 23497 36676 26302
rect 37002 26200 37058 27000
rect 37646 26200 37702 27000
rect 38290 26330 38346 27000
rect 38290 26302 38516 26330
rect 38290 26200 38346 26302
rect 36728 23656 36780 23662
rect 36728 23598 36780 23604
rect 36634 23488 36690 23497
rect 36634 23423 36690 23432
rect 36740 23050 36768 23598
rect 36728 23044 36780 23050
rect 36728 22986 36780 22992
rect 36360 22772 36412 22778
rect 36360 22714 36412 22720
rect 36450 22672 36506 22681
rect 36450 22607 36506 22616
rect 36464 22574 36492 22607
rect 36452 22568 36504 22574
rect 36452 22510 36504 22516
rect 37016 22438 37044 26200
rect 37556 24404 37608 24410
rect 37556 24346 37608 24352
rect 37568 24274 37596 24346
rect 37556 24268 37608 24274
rect 37556 24210 37608 24216
rect 37464 24064 37516 24070
rect 37464 24006 37516 24012
rect 37476 23866 37504 24006
rect 37464 23860 37516 23866
rect 37464 23802 37516 23808
rect 37372 23724 37424 23730
rect 37372 23666 37424 23672
rect 37094 23624 37150 23633
rect 37094 23559 37150 23568
rect 37004 22432 37056 22438
rect 37004 22374 37056 22380
rect 36544 21888 36596 21894
rect 36544 21830 36596 21836
rect 36268 21616 36320 21622
rect 36268 21558 36320 21564
rect 36176 21480 36228 21486
rect 36176 21422 36228 21428
rect 36556 21418 36584 21830
rect 37108 21554 37136 23559
rect 37280 23112 37332 23118
rect 37280 23054 37332 23060
rect 37188 23044 37240 23050
rect 37188 22986 37240 22992
rect 37200 22778 37228 22986
rect 37188 22772 37240 22778
rect 37188 22714 37240 22720
rect 37292 22574 37320 23054
rect 37280 22568 37332 22574
rect 37280 22510 37332 22516
rect 37292 22030 37320 22510
rect 37280 22024 37332 22030
rect 37280 21966 37332 21972
rect 37292 21554 37320 21966
rect 37096 21548 37148 21554
rect 37096 21490 37148 21496
rect 37280 21548 37332 21554
rect 37280 21490 37332 21496
rect 36912 21480 36964 21486
rect 36912 21422 36964 21428
rect 36544 21412 36596 21418
rect 36544 21354 36596 21360
rect 36176 21344 36228 21350
rect 36176 21286 36228 21292
rect 35900 21004 35952 21010
rect 35900 20946 35952 20952
rect 35808 20596 35860 20602
rect 35808 20538 35860 20544
rect 35912 20534 35940 20946
rect 35900 20528 35952 20534
rect 35900 20470 35952 20476
rect 36084 20460 36136 20466
rect 36084 20402 36136 20408
rect 35900 19712 35952 19718
rect 35900 19654 35952 19660
rect 35992 19712 36044 19718
rect 35992 19654 36044 19660
rect 35714 19544 35770 19553
rect 35714 19479 35770 19488
rect 35728 18358 35756 19479
rect 35912 19378 35940 19654
rect 35900 19372 35952 19378
rect 35900 19314 35952 19320
rect 36004 18970 36032 19654
rect 35992 18964 36044 18970
rect 35992 18906 36044 18912
rect 35716 18352 35768 18358
rect 35716 18294 35768 18300
rect 35728 17746 35756 18294
rect 35716 17740 35768 17746
rect 35716 17682 35768 17688
rect 35624 16720 35676 16726
rect 35624 16662 35676 16668
rect 35728 16658 35756 17682
rect 35992 17604 36044 17610
rect 35992 17546 36044 17552
rect 35716 16652 35768 16658
rect 35716 16594 35768 16600
rect 36004 16590 36032 17546
rect 36096 17066 36124 20402
rect 36188 19446 36216 21286
rect 36268 21140 36320 21146
rect 36268 21082 36320 21088
rect 36176 19440 36228 19446
rect 36176 19382 36228 19388
rect 36176 19236 36228 19242
rect 36176 19178 36228 19184
rect 36188 17746 36216 19178
rect 36280 18426 36308 21082
rect 36728 20052 36780 20058
rect 36728 19994 36780 20000
rect 36544 19712 36596 19718
rect 36544 19654 36596 19660
rect 36556 19514 36584 19654
rect 36544 19508 36596 19514
rect 36544 19450 36596 19456
rect 36636 19440 36688 19446
rect 36636 19382 36688 19388
rect 36544 18692 36596 18698
rect 36544 18634 36596 18640
rect 36556 18465 36584 18634
rect 36542 18456 36598 18465
rect 36268 18420 36320 18426
rect 36542 18391 36598 18400
rect 36268 18362 36320 18368
rect 36360 18216 36412 18222
rect 36360 18158 36412 18164
rect 36176 17740 36228 17746
rect 36176 17682 36228 17688
rect 36176 17128 36228 17134
rect 36176 17070 36228 17076
rect 36084 17060 36136 17066
rect 36084 17002 36136 17008
rect 35992 16584 36044 16590
rect 35992 16526 36044 16532
rect 35808 15904 35860 15910
rect 35808 15846 35860 15852
rect 35900 15904 35952 15910
rect 35900 15846 35952 15852
rect 35360 14742 35480 14770
rect 35716 14816 35768 14822
rect 35716 14758 35768 14764
rect 35360 14618 35388 14742
rect 35348 14612 35400 14618
rect 35348 14554 35400 14560
rect 35256 14340 35308 14346
rect 35256 14282 35308 14288
rect 35164 13388 35216 13394
rect 35164 13330 35216 13336
rect 35452 12102 35480 14742
rect 35532 13728 35584 13734
rect 35532 13670 35584 13676
rect 35544 13394 35572 13670
rect 35532 13388 35584 13394
rect 35532 13330 35584 13336
rect 35728 12986 35756 14758
rect 35820 14618 35848 15846
rect 35912 15366 35940 15846
rect 35900 15360 35952 15366
rect 35900 15302 35952 15308
rect 35808 14612 35860 14618
rect 35808 14554 35860 14560
rect 35992 13864 36044 13870
rect 35992 13806 36044 13812
rect 35808 13320 35860 13326
rect 35808 13262 35860 13268
rect 35716 12980 35768 12986
rect 35716 12922 35768 12928
rect 35820 12306 35848 13262
rect 35808 12300 35860 12306
rect 35808 12242 35860 12248
rect 35440 12096 35492 12102
rect 35440 12038 35492 12044
rect 35808 12096 35860 12102
rect 35808 12038 35860 12044
rect 35348 11076 35400 11082
rect 35348 11018 35400 11024
rect 35072 10804 35124 10810
rect 35072 10746 35124 10752
rect 35084 9994 35112 10746
rect 35360 10742 35388 11018
rect 35532 11008 35584 11014
rect 35532 10950 35584 10956
rect 35348 10736 35400 10742
rect 35348 10678 35400 10684
rect 35072 9988 35124 9994
rect 35360 9976 35388 10678
rect 35544 10470 35572 10950
rect 35820 10674 35848 12038
rect 36004 11558 36032 13806
rect 36188 11801 36216 17070
rect 36268 16448 36320 16454
rect 36268 16390 36320 16396
rect 36280 14006 36308 16390
rect 36372 15706 36400 18158
rect 36452 18148 36504 18154
rect 36452 18090 36504 18096
rect 36464 17338 36492 18090
rect 36556 17610 36584 18391
rect 36544 17604 36596 17610
rect 36544 17546 36596 17552
rect 36452 17332 36504 17338
rect 36452 17274 36504 17280
rect 36452 16108 36504 16114
rect 36556 16096 36584 17546
rect 36504 16068 36584 16096
rect 36452 16050 36504 16056
rect 36360 15700 36412 15706
rect 36360 15642 36412 15648
rect 36464 15434 36492 16050
rect 36452 15428 36504 15434
rect 36504 15388 36584 15416
rect 36452 15370 36504 15376
rect 36452 14952 36504 14958
rect 36452 14894 36504 14900
rect 36268 14000 36320 14006
rect 36268 13942 36320 13948
rect 36360 13184 36412 13190
rect 36360 13126 36412 13132
rect 36268 12844 36320 12850
rect 36268 12786 36320 12792
rect 36174 11792 36230 11801
rect 36174 11727 36230 11736
rect 35992 11552 36044 11558
rect 35992 11494 36044 11500
rect 36084 11552 36136 11558
rect 36084 11494 36136 11500
rect 36096 11218 36124 11494
rect 36188 11393 36216 11727
rect 36174 11384 36230 11393
rect 36174 11319 36230 11328
rect 36084 11212 36136 11218
rect 36084 11154 36136 11160
rect 35808 10668 35860 10674
rect 35808 10610 35860 10616
rect 35532 10464 35584 10470
rect 35532 10406 35584 10412
rect 35440 9988 35492 9994
rect 35360 9948 35440 9976
rect 35072 9930 35124 9936
rect 35440 9930 35492 9936
rect 35624 9988 35676 9994
rect 35624 9930 35676 9936
rect 35084 9466 35112 9930
rect 35636 9654 35664 9930
rect 35624 9648 35676 9654
rect 35624 9590 35676 9596
rect 35084 9450 35204 9466
rect 35084 9444 35216 9450
rect 35084 9438 35164 9444
rect 35164 9386 35216 9392
rect 35532 9376 35584 9382
rect 35532 9318 35584 9324
rect 34980 9104 35032 9110
rect 34980 9046 35032 9052
rect 35544 9042 35572 9318
rect 35624 9104 35676 9110
rect 35624 9046 35676 9052
rect 35532 9036 35584 9042
rect 35532 8978 35584 8984
rect 35636 8838 35664 9046
rect 34888 8832 34940 8838
rect 34888 8774 34940 8780
rect 35256 8832 35308 8838
rect 35256 8774 35308 8780
rect 35624 8832 35676 8838
rect 35624 8774 35676 8780
rect 34900 8566 34928 8774
rect 34888 8560 34940 8566
rect 34888 8502 34940 8508
rect 34704 8424 34756 8430
rect 34704 8366 34756 8372
rect 35268 8090 35296 8774
rect 35532 8424 35584 8430
rect 35532 8366 35584 8372
rect 35256 8084 35308 8090
rect 35256 8026 35308 8032
rect 34244 7404 34296 7410
rect 34244 7346 34296 7352
rect 35544 7342 35572 8366
rect 35820 7954 35848 10610
rect 36280 10606 36308 12786
rect 36372 12782 36400 13126
rect 36360 12776 36412 12782
rect 36360 12718 36412 12724
rect 36464 12102 36492 14894
rect 36556 14346 36584 15388
rect 36648 14890 36676 19382
rect 36740 15094 36768 19994
rect 36924 17898 36952 21422
rect 37292 21010 37320 21490
rect 37384 21146 37412 23666
rect 37568 22098 37596 24210
rect 37660 22098 37688 26200
rect 37922 24848 37978 24857
rect 37922 24783 37978 24792
rect 37936 24274 37964 24783
rect 37924 24268 37976 24274
rect 37924 24210 37976 24216
rect 38384 24268 38436 24274
rect 38384 24210 38436 24216
rect 37740 24132 37792 24138
rect 37740 24074 37792 24080
rect 37752 22710 37780 24074
rect 37950 23964 38258 23973
rect 37950 23962 37956 23964
rect 38012 23962 38036 23964
rect 38092 23962 38116 23964
rect 38172 23962 38196 23964
rect 38252 23962 38258 23964
rect 38012 23910 38014 23962
rect 38194 23910 38196 23962
rect 37950 23908 37956 23910
rect 38012 23908 38036 23910
rect 38092 23908 38116 23910
rect 38172 23908 38196 23910
rect 38252 23908 38258 23910
rect 37950 23899 38258 23908
rect 37832 23724 37884 23730
rect 37832 23666 37884 23672
rect 37740 22704 37792 22710
rect 37740 22646 37792 22652
rect 37740 22568 37792 22574
rect 37740 22510 37792 22516
rect 37752 22137 37780 22510
rect 37738 22128 37794 22137
rect 37556 22092 37608 22098
rect 37556 22034 37608 22040
rect 37648 22092 37700 22098
rect 37738 22063 37794 22072
rect 37648 22034 37700 22040
rect 37462 21856 37518 21865
rect 37462 21791 37518 21800
rect 37476 21321 37504 21791
rect 37752 21690 37780 22063
rect 37740 21684 37792 21690
rect 37740 21626 37792 21632
rect 37462 21312 37518 21321
rect 37462 21247 37518 21256
rect 37372 21140 37424 21146
rect 37372 21082 37424 21088
rect 37280 21004 37332 21010
rect 37280 20946 37332 20952
rect 37280 19916 37332 19922
rect 37280 19858 37332 19864
rect 37188 19372 37240 19378
rect 37188 19314 37240 19320
rect 37004 19168 37056 19174
rect 37004 19110 37056 19116
rect 37016 18970 37044 19110
rect 37004 18964 37056 18970
rect 37004 18906 37056 18912
rect 36832 17882 36952 17898
rect 37200 17882 37228 19314
rect 37292 18290 37320 19858
rect 37372 19848 37424 19854
rect 37372 19790 37424 19796
rect 37384 19689 37412 19790
rect 37370 19680 37426 19689
rect 37370 19615 37426 19624
rect 37476 18766 37504 21247
rect 37740 21004 37792 21010
rect 37740 20946 37792 20952
rect 37752 20466 37780 20946
rect 37556 20460 37608 20466
rect 37556 20402 37608 20408
rect 37740 20460 37792 20466
rect 37740 20402 37792 20408
rect 37464 18760 37516 18766
rect 37462 18728 37464 18737
rect 37516 18728 37518 18737
rect 37462 18663 37518 18672
rect 37568 18426 37596 20402
rect 37648 20392 37700 20398
rect 37648 20334 37700 20340
rect 37660 18698 37688 20334
rect 37752 19553 37780 20402
rect 37844 20058 37872 23666
rect 38292 23656 38344 23662
rect 38292 23598 38344 23604
rect 37950 22876 38258 22885
rect 37950 22874 37956 22876
rect 38012 22874 38036 22876
rect 38092 22874 38116 22876
rect 38172 22874 38196 22876
rect 38252 22874 38258 22876
rect 38012 22822 38014 22874
rect 38194 22822 38196 22874
rect 37950 22820 37956 22822
rect 38012 22820 38036 22822
rect 38092 22820 38116 22822
rect 38172 22820 38196 22822
rect 38252 22820 38258 22822
rect 37950 22811 38258 22820
rect 37950 21788 38258 21797
rect 37950 21786 37956 21788
rect 38012 21786 38036 21788
rect 38092 21786 38116 21788
rect 38172 21786 38196 21788
rect 38252 21786 38258 21788
rect 38012 21734 38014 21786
rect 38194 21734 38196 21786
rect 37950 21732 37956 21734
rect 38012 21732 38036 21734
rect 38092 21732 38116 21734
rect 38172 21732 38196 21734
rect 38252 21732 38258 21734
rect 37950 21723 38258 21732
rect 37924 21344 37976 21350
rect 37924 21286 37976 21292
rect 37936 20874 37964 21286
rect 37924 20868 37976 20874
rect 37924 20810 37976 20816
rect 38304 20806 38332 23598
rect 38396 23361 38424 24210
rect 38382 23352 38438 23361
rect 38382 23287 38438 23296
rect 38488 22001 38516 26302
rect 38934 26200 38990 27000
rect 39578 26200 39634 27000
rect 40222 26200 40278 27000
rect 42154 26200 42210 27000
rect 42798 26200 42854 27000
rect 43350 26344 43406 26353
rect 43350 26279 43406 26288
rect 38948 24818 38976 26200
rect 39212 24948 39264 24954
rect 39212 24890 39264 24896
rect 38936 24812 38988 24818
rect 38936 24754 38988 24760
rect 38658 24712 38714 24721
rect 38658 24647 38714 24656
rect 38568 24404 38620 24410
rect 38568 24346 38620 24352
rect 38580 23610 38608 24346
rect 38672 24274 38700 24647
rect 39224 24410 39252 24890
rect 39212 24404 39264 24410
rect 39212 24346 39264 24352
rect 38660 24268 38712 24274
rect 38660 24210 38712 24216
rect 39224 24206 39252 24346
rect 39120 24200 39172 24206
rect 39120 24142 39172 24148
rect 39212 24200 39264 24206
rect 39212 24142 39264 24148
rect 38752 23724 38804 23730
rect 38752 23666 38804 23672
rect 38580 23582 38700 23610
rect 38568 23520 38620 23526
rect 38568 23462 38620 23468
rect 38580 23322 38608 23462
rect 38672 23322 38700 23582
rect 38568 23316 38620 23322
rect 38568 23258 38620 23264
rect 38660 23316 38712 23322
rect 38660 23258 38712 23264
rect 38568 22976 38620 22982
rect 38568 22918 38620 22924
rect 38580 22166 38608 22918
rect 38568 22160 38620 22166
rect 38568 22102 38620 22108
rect 38474 21992 38530 22001
rect 38474 21927 38530 21936
rect 38764 21146 38792 23666
rect 38844 23248 38896 23254
rect 38844 23190 38896 23196
rect 38856 23050 38884 23190
rect 38844 23044 38896 23050
rect 38844 22986 38896 22992
rect 38856 22642 38884 22986
rect 39026 22808 39082 22817
rect 39026 22743 39082 22752
rect 38844 22636 38896 22642
rect 38844 22578 38896 22584
rect 38856 22234 38884 22578
rect 39040 22506 39068 22743
rect 39132 22506 39160 24142
rect 39592 23050 39620 26200
rect 39946 24848 40002 24857
rect 39946 24783 40002 24792
rect 39960 24342 39988 24783
rect 40040 24608 40092 24614
rect 40040 24550 40092 24556
rect 40052 24410 40080 24550
rect 40040 24404 40092 24410
rect 40040 24346 40092 24352
rect 39672 24336 39724 24342
rect 39672 24278 39724 24284
rect 39948 24336 40000 24342
rect 39948 24278 40000 24284
rect 39580 23044 39632 23050
rect 39580 22986 39632 22992
rect 39684 22778 39712 24278
rect 39856 24064 39908 24070
rect 39856 24006 39908 24012
rect 39868 23866 39896 24006
rect 39856 23860 39908 23866
rect 39856 23802 39908 23808
rect 39960 23662 39988 24278
rect 40040 23792 40092 23798
rect 40040 23734 40092 23740
rect 39948 23656 40000 23662
rect 39948 23598 40000 23604
rect 39764 23588 39816 23594
rect 39764 23530 39816 23536
rect 39672 22772 39724 22778
rect 39672 22714 39724 22720
rect 39028 22500 39080 22506
rect 39028 22442 39080 22448
rect 39120 22500 39172 22506
rect 39120 22442 39172 22448
rect 38844 22228 38896 22234
rect 38844 22170 38896 22176
rect 38856 22030 38884 22170
rect 38844 22024 38896 22030
rect 38844 21966 38896 21972
rect 39028 22024 39080 22030
rect 39028 21966 39080 21972
rect 39040 21622 39068 21966
rect 39776 21894 39804 23530
rect 40052 23322 40080 23734
rect 40236 23322 40264 26200
rect 41788 24812 41840 24818
rect 41788 24754 41840 24760
rect 40684 24744 40736 24750
rect 40684 24686 40736 24692
rect 40696 24410 40724 24686
rect 40684 24404 40736 24410
rect 40684 24346 40736 24352
rect 40960 24336 41012 24342
rect 40960 24278 41012 24284
rect 41234 24304 41290 24313
rect 40972 24138 41000 24278
rect 41234 24239 41290 24248
rect 40960 24132 41012 24138
rect 40960 24074 41012 24080
rect 41144 24132 41196 24138
rect 41144 24074 41196 24080
rect 40776 24064 40828 24070
rect 40776 24006 40828 24012
rect 40788 23633 40816 24006
rect 40774 23624 40830 23633
rect 40774 23559 40830 23568
rect 40500 23520 40552 23526
rect 40500 23462 40552 23468
rect 40040 23316 40092 23322
rect 40040 23258 40092 23264
rect 40224 23316 40276 23322
rect 40224 23258 40276 23264
rect 40316 23044 40368 23050
rect 40316 22986 40368 22992
rect 40224 22976 40276 22982
rect 40224 22918 40276 22924
rect 40132 22772 40184 22778
rect 40132 22714 40184 22720
rect 40040 22636 40092 22642
rect 40040 22578 40092 22584
rect 40052 22234 40080 22578
rect 40040 22228 40092 22234
rect 40040 22170 40092 22176
rect 39120 21888 39172 21894
rect 39120 21830 39172 21836
rect 39764 21888 39816 21894
rect 39764 21830 39816 21836
rect 39028 21616 39080 21622
rect 39028 21558 39080 21564
rect 39132 21486 39160 21830
rect 39488 21616 39540 21622
rect 39488 21558 39540 21564
rect 39120 21480 39172 21486
rect 39120 21422 39172 21428
rect 39212 21344 39264 21350
rect 39212 21286 39264 21292
rect 38752 21140 38804 21146
rect 38752 21082 38804 21088
rect 39224 21010 39252 21286
rect 39212 21004 39264 21010
rect 39212 20946 39264 20952
rect 39500 20942 39528 21558
rect 39672 21548 39724 21554
rect 39672 21490 39724 21496
rect 39684 21350 39712 21490
rect 39672 21344 39724 21350
rect 39670 21312 39672 21321
rect 39724 21312 39726 21321
rect 39670 21247 39726 21256
rect 39776 20942 39804 21830
rect 40144 21690 40172 22714
rect 40132 21684 40184 21690
rect 40132 21626 40184 21632
rect 40236 21162 40264 22918
rect 40328 22710 40356 22986
rect 40316 22704 40368 22710
rect 40316 22646 40368 22652
rect 40408 21480 40460 21486
rect 40408 21422 40460 21428
rect 39960 21134 40264 21162
rect 40316 21140 40368 21146
rect 39488 20936 39540 20942
rect 39488 20878 39540 20884
rect 39764 20936 39816 20942
rect 39764 20878 39816 20884
rect 38292 20800 38344 20806
rect 38292 20742 38344 20748
rect 37950 20700 38258 20709
rect 37950 20698 37956 20700
rect 38012 20698 38036 20700
rect 38092 20698 38116 20700
rect 38172 20698 38196 20700
rect 38252 20698 38258 20700
rect 38012 20646 38014 20698
rect 38194 20646 38196 20698
rect 37950 20644 37956 20646
rect 38012 20644 38036 20646
rect 38092 20644 38116 20646
rect 38172 20644 38196 20646
rect 38252 20644 38258 20646
rect 37950 20635 38258 20644
rect 38304 20534 38332 20742
rect 39500 20534 39528 20878
rect 39960 20874 39988 21134
rect 40316 21082 40368 21088
rect 39948 20868 40000 20874
rect 39948 20810 40000 20816
rect 37924 20528 37976 20534
rect 37924 20470 37976 20476
rect 38292 20528 38344 20534
rect 38292 20470 38344 20476
rect 39488 20528 39540 20534
rect 39488 20470 39540 20476
rect 37832 20052 37884 20058
rect 37832 19994 37884 20000
rect 37936 19922 37964 20470
rect 38660 20256 38712 20262
rect 38660 20198 38712 20204
rect 37924 19916 37976 19922
rect 37924 19858 37976 19864
rect 38384 19916 38436 19922
rect 38384 19858 38436 19864
rect 38568 19916 38620 19922
rect 38568 19858 38620 19864
rect 38396 19689 38424 19858
rect 38382 19680 38438 19689
rect 37950 19612 38258 19621
rect 38382 19615 38438 19624
rect 37950 19610 37956 19612
rect 38012 19610 38036 19612
rect 38092 19610 38116 19612
rect 38172 19610 38196 19612
rect 38252 19610 38258 19612
rect 38012 19558 38014 19610
rect 38194 19558 38196 19610
rect 37950 19556 37956 19558
rect 38012 19556 38036 19558
rect 38092 19556 38116 19558
rect 38172 19556 38196 19558
rect 38252 19556 38258 19558
rect 37738 19544 37794 19553
rect 37950 19547 38258 19556
rect 37738 19479 37794 19488
rect 37752 19378 37780 19479
rect 37740 19372 37792 19378
rect 37740 19314 37792 19320
rect 37832 19304 37884 19310
rect 37832 19246 37884 19252
rect 38382 19272 38438 19281
rect 37648 18692 37700 18698
rect 37648 18634 37700 18640
rect 37556 18420 37608 18426
rect 37556 18362 37608 18368
rect 37280 18284 37332 18290
rect 37280 18226 37332 18232
rect 36820 17876 36952 17882
rect 36872 17870 36952 17876
rect 36820 17818 36872 17824
rect 36820 16652 36872 16658
rect 36820 16594 36872 16600
rect 36728 15088 36780 15094
rect 36728 15030 36780 15036
rect 36636 14884 36688 14890
rect 36636 14826 36688 14832
rect 36832 14618 36860 16594
rect 36924 15978 36952 17870
rect 37188 17876 37240 17882
rect 37188 17818 37240 17824
rect 37292 17814 37320 18226
rect 37556 18216 37608 18222
rect 37556 18158 37608 18164
rect 37280 17808 37332 17814
rect 37280 17750 37332 17756
rect 37372 17672 37424 17678
rect 37372 17614 37424 17620
rect 37188 16652 37240 16658
rect 37188 16594 37240 16600
rect 36912 15972 36964 15978
rect 36912 15914 36964 15920
rect 37096 15496 37148 15502
rect 37096 15438 37148 15444
rect 37108 14958 37136 15438
rect 37200 15026 37228 16594
rect 37384 16046 37412 17614
rect 37568 17134 37596 18158
rect 37556 17128 37608 17134
rect 37556 17070 37608 17076
rect 37648 17128 37700 17134
rect 37648 17070 37700 17076
rect 37556 16992 37608 16998
rect 37556 16934 37608 16940
rect 37568 16250 37596 16934
rect 37556 16244 37608 16250
rect 37556 16186 37608 16192
rect 37372 16040 37424 16046
rect 37372 15982 37424 15988
rect 37384 15706 37412 15982
rect 37660 15706 37688 17070
rect 37740 17060 37792 17066
rect 37740 17002 37792 17008
rect 37752 16590 37780 17002
rect 37740 16584 37792 16590
rect 37740 16526 37792 16532
rect 37752 16046 37780 16526
rect 37844 16454 37872 19246
rect 38382 19207 38438 19216
rect 38292 18828 38344 18834
rect 38292 18770 38344 18776
rect 37950 18524 38258 18533
rect 37950 18522 37956 18524
rect 38012 18522 38036 18524
rect 38092 18522 38116 18524
rect 38172 18522 38196 18524
rect 38252 18522 38258 18524
rect 38012 18470 38014 18522
rect 38194 18470 38196 18522
rect 37950 18468 37956 18470
rect 38012 18468 38036 18470
rect 38092 18468 38116 18470
rect 38172 18468 38196 18470
rect 38252 18468 38258 18470
rect 37950 18459 38258 18468
rect 37950 17436 38258 17445
rect 37950 17434 37956 17436
rect 38012 17434 38036 17436
rect 38092 17434 38116 17436
rect 38172 17434 38196 17436
rect 38252 17434 38258 17436
rect 38012 17382 38014 17434
rect 38194 17382 38196 17434
rect 37950 17380 37956 17382
rect 38012 17380 38036 17382
rect 38092 17380 38116 17382
rect 38172 17380 38196 17382
rect 38252 17380 38258 17382
rect 37950 17371 38258 17380
rect 37832 16448 37884 16454
rect 37832 16390 37884 16396
rect 37844 16182 37872 16390
rect 37950 16348 38258 16357
rect 37950 16346 37956 16348
rect 38012 16346 38036 16348
rect 38092 16346 38116 16348
rect 38172 16346 38196 16348
rect 38252 16346 38258 16348
rect 38012 16294 38014 16346
rect 38194 16294 38196 16346
rect 37950 16292 37956 16294
rect 38012 16292 38036 16294
rect 38092 16292 38116 16294
rect 38172 16292 38196 16294
rect 38252 16292 38258 16294
rect 37950 16283 38258 16292
rect 37832 16176 37884 16182
rect 37832 16118 37884 16124
rect 37740 16040 37792 16046
rect 37740 15982 37792 15988
rect 37372 15700 37424 15706
rect 37372 15642 37424 15648
rect 37648 15700 37700 15706
rect 37648 15642 37700 15648
rect 37556 15428 37608 15434
rect 37556 15370 37608 15376
rect 37188 15020 37240 15026
rect 37188 14962 37240 14968
rect 37096 14952 37148 14958
rect 37096 14894 37148 14900
rect 36820 14612 36872 14618
rect 36820 14554 36872 14560
rect 36544 14340 36596 14346
rect 36544 14282 36596 14288
rect 36556 13190 36584 14282
rect 36832 13870 36860 14554
rect 37108 14482 37136 14894
rect 37280 14816 37332 14822
rect 37280 14758 37332 14764
rect 37096 14476 37148 14482
rect 37096 14418 37148 14424
rect 36636 13864 36688 13870
rect 36636 13806 36688 13812
rect 36820 13864 36872 13870
rect 36820 13806 36872 13812
rect 36648 13258 36676 13806
rect 36636 13252 36688 13258
rect 36636 13194 36688 13200
rect 36544 13184 36596 13190
rect 36544 13126 36596 13132
rect 36556 12170 36584 13126
rect 36544 12164 36596 12170
rect 36544 12106 36596 12112
rect 36452 12096 36504 12102
rect 36452 12038 36504 12044
rect 36556 11762 36584 12106
rect 36728 12096 36780 12102
rect 36728 12038 36780 12044
rect 36740 11762 36768 12038
rect 37292 11830 37320 14758
rect 37372 13932 37424 13938
rect 37372 13874 37424 13880
rect 37384 13138 37412 13874
rect 37568 13734 37596 15370
rect 37660 15094 37688 15642
rect 37752 15502 37780 15982
rect 38016 15972 38068 15978
rect 38016 15914 38068 15920
rect 37740 15496 37792 15502
rect 37740 15438 37792 15444
rect 38028 15434 38056 15914
rect 38016 15428 38068 15434
rect 38016 15370 38068 15376
rect 37950 15260 38258 15269
rect 37950 15258 37956 15260
rect 38012 15258 38036 15260
rect 38092 15258 38116 15260
rect 38172 15258 38196 15260
rect 38252 15258 38258 15260
rect 38012 15206 38014 15258
rect 38194 15206 38196 15258
rect 37950 15204 37956 15206
rect 38012 15204 38036 15206
rect 38092 15204 38116 15206
rect 38172 15204 38196 15206
rect 38252 15204 38258 15206
rect 37950 15195 38258 15204
rect 37648 15088 37700 15094
rect 37648 15030 37700 15036
rect 37832 15088 37884 15094
rect 37832 15030 37884 15036
rect 37844 14346 37872 15030
rect 38304 14958 38332 18770
rect 38396 18630 38424 19207
rect 38384 18624 38436 18630
rect 38384 18566 38436 18572
rect 38476 18080 38528 18086
rect 38476 18022 38528 18028
rect 38488 17746 38516 18022
rect 38476 17740 38528 17746
rect 38476 17682 38528 17688
rect 38384 17264 38436 17270
rect 38384 17206 38436 17212
rect 38292 14952 38344 14958
rect 38292 14894 38344 14900
rect 38108 14476 38160 14482
rect 38304 14464 38332 14894
rect 38160 14436 38332 14464
rect 38108 14418 38160 14424
rect 37832 14340 37884 14346
rect 37832 14282 37884 14288
rect 37950 14172 38258 14181
rect 37950 14170 37956 14172
rect 38012 14170 38036 14172
rect 38092 14170 38116 14172
rect 38172 14170 38196 14172
rect 38252 14170 38258 14172
rect 38012 14118 38014 14170
rect 38194 14118 38196 14170
rect 37950 14116 37956 14118
rect 38012 14116 38036 14118
rect 38092 14116 38116 14118
rect 38172 14116 38196 14118
rect 38252 14116 38258 14118
rect 37950 14107 38258 14116
rect 37832 13796 37884 13802
rect 37832 13738 37884 13744
rect 37556 13728 37608 13734
rect 37556 13670 37608 13676
rect 37844 13394 37872 13738
rect 38396 13530 38424 17206
rect 38580 15994 38608 19858
rect 38672 19310 38700 20198
rect 39118 20088 39174 20097
rect 39118 20023 39174 20032
rect 39132 19854 39160 20023
rect 39120 19848 39172 19854
rect 39120 19790 39172 19796
rect 39500 19446 39528 20470
rect 39960 20233 39988 20810
rect 40328 20466 40356 21082
rect 40420 20602 40448 21422
rect 40512 21010 40540 23462
rect 40590 23352 40646 23361
rect 40590 23287 40646 23296
rect 40604 23186 40632 23287
rect 40592 23180 40644 23186
rect 40592 23122 40644 23128
rect 41050 22672 41106 22681
rect 41050 22607 41106 22616
rect 41064 22574 41092 22607
rect 40960 22568 41012 22574
rect 40682 22536 40738 22545
rect 40960 22510 41012 22516
rect 41052 22568 41104 22574
rect 41052 22510 41104 22516
rect 40682 22471 40738 22480
rect 40592 21888 40644 21894
rect 40592 21830 40644 21836
rect 40604 21690 40632 21830
rect 40592 21684 40644 21690
rect 40592 21626 40644 21632
rect 40604 21298 40632 21626
rect 40696 21486 40724 22471
rect 40776 22160 40828 22166
rect 40774 22128 40776 22137
rect 40828 22128 40830 22137
rect 40774 22063 40830 22072
rect 40788 21486 40816 22063
rect 40972 21894 41000 22510
rect 41156 22094 41184 24074
rect 41248 23866 41276 24239
rect 41236 23860 41288 23866
rect 41236 23802 41288 23808
rect 41328 23792 41380 23798
rect 41328 23734 41380 23740
rect 41420 23792 41472 23798
rect 41420 23734 41472 23740
rect 41236 23656 41288 23662
rect 41236 23598 41288 23604
rect 41064 22066 41184 22094
rect 40960 21888 41012 21894
rect 40960 21830 41012 21836
rect 40684 21480 40736 21486
rect 40684 21422 40736 21428
rect 40776 21480 40828 21486
rect 40776 21422 40828 21428
rect 40604 21270 40724 21298
rect 40500 21004 40552 21010
rect 40500 20946 40552 20952
rect 40592 21004 40644 21010
rect 40592 20946 40644 20952
rect 40408 20596 40460 20602
rect 40408 20538 40460 20544
rect 40316 20460 40368 20466
rect 40316 20402 40368 20408
rect 40328 20369 40356 20402
rect 40500 20392 40552 20398
rect 40314 20360 40370 20369
rect 40132 20324 40184 20330
rect 40500 20334 40552 20340
rect 40314 20295 40370 20304
rect 40408 20324 40460 20330
rect 40132 20266 40184 20272
rect 40408 20266 40460 20272
rect 39946 20224 40002 20233
rect 39946 20159 40002 20168
rect 40144 20058 40172 20266
rect 40132 20052 40184 20058
rect 40132 19994 40184 20000
rect 40420 19825 40448 20266
rect 40406 19816 40462 19825
rect 39948 19780 40000 19786
rect 40406 19751 40462 19760
rect 39948 19722 40000 19728
rect 39960 19446 39988 19722
rect 40420 19514 40448 19751
rect 40408 19508 40460 19514
rect 40408 19450 40460 19456
rect 39488 19440 39540 19446
rect 39488 19382 39540 19388
rect 39948 19440 40000 19446
rect 39948 19382 40000 19388
rect 38660 19304 38712 19310
rect 38660 19246 38712 19252
rect 39212 19304 39264 19310
rect 39212 19246 39264 19252
rect 38660 18760 38712 18766
rect 38660 18702 38712 18708
rect 38672 18358 38700 18702
rect 38660 18352 38712 18358
rect 38660 18294 38712 18300
rect 39224 17270 39252 19246
rect 39500 18834 39528 19382
rect 40512 19242 40540 20334
rect 40604 19922 40632 20946
rect 40592 19916 40644 19922
rect 40592 19858 40644 19864
rect 40696 19802 40724 21270
rect 40868 20256 40920 20262
rect 40868 20198 40920 20204
rect 40604 19774 40724 19802
rect 40500 19236 40552 19242
rect 40500 19178 40552 19184
rect 39672 19168 39724 19174
rect 39672 19110 39724 19116
rect 40132 19168 40184 19174
rect 40132 19110 40184 19116
rect 39488 18828 39540 18834
rect 39488 18770 39540 18776
rect 39500 18290 39528 18770
rect 39488 18284 39540 18290
rect 39488 18226 39540 18232
rect 39212 17264 39264 17270
rect 39212 17206 39264 17212
rect 39500 17218 39528 18226
rect 39684 18222 39712 19110
rect 40040 18896 40092 18902
rect 40040 18838 40092 18844
rect 39856 18692 39908 18698
rect 39856 18634 39908 18640
rect 39868 18426 39896 18634
rect 39856 18420 39908 18426
rect 39856 18362 39908 18368
rect 39672 18216 39724 18222
rect 39672 18158 39724 18164
rect 39672 17264 39724 17270
rect 39500 17212 39672 17218
rect 39500 17206 39724 17212
rect 38844 17196 38896 17202
rect 39500 17190 39712 17206
rect 38844 17138 38896 17144
rect 38856 16250 38884 17138
rect 39592 16522 39620 17190
rect 39580 16516 39632 16522
rect 39580 16458 39632 16464
rect 38844 16244 38896 16250
rect 38844 16186 38896 16192
rect 39592 16114 39620 16458
rect 39580 16108 39632 16114
rect 39580 16050 39632 16056
rect 38580 15966 38700 15994
rect 38672 15910 38700 15966
rect 38660 15904 38712 15910
rect 38660 15846 38712 15852
rect 39592 15366 39620 16050
rect 39948 15904 40000 15910
rect 39948 15846 40000 15852
rect 39960 15434 39988 15846
rect 39948 15428 40000 15434
rect 39948 15370 40000 15376
rect 39580 15360 39632 15366
rect 39580 15302 39632 15308
rect 40052 15162 40080 18838
rect 40144 17746 40172 19110
rect 40132 17740 40184 17746
rect 40132 17682 40184 17688
rect 40604 17649 40632 19774
rect 40880 18426 40908 20198
rect 40960 19712 41012 19718
rect 40960 19654 41012 19660
rect 40868 18420 40920 18426
rect 40868 18362 40920 18368
rect 40868 17808 40920 17814
rect 40868 17750 40920 17756
rect 40684 17672 40736 17678
rect 40590 17640 40646 17649
rect 40684 17614 40736 17620
rect 40590 17575 40646 17584
rect 40696 16998 40724 17614
rect 40684 16992 40736 16998
rect 40684 16934 40736 16940
rect 40696 16658 40724 16934
rect 40684 16652 40736 16658
rect 40684 16594 40736 16600
rect 40040 15156 40092 15162
rect 40040 15098 40092 15104
rect 40880 15026 40908 17750
rect 40972 16250 41000 19654
rect 41064 19514 41092 22066
rect 41144 21888 41196 21894
rect 41144 21830 41196 21836
rect 41156 21622 41184 21830
rect 41144 21616 41196 21622
rect 41144 21558 41196 21564
rect 41144 19712 41196 19718
rect 41144 19654 41196 19660
rect 41052 19508 41104 19514
rect 41052 19450 41104 19456
rect 41156 19446 41184 19654
rect 41144 19440 41196 19446
rect 41144 19382 41196 19388
rect 41248 18329 41276 23598
rect 41340 23497 41368 23734
rect 41326 23488 41382 23497
rect 41326 23423 41382 23432
rect 41432 22982 41460 23734
rect 41604 23316 41656 23322
rect 41604 23258 41656 23264
rect 41616 22982 41644 23258
rect 41420 22976 41472 22982
rect 41420 22918 41472 22924
rect 41604 22976 41656 22982
rect 41604 22918 41656 22924
rect 41800 22642 41828 24754
rect 42168 24206 42196 26200
rect 42950 24508 43258 24517
rect 42950 24506 42956 24508
rect 43012 24506 43036 24508
rect 43092 24506 43116 24508
rect 43172 24506 43196 24508
rect 43252 24506 43258 24508
rect 43012 24454 43014 24506
rect 43194 24454 43196 24506
rect 42950 24452 42956 24454
rect 43012 24452 43036 24454
rect 43092 24452 43116 24454
rect 43172 24452 43196 24454
rect 43252 24452 43258 24454
rect 42950 24443 43258 24452
rect 42156 24200 42208 24206
rect 42156 24142 42208 24148
rect 43364 24154 43392 26279
rect 43442 26200 43498 27000
rect 44086 26200 44142 27000
rect 44730 26200 44786 27000
rect 45374 26330 45430 27000
rect 45374 26302 45508 26330
rect 45374 26200 45430 26302
rect 43536 24676 43588 24682
rect 43536 24618 43588 24624
rect 43364 24126 43484 24154
rect 43352 24064 43404 24070
rect 43352 24006 43404 24012
rect 42800 23520 42852 23526
rect 42800 23462 42852 23468
rect 42156 23044 42208 23050
rect 42156 22986 42208 22992
rect 41878 22808 41934 22817
rect 41878 22743 41934 22752
rect 41892 22642 41920 22743
rect 41512 22636 41564 22642
rect 41512 22578 41564 22584
rect 41788 22636 41840 22642
rect 41788 22578 41840 22584
rect 41880 22636 41932 22642
rect 41880 22578 41932 22584
rect 41328 22432 41380 22438
rect 41328 22374 41380 22380
rect 41340 21865 41368 22374
rect 41524 21962 41552 22578
rect 41604 22432 41656 22438
rect 41602 22400 41604 22409
rect 41696 22432 41748 22438
rect 41656 22400 41658 22409
rect 41696 22374 41748 22380
rect 41602 22335 41658 22344
rect 41512 21956 41564 21962
rect 41512 21898 41564 21904
rect 41326 21856 41382 21865
rect 41326 21791 41382 21800
rect 41328 21616 41380 21622
rect 41328 21558 41380 21564
rect 41602 21584 41658 21593
rect 41340 18970 41368 21558
rect 41602 21519 41658 21528
rect 41616 21350 41644 21519
rect 41604 21344 41656 21350
rect 41604 21286 41656 21292
rect 41616 19922 41644 21286
rect 41708 20369 41736 22374
rect 42168 22234 42196 22986
rect 42812 22982 42840 23462
rect 42950 23420 43258 23429
rect 42950 23418 42956 23420
rect 43012 23418 43036 23420
rect 43092 23418 43116 23420
rect 43172 23418 43196 23420
rect 43252 23418 43258 23420
rect 43012 23366 43014 23418
rect 43194 23366 43196 23418
rect 42950 23364 42956 23366
rect 43012 23364 43036 23366
rect 43092 23364 43116 23366
rect 43172 23364 43196 23366
rect 43252 23364 43258 23366
rect 42950 23355 43258 23364
rect 43364 23322 43392 24006
rect 43352 23316 43404 23322
rect 43352 23258 43404 23264
rect 43364 23050 43392 23258
rect 43352 23044 43404 23050
rect 43352 22986 43404 22992
rect 42616 22976 42668 22982
rect 42616 22918 42668 22924
rect 42800 22976 42852 22982
rect 42800 22918 42852 22924
rect 42156 22228 42208 22234
rect 42156 22170 42208 22176
rect 42628 22098 42656 22918
rect 42616 22092 42668 22098
rect 42616 22034 42668 22040
rect 42812 21457 42840 22918
rect 43456 22642 43484 24126
rect 43548 23662 43576 24618
rect 43536 23656 43588 23662
rect 43536 23598 43588 23604
rect 44100 23118 44128 26200
rect 44744 24206 44772 26200
rect 45480 24290 45508 26302
rect 46018 26200 46074 27000
rect 46662 26330 46718 27000
rect 46662 26302 46888 26330
rect 46662 26200 46718 26302
rect 45480 24262 45600 24290
rect 45572 24206 45600 24262
rect 46032 24206 46060 26200
rect 46754 25120 46810 25129
rect 46754 25055 46810 25064
rect 46662 24712 46718 24721
rect 46662 24647 46718 24656
rect 44732 24200 44784 24206
rect 44732 24142 44784 24148
rect 45560 24200 45612 24206
rect 45560 24142 45612 24148
rect 46020 24200 46072 24206
rect 46020 24142 46072 24148
rect 46112 24064 46164 24070
rect 46112 24006 46164 24012
rect 45466 23760 45522 23769
rect 45466 23695 45468 23704
rect 45520 23695 45522 23704
rect 45468 23666 45520 23672
rect 43996 23112 44048 23118
rect 43996 23054 44048 23060
rect 44088 23112 44140 23118
rect 44088 23054 44140 23060
rect 43628 23044 43680 23050
rect 43628 22986 43680 22992
rect 43812 23044 43864 23050
rect 43812 22986 43864 22992
rect 43640 22681 43668 22986
rect 43626 22672 43682 22681
rect 43444 22636 43496 22642
rect 43626 22607 43682 22616
rect 43444 22578 43496 22584
rect 43536 22568 43588 22574
rect 43536 22510 43588 22516
rect 42950 22332 43258 22341
rect 42950 22330 42956 22332
rect 43012 22330 43036 22332
rect 43092 22330 43116 22332
rect 43172 22330 43196 22332
rect 43252 22330 43258 22332
rect 43012 22278 43014 22330
rect 43194 22278 43196 22330
rect 42950 22276 42956 22278
rect 43012 22276 43036 22278
rect 43092 22276 43116 22278
rect 43172 22276 43196 22278
rect 43252 22276 43258 22278
rect 42950 22267 43258 22276
rect 43260 21888 43312 21894
rect 43260 21830 43312 21836
rect 42798 21448 42854 21457
rect 43272 21418 43300 21830
rect 42798 21383 42854 21392
rect 43260 21412 43312 21418
rect 43260 21354 43312 21360
rect 42950 21244 43258 21253
rect 42950 21242 42956 21244
rect 43012 21242 43036 21244
rect 43092 21242 43116 21244
rect 43172 21242 43196 21244
rect 43252 21242 43258 21244
rect 43012 21190 43014 21242
rect 43194 21190 43196 21242
rect 42950 21188 42956 21190
rect 43012 21188 43036 21190
rect 43092 21188 43116 21190
rect 43172 21188 43196 21190
rect 43252 21188 43258 21190
rect 42950 21179 43258 21188
rect 43548 20913 43576 22510
rect 43824 22001 43852 22986
rect 43810 21992 43866 22001
rect 43810 21927 43866 21936
rect 43628 21412 43680 21418
rect 43628 21354 43680 21360
rect 43640 21146 43668 21354
rect 43628 21140 43680 21146
rect 43628 21082 43680 21088
rect 44008 21049 44036 23054
rect 45192 22976 45244 22982
rect 45192 22918 45244 22924
rect 45376 22976 45428 22982
rect 45376 22918 45428 22924
rect 45468 22976 45520 22982
rect 45468 22918 45520 22924
rect 45204 22545 45232 22918
rect 45190 22536 45246 22545
rect 45190 22471 45246 22480
rect 44732 22432 44784 22438
rect 44732 22374 44784 22380
rect 44744 22137 44772 22374
rect 44730 22128 44786 22137
rect 44730 22063 44786 22072
rect 43994 21040 44050 21049
rect 43994 20975 44050 20984
rect 43534 20904 43590 20913
rect 43534 20839 43590 20848
rect 45388 20466 45416 22918
rect 45480 22098 45508 22918
rect 45468 22092 45520 22098
rect 45468 22034 45520 22040
rect 45376 20460 45428 20466
rect 45376 20402 45428 20408
rect 41694 20360 41750 20369
rect 41694 20295 41750 20304
rect 42950 20156 43258 20165
rect 42950 20154 42956 20156
rect 43012 20154 43036 20156
rect 43092 20154 43116 20156
rect 43172 20154 43196 20156
rect 43252 20154 43258 20156
rect 43012 20102 43014 20154
rect 43194 20102 43196 20154
rect 42950 20100 42956 20102
rect 43012 20100 43036 20102
rect 43092 20100 43116 20102
rect 43172 20100 43196 20102
rect 43252 20100 43258 20102
rect 41878 20088 41934 20097
rect 42950 20091 43258 20100
rect 41878 20023 41934 20032
rect 41892 19922 41920 20023
rect 41604 19916 41656 19922
rect 41604 19858 41656 19864
rect 41880 19916 41932 19922
rect 41880 19858 41932 19864
rect 46124 19689 46152 24006
rect 46294 23760 46350 23769
rect 46294 23695 46350 23704
rect 46308 23118 46336 23695
rect 46296 23112 46348 23118
rect 46296 23054 46348 23060
rect 46676 22094 46704 24647
rect 46768 22642 46796 25055
rect 46860 23798 46888 26302
rect 47306 26200 47362 27000
rect 47950 26330 48006 27000
rect 47872 26302 48006 26330
rect 47320 24206 47348 26200
rect 47308 24200 47360 24206
rect 47308 24142 47360 24148
rect 46940 24132 46992 24138
rect 46940 24074 46992 24080
rect 46848 23792 46900 23798
rect 46848 23734 46900 23740
rect 46848 23044 46900 23050
rect 46848 22986 46900 22992
rect 46756 22636 46808 22642
rect 46756 22578 46808 22584
rect 46676 22066 46796 22094
rect 46768 22030 46796 22066
rect 46756 22024 46808 22030
rect 46756 21966 46808 21972
rect 46860 21690 46888 22986
rect 46848 21684 46900 21690
rect 46848 21626 46900 21632
rect 46952 21554 46980 24074
rect 47872 23798 47900 26302
rect 47950 26200 48006 26302
rect 48594 26330 48650 27000
rect 48594 26302 48820 26330
rect 48594 26200 48650 26302
rect 48226 25528 48282 25537
rect 48226 25463 48282 25472
rect 48240 24274 48268 25463
rect 48318 24984 48374 24993
rect 48318 24919 48374 24928
rect 48332 24410 48360 24919
rect 48688 24880 48740 24886
rect 48688 24822 48740 24828
rect 48320 24404 48372 24410
rect 48320 24346 48372 24352
rect 48410 24304 48466 24313
rect 48228 24268 48280 24274
rect 48410 24239 48466 24248
rect 48228 24210 48280 24216
rect 47950 23964 48258 23973
rect 47950 23962 47956 23964
rect 48012 23962 48036 23964
rect 48092 23962 48116 23964
rect 48172 23962 48196 23964
rect 48252 23962 48258 23964
rect 48012 23910 48014 23962
rect 48194 23910 48196 23962
rect 47950 23908 47956 23910
rect 48012 23908 48036 23910
rect 48092 23908 48116 23910
rect 48172 23908 48196 23910
rect 48252 23908 48258 23910
rect 47950 23899 48258 23908
rect 47860 23792 47912 23798
rect 47860 23734 47912 23740
rect 47124 23520 47176 23526
rect 47124 23462 47176 23468
rect 47858 23488 47914 23497
rect 47136 21622 47164 23462
rect 47858 23423 47914 23432
rect 47872 23118 47900 23423
rect 47860 23112 47912 23118
rect 48320 23112 48372 23118
rect 47860 23054 47912 23060
rect 48318 23080 48320 23089
rect 48372 23080 48374 23089
rect 48318 23015 48374 23024
rect 47676 22976 47728 22982
rect 47676 22918 47728 22924
rect 47308 22500 47360 22506
rect 47308 22442 47360 22448
rect 47124 21616 47176 21622
rect 47124 21558 47176 21564
rect 46940 21548 46992 21554
rect 46940 21490 46992 21496
rect 46110 19680 46166 19689
rect 46110 19615 46166 19624
rect 41788 19236 41840 19242
rect 41788 19178 41840 19184
rect 41800 18970 41828 19178
rect 42950 19068 43258 19077
rect 42950 19066 42956 19068
rect 43012 19066 43036 19068
rect 43092 19066 43116 19068
rect 43172 19066 43196 19068
rect 43252 19066 43258 19068
rect 43012 19014 43014 19066
rect 43194 19014 43196 19066
rect 42950 19012 42956 19014
rect 43012 19012 43036 19014
rect 43092 19012 43116 19014
rect 43172 19012 43196 19014
rect 43252 19012 43258 19014
rect 42950 19003 43258 19012
rect 41328 18964 41380 18970
rect 41328 18906 41380 18912
rect 41788 18964 41840 18970
rect 41788 18906 41840 18912
rect 47320 18873 47348 22442
rect 47688 21962 47716 22918
rect 47950 22876 48258 22885
rect 47950 22874 47956 22876
rect 48012 22874 48036 22876
rect 48092 22874 48116 22876
rect 48172 22874 48196 22876
rect 48252 22874 48258 22876
rect 48012 22822 48014 22874
rect 48194 22822 48196 22874
rect 47950 22820 47956 22822
rect 48012 22820 48036 22822
rect 48092 22820 48116 22822
rect 48172 22820 48196 22822
rect 48252 22820 48258 22822
rect 47950 22811 48258 22820
rect 48424 22642 48452 24239
rect 48596 24200 48648 24206
rect 48594 24168 48596 24177
rect 48648 24168 48650 24177
rect 48594 24103 48650 24112
rect 48504 22976 48556 22982
rect 48504 22918 48556 22924
rect 48412 22636 48464 22642
rect 48412 22578 48464 22584
rect 47676 21956 47728 21962
rect 47676 21898 47728 21904
rect 48412 21888 48464 21894
rect 48412 21830 48464 21836
rect 47950 21788 48258 21797
rect 47950 21786 47956 21788
rect 48012 21786 48036 21788
rect 48092 21786 48116 21788
rect 48172 21786 48196 21788
rect 48252 21786 48258 21788
rect 48012 21734 48014 21786
rect 48194 21734 48196 21786
rect 47950 21732 47956 21734
rect 48012 21732 48036 21734
rect 48092 21732 48116 21734
rect 48172 21732 48196 21734
rect 48252 21732 48258 21734
rect 47950 21723 48258 21732
rect 48424 20874 48452 21830
rect 48412 20868 48464 20874
rect 48412 20810 48464 20816
rect 47950 20700 48258 20709
rect 47950 20698 47956 20700
rect 48012 20698 48036 20700
rect 48092 20698 48116 20700
rect 48172 20698 48196 20700
rect 48252 20698 48258 20700
rect 48012 20646 48014 20698
rect 48194 20646 48196 20698
rect 47950 20644 47956 20646
rect 48012 20644 48036 20646
rect 48092 20644 48116 20646
rect 48172 20644 48196 20646
rect 48252 20644 48258 20646
rect 47950 20635 48258 20644
rect 48412 20256 48464 20262
rect 48412 20198 48464 20204
rect 48424 19786 48452 20198
rect 48516 19961 48544 22918
rect 48700 22778 48728 24822
rect 48792 23730 48820 26302
rect 49238 26200 49294 27000
rect 48780 23724 48832 23730
rect 48780 23666 48832 23672
rect 49252 23186 49280 26200
rect 49240 23180 49292 23186
rect 49240 23122 49292 23128
rect 49148 23112 49200 23118
rect 49148 23054 49200 23060
rect 48688 22772 48740 22778
rect 48688 22714 48740 22720
rect 49160 22681 49188 23054
rect 49146 22672 49202 22681
rect 49056 22636 49108 22642
rect 49146 22607 49202 22616
rect 49056 22578 49108 22584
rect 49068 22273 49096 22578
rect 49054 22264 49110 22273
rect 49054 22199 49110 22208
rect 48596 22024 48648 22030
rect 48596 21966 48648 21972
rect 48608 21865 48636 21966
rect 49148 21956 49200 21962
rect 49148 21898 49200 21904
rect 48688 21888 48740 21894
rect 48594 21856 48650 21865
rect 48688 21830 48740 21836
rect 48594 21791 48650 21800
rect 48596 20460 48648 20466
rect 48596 20402 48648 20408
rect 48608 20233 48636 20402
rect 48594 20224 48650 20233
rect 48594 20159 48650 20168
rect 48502 19952 48558 19961
rect 48502 19887 48558 19896
rect 48412 19780 48464 19786
rect 48412 19722 48464 19728
rect 47950 19612 48258 19621
rect 47950 19610 47956 19612
rect 48012 19610 48036 19612
rect 48092 19610 48116 19612
rect 48172 19610 48196 19612
rect 48252 19610 48258 19612
rect 48012 19558 48014 19610
rect 48194 19558 48196 19610
rect 47950 19556 47956 19558
rect 48012 19556 48036 19558
rect 48092 19556 48116 19558
rect 48172 19556 48196 19558
rect 48252 19556 48258 19558
rect 47950 19547 48258 19556
rect 48700 19417 48728 21830
rect 49056 21548 49108 21554
rect 49056 21490 49108 21496
rect 48964 21412 49016 21418
rect 48964 21354 49016 21360
rect 48976 21146 49004 21354
rect 48964 21140 49016 21146
rect 48964 21082 49016 21088
rect 49068 21049 49096 21490
rect 49160 21457 49188 21898
rect 49146 21448 49202 21457
rect 49146 21383 49202 21392
rect 49054 21040 49110 21049
rect 49054 20975 49110 20984
rect 49056 20936 49108 20942
rect 49056 20878 49108 20884
rect 49068 20641 49096 20878
rect 49054 20632 49110 20641
rect 49054 20567 49110 20576
rect 49056 20460 49108 20466
rect 49056 20402 49108 20408
rect 49068 19825 49096 20402
rect 49054 19816 49110 19825
rect 49054 19751 49110 19760
rect 49332 19780 49384 19786
rect 49332 19722 49384 19728
rect 49344 19417 49372 19722
rect 48686 19408 48742 19417
rect 49330 19408 49386 19417
rect 48686 19343 48742 19352
rect 49148 19372 49200 19378
rect 49330 19343 49386 19352
rect 49148 19314 49200 19320
rect 47400 19168 47452 19174
rect 47400 19110 47452 19116
rect 47306 18864 47362 18873
rect 47306 18799 47362 18808
rect 47412 18630 47440 19110
rect 49160 19009 49188 19314
rect 49146 19000 49202 19009
rect 49146 18935 49202 18944
rect 48596 18760 48648 18766
rect 48596 18702 48648 18708
rect 49148 18760 49200 18766
rect 49148 18702 49200 18708
rect 47400 18624 47452 18630
rect 47400 18566 47452 18572
rect 48412 18624 48464 18630
rect 48608 18601 48636 18702
rect 48412 18566 48464 18572
rect 48594 18592 48650 18601
rect 47950 18524 48258 18533
rect 47950 18522 47956 18524
rect 48012 18522 48036 18524
rect 48092 18522 48116 18524
rect 48172 18522 48196 18524
rect 48252 18522 48258 18524
rect 48012 18470 48014 18522
rect 48194 18470 48196 18522
rect 47950 18468 47956 18470
rect 48012 18468 48036 18470
rect 48092 18468 48116 18470
rect 48172 18468 48196 18470
rect 48252 18468 48258 18470
rect 47950 18459 48258 18468
rect 41420 18420 41472 18426
rect 41420 18362 41472 18368
rect 41234 18320 41290 18329
rect 41234 18255 41290 18264
rect 41432 17241 41460 18362
rect 48424 18358 48452 18566
rect 48594 18527 48650 18536
rect 48412 18352 48464 18358
rect 48412 18294 48464 18300
rect 49056 18284 49108 18290
rect 49056 18226 49108 18232
rect 45560 18080 45612 18086
rect 45560 18022 45612 18028
rect 42950 17980 43258 17989
rect 42950 17978 42956 17980
rect 43012 17978 43036 17980
rect 43092 17978 43116 17980
rect 43172 17978 43196 17980
rect 43252 17978 43258 17980
rect 43012 17926 43014 17978
rect 43194 17926 43196 17978
rect 42950 17924 42956 17926
rect 43012 17924 43036 17926
rect 43092 17924 43116 17926
rect 43172 17924 43196 17926
rect 43252 17924 43258 17926
rect 42950 17915 43258 17924
rect 41418 17232 41474 17241
rect 41418 17167 41474 17176
rect 42950 16892 43258 16901
rect 42950 16890 42956 16892
rect 43012 16890 43036 16892
rect 43092 16890 43116 16892
rect 43172 16890 43196 16892
rect 43252 16890 43258 16892
rect 43012 16838 43014 16890
rect 43194 16838 43196 16890
rect 42950 16836 42956 16838
rect 43012 16836 43036 16838
rect 43092 16836 43116 16838
rect 43172 16836 43196 16838
rect 43252 16836 43258 16838
rect 42950 16827 43258 16836
rect 40960 16244 41012 16250
rect 40960 16186 41012 16192
rect 41788 16040 41840 16046
rect 41788 15982 41840 15988
rect 41800 15706 41828 15982
rect 42950 15804 43258 15813
rect 42950 15802 42956 15804
rect 43012 15802 43036 15804
rect 43092 15802 43116 15804
rect 43172 15802 43196 15804
rect 43252 15802 43258 15804
rect 43012 15750 43014 15802
rect 43194 15750 43196 15802
rect 42950 15748 42956 15750
rect 43012 15748 43036 15750
rect 43092 15748 43116 15750
rect 43172 15748 43196 15750
rect 43252 15748 43258 15750
rect 42950 15739 43258 15748
rect 41788 15700 41840 15706
rect 41788 15642 41840 15648
rect 45572 15609 45600 18022
rect 49068 17785 49096 18226
rect 49160 18193 49188 18702
rect 49240 18624 49292 18630
rect 49240 18566 49292 18572
rect 49252 18426 49280 18566
rect 49240 18420 49292 18426
rect 49240 18362 49292 18368
rect 49146 18184 49202 18193
rect 49146 18119 49202 18128
rect 49054 17776 49110 17785
rect 49054 17711 49110 17720
rect 49056 17672 49108 17678
rect 49056 17614 49108 17620
rect 48412 17604 48464 17610
rect 48412 17546 48464 17552
rect 47400 17536 47452 17542
rect 47400 17478 47452 17484
rect 47412 17066 47440 17478
rect 47950 17436 48258 17445
rect 47950 17434 47956 17436
rect 48012 17434 48036 17436
rect 48092 17434 48116 17436
rect 48172 17434 48196 17436
rect 48252 17434 48258 17436
rect 48012 17382 48014 17434
rect 48194 17382 48196 17434
rect 47950 17380 47956 17382
rect 48012 17380 48036 17382
rect 48092 17380 48116 17382
rect 48172 17380 48196 17382
rect 48252 17380 48258 17382
rect 47950 17371 48258 17380
rect 48424 17338 48452 17546
rect 49068 17377 49096 17614
rect 49054 17368 49110 17377
rect 48412 17332 48464 17338
rect 49054 17303 49110 17312
rect 48412 17274 48464 17280
rect 48228 17264 48280 17270
rect 48228 17206 48280 17212
rect 47400 17060 47452 17066
rect 47400 17002 47452 17008
rect 48240 16561 48268 17206
rect 48596 17196 48648 17202
rect 48596 17138 48648 17144
rect 48608 16969 48636 17138
rect 49240 16992 49292 16998
rect 48594 16960 48650 16969
rect 49240 16934 49292 16940
rect 48594 16895 48650 16904
rect 49252 16794 49280 16934
rect 49240 16788 49292 16794
rect 49240 16730 49292 16736
rect 49148 16584 49200 16590
rect 48226 16552 48282 16561
rect 49148 16526 49200 16532
rect 48226 16487 48282 16496
rect 47950 16348 48258 16357
rect 47950 16346 47956 16348
rect 48012 16346 48036 16348
rect 48092 16346 48116 16348
rect 48172 16346 48196 16348
rect 48252 16346 48258 16348
rect 48012 16294 48014 16346
rect 48194 16294 48196 16346
rect 47950 16292 47956 16294
rect 48012 16292 48036 16294
rect 48092 16292 48116 16294
rect 48172 16292 48196 16294
rect 48252 16292 48258 16294
rect 47950 16283 48258 16292
rect 49160 16153 49188 16526
rect 49240 16448 49292 16454
rect 49240 16390 49292 16396
rect 49146 16144 49202 16153
rect 48964 16108 49016 16114
rect 48964 16050 49016 16056
rect 49056 16108 49108 16114
rect 49146 16079 49202 16088
rect 49056 16050 49108 16056
rect 48688 15904 48740 15910
rect 48688 15846 48740 15852
rect 45558 15600 45614 15609
rect 45558 15535 45614 15544
rect 47950 15260 48258 15269
rect 47950 15258 47956 15260
rect 48012 15258 48036 15260
rect 48092 15258 48116 15260
rect 48172 15258 48196 15260
rect 48252 15258 48258 15260
rect 48012 15206 48014 15258
rect 48194 15206 48196 15258
rect 47950 15204 47956 15206
rect 48012 15204 48036 15206
rect 48092 15204 48116 15206
rect 48172 15204 48196 15206
rect 48252 15204 48258 15206
rect 47950 15195 48258 15204
rect 48502 15056 48558 15065
rect 40868 15020 40920 15026
rect 48502 14991 48558 15000
rect 40868 14962 40920 14968
rect 39304 14952 39356 14958
rect 48412 14952 48464 14958
rect 39304 14894 39356 14900
rect 48318 14920 48374 14929
rect 39316 14822 39344 14894
rect 48412 14894 48464 14900
rect 48318 14855 48320 14864
rect 48372 14855 48374 14864
rect 48320 14826 48372 14832
rect 38476 14816 38528 14822
rect 38476 14758 38528 14764
rect 39304 14816 39356 14822
rect 39304 14758 39356 14764
rect 45836 14816 45888 14822
rect 45836 14758 45888 14764
rect 38488 13977 38516 14758
rect 39316 14550 39344 14758
rect 42950 14716 43258 14725
rect 42950 14714 42956 14716
rect 43012 14714 43036 14716
rect 43092 14714 43116 14716
rect 43172 14714 43196 14716
rect 43252 14714 43258 14716
rect 43012 14662 43014 14714
rect 43194 14662 43196 14714
rect 42950 14660 42956 14662
rect 43012 14660 43036 14662
rect 43092 14660 43116 14662
rect 43172 14660 43196 14662
rect 43252 14660 43258 14662
rect 42950 14651 43258 14660
rect 39304 14544 39356 14550
rect 39304 14486 39356 14492
rect 45008 14272 45060 14278
rect 45008 14214 45060 14220
rect 41512 14068 41564 14074
rect 41512 14010 41564 14016
rect 38474 13968 38530 13977
rect 38474 13903 38530 13912
rect 38844 13728 38896 13734
rect 38844 13670 38896 13676
rect 38384 13524 38436 13530
rect 38384 13466 38436 13472
rect 38856 13462 38884 13670
rect 38844 13456 38896 13462
rect 38844 13398 38896 13404
rect 37832 13388 37884 13394
rect 37832 13330 37884 13336
rect 37384 13110 37780 13138
rect 37648 12096 37700 12102
rect 37648 12038 37700 12044
rect 37280 11824 37332 11830
rect 37280 11766 37332 11772
rect 36544 11756 36596 11762
rect 36544 11698 36596 11704
rect 36728 11756 36780 11762
rect 36728 11698 36780 11704
rect 36450 11112 36506 11121
rect 36556 11082 36584 11698
rect 37004 11620 37056 11626
rect 37004 11562 37056 11568
rect 36450 11047 36506 11056
rect 36544 11076 36596 11082
rect 36464 11014 36492 11047
rect 36544 11018 36596 11024
rect 36452 11008 36504 11014
rect 36452 10950 36504 10956
rect 36542 10976 36598 10985
rect 36464 10674 36492 10950
rect 36542 10911 36598 10920
rect 36556 10674 36584 10911
rect 37016 10810 37044 11562
rect 37464 11076 37516 11082
rect 37464 11018 37516 11024
rect 37004 10804 37056 10810
rect 37004 10746 37056 10752
rect 37280 10736 37332 10742
rect 37280 10678 37332 10684
rect 36452 10668 36504 10674
rect 36452 10610 36504 10616
rect 36544 10668 36596 10674
rect 36544 10610 36596 10616
rect 36268 10600 36320 10606
rect 36268 10542 36320 10548
rect 35808 7948 35860 7954
rect 35808 7890 35860 7896
rect 35532 7336 35584 7342
rect 35532 7278 35584 7284
rect 36556 4690 36584 10610
rect 37292 9178 37320 10678
rect 37476 9518 37504 11018
rect 37660 10606 37688 12038
rect 37648 10600 37700 10606
rect 37648 10542 37700 10548
rect 37752 10130 37780 13110
rect 37844 12306 37872 13330
rect 41524 13326 41552 14010
rect 45020 14006 45048 14214
rect 45008 14000 45060 14006
rect 45008 13942 45060 13948
rect 45848 13938 45876 14758
rect 47950 14172 48258 14181
rect 47950 14170 47956 14172
rect 48012 14170 48036 14172
rect 48092 14170 48116 14172
rect 48172 14170 48196 14172
rect 48252 14170 48258 14172
rect 48012 14118 48014 14170
rect 48194 14118 48196 14170
rect 47950 14116 47956 14118
rect 48012 14116 48036 14118
rect 48092 14116 48116 14118
rect 48172 14116 48196 14118
rect 48252 14116 48258 14118
rect 47950 14107 48258 14116
rect 48424 14074 48452 14894
rect 48516 14074 48544 14991
rect 47032 14068 47084 14074
rect 47032 14010 47084 14016
rect 48412 14068 48464 14074
rect 48412 14010 48464 14016
rect 48504 14068 48556 14074
rect 48504 14010 48556 14016
rect 46848 14000 46900 14006
rect 46848 13942 46900 13948
rect 45836 13932 45888 13938
rect 45836 13874 45888 13880
rect 46296 13864 46348 13870
rect 46296 13806 46348 13812
rect 42950 13628 43258 13637
rect 42950 13626 42956 13628
rect 43012 13626 43036 13628
rect 43092 13626 43116 13628
rect 43172 13626 43196 13628
rect 43252 13626 43258 13628
rect 43012 13574 43014 13626
rect 43194 13574 43196 13626
rect 42950 13572 42956 13574
rect 43012 13572 43036 13574
rect 43092 13572 43116 13574
rect 43172 13572 43196 13574
rect 43252 13572 43258 13574
rect 42950 13563 43258 13572
rect 46308 13326 46336 13806
rect 41512 13320 41564 13326
rect 41512 13262 41564 13268
rect 46296 13320 46348 13326
rect 46296 13262 46348 13268
rect 46112 13184 46164 13190
rect 46112 13126 46164 13132
rect 37950 13084 38258 13093
rect 37950 13082 37956 13084
rect 38012 13082 38036 13084
rect 38092 13082 38116 13084
rect 38172 13082 38196 13084
rect 38252 13082 38258 13084
rect 38012 13030 38014 13082
rect 38194 13030 38196 13082
rect 37950 13028 37956 13030
rect 38012 13028 38036 13030
rect 38092 13028 38116 13030
rect 38172 13028 38196 13030
rect 38252 13028 38258 13030
rect 37950 13019 38258 13028
rect 39948 12912 40000 12918
rect 39948 12854 40000 12860
rect 39304 12708 39356 12714
rect 39304 12650 39356 12656
rect 37832 12300 37884 12306
rect 37832 12242 37884 12248
rect 38292 12300 38344 12306
rect 38292 12242 38344 12248
rect 37950 11996 38258 12005
rect 37950 11994 37956 11996
rect 38012 11994 38036 11996
rect 38092 11994 38116 11996
rect 38172 11994 38196 11996
rect 38252 11994 38258 11996
rect 38012 11942 38014 11994
rect 38194 11942 38196 11994
rect 37950 11940 37956 11942
rect 38012 11940 38036 11942
rect 38092 11940 38116 11942
rect 38172 11940 38196 11942
rect 38252 11940 38258 11942
rect 37950 11931 38258 11940
rect 38304 11558 38332 12242
rect 39316 12238 39344 12650
rect 39396 12436 39448 12442
rect 39396 12378 39448 12384
rect 39304 12232 39356 12238
rect 39304 12174 39356 12180
rect 39408 11830 39436 12378
rect 39960 12238 39988 12854
rect 46124 12850 46152 13126
rect 46112 12844 46164 12850
rect 46112 12786 46164 12792
rect 46860 12753 46888 13942
rect 47044 12850 47072 14010
rect 48700 14006 48728 15846
rect 48976 15706 49004 16050
rect 49068 15745 49096 16050
rect 49054 15736 49110 15745
rect 48964 15700 49016 15706
rect 49054 15671 49110 15680
rect 48964 15642 49016 15648
rect 49252 15473 49280 16390
rect 49332 15496 49384 15502
rect 49238 15464 49294 15473
rect 49332 15438 49384 15444
rect 49238 15399 49294 15408
rect 49344 15337 49372 15438
rect 49330 15328 49386 15337
rect 49330 15263 49386 15272
rect 49056 15020 49108 15026
rect 49056 14962 49108 14968
rect 49068 14929 49096 14962
rect 49054 14920 49110 14929
rect 49054 14855 49110 14864
rect 49054 14512 49110 14521
rect 49054 14447 49110 14456
rect 49068 14414 49096 14447
rect 49056 14408 49108 14414
rect 49056 14350 49108 14356
rect 49238 14376 49294 14385
rect 49238 14311 49294 14320
rect 49252 14278 49280 14311
rect 49240 14272 49292 14278
rect 49240 14214 49292 14220
rect 49146 14104 49202 14113
rect 49146 14039 49202 14048
rect 49160 14006 49188 14039
rect 48688 14000 48740 14006
rect 48688 13942 48740 13948
rect 49148 14000 49200 14006
rect 49148 13942 49200 13948
rect 48228 13932 48280 13938
rect 48228 13874 48280 13880
rect 48240 13705 48268 13874
rect 48226 13696 48282 13705
rect 48226 13631 48282 13640
rect 49148 13320 49200 13326
rect 49146 13288 49148 13297
rect 49200 13288 49202 13297
rect 49146 13223 49202 13232
rect 47950 13084 48258 13093
rect 47950 13082 47956 13084
rect 48012 13082 48036 13084
rect 48092 13082 48116 13084
rect 48172 13082 48196 13084
rect 48252 13082 48258 13084
rect 48012 13030 48014 13082
rect 48194 13030 48196 13082
rect 47950 13028 47956 13030
rect 48012 13028 48036 13030
rect 48092 13028 48116 13030
rect 48172 13028 48196 13030
rect 48252 13028 48258 13030
rect 47950 13019 48258 13028
rect 49146 12880 49202 12889
rect 47032 12844 47084 12850
rect 49146 12815 49148 12824
rect 47032 12786 47084 12792
rect 49200 12815 49202 12824
rect 49148 12786 49200 12792
rect 46846 12744 46902 12753
rect 46846 12679 46902 12688
rect 42708 12640 42760 12646
rect 42708 12582 42760 12588
rect 47952 12640 48004 12646
rect 47952 12582 48004 12588
rect 39948 12232 40000 12238
rect 39948 12174 40000 12180
rect 40224 12096 40276 12102
rect 40224 12038 40276 12044
rect 40236 11830 40264 12038
rect 39396 11824 39448 11830
rect 39396 11766 39448 11772
rect 40224 11824 40276 11830
rect 40224 11766 40276 11772
rect 38384 11756 38436 11762
rect 38384 11698 38436 11704
rect 38292 11552 38344 11558
rect 38292 11494 38344 11500
rect 37950 10908 38258 10917
rect 37950 10906 37956 10908
rect 38012 10906 38036 10908
rect 38092 10906 38116 10908
rect 38172 10906 38196 10908
rect 38252 10906 38258 10908
rect 38012 10854 38014 10906
rect 38194 10854 38196 10906
rect 37950 10852 37956 10854
rect 38012 10852 38036 10854
rect 38092 10852 38116 10854
rect 38172 10852 38196 10854
rect 38252 10852 38258 10854
rect 37950 10843 38258 10852
rect 37832 10464 37884 10470
rect 37832 10406 37884 10412
rect 37740 10124 37792 10130
rect 37740 10066 37792 10072
rect 37844 10062 37872 10406
rect 37832 10056 37884 10062
rect 37832 9998 37884 10004
rect 37950 9820 38258 9829
rect 37950 9818 37956 9820
rect 38012 9818 38036 9820
rect 38092 9818 38116 9820
rect 38172 9818 38196 9820
rect 38252 9818 38258 9820
rect 38012 9766 38014 9818
rect 38194 9766 38196 9818
rect 37950 9764 37956 9766
rect 38012 9764 38036 9766
rect 38092 9764 38116 9766
rect 38172 9764 38196 9766
rect 38252 9764 38258 9766
rect 37950 9755 38258 9764
rect 37464 9512 37516 9518
rect 37464 9454 37516 9460
rect 37280 9172 37332 9178
rect 37280 9114 37332 9120
rect 37950 8732 38258 8741
rect 37950 8730 37956 8732
rect 38012 8730 38036 8732
rect 38092 8730 38116 8732
rect 38172 8730 38196 8732
rect 38252 8730 38258 8732
rect 38012 8678 38014 8730
rect 38194 8678 38196 8730
rect 37950 8676 37956 8678
rect 38012 8676 38036 8678
rect 38092 8676 38116 8678
rect 38172 8676 38196 8678
rect 38252 8676 38258 8678
rect 37950 8667 38258 8676
rect 38396 8022 38424 11698
rect 40130 11384 40186 11393
rect 40130 11319 40186 11328
rect 42616 11348 42668 11354
rect 39764 10668 39816 10674
rect 39764 10610 39816 10616
rect 39776 10169 39804 10610
rect 39762 10160 39818 10169
rect 39762 10095 39818 10104
rect 40144 9994 40172 11319
rect 42616 11290 42668 11296
rect 40960 11144 41012 11150
rect 40960 11086 41012 11092
rect 40972 10266 41000 11086
rect 40960 10260 41012 10266
rect 40960 10202 41012 10208
rect 42628 10062 42656 11290
rect 42720 11286 42748 12582
rect 42950 12540 43258 12549
rect 42950 12538 42956 12540
rect 43012 12538 43036 12540
rect 43092 12538 43116 12540
rect 43172 12538 43196 12540
rect 43252 12538 43258 12540
rect 43012 12486 43014 12538
rect 43194 12486 43196 12538
rect 42950 12484 42956 12486
rect 43012 12484 43036 12486
rect 43092 12484 43116 12486
rect 43172 12484 43196 12486
rect 43252 12484 43258 12486
rect 42950 12475 43258 12484
rect 47964 12238 47992 12582
rect 49146 12472 49202 12481
rect 49146 12407 49202 12416
rect 49160 12306 49188 12407
rect 49148 12300 49200 12306
rect 49148 12242 49200 12248
rect 47952 12232 48004 12238
rect 47952 12174 48004 12180
rect 47032 12164 47084 12170
rect 47032 12106 47084 12112
rect 45928 12096 45980 12102
rect 45928 12038 45980 12044
rect 45940 11762 45968 12038
rect 45928 11756 45980 11762
rect 45928 11698 45980 11704
rect 44180 11620 44232 11626
rect 44180 11562 44232 11568
rect 46664 11620 46716 11626
rect 46664 11562 46716 11568
rect 42950 11452 43258 11461
rect 42950 11450 42956 11452
rect 43012 11450 43036 11452
rect 43092 11450 43116 11452
rect 43172 11450 43196 11452
rect 43252 11450 43258 11452
rect 43012 11398 43014 11450
rect 43194 11398 43196 11450
rect 42950 11396 42956 11398
rect 43012 11396 43036 11398
rect 43092 11396 43116 11398
rect 43172 11396 43196 11398
rect 43252 11396 43258 11398
rect 42950 11387 43258 11396
rect 42708 11280 42760 11286
rect 42708 11222 42760 11228
rect 43720 10532 43772 10538
rect 43720 10474 43772 10480
rect 42950 10364 43258 10373
rect 42950 10362 42956 10364
rect 43012 10362 43036 10364
rect 43092 10362 43116 10364
rect 43172 10362 43196 10364
rect 43252 10362 43258 10364
rect 43012 10310 43014 10362
rect 43194 10310 43196 10362
rect 42950 10308 42956 10310
rect 43012 10308 43036 10310
rect 43092 10308 43116 10310
rect 43172 10308 43196 10310
rect 43252 10308 43258 10310
rect 42950 10299 43258 10308
rect 42616 10056 42668 10062
rect 42616 9998 42668 10004
rect 38752 9988 38804 9994
rect 38752 9930 38804 9936
rect 40132 9988 40184 9994
rect 40132 9930 40184 9936
rect 42708 9988 42760 9994
rect 42708 9930 42760 9936
rect 38764 9722 38792 9930
rect 38752 9716 38804 9722
rect 38752 9658 38804 9664
rect 38750 8936 38806 8945
rect 38750 8871 38806 8880
rect 38476 8288 38528 8294
rect 38476 8230 38528 8236
rect 38384 8016 38436 8022
rect 38384 7958 38436 7964
rect 37950 7644 38258 7653
rect 37950 7642 37956 7644
rect 38012 7642 38036 7644
rect 38092 7642 38116 7644
rect 38172 7642 38196 7644
rect 38252 7642 38258 7644
rect 38012 7590 38014 7642
rect 38194 7590 38196 7642
rect 37950 7588 37956 7590
rect 38012 7588 38036 7590
rect 38092 7588 38116 7590
rect 38172 7588 38196 7590
rect 38252 7588 38258 7590
rect 37950 7579 38258 7588
rect 37924 7200 37976 7206
rect 37924 7142 37976 7148
rect 37936 6934 37964 7142
rect 37924 6928 37976 6934
rect 37924 6870 37976 6876
rect 37740 6860 37792 6866
rect 37740 6802 37792 6808
rect 37648 6112 37700 6118
rect 37648 6054 37700 6060
rect 37660 5914 37688 6054
rect 37648 5908 37700 5914
rect 37648 5850 37700 5856
rect 37752 5302 37780 6802
rect 37950 6556 38258 6565
rect 37950 6554 37956 6556
rect 38012 6554 38036 6556
rect 38092 6554 38116 6556
rect 38172 6554 38196 6556
rect 38252 6554 38258 6556
rect 38012 6502 38014 6554
rect 38194 6502 38196 6554
rect 37950 6500 37956 6502
rect 38012 6500 38036 6502
rect 38092 6500 38116 6502
rect 38172 6500 38196 6502
rect 38252 6500 38258 6502
rect 37950 6491 38258 6500
rect 37950 5468 38258 5477
rect 37950 5466 37956 5468
rect 38012 5466 38036 5468
rect 38092 5466 38116 5468
rect 38172 5466 38196 5468
rect 38252 5466 38258 5468
rect 38012 5414 38014 5466
rect 38194 5414 38196 5466
rect 37950 5412 37956 5414
rect 38012 5412 38036 5414
rect 38092 5412 38116 5414
rect 38172 5412 38196 5414
rect 38252 5412 38258 5414
rect 37950 5403 38258 5412
rect 38488 5302 38516 8230
rect 38764 7886 38792 8871
rect 40224 8628 40276 8634
rect 40224 8570 40276 8576
rect 40132 8356 40184 8362
rect 40132 8298 40184 8304
rect 38752 7880 38804 7886
rect 38752 7822 38804 7828
rect 40040 7812 40092 7818
rect 40040 7754 40092 7760
rect 38660 7744 38712 7750
rect 38660 7686 38712 7692
rect 38672 7546 38700 7686
rect 38660 7540 38712 7546
rect 38660 7482 38712 7488
rect 40052 6798 40080 7754
rect 40144 7478 40172 8298
rect 40132 7472 40184 7478
rect 40132 7414 40184 7420
rect 40040 6792 40092 6798
rect 40040 6734 40092 6740
rect 40236 6390 40264 8570
rect 42720 8498 42748 9930
rect 42800 9920 42852 9926
rect 42800 9862 42852 9868
rect 42708 8492 42760 8498
rect 42708 8434 42760 8440
rect 42812 7410 42840 9862
rect 42950 9276 43258 9285
rect 42950 9274 42956 9276
rect 43012 9274 43036 9276
rect 43092 9274 43116 9276
rect 43172 9274 43196 9276
rect 43252 9274 43258 9276
rect 43012 9222 43014 9274
rect 43194 9222 43196 9274
rect 42950 9220 42956 9222
rect 43012 9220 43036 9222
rect 43092 9220 43116 9222
rect 43172 9220 43196 9222
rect 43252 9220 43258 9222
rect 42950 9211 43258 9220
rect 43628 8968 43680 8974
rect 43628 8910 43680 8916
rect 42950 8188 43258 8197
rect 42950 8186 42956 8188
rect 43012 8186 43036 8188
rect 43092 8186 43116 8188
rect 43172 8186 43196 8188
rect 43252 8186 43258 8188
rect 43012 8134 43014 8186
rect 43194 8134 43196 8186
rect 42950 8132 42956 8134
rect 43012 8132 43036 8134
rect 43092 8132 43116 8134
rect 43172 8132 43196 8134
rect 43252 8132 43258 8134
rect 42950 8123 43258 8132
rect 42800 7404 42852 7410
rect 42800 7346 42852 7352
rect 42950 7100 43258 7109
rect 42950 7098 42956 7100
rect 43012 7098 43036 7100
rect 43092 7098 43116 7100
rect 43172 7098 43196 7100
rect 43252 7098 43258 7100
rect 43012 7046 43014 7098
rect 43194 7046 43196 7098
rect 42950 7044 42956 7046
rect 43012 7044 43036 7046
rect 43092 7044 43116 7046
rect 43172 7044 43196 7046
rect 43252 7044 43258 7046
rect 42950 7035 43258 7044
rect 43640 6914 43668 8910
rect 43732 7886 43760 10474
rect 44192 8974 44220 11562
rect 45744 11076 45796 11082
rect 45744 11018 45796 11024
rect 45756 10062 45784 11018
rect 46676 10062 46704 11562
rect 46940 11076 46992 11082
rect 46940 11018 46992 11024
rect 46952 10674 46980 11018
rect 46940 10668 46992 10674
rect 46940 10610 46992 10616
rect 45744 10056 45796 10062
rect 45744 9998 45796 10004
rect 46664 10056 46716 10062
rect 46664 9998 46716 10004
rect 46756 9988 46808 9994
rect 46756 9930 46808 9936
rect 44180 8968 44232 8974
rect 44180 8910 44232 8916
rect 46572 8900 46624 8906
rect 46572 8842 46624 8848
rect 44272 8832 44324 8838
rect 44272 8774 44324 8780
rect 44284 8566 44312 8774
rect 44272 8560 44324 8566
rect 44272 8502 44324 8508
rect 43720 7880 43772 7886
rect 43720 7822 43772 7828
rect 45744 7268 45796 7274
rect 45744 7210 45796 7216
rect 43640 6886 43760 6914
rect 40224 6384 40276 6390
rect 40224 6326 40276 6332
rect 42950 6012 43258 6021
rect 42950 6010 42956 6012
rect 43012 6010 43036 6012
rect 43092 6010 43116 6012
rect 43172 6010 43196 6012
rect 43252 6010 43258 6012
rect 43012 5958 43014 6010
rect 43194 5958 43196 6010
rect 42950 5956 42956 5958
rect 43012 5956 43036 5958
rect 43092 5956 43116 5958
rect 43172 5956 43196 5958
rect 43252 5956 43258 5958
rect 42950 5947 43258 5956
rect 43732 5710 43760 6886
rect 45560 6112 45612 6118
rect 45560 6054 45612 6060
rect 43720 5704 43772 5710
rect 43720 5646 43772 5652
rect 37740 5296 37792 5302
rect 37740 5238 37792 5244
rect 38476 5296 38528 5302
rect 38476 5238 38528 5244
rect 40040 5092 40092 5098
rect 40040 5034 40092 5040
rect 37280 5024 37332 5030
rect 37280 4966 37332 4972
rect 37832 5024 37884 5030
rect 37832 4966 37884 4972
rect 36544 4684 36596 4690
rect 36544 4626 36596 4632
rect 37292 4554 37320 4966
rect 37844 4826 37872 4966
rect 37832 4820 37884 4826
rect 37832 4762 37884 4768
rect 37280 4548 37332 4554
rect 37280 4490 37332 4496
rect 39856 4548 39908 4554
rect 39856 4490 39908 4496
rect 37950 4380 38258 4389
rect 37950 4378 37956 4380
rect 38012 4378 38036 4380
rect 38092 4378 38116 4380
rect 38172 4378 38196 4380
rect 38252 4378 38258 4380
rect 38012 4326 38014 4378
rect 38194 4326 38196 4378
rect 37950 4324 37956 4326
rect 38012 4324 38036 4326
rect 38092 4324 38116 4326
rect 38172 4324 38196 4326
rect 38252 4324 38258 4326
rect 37950 4315 38258 4324
rect 36544 4140 36596 4146
rect 36544 4082 36596 4088
rect 34428 3936 34480 3942
rect 34428 3878 34480 3884
rect 32950 2748 33258 2757
rect 32950 2746 32956 2748
rect 33012 2746 33036 2748
rect 33092 2746 33116 2748
rect 33172 2746 33196 2748
rect 33252 2746 33258 2748
rect 34164 2746 34376 2774
rect 33012 2694 33014 2746
rect 33194 2694 33196 2746
rect 32950 2692 32956 2694
rect 33012 2692 33036 2694
rect 33092 2692 33116 2694
rect 33172 2692 33196 2694
rect 33252 2692 33258 2694
rect 32950 2683 33258 2692
rect 28908 2644 28960 2650
rect 28908 2586 28960 2592
rect 34348 2582 34376 2746
rect 34440 2650 34468 3878
rect 36556 3738 36584 4082
rect 36544 3732 36596 3738
rect 36544 3674 36596 3680
rect 39212 3392 39264 3398
rect 39212 3334 39264 3340
rect 37950 3292 38258 3301
rect 37950 3290 37956 3292
rect 38012 3290 38036 3292
rect 38092 3290 38116 3292
rect 38172 3290 38196 3292
rect 38252 3290 38258 3292
rect 38012 3238 38014 3290
rect 38194 3238 38196 3290
rect 37950 3236 37956 3238
rect 38012 3236 38036 3238
rect 38092 3236 38116 3238
rect 38172 3236 38196 3238
rect 38252 3236 38258 3238
rect 37950 3227 38258 3236
rect 36820 3188 36872 3194
rect 36820 3130 36872 3136
rect 34428 2644 34480 2650
rect 34428 2586 34480 2592
rect 34336 2576 34388 2582
rect 34336 2518 34388 2524
rect 36832 2514 36860 3130
rect 38108 2848 38160 2854
rect 38108 2790 38160 2796
rect 36820 2508 36872 2514
rect 36820 2450 36872 2456
rect 38120 2446 38148 2790
rect 30748 2440 30800 2446
rect 30748 2382 30800 2388
rect 32864 2440 32916 2446
rect 32864 2382 32916 2388
rect 34980 2440 35032 2446
rect 34980 2382 35032 2388
rect 37096 2440 37148 2446
rect 37096 2382 37148 2388
rect 38108 2440 38160 2446
rect 38108 2382 38160 2388
rect 28724 2304 28776 2310
rect 28724 2246 28776 2252
rect 30760 800 30788 2382
rect 32876 800 32904 2382
rect 34992 800 35020 2382
rect 37108 800 37136 2382
rect 37950 2204 38258 2213
rect 37950 2202 37956 2204
rect 38012 2202 38036 2204
rect 38092 2202 38116 2204
rect 38172 2202 38196 2204
rect 38252 2202 38258 2204
rect 38012 2150 38014 2202
rect 38194 2150 38196 2202
rect 37950 2148 37956 2150
rect 38012 2148 38036 2150
rect 38092 2148 38116 2150
rect 38172 2148 38196 2150
rect 38252 2148 38258 2150
rect 37950 2139 38258 2148
rect 39224 800 39252 3334
rect 39868 3058 39896 4490
rect 40052 3602 40080 5034
rect 42950 4924 43258 4933
rect 42950 4922 42956 4924
rect 43012 4922 43036 4924
rect 43092 4922 43116 4924
rect 43172 4922 43196 4924
rect 43252 4922 43258 4924
rect 43012 4870 43014 4922
rect 43194 4870 43196 4922
rect 42950 4868 42956 4870
rect 43012 4868 43036 4870
rect 43092 4868 43116 4870
rect 43172 4868 43196 4870
rect 43252 4868 43258 4870
rect 42950 4859 43258 4868
rect 44640 4480 44692 4486
rect 44640 4422 44692 4428
rect 42950 3836 43258 3845
rect 42950 3834 42956 3836
rect 43012 3834 43036 3836
rect 43092 3834 43116 3836
rect 43172 3834 43196 3836
rect 43252 3834 43258 3836
rect 43012 3782 43014 3834
rect 43194 3782 43196 3834
rect 42950 3780 42956 3782
rect 43012 3780 43036 3782
rect 43092 3780 43116 3782
rect 43172 3780 43196 3782
rect 43252 3780 43258 3782
rect 42950 3771 43258 3780
rect 40040 3596 40092 3602
rect 40040 3538 40092 3544
rect 39856 3052 39908 3058
rect 39856 2994 39908 3000
rect 42950 2748 43258 2757
rect 42950 2746 42956 2748
rect 43012 2746 43036 2748
rect 43092 2746 43116 2748
rect 43172 2746 43196 2748
rect 43252 2746 43258 2748
rect 43012 2694 43014 2746
rect 43194 2694 43196 2746
rect 42950 2692 42956 2694
rect 43012 2692 43036 2694
rect 43092 2692 43116 2694
rect 43172 2692 43196 2694
rect 43252 2692 43258 2694
rect 42950 2683 43258 2692
rect 41328 2508 41380 2514
rect 41328 2450 41380 2456
rect 41340 800 41368 2450
rect 44652 2446 44680 4422
rect 45572 3738 45600 6054
rect 45756 5234 45784 7210
rect 46584 6322 46612 8842
rect 46768 8498 46796 9930
rect 47044 9586 47072 12106
rect 49146 12064 49202 12073
rect 47950 11996 48258 12005
rect 49146 11999 49202 12008
rect 47950 11994 47956 11996
rect 48012 11994 48036 11996
rect 48092 11994 48116 11996
rect 48172 11994 48196 11996
rect 48252 11994 48258 11996
rect 48012 11942 48014 11994
rect 48194 11942 48196 11994
rect 47950 11940 47956 11942
rect 48012 11940 48036 11942
rect 48092 11940 48116 11942
rect 48172 11940 48196 11942
rect 48252 11940 48258 11942
rect 47950 11931 48258 11940
rect 49160 11830 49188 11999
rect 49148 11824 49200 11830
rect 49148 11766 49200 11772
rect 49146 11656 49202 11665
rect 49146 11591 49202 11600
rect 49160 11218 49188 11591
rect 49238 11248 49294 11257
rect 49148 11212 49200 11218
rect 49238 11183 49294 11192
rect 49148 11154 49200 11160
rect 47950 10908 48258 10917
rect 47950 10906 47956 10908
rect 48012 10906 48036 10908
rect 48092 10906 48116 10908
rect 48172 10906 48196 10908
rect 48252 10906 48258 10908
rect 48012 10854 48014 10906
rect 48194 10854 48196 10906
rect 47950 10852 47956 10854
rect 48012 10852 48036 10854
rect 48092 10852 48116 10854
rect 48172 10852 48196 10854
rect 48252 10852 48258 10854
rect 47950 10843 48258 10852
rect 49146 10840 49202 10849
rect 49146 10775 49202 10784
rect 49160 10130 49188 10775
rect 49252 10742 49280 11183
rect 49240 10736 49292 10742
rect 49240 10678 49292 10684
rect 49330 10432 49386 10441
rect 49330 10367 49386 10376
rect 49148 10124 49200 10130
rect 49148 10066 49200 10072
rect 49238 10024 49294 10033
rect 47308 9988 47360 9994
rect 49238 9959 49294 9968
rect 47308 9930 47360 9936
rect 47320 9625 47348 9930
rect 47950 9820 48258 9829
rect 47950 9818 47956 9820
rect 48012 9818 48036 9820
rect 48092 9818 48116 9820
rect 48172 9818 48196 9820
rect 48252 9818 48258 9820
rect 48012 9766 48014 9818
rect 48194 9766 48196 9818
rect 47950 9764 47956 9766
rect 48012 9764 48036 9766
rect 48092 9764 48116 9766
rect 48172 9764 48196 9766
rect 48252 9764 48258 9766
rect 47950 9755 48258 9764
rect 47306 9616 47362 9625
rect 47032 9580 47084 9586
rect 47306 9551 47362 9560
rect 47032 9522 47084 9528
rect 49146 9208 49202 9217
rect 49146 9143 49202 9152
rect 47950 8732 48258 8741
rect 47950 8730 47956 8732
rect 48012 8730 48036 8732
rect 48092 8730 48116 8732
rect 48172 8730 48196 8732
rect 48252 8730 48258 8732
rect 48012 8678 48014 8730
rect 48194 8678 48196 8730
rect 47950 8676 47956 8678
rect 48012 8676 48036 8678
rect 48092 8676 48116 8678
rect 48172 8676 48196 8678
rect 48252 8676 48258 8678
rect 47950 8667 48258 8676
rect 47676 8628 47728 8634
rect 47676 8570 47728 8576
rect 46756 8492 46808 8498
rect 46756 8434 46808 8440
rect 46848 8424 46900 8430
rect 46848 8366 46900 8372
rect 46860 7993 46888 8366
rect 46846 7984 46902 7993
rect 46846 7919 46902 7928
rect 47584 7540 47636 7546
rect 47584 7482 47636 7488
rect 46940 6928 46992 6934
rect 46940 6870 46992 6876
rect 46572 6316 46624 6322
rect 46572 6258 46624 6264
rect 45836 5636 45888 5642
rect 45836 5578 45888 5584
rect 45744 5228 45796 5234
rect 45744 5170 45796 5176
rect 45560 3732 45612 3738
rect 45560 3674 45612 3680
rect 45560 3528 45612 3534
rect 45560 3470 45612 3476
rect 43444 2440 43496 2446
rect 43444 2382 43496 2388
rect 44640 2440 44692 2446
rect 44640 2382 44692 2388
rect 43456 800 43484 2382
rect 45572 800 45600 3470
rect 45848 3058 45876 5578
rect 46952 4146 46980 6870
rect 47032 6180 47084 6186
rect 47032 6122 47084 6128
rect 46940 4140 46992 4146
rect 46940 4082 46992 4088
rect 46664 4072 46716 4078
rect 46664 4014 46716 4020
rect 45836 3052 45888 3058
rect 45836 2994 45888 3000
rect 46676 1465 46704 4014
rect 47044 3534 47072 6122
rect 47216 5908 47268 5914
rect 47216 5850 47268 5856
rect 47124 4820 47176 4826
rect 47124 4762 47176 4768
rect 47032 3528 47084 3534
rect 47032 3470 47084 3476
rect 46756 2984 46808 2990
rect 46756 2926 46808 2932
rect 46848 2984 46900 2990
rect 46848 2926 46900 2932
rect 46768 1873 46796 2926
rect 46860 2689 46888 2926
rect 46846 2680 46902 2689
rect 46846 2615 46902 2624
rect 47136 2446 47164 4762
rect 47228 3058 47256 5850
rect 47596 4622 47624 7482
rect 47688 5710 47716 8570
rect 49160 8566 49188 9143
rect 49252 9042 49280 9959
rect 49344 9654 49372 10367
rect 49332 9648 49384 9654
rect 49332 9590 49384 9596
rect 49240 9036 49292 9042
rect 49240 8978 49292 8984
rect 49238 8800 49294 8809
rect 49238 8735 49294 8744
rect 49148 8560 49200 8566
rect 49148 8502 49200 8508
rect 47860 8356 47912 8362
rect 47860 8298 47912 8304
rect 47768 7200 47820 7206
rect 47768 7142 47820 7148
rect 47676 5704 47728 5710
rect 47676 5646 47728 5652
rect 47780 5234 47808 7142
rect 47872 6798 47900 8298
rect 49252 7954 49280 8735
rect 49330 8392 49386 8401
rect 49330 8327 49386 8336
rect 49240 7948 49292 7954
rect 49240 7890 49292 7896
rect 47950 7644 48258 7653
rect 47950 7642 47956 7644
rect 48012 7642 48036 7644
rect 48092 7642 48116 7644
rect 48172 7642 48196 7644
rect 48252 7642 48258 7644
rect 48012 7590 48014 7642
rect 48194 7590 48196 7642
rect 47950 7588 47956 7590
rect 48012 7588 48036 7590
rect 48092 7588 48116 7590
rect 48172 7588 48196 7590
rect 48252 7588 48258 7590
rect 47950 7579 48258 7588
rect 49146 7576 49202 7585
rect 49146 7511 49202 7520
rect 49160 6866 49188 7511
rect 49344 7478 49372 8327
rect 49332 7472 49384 7478
rect 49332 7414 49384 7420
rect 49238 7168 49294 7177
rect 49238 7103 49294 7112
rect 49148 6860 49200 6866
rect 49148 6802 49200 6808
rect 47860 6792 47912 6798
rect 47860 6734 47912 6740
rect 48872 6724 48924 6730
rect 48872 6666 48924 6672
rect 47950 6556 48258 6565
rect 47950 6554 47956 6556
rect 48012 6554 48036 6556
rect 48092 6554 48116 6556
rect 48172 6554 48196 6556
rect 48252 6554 48258 6556
rect 48012 6502 48014 6554
rect 48194 6502 48196 6554
rect 47950 6500 47956 6502
rect 48012 6500 48036 6502
rect 48092 6500 48116 6502
rect 48172 6500 48196 6502
rect 48252 6500 48258 6502
rect 47950 6491 48258 6500
rect 48884 6361 48912 6666
rect 49252 6390 49280 7103
rect 49422 6760 49478 6769
rect 49422 6695 49478 6704
rect 49240 6384 49292 6390
rect 48870 6352 48926 6361
rect 49240 6326 49292 6332
rect 48870 6287 48926 6296
rect 49146 5944 49202 5953
rect 49146 5879 49202 5888
rect 47950 5468 48258 5477
rect 47950 5466 47956 5468
rect 48012 5466 48036 5468
rect 48092 5466 48116 5468
rect 48172 5466 48196 5468
rect 48252 5466 48258 5468
rect 48012 5414 48014 5466
rect 48194 5414 48196 5466
rect 47950 5412 47956 5414
rect 48012 5412 48036 5414
rect 48092 5412 48116 5414
rect 48172 5412 48196 5414
rect 48252 5412 48258 5414
rect 47950 5403 48258 5412
rect 49160 5302 49188 5879
rect 49436 5778 49464 6695
rect 49424 5772 49476 5778
rect 49424 5714 49476 5720
rect 49422 5536 49478 5545
rect 49422 5471 49478 5480
rect 49148 5296 49200 5302
rect 49148 5238 49200 5244
rect 47768 5228 47820 5234
rect 47768 5170 47820 5176
rect 48320 5160 48372 5166
rect 48320 5102 48372 5108
rect 49330 5128 49386 5137
rect 48332 4729 48360 5102
rect 49330 5063 49386 5072
rect 48318 4720 48374 4729
rect 48318 4655 48374 4664
rect 47584 4616 47636 4622
rect 47584 4558 47636 4564
rect 47676 4548 47728 4554
rect 47676 4490 47728 4496
rect 47216 3052 47268 3058
rect 47216 2994 47268 3000
rect 47124 2440 47176 2446
rect 47124 2382 47176 2388
rect 46754 1864 46810 1873
rect 46754 1799 46810 1808
rect 46662 1456 46718 1465
rect 46662 1391 46718 1400
rect 47688 800 47716 4490
rect 47950 4380 48258 4389
rect 47950 4378 47956 4380
rect 48012 4378 48036 4380
rect 48092 4378 48116 4380
rect 48172 4378 48196 4380
rect 48252 4378 48258 4380
rect 48012 4326 48014 4378
rect 48194 4326 48196 4378
rect 47950 4324 47956 4326
rect 48012 4324 48036 4326
rect 48092 4324 48116 4326
rect 48172 4324 48196 4326
rect 48252 4324 48258 4326
rect 47950 4315 48258 4324
rect 49146 4312 49202 4321
rect 49146 4247 49202 4256
rect 49160 3602 49188 4247
rect 49344 4146 49372 5063
rect 49436 4690 49464 5471
rect 49424 4684 49476 4690
rect 49424 4626 49476 4632
rect 49792 4480 49844 4486
rect 49792 4422 49844 4428
rect 49332 4140 49384 4146
rect 49332 4082 49384 4088
rect 49238 3904 49294 3913
rect 49238 3839 49294 3848
rect 49148 3596 49200 3602
rect 49148 3538 49200 3544
rect 49146 3496 49202 3505
rect 48688 3460 48740 3466
rect 49146 3431 49202 3440
rect 48688 3402 48740 3408
rect 47950 3292 48258 3301
rect 47950 3290 47956 3292
rect 48012 3290 48036 3292
rect 48092 3290 48116 3292
rect 48172 3290 48196 3292
rect 48252 3290 48258 3292
rect 48012 3238 48014 3290
rect 48194 3238 48196 3290
rect 47950 3236 47956 3238
rect 48012 3236 48036 3238
rect 48092 3236 48116 3238
rect 48172 3236 48196 3238
rect 48252 3236 48258 3238
rect 47950 3227 48258 3236
rect 48700 3097 48728 3402
rect 48686 3088 48742 3097
rect 48686 3023 48742 3032
rect 49160 2514 49188 3431
rect 49252 3126 49280 3839
rect 49240 3120 49292 3126
rect 49240 3062 49292 3068
rect 49148 2508 49200 2514
rect 49148 2450 49200 2456
rect 48504 2372 48556 2378
rect 48504 2314 48556 2320
rect 48516 2281 48544 2314
rect 48502 2272 48558 2281
rect 47950 2204 48258 2213
rect 48502 2207 48558 2216
rect 47950 2202 47956 2204
rect 48012 2202 48036 2204
rect 48092 2202 48116 2204
rect 48172 2202 48196 2204
rect 48252 2202 48258 2204
rect 48012 2150 48014 2202
rect 48194 2150 48196 2202
rect 47950 2148 47956 2150
rect 48012 2148 48036 2150
rect 48092 2148 48116 2150
rect 48172 2148 48196 2150
rect 48252 2148 48258 2150
rect 47950 2139 48258 2148
rect 49804 800 49832 4422
rect 18156 734 18460 762
rect 20166 0 20222 800
rect 22282 0 22338 800
rect 24398 0 24454 800
rect 26514 0 26570 800
rect 28630 0 28686 800
rect 30746 0 30802 800
rect 32862 0 32918 800
rect 34978 0 35034 800
rect 37094 0 37150 800
rect 39210 0 39266 800
rect 41326 0 41382 800
rect 43442 0 43498 800
rect 45558 0 45614 800
rect 47674 0 47730 800
rect 49790 0 49846 800
<< via2 >>
rect 2778 24404 2834 24440
rect 2778 24384 2780 24404
rect 2780 24384 2832 24404
rect 2832 24384 2834 24404
rect 1306 20712 1362 20768
rect 3422 25608 3478 25664
rect 3330 25200 3386 25256
rect 3146 24792 3202 24848
rect 2956 24506 3012 24508
rect 3036 24506 3092 24508
rect 3116 24506 3172 24508
rect 3196 24506 3252 24508
rect 2956 24454 3002 24506
rect 3002 24454 3012 24506
rect 3036 24454 3066 24506
rect 3066 24454 3078 24506
rect 3078 24454 3092 24506
rect 3116 24454 3130 24506
rect 3130 24454 3142 24506
rect 3142 24454 3172 24506
rect 3196 24454 3206 24506
rect 3206 24454 3252 24506
rect 2956 24452 3012 24454
rect 3036 24452 3092 24454
rect 3116 24452 3172 24454
rect 3196 24452 3252 24454
rect 3698 23976 3754 24032
rect 3422 23588 3478 23624
rect 3422 23568 3424 23588
rect 3424 23568 3476 23588
rect 3476 23568 3478 23588
rect 2956 23418 3012 23420
rect 3036 23418 3092 23420
rect 3116 23418 3172 23420
rect 3196 23418 3252 23420
rect 2956 23366 3002 23418
rect 3002 23366 3012 23418
rect 3036 23366 3066 23418
rect 3066 23366 3078 23418
rect 3078 23366 3092 23418
rect 3116 23366 3130 23418
rect 3130 23366 3142 23418
rect 3142 23366 3172 23418
rect 3196 23366 3206 23418
rect 3206 23366 3252 23418
rect 2956 23364 3012 23366
rect 3036 23364 3092 23366
rect 3116 23364 3172 23366
rect 3196 23364 3252 23366
rect 3330 23160 3386 23216
rect 3422 22752 3478 22808
rect 2686 21528 2742 21584
rect 2778 21120 2834 21176
rect 2956 22330 3012 22332
rect 3036 22330 3092 22332
rect 3116 22330 3172 22332
rect 3196 22330 3252 22332
rect 2956 22278 3002 22330
rect 3002 22278 3012 22330
rect 3036 22278 3066 22330
rect 3066 22278 3078 22330
rect 3078 22278 3092 22330
rect 3116 22278 3130 22330
rect 3130 22278 3142 22330
rect 3142 22278 3172 22330
rect 3196 22278 3206 22330
rect 3206 22278 3252 22330
rect 2956 22276 3012 22278
rect 3036 22276 3092 22278
rect 3116 22276 3172 22278
rect 3196 22276 3252 22278
rect 2956 21242 3012 21244
rect 3036 21242 3092 21244
rect 3116 21242 3172 21244
rect 3196 21242 3252 21244
rect 2956 21190 3002 21242
rect 3002 21190 3012 21242
rect 3036 21190 3066 21242
rect 3066 21190 3078 21242
rect 3078 21190 3092 21242
rect 3116 21190 3130 21242
rect 3130 21190 3142 21242
rect 3142 21190 3172 21242
rect 3196 21190 3206 21242
rect 3206 21190 3252 21242
rect 2956 21188 3012 21190
rect 3036 21188 3092 21190
rect 3116 21188 3172 21190
rect 3196 21188 3252 21190
rect 2686 19488 2742 19544
rect 2956 20154 3012 20156
rect 3036 20154 3092 20156
rect 3116 20154 3172 20156
rect 3196 20154 3252 20156
rect 2956 20102 3002 20154
rect 3002 20102 3012 20154
rect 3036 20102 3066 20154
rect 3066 20102 3078 20154
rect 3078 20102 3092 20154
rect 3116 20102 3130 20154
rect 3130 20102 3142 20154
rect 3142 20102 3172 20154
rect 3196 20102 3206 20154
rect 3206 20102 3252 20154
rect 2956 20100 3012 20102
rect 3036 20100 3092 20102
rect 3116 20100 3172 20102
rect 3196 20100 3252 20102
rect 3330 19896 3386 19952
rect 2778 18808 2834 18864
rect 1766 18672 1822 18728
rect 2962 19216 3018 19272
rect 2956 19066 3012 19068
rect 3036 19066 3092 19068
rect 3116 19066 3172 19068
rect 3196 19066 3252 19068
rect 2956 19014 3002 19066
rect 3002 19014 3012 19066
rect 3036 19014 3066 19066
rect 3066 19014 3078 19066
rect 3078 19014 3092 19066
rect 3116 19014 3130 19066
rect 3130 19014 3142 19066
rect 3142 19014 3172 19066
rect 3196 19014 3206 19066
rect 3206 19014 3252 19066
rect 2956 19012 3012 19014
rect 3036 19012 3092 19014
rect 3116 19012 3172 19014
rect 3196 19012 3252 19014
rect 2870 18264 2926 18320
rect 3790 21936 3846 21992
rect 4250 22480 4306 22536
rect 3882 20340 3884 20360
rect 3884 20340 3936 20360
rect 3936 20340 3938 20360
rect 3882 20304 3938 20340
rect 2686 17856 2742 17912
rect 2956 17978 3012 17980
rect 3036 17978 3092 17980
rect 3116 17978 3172 17980
rect 3196 17978 3252 17980
rect 2956 17926 3002 17978
rect 3002 17926 3012 17978
rect 3036 17926 3066 17978
rect 3066 17926 3078 17978
rect 3078 17926 3092 17978
rect 3116 17926 3130 17978
rect 3130 17926 3142 17978
rect 3142 17926 3172 17978
rect 3196 17926 3206 17978
rect 3206 17926 3252 17978
rect 2956 17924 3012 17926
rect 3036 17924 3092 17926
rect 3116 17924 3172 17926
rect 3196 17924 3252 17926
rect 2778 17448 2834 17504
rect 1214 17040 1270 17096
rect 2956 16890 3012 16892
rect 3036 16890 3092 16892
rect 3116 16890 3172 16892
rect 3196 16890 3252 16892
rect 2956 16838 3002 16890
rect 3002 16838 3012 16890
rect 3036 16838 3066 16890
rect 3066 16838 3078 16890
rect 3078 16838 3092 16890
rect 3116 16838 3130 16890
rect 3130 16838 3142 16890
rect 3142 16838 3172 16890
rect 3196 16838 3206 16890
rect 3206 16838 3252 16890
rect 2956 16836 3012 16838
rect 3036 16836 3092 16838
rect 3116 16836 3172 16838
rect 3196 16836 3252 16838
rect 1306 16632 1362 16688
rect 1306 16224 1362 16280
rect 1306 15816 1362 15872
rect 2956 15802 3012 15804
rect 3036 15802 3092 15804
rect 3116 15802 3172 15804
rect 3196 15802 3252 15804
rect 2956 15750 3002 15802
rect 3002 15750 3012 15802
rect 3036 15750 3066 15802
rect 3066 15750 3078 15802
rect 3078 15750 3092 15802
rect 3116 15750 3130 15802
rect 3130 15750 3142 15802
rect 3142 15750 3172 15802
rect 3196 15750 3206 15802
rect 3206 15750 3252 15802
rect 2956 15748 3012 15750
rect 3036 15748 3092 15750
rect 3116 15748 3172 15750
rect 3196 15748 3252 15750
rect 1306 15408 1362 15464
rect 1306 15000 1362 15056
rect 1306 14592 1362 14648
rect 1306 14184 1362 14240
rect 938 12960 994 13016
rect 1306 12552 1362 12608
rect 1030 12144 1086 12200
rect 938 11736 994 11792
rect 938 11328 994 11384
rect 1582 10920 1638 10976
rect 938 10512 994 10568
rect 1214 10104 1270 10160
rect 938 9696 994 9752
rect 1766 9444 1822 9480
rect 1766 9424 1768 9444
rect 1768 9424 1820 9444
rect 1820 9424 1822 9444
rect 938 9288 994 9344
rect 938 8916 940 8936
rect 940 8916 992 8936
rect 992 8916 994 8936
rect 938 8880 994 8916
rect 1214 8472 1270 8528
rect 1582 8064 1638 8120
rect 938 7656 994 7712
rect 938 7248 994 7304
rect 938 6840 994 6896
rect 2956 14714 3012 14716
rect 3036 14714 3092 14716
rect 3116 14714 3172 14716
rect 3196 14714 3252 14716
rect 2956 14662 3002 14714
rect 3002 14662 3012 14714
rect 3036 14662 3066 14714
rect 3066 14662 3078 14714
rect 3078 14662 3092 14714
rect 3116 14662 3130 14714
rect 3130 14662 3142 14714
rect 3142 14662 3172 14714
rect 3196 14662 3206 14714
rect 3206 14662 3252 14714
rect 2956 14660 3012 14662
rect 3036 14660 3092 14662
rect 3116 14660 3172 14662
rect 3196 14660 3252 14662
rect 2778 13776 2834 13832
rect 2956 13626 3012 13628
rect 3036 13626 3092 13628
rect 3116 13626 3172 13628
rect 3196 13626 3252 13628
rect 2956 13574 3002 13626
rect 3002 13574 3012 13626
rect 3036 13574 3066 13626
rect 3066 13574 3078 13626
rect 3078 13574 3092 13626
rect 3116 13574 3130 13626
rect 3130 13574 3142 13626
rect 3142 13574 3172 13626
rect 3196 13574 3206 13626
rect 3206 13574 3252 13626
rect 2956 13572 3012 13574
rect 3036 13572 3092 13574
rect 3116 13572 3172 13574
rect 3196 13572 3252 13574
rect 3514 13368 3570 13424
rect 2956 12538 3012 12540
rect 3036 12538 3092 12540
rect 3116 12538 3172 12540
rect 3196 12538 3252 12540
rect 2956 12486 3002 12538
rect 3002 12486 3012 12538
rect 3036 12486 3066 12538
rect 3066 12486 3078 12538
rect 3078 12486 3092 12538
rect 3116 12486 3130 12538
rect 3130 12486 3142 12538
rect 3142 12486 3172 12538
rect 3196 12486 3206 12538
rect 3206 12486 3252 12538
rect 2956 12484 3012 12486
rect 3036 12484 3092 12486
rect 3116 12484 3172 12486
rect 3196 12484 3252 12486
rect 7470 24656 7526 24712
rect 7956 23962 8012 23964
rect 8036 23962 8092 23964
rect 8116 23962 8172 23964
rect 8196 23962 8252 23964
rect 7956 23910 8002 23962
rect 8002 23910 8012 23962
rect 8036 23910 8066 23962
rect 8066 23910 8078 23962
rect 8078 23910 8092 23962
rect 8116 23910 8130 23962
rect 8130 23910 8142 23962
rect 8142 23910 8172 23962
rect 8196 23910 8206 23962
rect 8206 23910 8252 23962
rect 7956 23908 8012 23910
rect 8036 23908 8092 23910
rect 8116 23908 8172 23910
rect 8196 23908 8252 23910
rect 7956 22874 8012 22876
rect 8036 22874 8092 22876
rect 8116 22874 8172 22876
rect 8196 22874 8252 22876
rect 7956 22822 8002 22874
rect 8002 22822 8012 22874
rect 8036 22822 8066 22874
rect 8066 22822 8078 22874
rect 8078 22822 8092 22874
rect 8116 22822 8130 22874
rect 8130 22822 8142 22874
rect 8142 22822 8172 22874
rect 8196 22822 8206 22874
rect 8206 22822 8252 22874
rect 7956 22820 8012 22822
rect 8036 22820 8092 22822
rect 8116 22820 8172 22822
rect 8196 22820 8252 22822
rect 7956 21786 8012 21788
rect 8036 21786 8092 21788
rect 8116 21786 8172 21788
rect 8196 21786 8252 21788
rect 7956 21734 8002 21786
rect 8002 21734 8012 21786
rect 8036 21734 8066 21786
rect 8066 21734 8078 21786
rect 8078 21734 8092 21786
rect 8116 21734 8130 21786
rect 8130 21734 8142 21786
rect 8142 21734 8172 21786
rect 8196 21734 8206 21786
rect 8206 21734 8252 21786
rect 7956 21732 8012 21734
rect 8036 21732 8092 21734
rect 8116 21732 8172 21734
rect 8196 21732 8252 21734
rect 7956 20698 8012 20700
rect 8036 20698 8092 20700
rect 8116 20698 8172 20700
rect 8196 20698 8252 20700
rect 7956 20646 8002 20698
rect 8002 20646 8012 20698
rect 8036 20646 8066 20698
rect 8066 20646 8078 20698
rect 8078 20646 8092 20698
rect 8116 20646 8130 20698
rect 8130 20646 8142 20698
rect 8142 20646 8172 20698
rect 8196 20646 8206 20698
rect 8206 20646 8252 20698
rect 7956 20644 8012 20646
rect 8036 20644 8092 20646
rect 8116 20644 8172 20646
rect 8196 20644 8252 20646
rect 7956 19610 8012 19612
rect 8036 19610 8092 19612
rect 8116 19610 8172 19612
rect 8196 19610 8252 19612
rect 7956 19558 8002 19610
rect 8002 19558 8012 19610
rect 8036 19558 8066 19610
rect 8066 19558 8078 19610
rect 8078 19558 8092 19610
rect 8116 19558 8130 19610
rect 8130 19558 8142 19610
rect 8142 19558 8172 19610
rect 8196 19558 8206 19610
rect 8206 19558 8252 19610
rect 7956 19556 8012 19558
rect 8036 19556 8092 19558
rect 8116 19556 8172 19558
rect 8196 19556 8252 19558
rect 7956 18522 8012 18524
rect 8036 18522 8092 18524
rect 8116 18522 8172 18524
rect 8196 18522 8252 18524
rect 7956 18470 8002 18522
rect 8002 18470 8012 18522
rect 8036 18470 8066 18522
rect 8066 18470 8078 18522
rect 8078 18470 8092 18522
rect 8116 18470 8130 18522
rect 8130 18470 8142 18522
rect 8142 18470 8172 18522
rect 8196 18470 8206 18522
rect 8206 18470 8252 18522
rect 7956 18468 8012 18470
rect 8036 18468 8092 18470
rect 8116 18468 8172 18470
rect 8196 18468 8252 18470
rect 7956 17434 8012 17436
rect 8036 17434 8092 17436
rect 8116 17434 8172 17436
rect 8196 17434 8252 17436
rect 7956 17382 8002 17434
rect 8002 17382 8012 17434
rect 8036 17382 8066 17434
rect 8066 17382 8078 17434
rect 8078 17382 8092 17434
rect 8116 17382 8130 17434
rect 8130 17382 8142 17434
rect 8142 17382 8172 17434
rect 8196 17382 8206 17434
rect 8206 17382 8252 17434
rect 7956 17380 8012 17382
rect 8036 17380 8092 17382
rect 8116 17380 8172 17382
rect 8196 17380 8252 17382
rect 7956 16346 8012 16348
rect 8036 16346 8092 16348
rect 8116 16346 8172 16348
rect 8196 16346 8252 16348
rect 7956 16294 8002 16346
rect 8002 16294 8012 16346
rect 8036 16294 8066 16346
rect 8066 16294 8078 16346
rect 8078 16294 8092 16346
rect 8116 16294 8130 16346
rect 8130 16294 8142 16346
rect 8142 16294 8172 16346
rect 8196 16294 8206 16346
rect 8206 16294 8252 16346
rect 7956 16292 8012 16294
rect 8036 16292 8092 16294
rect 8116 16292 8172 16294
rect 8196 16292 8252 16294
rect 7956 15258 8012 15260
rect 8036 15258 8092 15260
rect 8116 15258 8172 15260
rect 8196 15258 8252 15260
rect 7956 15206 8002 15258
rect 8002 15206 8012 15258
rect 8036 15206 8066 15258
rect 8066 15206 8078 15258
rect 8078 15206 8092 15258
rect 8116 15206 8130 15258
rect 8130 15206 8142 15258
rect 8142 15206 8172 15258
rect 8196 15206 8206 15258
rect 8206 15206 8252 15258
rect 7956 15204 8012 15206
rect 8036 15204 8092 15206
rect 8116 15204 8172 15206
rect 8196 15204 8252 15206
rect 7956 14170 8012 14172
rect 8036 14170 8092 14172
rect 8116 14170 8172 14172
rect 8196 14170 8252 14172
rect 7956 14118 8002 14170
rect 8002 14118 8012 14170
rect 8036 14118 8066 14170
rect 8066 14118 8078 14170
rect 8078 14118 8092 14170
rect 8116 14118 8130 14170
rect 8130 14118 8142 14170
rect 8142 14118 8172 14170
rect 8196 14118 8206 14170
rect 8206 14118 8252 14170
rect 7956 14116 8012 14118
rect 8036 14116 8092 14118
rect 8116 14116 8172 14118
rect 8196 14116 8252 14118
rect 12070 22616 12126 22672
rect 12956 24506 13012 24508
rect 13036 24506 13092 24508
rect 13116 24506 13172 24508
rect 13196 24506 13252 24508
rect 12956 24454 13002 24506
rect 13002 24454 13012 24506
rect 13036 24454 13066 24506
rect 13066 24454 13078 24506
rect 13078 24454 13092 24506
rect 13116 24454 13130 24506
rect 13130 24454 13142 24506
rect 13142 24454 13172 24506
rect 13196 24454 13206 24506
rect 13206 24454 13252 24506
rect 12956 24452 13012 24454
rect 13036 24452 13092 24454
rect 13116 24452 13172 24454
rect 13196 24452 13252 24454
rect 12070 21972 12072 21992
rect 12072 21972 12124 21992
rect 12124 21972 12126 21992
rect 11150 20984 11206 21040
rect 10138 14184 10194 14240
rect 7956 13082 8012 13084
rect 8036 13082 8092 13084
rect 8116 13082 8172 13084
rect 8196 13082 8252 13084
rect 7956 13030 8002 13082
rect 8002 13030 8012 13082
rect 8036 13030 8066 13082
rect 8066 13030 8078 13082
rect 8078 13030 8092 13082
rect 8116 13030 8130 13082
rect 8130 13030 8142 13082
rect 8142 13030 8172 13082
rect 8196 13030 8206 13082
rect 8206 13030 8252 13082
rect 7956 13028 8012 13030
rect 8036 13028 8092 13030
rect 8116 13028 8172 13030
rect 8196 13028 8252 13030
rect 11702 20712 11758 20768
rect 10322 13232 10378 13288
rect 11334 15952 11390 16008
rect 11150 14340 11206 14376
rect 11150 14320 11152 14340
rect 11152 14320 11204 14340
rect 11204 14320 11206 14340
rect 12070 21936 12126 21972
rect 12438 20848 12494 20904
rect 12070 17720 12126 17776
rect 11886 16088 11942 16144
rect 12956 23418 13012 23420
rect 13036 23418 13092 23420
rect 13116 23418 13172 23420
rect 13196 23418 13252 23420
rect 12956 23366 13002 23418
rect 13002 23366 13012 23418
rect 13036 23366 13066 23418
rect 13066 23366 13078 23418
rect 13078 23366 13092 23418
rect 13116 23366 13130 23418
rect 13130 23366 13142 23418
rect 13142 23366 13172 23418
rect 13196 23366 13206 23418
rect 13206 23366 13252 23418
rect 12956 23364 13012 23366
rect 13036 23364 13092 23366
rect 13116 23364 13172 23366
rect 13196 23364 13252 23366
rect 12956 22330 13012 22332
rect 13036 22330 13092 22332
rect 13116 22330 13172 22332
rect 13196 22330 13252 22332
rect 12956 22278 13002 22330
rect 13002 22278 13012 22330
rect 13036 22278 13066 22330
rect 13066 22278 13078 22330
rect 13078 22278 13092 22330
rect 13116 22278 13130 22330
rect 13130 22278 13142 22330
rect 13142 22278 13172 22330
rect 13196 22278 13206 22330
rect 13206 22278 13252 22330
rect 12956 22276 13012 22278
rect 13036 22276 13092 22278
rect 13116 22276 13172 22278
rect 13196 22276 13252 22278
rect 12714 19236 12770 19272
rect 12714 19216 12716 19236
rect 12716 19216 12768 19236
rect 12768 19216 12770 19236
rect 12956 21242 13012 21244
rect 13036 21242 13092 21244
rect 13116 21242 13172 21244
rect 13196 21242 13252 21244
rect 12956 21190 13002 21242
rect 13002 21190 13012 21242
rect 13036 21190 13066 21242
rect 13066 21190 13078 21242
rect 13078 21190 13092 21242
rect 13116 21190 13130 21242
rect 13130 21190 13142 21242
rect 13142 21190 13172 21242
rect 13196 21190 13206 21242
rect 13206 21190 13252 21242
rect 12956 21188 13012 21190
rect 13036 21188 13092 21190
rect 13116 21188 13172 21190
rect 13196 21188 13252 21190
rect 12956 20154 13012 20156
rect 13036 20154 13092 20156
rect 13116 20154 13172 20156
rect 13196 20154 13252 20156
rect 12956 20102 13002 20154
rect 13002 20102 13012 20154
rect 13036 20102 13066 20154
rect 13066 20102 13078 20154
rect 13078 20102 13092 20154
rect 13116 20102 13130 20154
rect 13130 20102 13142 20154
rect 13142 20102 13172 20154
rect 13196 20102 13206 20154
rect 13206 20102 13252 20154
rect 12956 20100 13012 20102
rect 13036 20100 13092 20102
rect 13116 20100 13172 20102
rect 13196 20100 13252 20102
rect 12956 19066 13012 19068
rect 13036 19066 13092 19068
rect 13116 19066 13172 19068
rect 13196 19066 13252 19068
rect 12956 19014 13002 19066
rect 13002 19014 13012 19066
rect 13036 19014 13066 19066
rect 13066 19014 13078 19066
rect 13078 19014 13092 19066
rect 13116 19014 13130 19066
rect 13130 19014 13142 19066
rect 13142 19014 13172 19066
rect 13196 19014 13206 19066
rect 13206 19014 13252 19066
rect 12956 19012 13012 19014
rect 13036 19012 13092 19014
rect 13116 19012 13172 19014
rect 13196 19012 13252 19014
rect 13634 20460 13690 20496
rect 13634 20440 13636 20460
rect 13636 20440 13688 20460
rect 13688 20440 13690 20460
rect 12956 17978 13012 17980
rect 13036 17978 13092 17980
rect 13116 17978 13172 17980
rect 13196 17978 13252 17980
rect 12956 17926 13002 17978
rect 13002 17926 13012 17978
rect 13036 17926 13066 17978
rect 13066 17926 13078 17978
rect 13078 17926 13092 17978
rect 13116 17926 13130 17978
rect 13130 17926 13142 17978
rect 13142 17926 13172 17978
rect 13196 17926 13206 17978
rect 13206 17926 13252 17978
rect 12956 17924 13012 17926
rect 13036 17924 13092 17926
rect 13116 17924 13172 17926
rect 13196 17924 13252 17926
rect 12956 16890 13012 16892
rect 13036 16890 13092 16892
rect 13116 16890 13172 16892
rect 13196 16890 13252 16892
rect 12956 16838 13002 16890
rect 13002 16838 13012 16890
rect 13036 16838 13066 16890
rect 13066 16838 13078 16890
rect 13078 16838 13092 16890
rect 13116 16838 13130 16890
rect 13130 16838 13142 16890
rect 13142 16838 13172 16890
rect 13196 16838 13206 16890
rect 13206 16838 13252 16890
rect 12956 16836 13012 16838
rect 13036 16836 13092 16838
rect 13116 16836 13172 16838
rect 13196 16836 13252 16838
rect 11334 12280 11390 12336
rect 11058 12144 11114 12200
rect 7956 11994 8012 11996
rect 8036 11994 8092 11996
rect 8116 11994 8172 11996
rect 8196 11994 8252 11996
rect 7956 11942 8002 11994
rect 8002 11942 8012 11994
rect 8036 11942 8066 11994
rect 8066 11942 8078 11994
rect 8078 11942 8092 11994
rect 8116 11942 8130 11994
rect 8130 11942 8142 11994
rect 8142 11942 8172 11994
rect 8196 11942 8206 11994
rect 8206 11942 8252 11994
rect 7956 11940 8012 11942
rect 8036 11940 8092 11942
rect 8116 11940 8172 11942
rect 8196 11940 8252 11942
rect 2956 11450 3012 11452
rect 3036 11450 3092 11452
rect 3116 11450 3172 11452
rect 3196 11450 3252 11452
rect 2956 11398 3002 11450
rect 3002 11398 3012 11450
rect 3036 11398 3066 11450
rect 3066 11398 3078 11450
rect 3078 11398 3092 11450
rect 3116 11398 3130 11450
rect 3130 11398 3142 11450
rect 3142 11398 3172 11450
rect 3196 11398 3206 11450
rect 3206 11398 3252 11450
rect 2956 11396 3012 11398
rect 3036 11396 3092 11398
rect 3116 11396 3172 11398
rect 3196 11396 3252 11398
rect 7956 10906 8012 10908
rect 8036 10906 8092 10908
rect 8116 10906 8172 10908
rect 8196 10906 8252 10908
rect 7956 10854 8002 10906
rect 8002 10854 8012 10906
rect 8036 10854 8066 10906
rect 8066 10854 8078 10906
rect 8078 10854 8092 10906
rect 8116 10854 8130 10906
rect 8130 10854 8142 10906
rect 8142 10854 8172 10906
rect 8196 10854 8206 10906
rect 8206 10854 8252 10906
rect 7956 10852 8012 10854
rect 8036 10852 8092 10854
rect 8116 10852 8172 10854
rect 8196 10852 8252 10854
rect 2956 10362 3012 10364
rect 3036 10362 3092 10364
rect 3116 10362 3172 10364
rect 3196 10362 3252 10364
rect 2956 10310 3002 10362
rect 3002 10310 3012 10362
rect 3036 10310 3066 10362
rect 3066 10310 3078 10362
rect 3078 10310 3092 10362
rect 3116 10310 3130 10362
rect 3130 10310 3142 10362
rect 3142 10310 3172 10362
rect 3196 10310 3206 10362
rect 3206 10310 3252 10362
rect 2956 10308 3012 10310
rect 3036 10308 3092 10310
rect 3116 10308 3172 10310
rect 3196 10308 3252 10310
rect 7956 9818 8012 9820
rect 8036 9818 8092 9820
rect 8116 9818 8172 9820
rect 8196 9818 8252 9820
rect 7956 9766 8002 9818
rect 8002 9766 8012 9818
rect 8036 9766 8066 9818
rect 8066 9766 8078 9818
rect 8078 9766 8092 9818
rect 8116 9766 8130 9818
rect 8130 9766 8142 9818
rect 8142 9766 8172 9818
rect 8196 9766 8206 9818
rect 8206 9766 8252 9818
rect 7956 9764 8012 9766
rect 8036 9764 8092 9766
rect 8116 9764 8172 9766
rect 8196 9764 8252 9766
rect 13726 19216 13782 19272
rect 14186 17992 14242 18048
rect 12956 15802 13012 15804
rect 13036 15802 13092 15804
rect 13116 15802 13172 15804
rect 13196 15802 13252 15804
rect 12956 15750 13002 15802
rect 13002 15750 13012 15802
rect 13036 15750 13066 15802
rect 13066 15750 13078 15802
rect 13078 15750 13092 15802
rect 13116 15750 13130 15802
rect 13130 15750 13142 15802
rect 13142 15750 13172 15802
rect 13196 15750 13206 15802
rect 13206 15750 13252 15802
rect 12956 15748 13012 15750
rect 13036 15748 13092 15750
rect 13116 15748 13172 15750
rect 13196 15748 13252 15750
rect 13174 15020 13230 15056
rect 13174 15000 13176 15020
rect 13176 15000 13228 15020
rect 13228 15000 13230 15020
rect 12956 14714 13012 14716
rect 13036 14714 13092 14716
rect 13116 14714 13172 14716
rect 13196 14714 13252 14716
rect 12956 14662 13002 14714
rect 13002 14662 13012 14714
rect 13036 14662 13066 14714
rect 13066 14662 13078 14714
rect 13078 14662 13092 14714
rect 13116 14662 13130 14714
rect 13130 14662 13142 14714
rect 13142 14662 13172 14714
rect 13196 14662 13206 14714
rect 13206 14662 13252 14714
rect 12956 14660 13012 14662
rect 13036 14660 13092 14662
rect 13116 14660 13172 14662
rect 13196 14660 13252 14662
rect 12956 13626 13012 13628
rect 13036 13626 13092 13628
rect 13116 13626 13172 13628
rect 13196 13626 13252 13628
rect 12956 13574 13002 13626
rect 13002 13574 13012 13626
rect 13036 13574 13066 13626
rect 13066 13574 13078 13626
rect 13078 13574 13092 13626
rect 13116 13574 13130 13626
rect 13130 13574 13142 13626
rect 13142 13574 13172 13626
rect 13196 13574 13206 13626
rect 13206 13574 13252 13626
rect 12956 13572 13012 13574
rect 13036 13572 13092 13574
rect 13116 13572 13172 13574
rect 13196 13572 13252 13574
rect 12956 12538 13012 12540
rect 13036 12538 13092 12540
rect 13116 12538 13172 12540
rect 13196 12538 13252 12540
rect 12956 12486 13002 12538
rect 13002 12486 13012 12538
rect 13036 12486 13066 12538
rect 13066 12486 13078 12538
rect 13078 12486 13092 12538
rect 13116 12486 13130 12538
rect 13130 12486 13142 12538
rect 13142 12486 13172 12538
rect 13196 12486 13206 12538
rect 13206 12486 13252 12538
rect 12956 12484 13012 12486
rect 13036 12484 13092 12486
rect 13116 12484 13172 12486
rect 13196 12484 13252 12486
rect 14646 19896 14702 19952
rect 14186 17212 14188 17232
rect 14188 17212 14240 17232
rect 14240 17212 14242 17232
rect 14186 17176 14242 17212
rect 14370 16124 14372 16144
rect 14372 16124 14424 16144
rect 14424 16124 14426 16144
rect 14370 16088 14426 16124
rect 14002 14864 14058 14920
rect 13542 12552 13598 12608
rect 12956 11450 13012 11452
rect 13036 11450 13092 11452
rect 13116 11450 13172 11452
rect 13196 11450 13252 11452
rect 12956 11398 13002 11450
rect 13002 11398 13012 11450
rect 13036 11398 13066 11450
rect 13066 11398 13078 11450
rect 13078 11398 13092 11450
rect 13116 11398 13130 11450
rect 13130 11398 13142 11450
rect 13142 11398 13172 11450
rect 13196 11398 13206 11450
rect 13206 11398 13252 11450
rect 12956 11396 13012 11398
rect 13036 11396 13092 11398
rect 13116 11396 13172 11398
rect 13196 11396 13252 11398
rect 12956 10362 13012 10364
rect 13036 10362 13092 10364
rect 13116 10362 13172 10364
rect 13196 10362 13252 10364
rect 12956 10310 13002 10362
rect 13002 10310 13012 10362
rect 13036 10310 13066 10362
rect 13066 10310 13078 10362
rect 13078 10310 13092 10362
rect 13116 10310 13130 10362
rect 13130 10310 13142 10362
rect 13142 10310 13172 10362
rect 13196 10310 13206 10362
rect 13206 10310 13252 10362
rect 12956 10308 13012 10310
rect 13036 10308 13092 10310
rect 13116 10308 13172 10310
rect 13196 10308 13252 10310
rect 13266 10004 13268 10024
rect 13268 10004 13320 10024
rect 13320 10004 13322 10024
rect 13266 9968 13322 10004
rect 2956 9274 3012 9276
rect 3036 9274 3092 9276
rect 3116 9274 3172 9276
rect 3196 9274 3252 9276
rect 2956 9222 3002 9274
rect 3002 9222 3012 9274
rect 3036 9222 3066 9274
rect 3066 9222 3078 9274
rect 3078 9222 3092 9274
rect 3116 9222 3130 9274
rect 3130 9222 3142 9274
rect 3142 9222 3172 9274
rect 3196 9222 3206 9274
rect 3206 9222 3252 9274
rect 2956 9220 3012 9222
rect 3036 9220 3092 9222
rect 3116 9220 3172 9222
rect 3196 9220 3252 9222
rect 7956 8730 8012 8732
rect 8036 8730 8092 8732
rect 8116 8730 8172 8732
rect 8196 8730 8252 8732
rect 7956 8678 8002 8730
rect 8002 8678 8012 8730
rect 8036 8678 8066 8730
rect 8066 8678 8078 8730
rect 8078 8678 8092 8730
rect 8116 8678 8130 8730
rect 8130 8678 8142 8730
rect 8142 8678 8172 8730
rect 8196 8678 8206 8730
rect 8206 8678 8252 8730
rect 7956 8676 8012 8678
rect 8036 8676 8092 8678
rect 8116 8676 8172 8678
rect 8196 8676 8252 8678
rect 2956 8186 3012 8188
rect 3036 8186 3092 8188
rect 3116 8186 3172 8188
rect 3196 8186 3252 8188
rect 2956 8134 3002 8186
rect 3002 8134 3012 8186
rect 3036 8134 3066 8186
rect 3066 8134 3078 8186
rect 3078 8134 3092 8186
rect 3116 8134 3130 8186
rect 3130 8134 3142 8186
rect 3142 8134 3172 8186
rect 3196 8134 3206 8186
rect 3206 8134 3252 8186
rect 2956 8132 3012 8134
rect 3036 8132 3092 8134
rect 3116 8132 3172 8134
rect 3196 8132 3252 8134
rect 12956 9274 13012 9276
rect 13036 9274 13092 9276
rect 13116 9274 13172 9276
rect 13196 9274 13252 9276
rect 12956 9222 13002 9274
rect 13002 9222 13012 9274
rect 13036 9222 13066 9274
rect 13066 9222 13078 9274
rect 13078 9222 13092 9274
rect 13116 9222 13130 9274
rect 13130 9222 13142 9274
rect 13142 9222 13172 9274
rect 13196 9222 13206 9274
rect 13206 9222 13252 9274
rect 12956 9220 13012 9222
rect 13036 9220 13092 9222
rect 13116 9220 13172 9222
rect 13196 9220 13252 9222
rect 12956 8186 13012 8188
rect 13036 8186 13092 8188
rect 13116 8186 13172 8188
rect 13196 8186 13252 8188
rect 12956 8134 13002 8186
rect 13002 8134 13012 8186
rect 13036 8134 13066 8186
rect 13066 8134 13078 8186
rect 13078 8134 13092 8186
rect 13116 8134 13130 8186
rect 13130 8134 13142 8186
rect 13142 8134 13172 8186
rect 13196 8134 13206 8186
rect 13206 8134 13252 8186
rect 12956 8132 13012 8134
rect 13036 8132 13092 8134
rect 13116 8132 13172 8134
rect 13196 8132 13252 8134
rect 7956 7642 8012 7644
rect 8036 7642 8092 7644
rect 8116 7642 8172 7644
rect 8196 7642 8252 7644
rect 7956 7590 8002 7642
rect 8002 7590 8012 7642
rect 8036 7590 8066 7642
rect 8066 7590 8078 7642
rect 8078 7590 8092 7642
rect 8116 7590 8130 7642
rect 8130 7590 8142 7642
rect 8142 7590 8172 7642
rect 8196 7590 8206 7642
rect 8206 7590 8252 7642
rect 7956 7588 8012 7590
rect 8036 7588 8092 7590
rect 8116 7588 8172 7590
rect 8196 7588 8252 7590
rect 2956 7098 3012 7100
rect 3036 7098 3092 7100
rect 3116 7098 3172 7100
rect 3196 7098 3252 7100
rect 2956 7046 3002 7098
rect 3002 7046 3012 7098
rect 3036 7046 3066 7098
rect 3066 7046 3078 7098
rect 3078 7046 3092 7098
rect 3116 7046 3130 7098
rect 3130 7046 3142 7098
rect 3142 7046 3172 7098
rect 3196 7046 3206 7098
rect 3206 7046 3252 7098
rect 2956 7044 3012 7046
rect 3036 7044 3092 7046
rect 3116 7044 3172 7046
rect 3196 7044 3252 7046
rect 12956 7098 13012 7100
rect 13036 7098 13092 7100
rect 13116 7098 13172 7100
rect 13196 7098 13252 7100
rect 12956 7046 13002 7098
rect 13002 7046 13012 7098
rect 13036 7046 13066 7098
rect 13066 7046 13078 7098
rect 13078 7046 13092 7098
rect 13116 7046 13130 7098
rect 13130 7046 13142 7098
rect 13142 7046 13172 7098
rect 13196 7046 13206 7098
rect 13206 7046 13252 7098
rect 12956 7044 13012 7046
rect 13036 7044 13092 7046
rect 13116 7044 13172 7046
rect 13196 7044 13252 7046
rect 7956 6554 8012 6556
rect 8036 6554 8092 6556
rect 8116 6554 8172 6556
rect 8196 6554 8252 6556
rect 7956 6502 8002 6554
rect 8002 6502 8012 6554
rect 8036 6502 8066 6554
rect 8066 6502 8078 6554
rect 8078 6502 8092 6554
rect 8116 6502 8130 6554
rect 8130 6502 8142 6554
rect 8142 6502 8172 6554
rect 8196 6502 8206 6554
rect 8206 6502 8252 6554
rect 7956 6500 8012 6502
rect 8036 6500 8092 6502
rect 8116 6500 8172 6502
rect 8196 6500 8252 6502
rect 1306 6432 1362 6488
rect 938 6024 994 6080
rect 938 5652 940 5672
rect 940 5652 992 5672
rect 992 5652 994 5672
rect 938 5616 994 5652
rect 938 4800 994 4856
rect 938 4392 994 4448
rect 2956 6010 3012 6012
rect 3036 6010 3092 6012
rect 3116 6010 3172 6012
rect 3196 6010 3252 6012
rect 2956 5958 3002 6010
rect 3002 5958 3012 6010
rect 3036 5958 3066 6010
rect 3066 5958 3078 6010
rect 3078 5958 3092 6010
rect 3116 5958 3130 6010
rect 3130 5958 3142 6010
rect 3142 5958 3172 6010
rect 3196 5958 3206 6010
rect 3206 5958 3252 6010
rect 2956 5956 3012 5958
rect 3036 5956 3092 5958
rect 3116 5956 3172 5958
rect 3196 5956 3252 5958
rect 12956 6010 13012 6012
rect 13036 6010 13092 6012
rect 13116 6010 13172 6012
rect 13196 6010 13252 6012
rect 12956 5958 13002 6010
rect 13002 5958 13012 6010
rect 13036 5958 13066 6010
rect 13066 5958 13078 6010
rect 13078 5958 13092 6010
rect 13116 5958 13130 6010
rect 13130 5958 13142 6010
rect 13142 5958 13172 6010
rect 13196 5958 13206 6010
rect 13206 5958 13252 6010
rect 12956 5956 13012 5958
rect 13036 5956 13092 5958
rect 13116 5956 13172 5958
rect 13196 5956 13252 5958
rect 7956 5466 8012 5468
rect 8036 5466 8092 5468
rect 8116 5466 8172 5468
rect 8196 5466 8252 5468
rect 7956 5414 8002 5466
rect 8002 5414 8012 5466
rect 8036 5414 8066 5466
rect 8066 5414 8078 5466
rect 8078 5414 8092 5466
rect 8116 5414 8130 5466
rect 8130 5414 8142 5466
rect 8142 5414 8172 5466
rect 8196 5414 8206 5466
rect 8206 5414 8252 5466
rect 7956 5412 8012 5414
rect 8036 5412 8092 5414
rect 8116 5412 8172 5414
rect 8196 5412 8252 5414
rect 2318 5208 2374 5264
rect 2956 4922 3012 4924
rect 3036 4922 3092 4924
rect 3116 4922 3172 4924
rect 3196 4922 3252 4924
rect 2956 4870 3002 4922
rect 3002 4870 3012 4922
rect 3036 4870 3066 4922
rect 3066 4870 3078 4922
rect 3078 4870 3092 4922
rect 3116 4870 3130 4922
rect 3130 4870 3142 4922
rect 3142 4870 3172 4922
rect 3196 4870 3206 4922
rect 3206 4870 3252 4922
rect 2956 4868 3012 4870
rect 3036 4868 3092 4870
rect 3116 4868 3172 4870
rect 3196 4868 3252 4870
rect 12956 4922 13012 4924
rect 13036 4922 13092 4924
rect 13116 4922 13172 4924
rect 13196 4922 13252 4924
rect 12956 4870 13002 4922
rect 13002 4870 13012 4922
rect 13036 4870 13066 4922
rect 13066 4870 13078 4922
rect 13078 4870 13092 4922
rect 13116 4870 13130 4922
rect 13130 4870 13142 4922
rect 13142 4870 13172 4922
rect 13196 4870 13206 4922
rect 13206 4870 13252 4922
rect 12956 4868 13012 4870
rect 13036 4868 13092 4870
rect 13116 4868 13172 4870
rect 13196 4868 13252 4870
rect 7956 4378 8012 4380
rect 8036 4378 8092 4380
rect 8116 4378 8172 4380
rect 8196 4378 8252 4380
rect 7956 4326 8002 4378
rect 8002 4326 8012 4378
rect 8036 4326 8066 4378
rect 8066 4326 8078 4378
rect 8078 4326 8092 4378
rect 8116 4326 8130 4378
rect 8130 4326 8142 4378
rect 8142 4326 8172 4378
rect 8196 4326 8206 4378
rect 8206 4326 8252 4378
rect 7956 4324 8012 4326
rect 8036 4324 8092 4326
rect 8116 4324 8172 4326
rect 8196 4324 8252 4326
rect 1674 3984 1730 4040
rect 2956 3834 3012 3836
rect 3036 3834 3092 3836
rect 3116 3834 3172 3836
rect 3196 3834 3252 3836
rect 2956 3782 3002 3834
rect 3002 3782 3012 3834
rect 3036 3782 3066 3834
rect 3066 3782 3078 3834
rect 3078 3782 3092 3834
rect 3116 3782 3130 3834
rect 3130 3782 3142 3834
rect 3142 3782 3172 3834
rect 3196 3782 3206 3834
rect 3206 3782 3252 3834
rect 2956 3780 3012 3782
rect 3036 3780 3092 3782
rect 3116 3780 3172 3782
rect 3196 3780 3252 3782
rect 12956 3834 13012 3836
rect 13036 3834 13092 3836
rect 13116 3834 13172 3836
rect 13196 3834 13252 3836
rect 12956 3782 13002 3834
rect 13002 3782 13012 3834
rect 13036 3782 13066 3834
rect 13066 3782 13078 3834
rect 13078 3782 13092 3834
rect 13116 3782 13130 3834
rect 13130 3782 13142 3834
rect 13142 3782 13172 3834
rect 13196 3782 13206 3834
rect 13206 3782 13252 3834
rect 12956 3780 13012 3782
rect 13036 3780 13092 3782
rect 13116 3780 13172 3782
rect 13196 3780 13252 3782
rect 938 3576 994 3632
rect 5354 3576 5410 3632
rect 1122 3440 1178 3496
rect 938 3168 994 3224
rect 938 2760 994 2816
rect 938 2388 940 2408
rect 940 2388 992 2408
rect 992 2388 994 2408
rect 938 2352 994 2388
rect 2956 2746 3012 2748
rect 3036 2746 3092 2748
rect 3116 2746 3172 2748
rect 3196 2746 3252 2748
rect 2956 2694 3002 2746
rect 3002 2694 3012 2746
rect 3036 2694 3066 2746
rect 3066 2694 3078 2746
rect 3078 2694 3092 2746
rect 3116 2694 3130 2746
rect 3130 2694 3142 2746
rect 3142 2694 3172 2746
rect 3196 2694 3206 2746
rect 3206 2694 3252 2746
rect 2956 2692 3012 2694
rect 3036 2692 3092 2694
rect 3116 2692 3172 2694
rect 3196 2692 3252 2694
rect 1214 1944 1270 2000
rect 1306 1536 1362 1592
rect 7956 3290 8012 3292
rect 8036 3290 8092 3292
rect 8116 3290 8172 3292
rect 8196 3290 8252 3292
rect 7956 3238 8002 3290
rect 8002 3238 8012 3290
rect 8036 3238 8066 3290
rect 8066 3238 8078 3290
rect 8078 3238 8092 3290
rect 8116 3238 8130 3290
rect 8130 3238 8142 3290
rect 8142 3238 8172 3290
rect 8196 3238 8206 3290
rect 8206 3238 8252 3290
rect 7956 3236 8012 3238
rect 8036 3236 8092 3238
rect 8116 3236 8172 3238
rect 8196 3236 8252 3238
rect 7956 2202 8012 2204
rect 8036 2202 8092 2204
rect 8116 2202 8172 2204
rect 8196 2202 8252 2204
rect 7956 2150 8002 2202
rect 8002 2150 8012 2202
rect 8036 2150 8066 2202
rect 8066 2150 8078 2202
rect 8078 2150 8092 2202
rect 8116 2150 8130 2202
rect 8130 2150 8142 2202
rect 8142 2150 8172 2202
rect 8196 2150 8206 2202
rect 8206 2150 8252 2202
rect 7956 2148 8012 2150
rect 8036 2148 8092 2150
rect 8116 2148 8172 2150
rect 8196 2148 8252 2150
rect 12956 2746 13012 2748
rect 13036 2746 13092 2748
rect 13116 2746 13172 2748
rect 13196 2746 13252 2748
rect 12956 2694 13002 2746
rect 13002 2694 13012 2746
rect 13036 2694 13066 2746
rect 13066 2694 13078 2746
rect 13078 2694 13092 2746
rect 13116 2694 13130 2746
rect 13130 2694 13142 2746
rect 13142 2694 13172 2746
rect 13196 2694 13206 2746
rect 13206 2694 13252 2746
rect 12956 2692 13012 2694
rect 13036 2692 13092 2694
rect 13116 2692 13172 2694
rect 13196 2692 13252 2694
rect 14830 18128 14886 18184
rect 15382 20304 15438 20360
rect 15658 18808 15714 18864
rect 14922 16360 14978 16416
rect 14738 15136 14794 15192
rect 15106 15136 15162 15192
rect 14462 10668 14518 10704
rect 14462 10648 14464 10668
rect 14464 10648 14516 10668
rect 14516 10648 14518 10668
rect 15106 13640 15162 13696
rect 15014 12144 15070 12200
rect 15658 13776 15714 13832
rect 15566 12552 15622 12608
rect 15474 12280 15530 12336
rect 16578 23568 16634 23624
rect 16486 20748 16488 20768
rect 16488 20748 16540 20768
rect 16540 20748 16542 20768
rect 16486 20712 16542 20748
rect 16210 18672 16266 18728
rect 16670 19780 16726 19816
rect 16670 19760 16672 19780
rect 16672 19760 16724 19780
rect 16724 19760 16726 19780
rect 16486 18264 16542 18320
rect 16026 16532 16028 16552
rect 16028 16532 16080 16552
rect 16080 16532 16082 16552
rect 16026 16496 16082 16532
rect 16302 15408 16358 15464
rect 15842 12844 15898 12880
rect 15842 12824 15844 12844
rect 15844 12824 15896 12844
rect 15896 12824 15898 12844
rect 16210 14476 16266 14512
rect 16210 14456 16212 14476
rect 16212 14456 16264 14476
rect 16264 14456 16266 14476
rect 16578 17040 16634 17096
rect 16486 16360 16542 16416
rect 16302 12960 16358 13016
rect 16302 12824 16358 12880
rect 15474 9560 15530 9616
rect 14830 9036 14886 9072
rect 14830 9016 14832 9036
rect 14832 9016 14884 9036
rect 14884 9016 14886 9036
rect 16486 12960 16542 13016
rect 17956 23962 18012 23964
rect 18036 23962 18092 23964
rect 18116 23962 18172 23964
rect 18196 23962 18252 23964
rect 17956 23910 18002 23962
rect 18002 23910 18012 23962
rect 18036 23910 18066 23962
rect 18066 23910 18078 23962
rect 18078 23910 18092 23962
rect 18116 23910 18130 23962
rect 18130 23910 18142 23962
rect 18142 23910 18172 23962
rect 18196 23910 18206 23962
rect 18206 23910 18252 23962
rect 17956 23908 18012 23910
rect 18036 23908 18092 23910
rect 18116 23908 18172 23910
rect 18196 23908 18252 23910
rect 17956 22874 18012 22876
rect 18036 22874 18092 22876
rect 18116 22874 18172 22876
rect 18196 22874 18252 22876
rect 17956 22822 18002 22874
rect 18002 22822 18012 22874
rect 18036 22822 18066 22874
rect 18066 22822 18078 22874
rect 18078 22822 18092 22874
rect 18116 22822 18130 22874
rect 18130 22822 18142 22874
rect 18142 22822 18172 22874
rect 18196 22822 18206 22874
rect 18206 22822 18252 22874
rect 17956 22820 18012 22822
rect 18036 22820 18092 22822
rect 18116 22820 18172 22822
rect 18196 22820 18252 22822
rect 17956 21786 18012 21788
rect 18036 21786 18092 21788
rect 18116 21786 18172 21788
rect 18196 21786 18252 21788
rect 17956 21734 18002 21786
rect 18002 21734 18012 21786
rect 18036 21734 18066 21786
rect 18066 21734 18078 21786
rect 18078 21734 18092 21786
rect 18116 21734 18130 21786
rect 18130 21734 18142 21786
rect 18142 21734 18172 21786
rect 18196 21734 18206 21786
rect 18206 21734 18252 21786
rect 17956 21732 18012 21734
rect 18036 21732 18092 21734
rect 18116 21732 18172 21734
rect 18196 21732 18252 21734
rect 17956 20698 18012 20700
rect 18036 20698 18092 20700
rect 18116 20698 18172 20700
rect 18196 20698 18252 20700
rect 17956 20646 18002 20698
rect 18002 20646 18012 20698
rect 18036 20646 18066 20698
rect 18066 20646 18078 20698
rect 18078 20646 18092 20698
rect 18116 20646 18130 20698
rect 18130 20646 18142 20698
rect 18142 20646 18172 20698
rect 18196 20646 18206 20698
rect 18206 20646 18252 20698
rect 17956 20644 18012 20646
rect 18036 20644 18092 20646
rect 18116 20644 18172 20646
rect 18196 20644 18252 20646
rect 20534 22752 20590 22808
rect 17956 19610 18012 19612
rect 18036 19610 18092 19612
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 17956 19558 18002 19610
rect 18002 19558 18012 19610
rect 18036 19558 18066 19610
rect 18066 19558 18078 19610
rect 18078 19558 18092 19610
rect 18116 19558 18130 19610
rect 18130 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 17956 19556 18012 19558
rect 18036 19556 18092 19558
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 17406 19352 17462 19408
rect 18418 19624 18474 19680
rect 18418 18672 18474 18728
rect 17956 18522 18012 18524
rect 18036 18522 18092 18524
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 17956 18470 18002 18522
rect 18002 18470 18012 18522
rect 18036 18470 18066 18522
rect 18066 18470 18078 18522
rect 18078 18470 18092 18522
rect 18116 18470 18130 18522
rect 18130 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 17956 18468 18012 18470
rect 18036 18468 18092 18470
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 16854 14864 16910 14920
rect 16762 14220 16764 14240
rect 16764 14220 16816 14240
rect 16816 14220 16818 14240
rect 16762 14184 16818 14220
rect 17956 17434 18012 17436
rect 18036 17434 18092 17436
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 17956 17382 18002 17434
rect 18002 17382 18012 17434
rect 18036 17382 18066 17434
rect 18066 17382 18078 17434
rect 18078 17382 18092 17434
rect 18116 17382 18130 17434
rect 18130 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 17956 17380 18012 17382
rect 18036 17380 18092 17382
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 17406 15136 17462 15192
rect 17222 14456 17278 14512
rect 17222 12144 17278 12200
rect 17222 11192 17278 11248
rect 17956 16346 18012 16348
rect 18036 16346 18092 16348
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 17956 16294 18002 16346
rect 18002 16294 18012 16346
rect 18036 16294 18066 16346
rect 18066 16294 18078 16346
rect 18078 16294 18092 16346
rect 18116 16294 18130 16346
rect 18130 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 17956 16292 18012 16294
rect 18036 16292 18092 16294
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 18878 19624 18934 19680
rect 18786 17992 18842 18048
rect 17956 15258 18012 15260
rect 18036 15258 18092 15260
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 17956 15206 18002 15258
rect 18002 15206 18012 15258
rect 18036 15206 18066 15258
rect 18066 15206 18078 15258
rect 18078 15206 18092 15258
rect 18116 15206 18130 15258
rect 18130 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 17956 15204 18012 15206
rect 18036 15204 18092 15206
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 17958 14456 18014 14512
rect 17956 14170 18012 14172
rect 18036 14170 18092 14172
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 17956 14118 18002 14170
rect 18002 14118 18012 14170
rect 18036 14118 18066 14170
rect 18066 14118 18078 14170
rect 18078 14118 18092 14170
rect 18116 14118 18130 14170
rect 18130 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 17956 14116 18012 14118
rect 18036 14116 18092 14118
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 17958 13232 18014 13288
rect 17956 13082 18012 13084
rect 18036 13082 18092 13084
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 17956 13030 18002 13082
rect 18002 13030 18012 13082
rect 18036 13030 18066 13082
rect 18066 13030 18078 13082
rect 18078 13030 18092 13082
rect 18116 13030 18130 13082
rect 18130 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 17956 13028 18012 13030
rect 18036 13028 18092 13030
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 17774 12180 17776 12200
rect 17776 12180 17828 12200
rect 17828 12180 17830 12200
rect 17774 12144 17830 12180
rect 17956 11994 18012 11996
rect 18036 11994 18092 11996
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 17956 11942 18002 11994
rect 18002 11942 18012 11994
rect 18036 11942 18066 11994
rect 18066 11942 18078 11994
rect 18078 11942 18092 11994
rect 18116 11942 18130 11994
rect 18130 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 17956 11940 18012 11942
rect 18036 11940 18092 11942
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 19154 20596 19210 20632
rect 19154 20576 19156 20596
rect 19156 20576 19208 20596
rect 19208 20576 19210 20596
rect 22956 24506 23012 24508
rect 23036 24506 23092 24508
rect 23116 24506 23172 24508
rect 23196 24506 23252 24508
rect 22956 24454 23002 24506
rect 23002 24454 23012 24506
rect 23036 24454 23066 24506
rect 23066 24454 23078 24506
rect 23078 24454 23092 24506
rect 23116 24454 23130 24506
rect 23130 24454 23142 24506
rect 23142 24454 23172 24506
rect 23196 24454 23206 24506
rect 23206 24454 23252 24506
rect 22956 24452 23012 24454
rect 23036 24452 23092 24454
rect 23116 24452 23172 24454
rect 23196 24452 23252 24454
rect 22956 23418 23012 23420
rect 23036 23418 23092 23420
rect 23116 23418 23172 23420
rect 23196 23418 23252 23420
rect 22956 23366 23002 23418
rect 23002 23366 23012 23418
rect 23036 23366 23066 23418
rect 23066 23366 23078 23418
rect 23078 23366 23092 23418
rect 23116 23366 23130 23418
rect 23130 23366 23142 23418
rect 23142 23366 23172 23418
rect 23196 23366 23206 23418
rect 23206 23366 23252 23418
rect 22956 23364 23012 23366
rect 23036 23364 23092 23366
rect 23116 23364 23172 23366
rect 23196 23364 23252 23366
rect 19338 19896 19394 19952
rect 19338 18536 19394 18592
rect 19246 18400 19302 18456
rect 19246 17720 19302 17776
rect 18878 15408 18934 15464
rect 18602 14456 18658 14512
rect 17956 10906 18012 10908
rect 18036 10906 18092 10908
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 17956 10854 18002 10906
rect 18002 10854 18012 10906
rect 18036 10854 18066 10906
rect 18066 10854 18078 10906
rect 18078 10854 18092 10906
rect 18116 10854 18130 10906
rect 18130 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 17956 10852 18012 10854
rect 18036 10852 18092 10854
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 17956 9818 18012 9820
rect 18036 9818 18092 9820
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 17956 9766 18002 9818
rect 18002 9766 18012 9818
rect 18036 9766 18066 9818
rect 18066 9766 18078 9818
rect 18078 9766 18092 9818
rect 18116 9766 18130 9818
rect 18130 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 17956 9764 18012 9766
rect 18036 9764 18092 9766
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 17956 8730 18012 8732
rect 18036 8730 18092 8732
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 17956 8678 18002 8730
rect 18002 8678 18012 8730
rect 18036 8678 18066 8730
rect 18066 8678 18078 8730
rect 18078 8678 18092 8730
rect 18116 8678 18130 8730
rect 18130 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 17956 8676 18012 8678
rect 18036 8676 18092 8678
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 18786 13232 18842 13288
rect 18418 9016 18474 9072
rect 17956 7642 18012 7644
rect 18036 7642 18092 7644
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 17956 7590 18002 7642
rect 18002 7590 18012 7642
rect 18036 7590 18066 7642
rect 18066 7590 18078 7642
rect 18078 7590 18092 7642
rect 18116 7590 18130 7642
rect 18130 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 17956 7588 18012 7590
rect 18036 7588 18092 7590
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 17956 6554 18012 6556
rect 18036 6554 18092 6556
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 17956 6502 18002 6554
rect 18002 6502 18012 6554
rect 18036 6502 18066 6554
rect 18066 6502 18078 6554
rect 18078 6502 18092 6554
rect 18116 6502 18130 6554
rect 18130 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 17956 6500 18012 6502
rect 18036 6500 18092 6502
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 17956 5466 18012 5468
rect 18036 5466 18092 5468
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 17956 5414 18002 5466
rect 18002 5414 18012 5466
rect 18036 5414 18066 5466
rect 18066 5414 18078 5466
rect 18078 5414 18092 5466
rect 18116 5414 18130 5466
rect 18130 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 17956 5412 18012 5414
rect 18036 5412 18092 5414
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 17956 4378 18012 4380
rect 18036 4378 18092 4380
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 17956 4326 18002 4378
rect 18002 4326 18012 4378
rect 18036 4326 18066 4378
rect 18066 4326 18078 4378
rect 18078 4326 18092 4378
rect 18116 4326 18130 4378
rect 18130 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 17956 4324 18012 4326
rect 18036 4324 18092 4326
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 19706 18536 19762 18592
rect 19982 17312 20038 17368
rect 19338 10668 19394 10704
rect 19338 10648 19340 10668
rect 19340 10648 19392 10668
rect 19392 10648 19394 10668
rect 20534 18944 20590 19000
rect 21178 20440 21234 20496
rect 21454 19216 21510 19272
rect 20626 17448 20682 17504
rect 20994 17312 21050 17368
rect 20074 14048 20130 14104
rect 20902 15544 20958 15600
rect 21270 18400 21326 18456
rect 21178 16224 21234 16280
rect 21178 13640 21234 13696
rect 22282 22752 22338 22808
rect 22282 21800 22338 21856
rect 22190 20984 22246 21040
rect 22282 18944 22338 19000
rect 22374 18400 22430 18456
rect 22190 17720 22246 17776
rect 20994 11736 21050 11792
rect 20626 10648 20682 10704
rect 21730 15156 21786 15192
rect 21730 15136 21732 15156
rect 21732 15136 21784 15156
rect 21784 15136 21786 15156
rect 17956 3290 18012 3292
rect 18036 3290 18092 3292
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 17956 3238 18002 3290
rect 18002 3238 18012 3290
rect 18036 3238 18066 3290
rect 18066 3238 18078 3290
rect 18078 3238 18092 3290
rect 18116 3238 18130 3290
rect 18130 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 17956 3236 18012 3238
rect 18036 3236 18092 3238
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 17956 2202 18012 2204
rect 18036 2202 18092 2204
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 17956 2150 18002 2202
rect 18002 2150 18012 2202
rect 18036 2150 18066 2202
rect 18066 2150 18078 2202
rect 18078 2150 18092 2202
rect 18116 2150 18130 2202
rect 18130 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 17956 2148 18012 2150
rect 18036 2148 18092 2150
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 22282 15544 22338 15600
rect 22956 22330 23012 22332
rect 23036 22330 23092 22332
rect 23116 22330 23172 22332
rect 23196 22330 23252 22332
rect 22956 22278 23002 22330
rect 23002 22278 23012 22330
rect 23036 22278 23066 22330
rect 23066 22278 23078 22330
rect 23078 22278 23092 22330
rect 23116 22278 23130 22330
rect 23130 22278 23142 22330
rect 23142 22278 23172 22330
rect 23196 22278 23206 22330
rect 23206 22278 23252 22330
rect 22956 22276 23012 22278
rect 23036 22276 23092 22278
rect 23116 22276 23172 22278
rect 23196 22276 23252 22278
rect 23386 21936 23442 21992
rect 22956 21242 23012 21244
rect 23036 21242 23092 21244
rect 23116 21242 23172 21244
rect 23196 21242 23252 21244
rect 22956 21190 23002 21242
rect 23002 21190 23012 21242
rect 23036 21190 23066 21242
rect 23066 21190 23078 21242
rect 23078 21190 23092 21242
rect 23116 21190 23130 21242
rect 23130 21190 23142 21242
rect 23142 21190 23172 21242
rect 23196 21190 23206 21242
rect 23206 21190 23252 21242
rect 22956 21188 23012 21190
rect 23036 21188 23092 21190
rect 23116 21188 23172 21190
rect 23196 21188 23252 21190
rect 22956 20154 23012 20156
rect 23036 20154 23092 20156
rect 23116 20154 23172 20156
rect 23196 20154 23252 20156
rect 22956 20102 23002 20154
rect 23002 20102 23012 20154
rect 23036 20102 23066 20154
rect 23066 20102 23078 20154
rect 23078 20102 23092 20154
rect 23116 20102 23130 20154
rect 23130 20102 23142 20154
rect 23142 20102 23172 20154
rect 23196 20102 23206 20154
rect 23206 20102 23252 20154
rect 22956 20100 23012 20102
rect 23036 20100 23092 20102
rect 23116 20100 23172 20102
rect 23196 20100 23252 20102
rect 22742 18808 22798 18864
rect 24950 24112 25006 24168
rect 26054 24792 26110 24848
rect 26330 24656 26386 24712
rect 24766 23296 24822 23352
rect 24950 23160 25006 23216
rect 24674 22344 24730 22400
rect 26238 23568 26294 23624
rect 22956 19066 23012 19068
rect 23036 19066 23092 19068
rect 23116 19066 23172 19068
rect 23196 19066 23252 19068
rect 22956 19014 23002 19066
rect 23002 19014 23012 19066
rect 23036 19014 23066 19066
rect 23066 19014 23078 19066
rect 23078 19014 23092 19066
rect 23116 19014 23130 19066
rect 23130 19014 23142 19066
rect 23142 19014 23172 19066
rect 23196 19014 23206 19066
rect 23206 19014 23252 19066
rect 22956 19012 23012 19014
rect 23036 19012 23092 19014
rect 23116 19012 23172 19014
rect 23196 19012 23252 19014
rect 22956 17978 23012 17980
rect 23036 17978 23092 17980
rect 23116 17978 23172 17980
rect 23196 17978 23252 17980
rect 22956 17926 23002 17978
rect 23002 17926 23012 17978
rect 23036 17926 23066 17978
rect 23066 17926 23078 17978
rect 23078 17926 23092 17978
rect 23116 17926 23130 17978
rect 23130 17926 23142 17978
rect 23142 17926 23172 17978
rect 23196 17926 23206 17978
rect 23206 17926 23252 17978
rect 22956 17924 23012 17926
rect 23036 17924 23092 17926
rect 23116 17924 23172 17926
rect 23196 17924 23252 17926
rect 22374 14320 22430 14376
rect 22558 14320 22614 14376
rect 22374 12688 22430 12744
rect 22956 16890 23012 16892
rect 23036 16890 23092 16892
rect 23116 16890 23172 16892
rect 23196 16890 23252 16892
rect 22956 16838 23002 16890
rect 23002 16838 23012 16890
rect 23036 16838 23066 16890
rect 23066 16838 23078 16890
rect 23078 16838 23092 16890
rect 23116 16838 23130 16890
rect 23130 16838 23142 16890
rect 23142 16838 23172 16890
rect 23196 16838 23206 16890
rect 23206 16838 23252 16890
rect 22956 16836 23012 16838
rect 23036 16836 23092 16838
rect 23116 16836 23172 16838
rect 23196 16836 23252 16838
rect 22956 15802 23012 15804
rect 23036 15802 23092 15804
rect 23116 15802 23172 15804
rect 23196 15802 23252 15804
rect 22956 15750 23002 15802
rect 23002 15750 23012 15802
rect 23036 15750 23066 15802
rect 23066 15750 23078 15802
rect 23078 15750 23092 15802
rect 23116 15750 23130 15802
rect 23130 15750 23142 15802
rect 23142 15750 23172 15802
rect 23196 15750 23206 15802
rect 23206 15750 23252 15802
rect 22956 15748 23012 15750
rect 23036 15748 23092 15750
rect 23116 15748 23172 15750
rect 23196 15748 23252 15750
rect 22956 14714 23012 14716
rect 23036 14714 23092 14716
rect 23116 14714 23172 14716
rect 23196 14714 23252 14716
rect 22956 14662 23002 14714
rect 23002 14662 23012 14714
rect 23036 14662 23066 14714
rect 23066 14662 23078 14714
rect 23078 14662 23092 14714
rect 23116 14662 23130 14714
rect 23130 14662 23142 14714
rect 23142 14662 23172 14714
rect 23196 14662 23206 14714
rect 23206 14662 23252 14714
rect 22956 14660 23012 14662
rect 23036 14660 23092 14662
rect 23116 14660 23172 14662
rect 23196 14660 23252 14662
rect 22956 13626 23012 13628
rect 23036 13626 23092 13628
rect 23116 13626 23172 13628
rect 23196 13626 23252 13628
rect 22956 13574 23002 13626
rect 23002 13574 23012 13626
rect 23036 13574 23066 13626
rect 23066 13574 23078 13626
rect 23078 13574 23092 13626
rect 23116 13574 23130 13626
rect 23130 13574 23142 13626
rect 23142 13574 23172 13626
rect 23196 13574 23206 13626
rect 23206 13574 23252 13626
rect 22956 13572 23012 13574
rect 23036 13572 23092 13574
rect 23116 13572 23172 13574
rect 23196 13572 23252 13574
rect 22466 12008 22522 12064
rect 22956 12538 23012 12540
rect 23036 12538 23092 12540
rect 23116 12538 23172 12540
rect 23196 12538 23252 12540
rect 22956 12486 23002 12538
rect 23002 12486 23012 12538
rect 23036 12486 23066 12538
rect 23066 12486 23078 12538
rect 23078 12486 23092 12538
rect 23116 12486 23130 12538
rect 23130 12486 23142 12538
rect 23142 12486 23172 12538
rect 23196 12486 23206 12538
rect 23206 12486 23252 12538
rect 22956 12484 23012 12486
rect 23036 12484 23092 12486
rect 23116 12484 23172 12486
rect 23196 12484 23252 12486
rect 24214 20712 24270 20768
rect 23662 14048 23718 14104
rect 22956 11450 23012 11452
rect 23036 11450 23092 11452
rect 23116 11450 23172 11452
rect 23196 11450 23252 11452
rect 22956 11398 23002 11450
rect 23002 11398 23012 11450
rect 23036 11398 23066 11450
rect 23066 11398 23078 11450
rect 23078 11398 23092 11450
rect 23116 11398 23130 11450
rect 23130 11398 23142 11450
rect 23142 11398 23172 11450
rect 23196 11398 23206 11450
rect 23206 11398 23252 11450
rect 22956 11396 23012 11398
rect 23036 11396 23092 11398
rect 23116 11396 23172 11398
rect 23196 11396 23252 11398
rect 23294 11212 23350 11248
rect 23294 11192 23296 11212
rect 23296 11192 23348 11212
rect 23348 11192 23350 11212
rect 22956 10362 23012 10364
rect 23036 10362 23092 10364
rect 23116 10362 23172 10364
rect 23196 10362 23252 10364
rect 22956 10310 23002 10362
rect 23002 10310 23012 10362
rect 23036 10310 23066 10362
rect 23066 10310 23078 10362
rect 23078 10310 23092 10362
rect 23116 10310 23130 10362
rect 23130 10310 23142 10362
rect 23142 10310 23172 10362
rect 23196 10310 23206 10362
rect 23206 10310 23252 10362
rect 22956 10308 23012 10310
rect 23036 10308 23092 10310
rect 23116 10308 23172 10310
rect 23196 10308 23252 10310
rect 25134 21392 25190 21448
rect 25042 20884 25044 20904
rect 25044 20884 25096 20904
rect 25096 20884 25098 20904
rect 25042 20848 25098 20884
rect 24674 19216 24730 19272
rect 24306 17720 24362 17776
rect 24674 17992 24730 18048
rect 24490 16124 24492 16144
rect 24492 16124 24544 16144
rect 24544 16124 24546 16144
rect 24490 16088 24546 16124
rect 25134 20440 25190 20496
rect 25594 22616 25650 22672
rect 25042 19080 25098 19136
rect 26698 23024 26754 23080
rect 26422 22208 26478 22264
rect 26606 21836 26608 21856
rect 26608 21836 26660 21856
rect 26660 21836 26662 21856
rect 26422 20984 26478 21040
rect 25870 20440 25926 20496
rect 26146 20304 26202 20360
rect 25962 20168 26018 20224
rect 25962 19352 26018 19408
rect 25042 18536 25098 18592
rect 24950 18128 25006 18184
rect 24858 15952 24914 16008
rect 24858 15564 24914 15600
rect 24858 15544 24860 15564
rect 24860 15544 24912 15564
rect 24912 15544 24914 15564
rect 23754 12044 23756 12064
rect 23756 12044 23808 12064
rect 23808 12044 23810 12064
rect 23754 12008 23810 12044
rect 22956 9274 23012 9276
rect 23036 9274 23092 9276
rect 23116 9274 23172 9276
rect 23196 9274 23252 9276
rect 22956 9222 23002 9274
rect 23002 9222 23012 9274
rect 23036 9222 23066 9274
rect 23066 9222 23078 9274
rect 23078 9222 23092 9274
rect 23116 9222 23130 9274
rect 23130 9222 23142 9274
rect 23142 9222 23172 9274
rect 23196 9222 23206 9274
rect 23206 9222 23252 9274
rect 22956 9220 23012 9222
rect 23036 9220 23092 9222
rect 23116 9220 23172 9222
rect 23196 9220 23252 9222
rect 22956 8186 23012 8188
rect 23036 8186 23092 8188
rect 23116 8186 23172 8188
rect 23196 8186 23252 8188
rect 22956 8134 23002 8186
rect 23002 8134 23012 8186
rect 23036 8134 23066 8186
rect 23066 8134 23078 8186
rect 23078 8134 23092 8186
rect 23116 8134 23130 8186
rect 23130 8134 23142 8186
rect 23142 8134 23172 8186
rect 23196 8134 23206 8186
rect 23206 8134 23252 8186
rect 22956 8132 23012 8134
rect 23036 8132 23092 8134
rect 23116 8132 23172 8134
rect 23196 8132 23252 8134
rect 22190 3440 22246 3496
rect 22956 7098 23012 7100
rect 23036 7098 23092 7100
rect 23116 7098 23172 7100
rect 23196 7098 23252 7100
rect 22956 7046 23002 7098
rect 23002 7046 23012 7098
rect 23036 7046 23066 7098
rect 23066 7046 23078 7098
rect 23078 7046 23092 7098
rect 23116 7046 23130 7098
rect 23130 7046 23142 7098
rect 23142 7046 23172 7098
rect 23196 7046 23206 7098
rect 23206 7046 23252 7098
rect 22956 7044 23012 7046
rect 23036 7044 23092 7046
rect 23116 7044 23172 7046
rect 23196 7044 23252 7046
rect 22956 6010 23012 6012
rect 23036 6010 23092 6012
rect 23116 6010 23172 6012
rect 23196 6010 23252 6012
rect 22956 5958 23002 6010
rect 23002 5958 23012 6010
rect 23036 5958 23066 6010
rect 23066 5958 23078 6010
rect 23078 5958 23092 6010
rect 23116 5958 23130 6010
rect 23130 5958 23142 6010
rect 23142 5958 23172 6010
rect 23196 5958 23206 6010
rect 23206 5958 23252 6010
rect 22956 5956 23012 5958
rect 23036 5956 23092 5958
rect 23116 5956 23172 5958
rect 23196 5956 23252 5958
rect 22956 4922 23012 4924
rect 23036 4922 23092 4924
rect 23116 4922 23172 4924
rect 23196 4922 23252 4924
rect 22956 4870 23002 4922
rect 23002 4870 23012 4922
rect 23036 4870 23066 4922
rect 23066 4870 23078 4922
rect 23078 4870 23092 4922
rect 23116 4870 23130 4922
rect 23130 4870 23142 4922
rect 23142 4870 23172 4922
rect 23196 4870 23206 4922
rect 23206 4870 23252 4922
rect 22956 4868 23012 4870
rect 23036 4868 23092 4870
rect 23116 4868 23172 4870
rect 23196 4868 23252 4870
rect 22956 3834 23012 3836
rect 23036 3834 23092 3836
rect 23116 3834 23172 3836
rect 23196 3834 23252 3836
rect 22956 3782 23002 3834
rect 23002 3782 23012 3834
rect 23036 3782 23066 3834
rect 23066 3782 23078 3834
rect 23078 3782 23092 3834
rect 23116 3782 23130 3834
rect 23130 3782 23142 3834
rect 23142 3782 23172 3834
rect 23196 3782 23206 3834
rect 23206 3782 23252 3834
rect 22956 3780 23012 3782
rect 23036 3780 23092 3782
rect 23116 3780 23172 3782
rect 23196 3780 23252 3782
rect 24674 13948 24676 13968
rect 24676 13948 24728 13968
rect 24728 13948 24730 13968
rect 24674 13912 24730 13948
rect 25686 17604 25742 17640
rect 26146 19388 26148 19408
rect 26148 19388 26200 19408
rect 26200 19388 26202 19408
rect 26146 19352 26202 19388
rect 25686 17584 25688 17604
rect 25688 17584 25740 17604
rect 25740 17584 25742 17604
rect 25594 17176 25650 17232
rect 25410 15428 25466 15464
rect 25410 15408 25412 15428
rect 25412 15408 25464 15428
rect 25464 15408 25466 15428
rect 25318 12824 25374 12880
rect 26054 18028 26056 18048
rect 26056 18028 26108 18048
rect 26108 18028 26110 18048
rect 26054 17992 26110 18028
rect 26606 21800 26662 21836
rect 26330 17448 26386 17504
rect 26054 16496 26110 16552
rect 26330 16244 26386 16280
rect 26330 16224 26332 16244
rect 26332 16224 26384 16244
rect 26384 16224 26386 16244
rect 26146 15952 26202 16008
rect 26606 17448 26662 17504
rect 26238 15544 26294 15600
rect 26146 15000 26202 15056
rect 26146 14900 26148 14920
rect 26148 14900 26200 14920
rect 26200 14900 26202 14920
rect 26146 14864 26202 14900
rect 25778 13948 25780 13968
rect 25780 13948 25832 13968
rect 25832 13948 25834 13968
rect 25778 13912 25834 13948
rect 26238 12824 26294 12880
rect 22956 2746 23012 2748
rect 23036 2746 23092 2748
rect 23116 2746 23172 2748
rect 23196 2746 23252 2748
rect 22956 2694 23002 2746
rect 23002 2694 23012 2746
rect 23036 2694 23066 2746
rect 23066 2694 23078 2746
rect 23078 2694 23092 2746
rect 23116 2694 23130 2746
rect 23130 2694 23142 2746
rect 23142 2694 23172 2746
rect 23196 2694 23206 2746
rect 23206 2694 23252 2746
rect 22956 2692 23012 2694
rect 23036 2692 23092 2694
rect 23116 2692 23172 2694
rect 23196 2692 23252 2694
rect 24398 3576 24454 3632
rect 26790 19780 26846 19816
rect 26790 19760 26792 19780
rect 26792 19760 26844 19780
rect 26844 19760 26846 19780
rect 27618 22072 27674 22128
rect 27956 23962 28012 23964
rect 28036 23962 28092 23964
rect 28116 23962 28172 23964
rect 28196 23962 28252 23964
rect 27956 23910 28002 23962
rect 28002 23910 28012 23962
rect 28036 23910 28066 23962
rect 28066 23910 28078 23962
rect 28078 23910 28092 23962
rect 28116 23910 28130 23962
rect 28130 23910 28142 23962
rect 28142 23910 28172 23962
rect 28196 23910 28206 23962
rect 28206 23910 28252 23962
rect 27956 23908 28012 23910
rect 28036 23908 28092 23910
rect 28116 23908 28172 23910
rect 28196 23908 28252 23910
rect 27894 23316 27950 23352
rect 27894 23296 27896 23316
rect 27896 23296 27948 23316
rect 27948 23296 27950 23316
rect 27956 22874 28012 22876
rect 28036 22874 28092 22876
rect 28116 22874 28172 22876
rect 28196 22874 28252 22876
rect 27956 22822 28002 22874
rect 28002 22822 28012 22874
rect 28036 22822 28066 22874
rect 28066 22822 28078 22874
rect 28078 22822 28092 22874
rect 28116 22822 28130 22874
rect 28130 22822 28142 22874
rect 28142 22822 28172 22874
rect 28196 22822 28206 22874
rect 28206 22822 28252 22874
rect 27956 22820 28012 22822
rect 28036 22820 28092 22822
rect 28116 22820 28172 22822
rect 28196 22820 28252 22822
rect 27802 22072 27858 22128
rect 27956 21786 28012 21788
rect 28036 21786 28092 21788
rect 28116 21786 28172 21788
rect 28196 21786 28252 21788
rect 27956 21734 28002 21786
rect 28002 21734 28012 21786
rect 28036 21734 28066 21786
rect 28066 21734 28078 21786
rect 28078 21734 28092 21786
rect 28116 21734 28130 21786
rect 28130 21734 28142 21786
rect 28142 21734 28172 21786
rect 28196 21734 28206 21786
rect 28206 21734 28252 21786
rect 27956 21732 28012 21734
rect 28036 21732 28092 21734
rect 28116 21732 28172 21734
rect 28196 21732 28252 21734
rect 27342 21120 27398 21176
rect 27710 21528 27766 21584
rect 27618 20848 27674 20904
rect 27710 20712 27766 20768
rect 28446 21800 28502 21856
rect 28998 23160 29054 23216
rect 28538 21256 28594 21312
rect 28354 20848 28410 20904
rect 28814 21800 28870 21856
rect 27956 20698 28012 20700
rect 28036 20698 28092 20700
rect 28116 20698 28172 20700
rect 28196 20698 28252 20700
rect 27956 20646 28002 20698
rect 28002 20646 28012 20698
rect 28036 20646 28066 20698
rect 28066 20646 28078 20698
rect 28078 20646 28092 20698
rect 28116 20646 28130 20698
rect 28130 20646 28142 20698
rect 28142 20646 28172 20698
rect 28196 20646 28206 20698
rect 28206 20646 28252 20698
rect 27956 20644 28012 20646
rect 28036 20644 28092 20646
rect 28116 20644 28172 20646
rect 28196 20644 28252 20646
rect 28262 19896 28318 19952
rect 28538 20304 28594 20360
rect 28446 20168 28502 20224
rect 27956 19610 28012 19612
rect 28036 19610 28092 19612
rect 28116 19610 28172 19612
rect 28196 19610 28252 19612
rect 27956 19558 28002 19610
rect 28002 19558 28012 19610
rect 28036 19558 28066 19610
rect 28066 19558 28078 19610
rect 28078 19558 28092 19610
rect 28116 19558 28130 19610
rect 28130 19558 28142 19610
rect 28142 19558 28172 19610
rect 28196 19558 28206 19610
rect 28206 19558 28252 19610
rect 27956 19556 28012 19558
rect 28036 19556 28092 19558
rect 28116 19556 28172 19558
rect 28196 19556 28252 19558
rect 28354 18944 28410 19000
rect 27956 18522 28012 18524
rect 28036 18522 28092 18524
rect 28116 18522 28172 18524
rect 28196 18522 28252 18524
rect 27956 18470 28002 18522
rect 28002 18470 28012 18522
rect 28036 18470 28066 18522
rect 28066 18470 28078 18522
rect 28078 18470 28092 18522
rect 28116 18470 28130 18522
rect 28130 18470 28142 18522
rect 28142 18470 28172 18522
rect 28196 18470 28206 18522
rect 28206 18470 28252 18522
rect 27956 18468 28012 18470
rect 28036 18468 28092 18470
rect 28116 18468 28172 18470
rect 28196 18468 28252 18470
rect 27802 17448 27858 17504
rect 27956 17434 28012 17436
rect 28036 17434 28092 17436
rect 28116 17434 28172 17436
rect 28196 17434 28252 17436
rect 27956 17382 28002 17434
rect 28002 17382 28012 17434
rect 28036 17382 28066 17434
rect 28066 17382 28078 17434
rect 28078 17382 28092 17434
rect 28116 17382 28130 17434
rect 28130 17382 28142 17434
rect 28142 17382 28172 17434
rect 28196 17382 28206 17434
rect 28206 17382 28252 17434
rect 27956 17380 28012 17382
rect 28036 17380 28092 17382
rect 28116 17380 28172 17382
rect 28196 17380 28252 17382
rect 27710 17196 27766 17232
rect 27710 17176 27712 17196
rect 27712 17176 27764 17196
rect 27764 17176 27766 17196
rect 27802 17076 27804 17096
rect 27804 17076 27856 17096
rect 27856 17076 27858 17096
rect 27802 17040 27858 17076
rect 27526 15020 27582 15056
rect 27526 15000 27528 15020
rect 27528 15000 27580 15020
rect 27580 15000 27582 15020
rect 27710 16088 27766 16144
rect 27956 16346 28012 16348
rect 28036 16346 28092 16348
rect 28116 16346 28172 16348
rect 28196 16346 28252 16348
rect 27956 16294 28002 16346
rect 28002 16294 28012 16346
rect 28036 16294 28066 16346
rect 28066 16294 28078 16346
rect 28078 16294 28092 16346
rect 28116 16294 28130 16346
rect 28130 16294 28142 16346
rect 28142 16294 28172 16346
rect 28196 16294 28206 16346
rect 28206 16294 28252 16346
rect 27956 16292 28012 16294
rect 28036 16292 28092 16294
rect 28116 16292 28172 16294
rect 28196 16292 28252 16294
rect 28538 20032 28594 20088
rect 28538 19624 28594 19680
rect 29090 22480 29146 22536
rect 29458 20984 29514 21040
rect 29458 20712 29514 20768
rect 27956 15258 28012 15260
rect 28036 15258 28092 15260
rect 28116 15258 28172 15260
rect 28196 15258 28252 15260
rect 27956 15206 28002 15258
rect 28002 15206 28012 15258
rect 28036 15206 28066 15258
rect 28066 15206 28078 15258
rect 28078 15206 28092 15258
rect 28116 15206 28130 15258
rect 28130 15206 28142 15258
rect 28142 15206 28172 15258
rect 28196 15206 28206 15258
rect 28206 15206 28252 15258
rect 27956 15204 28012 15206
rect 28036 15204 28092 15206
rect 28116 15204 28172 15206
rect 28196 15204 28252 15206
rect 26146 9580 26202 9616
rect 26146 9560 26148 9580
rect 26148 9560 26200 9580
rect 26200 9560 26202 9580
rect 27434 11736 27490 11792
rect 27956 14170 28012 14172
rect 28036 14170 28092 14172
rect 28116 14170 28172 14172
rect 28196 14170 28252 14172
rect 27956 14118 28002 14170
rect 28002 14118 28012 14170
rect 28036 14118 28066 14170
rect 28066 14118 28078 14170
rect 28078 14118 28092 14170
rect 28116 14118 28130 14170
rect 28130 14118 28142 14170
rect 28142 14118 28172 14170
rect 28196 14118 28206 14170
rect 28206 14118 28252 14170
rect 27956 14116 28012 14118
rect 28036 14116 28092 14118
rect 28116 14116 28172 14118
rect 28196 14116 28252 14118
rect 27956 13082 28012 13084
rect 28036 13082 28092 13084
rect 28116 13082 28172 13084
rect 28196 13082 28252 13084
rect 27956 13030 28002 13082
rect 28002 13030 28012 13082
rect 28036 13030 28066 13082
rect 28066 13030 28078 13082
rect 28078 13030 28092 13082
rect 28116 13030 28130 13082
rect 28130 13030 28142 13082
rect 28142 13030 28172 13082
rect 28196 13030 28206 13082
rect 28206 13030 28252 13082
rect 27956 13028 28012 13030
rect 28036 13028 28092 13030
rect 28116 13028 28172 13030
rect 28196 13028 28252 13030
rect 27710 12008 27766 12064
rect 27956 11994 28012 11996
rect 28036 11994 28092 11996
rect 28116 11994 28172 11996
rect 28196 11994 28252 11996
rect 27956 11942 28002 11994
rect 28002 11942 28012 11994
rect 28036 11942 28066 11994
rect 28066 11942 28078 11994
rect 28078 11942 28092 11994
rect 28116 11942 28130 11994
rect 28130 11942 28142 11994
rect 28142 11942 28172 11994
rect 28196 11942 28206 11994
rect 28206 11942 28252 11994
rect 27956 11940 28012 11942
rect 28036 11940 28092 11942
rect 28116 11940 28172 11942
rect 28196 11940 28252 11942
rect 27956 10906 28012 10908
rect 28036 10906 28092 10908
rect 28116 10906 28172 10908
rect 28196 10906 28252 10908
rect 27956 10854 28002 10906
rect 28002 10854 28012 10906
rect 28036 10854 28066 10906
rect 28066 10854 28078 10906
rect 28078 10854 28092 10906
rect 28116 10854 28130 10906
rect 28130 10854 28142 10906
rect 28142 10854 28172 10906
rect 28196 10854 28206 10906
rect 28206 10854 28252 10906
rect 27956 10852 28012 10854
rect 28036 10852 28092 10854
rect 28116 10852 28172 10854
rect 28196 10852 28252 10854
rect 28814 13368 28870 13424
rect 29642 20304 29698 20360
rect 29918 21936 29974 21992
rect 29918 21256 29974 21312
rect 29918 20984 29974 21040
rect 30286 22208 30342 22264
rect 34518 26288 34574 26344
rect 31114 22616 31170 22672
rect 30746 22072 30802 22128
rect 31482 22380 31484 22400
rect 31484 22380 31536 22400
rect 31536 22380 31538 22400
rect 31482 22344 31538 22380
rect 31666 22752 31722 22808
rect 30286 21140 30342 21176
rect 30286 21120 30288 21140
rect 30288 21120 30340 21140
rect 30340 21120 30342 21140
rect 30102 20340 30104 20360
rect 30104 20340 30156 20360
rect 30156 20340 30158 20360
rect 30102 20304 30158 20340
rect 30010 19624 30066 19680
rect 29734 17720 29790 17776
rect 29458 14728 29514 14784
rect 29550 14184 29606 14240
rect 30194 19216 30250 19272
rect 30010 18264 30066 18320
rect 30194 18264 30250 18320
rect 27956 9818 28012 9820
rect 28036 9818 28092 9820
rect 28116 9818 28172 9820
rect 28196 9818 28252 9820
rect 27956 9766 28002 9818
rect 28002 9766 28012 9818
rect 28036 9766 28066 9818
rect 28066 9766 28078 9818
rect 28078 9766 28092 9818
rect 28116 9766 28130 9818
rect 28130 9766 28142 9818
rect 28142 9766 28172 9818
rect 28196 9766 28206 9818
rect 28206 9766 28252 9818
rect 27956 9764 28012 9766
rect 28036 9764 28092 9766
rect 28116 9764 28172 9766
rect 28196 9764 28252 9766
rect 28630 8880 28686 8936
rect 27956 8730 28012 8732
rect 28036 8730 28092 8732
rect 28116 8730 28172 8732
rect 28196 8730 28252 8732
rect 27956 8678 28002 8730
rect 28002 8678 28012 8730
rect 28036 8678 28066 8730
rect 28066 8678 28078 8730
rect 28078 8678 28092 8730
rect 28116 8678 28130 8730
rect 28130 8678 28142 8730
rect 28142 8678 28172 8730
rect 28196 8678 28206 8730
rect 28206 8678 28252 8730
rect 27956 8676 28012 8678
rect 28036 8676 28092 8678
rect 28116 8676 28172 8678
rect 28196 8676 28252 8678
rect 30838 19896 30894 19952
rect 30746 19080 30802 19136
rect 30654 18536 30710 18592
rect 31114 20848 31170 20904
rect 31114 20596 31170 20632
rect 31114 20576 31116 20596
rect 31116 20576 31168 20596
rect 31168 20576 31170 20596
rect 32310 24248 32366 24304
rect 27956 7642 28012 7644
rect 28036 7642 28092 7644
rect 28116 7642 28172 7644
rect 28196 7642 28252 7644
rect 27956 7590 28002 7642
rect 28002 7590 28012 7642
rect 28036 7590 28066 7642
rect 28066 7590 28078 7642
rect 28078 7590 28092 7642
rect 28116 7590 28130 7642
rect 28130 7590 28142 7642
rect 28142 7590 28172 7642
rect 28196 7590 28206 7642
rect 28206 7590 28252 7642
rect 27956 7588 28012 7590
rect 28036 7588 28092 7590
rect 28116 7588 28172 7590
rect 28196 7588 28252 7590
rect 27956 6554 28012 6556
rect 28036 6554 28092 6556
rect 28116 6554 28172 6556
rect 28196 6554 28252 6556
rect 27956 6502 28002 6554
rect 28002 6502 28012 6554
rect 28036 6502 28066 6554
rect 28066 6502 28078 6554
rect 28078 6502 28092 6554
rect 28116 6502 28130 6554
rect 28130 6502 28142 6554
rect 28142 6502 28172 6554
rect 28196 6502 28206 6554
rect 28206 6502 28252 6554
rect 27956 6500 28012 6502
rect 28036 6500 28092 6502
rect 28116 6500 28172 6502
rect 28196 6500 28252 6502
rect 27956 5466 28012 5468
rect 28036 5466 28092 5468
rect 28116 5466 28172 5468
rect 28196 5466 28252 5468
rect 27956 5414 28002 5466
rect 28002 5414 28012 5466
rect 28036 5414 28066 5466
rect 28066 5414 28078 5466
rect 28078 5414 28092 5466
rect 28116 5414 28130 5466
rect 28130 5414 28142 5466
rect 28142 5414 28172 5466
rect 28196 5414 28206 5466
rect 28206 5414 28252 5466
rect 27956 5412 28012 5414
rect 28036 5412 28092 5414
rect 28116 5412 28172 5414
rect 28196 5412 28252 5414
rect 27956 4378 28012 4380
rect 28036 4378 28092 4380
rect 28116 4378 28172 4380
rect 28196 4378 28252 4380
rect 27956 4326 28002 4378
rect 28002 4326 28012 4378
rect 28036 4326 28066 4378
rect 28066 4326 28078 4378
rect 28078 4326 28092 4378
rect 28116 4326 28130 4378
rect 28130 4326 28142 4378
rect 28142 4326 28172 4378
rect 28196 4326 28206 4378
rect 28206 4326 28252 4378
rect 27956 4324 28012 4326
rect 28036 4324 28092 4326
rect 28116 4324 28172 4326
rect 28196 4324 28252 4326
rect 27618 3440 27674 3496
rect 27956 3290 28012 3292
rect 28036 3290 28092 3292
rect 28116 3290 28172 3292
rect 28196 3290 28252 3292
rect 27956 3238 28002 3290
rect 28002 3238 28012 3290
rect 28036 3238 28066 3290
rect 28066 3238 28078 3290
rect 28078 3238 28092 3290
rect 28116 3238 28130 3290
rect 28130 3238 28142 3290
rect 28142 3238 28172 3290
rect 28196 3238 28206 3290
rect 28206 3238 28252 3290
rect 27956 3236 28012 3238
rect 28036 3236 28092 3238
rect 28116 3236 28172 3238
rect 28196 3236 28252 3238
rect 27956 2202 28012 2204
rect 28036 2202 28092 2204
rect 28116 2202 28172 2204
rect 28196 2202 28252 2204
rect 27956 2150 28002 2202
rect 28002 2150 28012 2202
rect 28036 2150 28066 2202
rect 28066 2150 28078 2202
rect 28078 2150 28092 2202
rect 28116 2150 28130 2202
rect 28130 2150 28142 2202
rect 28142 2150 28172 2202
rect 28196 2150 28206 2202
rect 28206 2150 28252 2202
rect 27956 2148 28012 2150
rect 28036 2148 28092 2150
rect 28116 2148 28172 2150
rect 28196 2148 28252 2150
rect 32126 23044 32182 23080
rect 32126 23024 32128 23044
rect 32128 23024 32180 23044
rect 32180 23024 32182 23044
rect 32218 20032 32274 20088
rect 32586 22888 32642 22944
rect 33138 24656 33194 24712
rect 32956 24506 33012 24508
rect 33036 24506 33092 24508
rect 33116 24506 33172 24508
rect 33196 24506 33252 24508
rect 32956 24454 33002 24506
rect 33002 24454 33012 24506
rect 33036 24454 33066 24506
rect 33066 24454 33078 24506
rect 33078 24454 33092 24506
rect 33116 24454 33130 24506
rect 33130 24454 33142 24506
rect 33142 24454 33172 24506
rect 33196 24454 33206 24506
rect 33206 24454 33252 24506
rect 32956 24452 33012 24454
rect 33036 24452 33092 24454
rect 33116 24452 33172 24454
rect 33196 24452 33252 24454
rect 32770 23568 32826 23624
rect 32494 21800 32550 21856
rect 32586 20168 32642 20224
rect 32218 14728 32274 14784
rect 31942 12416 31998 12472
rect 32956 23418 33012 23420
rect 33036 23418 33092 23420
rect 33116 23418 33172 23420
rect 33196 23418 33252 23420
rect 32956 23366 33002 23418
rect 33002 23366 33012 23418
rect 33036 23366 33066 23418
rect 33066 23366 33078 23418
rect 33078 23366 33092 23418
rect 33116 23366 33130 23418
rect 33130 23366 33142 23418
rect 33142 23366 33172 23418
rect 33196 23366 33206 23418
rect 33206 23366 33252 23418
rect 32956 23364 33012 23366
rect 33036 23364 33092 23366
rect 33116 23364 33172 23366
rect 33196 23364 33252 23366
rect 33690 23024 33746 23080
rect 32956 22330 33012 22332
rect 33036 22330 33092 22332
rect 33116 22330 33172 22332
rect 33196 22330 33252 22332
rect 32956 22278 33002 22330
rect 33002 22278 33012 22330
rect 33036 22278 33066 22330
rect 33066 22278 33078 22330
rect 33078 22278 33092 22330
rect 33116 22278 33130 22330
rect 33130 22278 33142 22330
rect 33142 22278 33172 22330
rect 33196 22278 33206 22330
rect 33206 22278 33252 22330
rect 32956 22276 33012 22278
rect 33036 22276 33092 22278
rect 33116 22276 33172 22278
rect 33196 22276 33252 22278
rect 34702 23316 34758 23352
rect 34702 23296 34704 23316
rect 34704 23296 34756 23316
rect 34756 23296 34758 23316
rect 34334 23024 34390 23080
rect 34150 21972 34152 21992
rect 34152 21972 34204 21992
rect 34204 21972 34206 21992
rect 34150 21936 34206 21972
rect 32956 21242 33012 21244
rect 33036 21242 33092 21244
rect 33116 21242 33172 21244
rect 33196 21242 33252 21244
rect 32956 21190 33002 21242
rect 33002 21190 33012 21242
rect 33036 21190 33066 21242
rect 33066 21190 33078 21242
rect 33078 21190 33092 21242
rect 33116 21190 33130 21242
rect 33130 21190 33142 21242
rect 33142 21190 33172 21242
rect 33196 21190 33206 21242
rect 33206 21190 33252 21242
rect 32956 21188 33012 21190
rect 33036 21188 33092 21190
rect 33116 21188 33172 21190
rect 33196 21188 33252 21190
rect 33782 21392 33838 21448
rect 33598 20168 33654 20224
rect 32956 20154 33012 20156
rect 33036 20154 33092 20156
rect 33116 20154 33172 20156
rect 33196 20154 33252 20156
rect 32956 20102 33002 20154
rect 33002 20102 33012 20154
rect 33036 20102 33066 20154
rect 33066 20102 33078 20154
rect 33078 20102 33092 20154
rect 33116 20102 33130 20154
rect 33130 20102 33142 20154
rect 33142 20102 33172 20154
rect 33196 20102 33206 20154
rect 33206 20102 33252 20154
rect 32956 20100 33012 20102
rect 33036 20100 33092 20102
rect 33116 20100 33172 20102
rect 33196 20100 33252 20102
rect 32956 19066 33012 19068
rect 33036 19066 33092 19068
rect 33116 19066 33172 19068
rect 33196 19066 33252 19068
rect 32956 19014 33002 19066
rect 33002 19014 33012 19066
rect 33036 19014 33066 19066
rect 33066 19014 33078 19066
rect 33078 19014 33092 19066
rect 33116 19014 33130 19066
rect 33130 19014 33142 19066
rect 33142 19014 33172 19066
rect 33196 19014 33206 19066
rect 33206 19014 33252 19066
rect 32956 19012 33012 19014
rect 33036 19012 33092 19014
rect 33116 19012 33172 19014
rect 33196 19012 33252 19014
rect 33046 18828 33102 18864
rect 33046 18808 33048 18828
rect 33048 18808 33100 18828
rect 33100 18808 33102 18828
rect 33046 18536 33102 18592
rect 32956 17978 33012 17980
rect 33036 17978 33092 17980
rect 33116 17978 33172 17980
rect 33196 17978 33252 17980
rect 32956 17926 33002 17978
rect 33002 17926 33012 17978
rect 33036 17926 33066 17978
rect 33066 17926 33078 17978
rect 33078 17926 33092 17978
rect 33116 17926 33130 17978
rect 33130 17926 33142 17978
rect 33142 17926 33172 17978
rect 33196 17926 33206 17978
rect 33206 17926 33252 17978
rect 32956 17924 33012 17926
rect 33036 17924 33092 17926
rect 33116 17924 33172 17926
rect 33196 17924 33252 17926
rect 32956 16890 33012 16892
rect 33036 16890 33092 16892
rect 33116 16890 33172 16892
rect 33196 16890 33252 16892
rect 32956 16838 33002 16890
rect 33002 16838 33012 16890
rect 33036 16838 33066 16890
rect 33066 16838 33078 16890
rect 33078 16838 33092 16890
rect 33116 16838 33130 16890
rect 33130 16838 33142 16890
rect 33142 16838 33172 16890
rect 33196 16838 33206 16890
rect 33206 16838 33252 16890
rect 32956 16836 33012 16838
rect 33036 16836 33092 16838
rect 33116 16836 33172 16838
rect 33196 16836 33252 16838
rect 32956 15802 33012 15804
rect 33036 15802 33092 15804
rect 33116 15802 33172 15804
rect 33196 15802 33252 15804
rect 32956 15750 33002 15802
rect 33002 15750 33012 15802
rect 33036 15750 33066 15802
rect 33066 15750 33078 15802
rect 33078 15750 33092 15802
rect 33116 15750 33130 15802
rect 33130 15750 33142 15802
rect 33142 15750 33172 15802
rect 33196 15750 33206 15802
rect 33206 15750 33252 15802
rect 32956 15748 33012 15750
rect 33036 15748 33092 15750
rect 33116 15748 33172 15750
rect 33196 15748 33252 15750
rect 32494 14456 32550 14512
rect 32034 11872 32090 11928
rect 31482 10920 31538 10976
rect 31850 8880 31906 8936
rect 32310 12416 32366 12472
rect 32586 13912 32642 13968
rect 32494 12280 32550 12336
rect 32494 12164 32550 12200
rect 32494 12144 32496 12164
rect 32496 12144 32548 12164
rect 32548 12144 32550 12164
rect 32310 11872 32366 11928
rect 32956 14714 33012 14716
rect 33036 14714 33092 14716
rect 33116 14714 33172 14716
rect 33196 14714 33252 14716
rect 32956 14662 33002 14714
rect 33002 14662 33012 14714
rect 33036 14662 33066 14714
rect 33066 14662 33078 14714
rect 33078 14662 33092 14714
rect 33116 14662 33130 14714
rect 33130 14662 33142 14714
rect 33142 14662 33172 14714
rect 33196 14662 33206 14714
rect 33206 14662 33252 14714
rect 32956 14660 33012 14662
rect 33036 14660 33092 14662
rect 33116 14660 33172 14662
rect 33196 14660 33252 14662
rect 34794 22480 34850 22536
rect 34518 20576 34574 20632
rect 33966 19352 34022 19408
rect 32956 13626 33012 13628
rect 33036 13626 33092 13628
rect 33116 13626 33172 13628
rect 33196 13626 33252 13628
rect 32956 13574 33002 13626
rect 33002 13574 33012 13626
rect 33036 13574 33066 13626
rect 33066 13574 33078 13626
rect 33078 13574 33092 13626
rect 33116 13574 33130 13626
rect 33130 13574 33142 13626
rect 33142 13574 33172 13626
rect 33196 13574 33206 13626
rect 33206 13574 33252 13626
rect 32956 13572 33012 13574
rect 33036 13572 33092 13574
rect 33116 13572 33172 13574
rect 33196 13572 33252 13574
rect 32956 12538 33012 12540
rect 33036 12538 33092 12540
rect 33116 12538 33172 12540
rect 33196 12538 33252 12540
rect 32956 12486 33002 12538
rect 33002 12486 33012 12538
rect 33036 12486 33066 12538
rect 33066 12486 33078 12538
rect 33078 12486 33092 12538
rect 33116 12486 33130 12538
rect 33130 12486 33142 12538
rect 33142 12486 33172 12538
rect 33196 12486 33206 12538
rect 33206 12486 33252 12538
rect 32956 12484 33012 12486
rect 33036 12484 33092 12486
rect 33116 12484 33172 12486
rect 33196 12484 33252 12486
rect 32954 12280 33010 12336
rect 32770 12144 32826 12200
rect 33322 12144 33378 12200
rect 32956 11450 33012 11452
rect 33036 11450 33092 11452
rect 33116 11450 33172 11452
rect 33196 11450 33252 11452
rect 32956 11398 33002 11450
rect 33002 11398 33012 11450
rect 33036 11398 33066 11450
rect 33066 11398 33078 11450
rect 33078 11398 33092 11450
rect 33116 11398 33130 11450
rect 33130 11398 33142 11450
rect 33142 11398 33172 11450
rect 33196 11398 33206 11450
rect 33206 11398 33252 11450
rect 32956 11396 33012 11398
rect 33036 11396 33092 11398
rect 33116 11396 33172 11398
rect 33196 11396 33252 11398
rect 32956 10362 33012 10364
rect 33036 10362 33092 10364
rect 33116 10362 33172 10364
rect 33196 10362 33252 10364
rect 32956 10310 33002 10362
rect 33002 10310 33012 10362
rect 33036 10310 33066 10362
rect 33066 10310 33078 10362
rect 33078 10310 33092 10362
rect 33116 10310 33130 10362
rect 33130 10310 33142 10362
rect 33142 10310 33172 10362
rect 33196 10310 33206 10362
rect 33206 10310 33252 10362
rect 32956 10308 33012 10310
rect 33036 10308 33092 10310
rect 33116 10308 33172 10310
rect 33196 10308 33252 10310
rect 33874 13388 33930 13424
rect 33874 13368 33876 13388
rect 33876 13368 33928 13388
rect 33928 13368 33930 13388
rect 33690 12164 33746 12200
rect 33690 12144 33692 12164
rect 33692 12144 33744 12164
rect 33744 12144 33746 12164
rect 33598 10104 33654 10160
rect 32956 9274 33012 9276
rect 33036 9274 33092 9276
rect 33116 9274 33172 9276
rect 33196 9274 33252 9276
rect 32956 9222 33002 9274
rect 33002 9222 33012 9274
rect 33036 9222 33066 9274
rect 33066 9222 33078 9274
rect 33078 9222 33092 9274
rect 33116 9222 33130 9274
rect 33130 9222 33142 9274
rect 33142 9222 33172 9274
rect 33196 9222 33206 9274
rect 33206 9222 33252 9274
rect 32956 9220 33012 9222
rect 33036 9220 33092 9222
rect 33116 9220 33172 9222
rect 33196 9220 33252 9222
rect 33782 10920 33838 10976
rect 33966 9968 34022 10024
rect 33598 9424 33654 9480
rect 32956 8186 33012 8188
rect 33036 8186 33092 8188
rect 33116 8186 33172 8188
rect 33196 8186 33252 8188
rect 32956 8134 33002 8186
rect 33002 8134 33012 8186
rect 33036 8134 33066 8186
rect 33066 8134 33078 8186
rect 33078 8134 33092 8186
rect 33116 8134 33130 8186
rect 33130 8134 33142 8186
rect 33142 8134 33172 8186
rect 33196 8134 33206 8186
rect 33206 8134 33252 8186
rect 32956 8132 33012 8134
rect 33036 8132 33092 8134
rect 33116 8132 33172 8134
rect 33196 8132 33252 8134
rect 32956 7098 33012 7100
rect 33036 7098 33092 7100
rect 33116 7098 33172 7100
rect 33196 7098 33252 7100
rect 32956 7046 33002 7098
rect 33002 7046 33012 7098
rect 33036 7046 33066 7098
rect 33066 7046 33078 7098
rect 33078 7046 33092 7098
rect 33116 7046 33130 7098
rect 33130 7046 33142 7098
rect 33142 7046 33172 7098
rect 33196 7046 33206 7098
rect 33206 7046 33252 7098
rect 32956 7044 33012 7046
rect 33036 7044 33092 7046
rect 33116 7044 33172 7046
rect 33196 7044 33252 7046
rect 32956 6010 33012 6012
rect 33036 6010 33092 6012
rect 33116 6010 33172 6012
rect 33196 6010 33252 6012
rect 32956 5958 33002 6010
rect 33002 5958 33012 6010
rect 33036 5958 33066 6010
rect 33066 5958 33078 6010
rect 33078 5958 33092 6010
rect 33116 5958 33130 6010
rect 33130 5958 33142 6010
rect 33142 5958 33172 6010
rect 33196 5958 33206 6010
rect 33206 5958 33252 6010
rect 32956 5956 33012 5958
rect 33036 5956 33092 5958
rect 33116 5956 33172 5958
rect 33196 5956 33252 5958
rect 32956 4922 33012 4924
rect 33036 4922 33092 4924
rect 33116 4922 33172 4924
rect 33196 4922 33252 4924
rect 32956 4870 33002 4922
rect 33002 4870 33012 4922
rect 33036 4870 33066 4922
rect 33066 4870 33078 4922
rect 33078 4870 33092 4922
rect 33116 4870 33130 4922
rect 33130 4870 33142 4922
rect 33142 4870 33172 4922
rect 33196 4870 33206 4922
rect 33206 4870 33252 4922
rect 32956 4868 33012 4870
rect 33036 4868 33092 4870
rect 33116 4868 33172 4870
rect 33196 4868 33252 4870
rect 32956 3834 33012 3836
rect 33036 3834 33092 3836
rect 33116 3834 33172 3836
rect 33196 3834 33252 3836
rect 32956 3782 33002 3834
rect 33002 3782 33012 3834
rect 33036 3782 33066 3834
rect 33066 3782 33078 3834
rect 33078 3782 33092 3834
rect 33116 3782 33130 3834
rect 33130 3782 33142 3834
rect 33142 3782 33172 3834
rect 33196 3782 33206 3834
rect 33206 3782 33252 3834
rect 32956 3780 33012 3782
rect 33036 3780 33092 3782
rect 33116 3780 33172 3782
rect 33196 3780 33252 3782
rect 34242 10920 34298 10976
rect 34426 18400 34482 18456
rect 36174 23160 36230 23216
rect 35806 23044 35862 23080
rect 35806 23024 35808 23044
rect 35808 23024 35860 23044
rect 35860 23024 35862 23044
rect 35438 22752 35494 22808
rect 35254 22380 35256 22400
rect 35256 22380 35308 22400
rect 35308 22380 35310 22400
rect 35254 22344 35310 22380
rect 35070 17720 35126 17776
rect 35254 18400 35310 18456
rect 34886 14184 34942 14240
rect 34702 13252 34758 13288
rect 34702 13232 34704 13252
rect 34704 13232 34756 13252
rect 34756 13232 34758 13252
rect 34334 10104 34390 10160
rect 36266 22888 36322 22944
rect 36174 22516 36176 22536
rect 36176 22516 36228 22536
rect 36228 22516 36230 22536
rect 36174 22480 36230 22516
rect 36174 22208 36230 22264
rect 36082 21800 36138 21856
rect 36542 23604 36544 23624
rect 36544 23604 36596 23624
rect 36596 23604 36598 23624
rect 36542 23568 36598 23604
rect 36634 23432 36690 23488
rect 36450 22616 36506 22672
rect 37094 23568 37150 23624
rect 35714 19488 35770 19544
rect 36542 18400 36598 18456
rect 36174 11736 36230 11792
rect 36174 11328 36230 11384
rect 37922 24792 37978 24848
rect 37956 23962 38012 23964
rect 38036 23962 38092 23964
rect 38116 23962 38172 23964
rect 38196 23962 38252 23964
rect 37956 23910 38002 23962
rect 38002 23910 38012 23962
rect 38036 23910 38066 23962
rect 38066 23910 38078 23962
rect 38078 23910 38092 23962
rect 38116 23910 38130 23962
rect 38130 23910 38142 23962
rect 38142 23910 38172 23962
rect 38196 23910 38206 23962
rect 38206 23910 38252 23962
rect 37956 23908 38012 23910
rect 38036 23908 38092 23910
rect 38116 23908 38172 23910
rect 38196 23908 38252 23910
rect 37738 22072 37794 22128
rect 37462 21800 37518 21856
rect 37462 21256 37518 21312
rect 37370 19624 37426 19680
rect 37462 18708 37464 18728
rect 37464 18708 37516 18728
rect 37516 18708 37518 18728
rect 37462 18672 37518 18708
rect 37956 22874 38012 22876
rect 38036 22874 38092 22876
rect 38116 22874 38172 22876
rect 38196 22874 38252 22876
rect 37956 22822 38002 22874
rect 38002 22822 38012 22874
rect 38036 22822 38066 22874
rect 38066 22822 38078 22874
rect 38078 22822 38092 22874
rect 38116 22822 38130 22874
rect 38130 22822 38142 22874
rect 38142 22822 38172 22874
rect 38196 22822 38206 22874
rect 38206 22822 38252 22874
rect 37956 22820 38012 22822
rect 38036 22820 38092 22822
rect 38116 22820 38172 22822
rect 38196 22820 38252 22822
rect 37956 21786 38012 21788
rect 38036 21786 38092 21788
rect 38116 21786 38172 21788
rect 38196 21786 38252 21788
rect 37956 21734 38002 21786
rect 38002 21734 38012 21786
rect 38036 21734 38066 21786
rect 38066 21734 38078 21786
rect 38078 21734 38092 21786
rect 38116 21734 38130 21786
rect 38130 21734 38142 21786
rect 38142 21734 38172 21786
rect 38196 21734 38206 21786
rect 38206 21734 38252 21786
rect 37956 21732 38012 21734
rect 38036 21732 38092 21734
rect 38116 21732 38172 21734
rect 38196 21732 38252 21734
rect 38382 23296 38438 23352
rect 43350 26288 43406 26344
rect 38658 24656 38714 24712
rect 38474 21936 38530 21992
rect 39026 22752 39082 22808
rect 39946 24792 40002 24848
rect 41234 24248 41290 24304
rect 40774 23568 40830 23624
rect 39670 21292 39672 21312
rect 39672 21292 39724 21312
rect 39724 21292 39726 21312
rect 39670 21256 39726 21292
rect 37956 20698 38012 20700
rect 38036 20698 38092 20700
rect 38116 20698 38172 20700
rect 38196 20698 38252 20700
rect 37956 20646 38002 20698
rect 38002 20646 38012 20698
rect 38036 20646 38066 20698
rect 38066 20646 38078 20698
rect 38078 20646 38092 20698
rect 38116 20646 38130 20698
rect 38130 20646 38142 20698
rect 38142 20646 38172 20698
rect 38196 20646 38206 20698
rect 38206 20646 38252 20698
rect 37956 20644 38012 20646
rect 38036 20644 38092 20646
rect 38116 20644 38172 20646
rect 38196 20644 38252 20646
rect 38382 19624 38438 19680
rect 37956 19610 38012 19612
rect 38036 19610 38092 19612
rect 38116 19610 38172 19612
rect 38196 19610 38252 19612
rect 37956 19558 38002 19610
rect 38002 19558 38012 19610
rect 38036 19558 38066 19610
rect 38066 19558 38078 19610
rect 38078 19558 38092 19610
rect 38116 19558 38130 19610
rect 38130 19558 38142 19610
rect 38142 19558 38172 19610
rect 38196 19558 38206 19610
rect 38206 19558 38252 19610
rect 37956 19556 38012 19558
rect 38036 19556 38092 19558
rect 38116 19556 38172 19558
rect 38196 19556 38252 19558
rect 37738 19488 37794 19544
rect 38382 19216 38438 19272
rect 37956 18522 38012 18524
rect 38036 18522 38092 18524
rect 38116 18522 38172 18524
rect 38196 18522 38252 18524
rect 37956 18470 38002 18522
rect 38002 18470 38012 18522
rect 38036 18470 38066 18522
rect 38066 18470 38078 18522
rect 38078 18470 38092 18522
rect 38116 18470 38130 18522
rect 38130 18470 38142 18522
rect 38142 18470 38172 18522
rect 38196 18470 38206 18522
rect 38206 18470 38252 18522
rect 37956 18468 38012 18470
rect 38036 18468 38092 18470
rect 38116 18468 38172 18470
rect 38196 18468 38252 18470
rect 37956 17434 38012 17436
rect 38036 17434 38092 17436
rect 38116 17434 38172 17436
rect 38196 17434 38252 17436
rect 37956 17382 38002 17434
rect 38002 17382 38012 17434
rect 38036 17382 38066 17434
rect 38066 17382 38078 17434
rect 38078 17382 38092 17434
rect 38116 17382 38130 17434
rect 38130 17382 38142 17434
rect 38142 17382 38172 17434
rect 38196 17382 38206 17434
rect 38206 17382 38252 17434
rect 37956 17380 38012 17382
rect 38036 17380 38092 17382
rect 38116 17380 38172 17382
rect 38196 17380 38252 17382
rect 37956 16346 38012 16348
rect 38036 16346 38092 16348
rect 38116 16346 38172 16348
rect 38196 16346 38252 16348
rect 37956 16294 38002 16346
rect 38002 16294 38012 16346
rect 38036 16294 38066 16346
rect 38066 16294 38078 16346
rect 38078 16294 38092 16346
rect 38116 16294 38130 16346
rect 38130 16294 38142 16346
rect 38142 16294 38172 16346
rect 38196 16294 38206 16346
rect 38206 16294 38252 16346
rect 37956 16292 38012 16294
rect 38036 16292 38092 16294
rect 38116 16292 38172 16294
rect 38196 16292 38252 16294
rect 37956 15258 38012 15260
rect 38036 15258 38092 15260
rect 38116 15258 38172 15260
rect 38196 15258 38252 15260
rect 37956 15206 38002 15258
rect 38002 15206 38012 15258
rect 38036 15206 38066 15258
rect 38066 15206 38078 15258
rect 38078 15206 38092 15258
rect 38116 15206 38130 15258
rect 38130 15206 38142 15258
rect 38142 15206 38172 15258
rect 38196 15206 38206 15258
rect 38206 15206 38252 15258
rect 37956 15204 38012 15206
rect 38036 15204 38092 15206
rect 38116 15204 38172 15206
rect 38196 15204 38252 15206
rect 37956 14170 38012 14172
rect 38036 14170 38092 14172
rect 38116 14170 38172 14172
rect 38196 14170 38252 14172
rect 37956 14118 38002 14170
rect 38002 14118 38012 14170
rect 38036 14118 38066 14170
rect 38066 14118 38078 14170
rect 38078 14118 38092 14170
rect 38116 14118 38130 14170
rect 38130 14118 38142 14170
rect 38142 14118 38172 14170
rect 38196 14118 38206 14170
rect 38206 14118 38252 14170
rect 37956 14116 38012 14118
rect 38036 14116 38092 14118
rect 38116 14116 38172 14118
rect 38196 14116 38252 14118
rect 39118 20032 39174 20088
rect 40590 23296 40646 23352
rect 41050 22616 41106 22672
rect 40682 22480 40738 22536
rect 40774 22108 40776 22128
rect 40776 22108 40828 22128
rect 40828 22108 40830 22128
rect 40774 22072 40830 22108
rect 40314 20304 40370 20360
rect 39946 20168 40002 20224
rect 40406 19760 40462 19816
rect 40590 17584 40646 17640
rect 41326 23432 41382 23488
rect 42956 24506 43012 24508
rect 43036 24506 43092 24508
rect 43116 24506 43172 24508
rect 43196 24506 43252 24508
rect 42956 24454 43002 24506
rect 43002 24454 43012 24506
rect 43036 24454 43066 24506
rect 43066 24454 43078 24506
rect 43078 24454 43092 24506
rect 43116 24454 43130 24506
rect 43130 24454 43142 24506
rect 43142 24454 43172 24506
rect 43196 24454 43206 24506
rect 43206 24454 43252 24506
rect 42956 24452 43012 24454
rect 43036 24452 43092 24454
rect 43116 24452 43172 24454
rect 43196 24452 43252 24454
rect 41878 22752 41934 22808
rect 41602 22380 41604 22400
rect 41604 22380 41656 22400
rect 41656 22380 41658 22400
rect 41602 22344 41658 22380
rect 41326 21800 41382 21856
rect 41602 21528 41658 21584
rect 42956 23418 43012 23420
rect 43036 23418 43092 23420
rect 43116 23418 43172 23420
rect 43196 23418 43252 23420
rect 42956 23366 43002 23418
rect 43002 23366 43012 23418
rect 43036 23366 43066 23418
rect 43066 23366 43078 23418
rect 43078 23366 43092 23418
rect 43116 23366 43130 23418
rect 43130 23366 43142 23418
rect 43142 23366 43172 23418
rect 43196 23366 43206 23418
rect 43206 23366 43252 23418
rect 42956 23364 43012 23366
rect 43036 23364 43092 23366
rect 43116 23364 43172 23366
rect 43196 23364 43252 23366
rect 46754 25064 46810 25120
rect 46662 24656 46718 24712
rect 45466 23724 45522 23760
rect 45466 23704 45468 23724
rect 45468 23704 45520 23724
rect 45520 23704 45522 23724
rect 43626 22616 43682 22672
rect 42956 22330 43012 22332
rect 43036 22330 43092 22332
rect 43116 22330 43172 22332
rect 43196 22330 43252 22332
rect 42956 22278 43002 22330
rect 43002 22278 43012 22330
rect 43036 22278 43066 22330
rect 43066 22278 43078 22330
rect 43078 22278 43092 22330
rect 43116 22278 43130 22330
rect 43130 22278 43142 22330
rect 43142 22278 43172 22330
rect 43196 22278 43206 22330
rect 43206 22278 43252 22330
rect 42956 22276 43012 22278
rect 43036 22276 43092 22278
rect 43116 22276 43172 22278
rect 43196 22276 43252 22278
rect 42798 21392 42854 21448
rect 42956 21242 43012 21244
rect 43036 21242 43092 21244
rect 43116 21242 43172 21244
rect 43196 21242 43252 21244
rect 42956 21190 43002 21242
rect 43002 21190 43012 21242
rect 43036 21190 43066 21242
rect 43066 21190 43078 21242
rect 43078 21190 43092 21242
rect 43116 21190 43130 21242
rect 43130 21190 43142 21242
rect 43142 21190 43172 21242
rect 43196 21190 43206 21242
rect 43206 21190 43252 21242
rect 42956 21188 43012 21190
rect 43036 21188 43092 21190
rect 43116 21188 43172 21190
rect 43196 21188 43252 21190
rect 43810 21936 43866 21992
rect 45190 22480 45246 22536
rect 44730 22072 44786 22128
rect 43994 20984 44050 21040
rect 43534 20848 43590 20904
rect 41694 20304 41750 20360
rect 42956 20154 43012 20156
rect 43036 20154 43092 20156
rect 43116 20154 43172 20156
rect 43196 20154 43252 20156
rect 42956 20102 43002 20154
rect 43002 20102 43012 20154
rect 43036 20102 43066 20154
rect 43066 20102 43078 20154
rect 43078 20102 43092 20154
rect 43116 20102 43130 20154
rect 43130 20102 43142 20154
rect 43142 20102 43172 20154
rect 43196 20102 43206 20154
rect 43206 20102 43252 20154
rect 42956 20100 43012 20102
rect 43036 20100 43092 20102
rect 43116 20100 43172 20102
rect 43196 20100 43252 20102
rect 41878 20032 41934 20088
rect 46294 23704 46350 23760
rect 48226 25472 48282 25528
rect 48318 24928 48374 24984
rect 48410 24248 48466 24304
rect 47956 23962 48012 23964
rect 48036 23962 48092 23964
rect 48116 23962 48172 23964
rect 48196 23962 48252 23964
rect 47956 23910 48002 23962
rect 48002 23910 48012 23962
rect 48036 23910 48066 23962
rect 48066 23910 48078 23962
rect 48078 23910 48092 23962
rect 48116 23910 48130 23962
rect 48130 23910 48142 23962
rect 48142 23910 48172 23962
rect 48196 23910 48206 23962
rect 48206 23910 48252 23962
rect 47956 23908 48012 23910
rect 48036 23908 48092 23910
rect 48116 23908 48172 23910
rect 48196 23908 48252 23910
rect 47858 23432 47914 23488
rect 48318 23060 48320 23080
rect 48320 23060 48372 23080
rect 48372 23060 48374 23080
rect 48318 23024 48374 23060
rect 46110 19624 46166 19680
rect 42956 19066 43012 19068
rect 43036 19066 43092 19068
rect 43116 19066 43172 19068
rect 43196 19066 43252 19068
rect 42956 19014 43002 19066
rect 43002 19014 43012 19066
rect 43036 19014 43066 19066
rect 43066 19014 43078 19066
rect 43078 19014 43092 19066
rect 43116 19014 43130 19066
rect 43130 19014 43142 19066
rect 43142 19014 43172 19066
rect 43196 19014 43206 19066
rect 43206 19014 43252 19066
rect 42956 19012 43012 19014
rect 43036 19012 43092 19014
rect 43116 19012 43172 19014
rect 43196 19012 43252 19014
rect 47956 22874 48012 22876
rect 48036 22874 48092 22876
rect 48116 22874 48172 22876
rect 48196 22874 48252 22876
rect 47956 22822 48002 22874
rect 48002 22822 48012 22874
rect 48036 22822 48066 22874
rect 48066 22822 48078 22874
rect 48078 22822 48092 22874
rect 48116 22822 48130 22874
rect 48130 22822 48142 22874
rect 48142 22822 48172 22874
rect 48196 22822 48206 22874
rect 48206 22822 48252 22874
rect 47956 22820 48012 22822
rect 48036 22820 48092 22822
rect 48116 22820 48172 22822
rect 48196 22820 48252 22822
rect 48594 24148 48596 24168
rect 48596 24148 48648 24168
rect 48648 24148 48650 24168
rect 48594 24112 48650 24148
rect 47956 21786 48012 21788
rect 48036 21786 48092 21788
rect 48116 21786 48172 21788
rect 48196 21786 48252 21788
rect 47956 21734 48002 21786
rect 48002 21734 48012 21786
rect 48036 21734 48066 21786
rect 48066 21734 48078 21786
rect 48078 21734 48092 21786
rect 48116 21734 48130 21786
rect 48130 21734 48142 21786
rect 48142 21734 48172 21786
rect 48196 21734 48206 21786
rect 48206 21734 48252 21786
rect 47956 21732 48012 21734
rect 48036 21732 48092 21734
rect 48116 21732 48172 21734
rect 48196 21732 48252 21734
rect 47956 20698 48012 20700
rect 48036 20698 48092 20700
rect 48116 20698 48172 20700
rect 48196 20698 48252 20700
rect 47956 20646 48002 20698
rect 48002 20646 48012 20698
rect 48036 20646 48066 20698
rect 48066 20646 48078 20698
rect 48078 20646 48092 20698
rect 48116 20646 48130 20698
rect 48130 20646 48142 20698
rect 48142 20646 48172 20698
rect 48196 20646 48206 20698
rect 48206 20646 48252 20698
rect 47956 20644 48012 20646
rect 48036 20644 48092 20646
rect 48116 20644 48172 20646
rect 48196 20644 48252 20646
rect 49146 22616 49202 22672
rect 49054 22208 49110 22264
rect 48594 21800 48650 21856
rect 48594 20168 48650 20224
rect 48502 19896 48558 19952
rect 47956 19610 48012 19612
rect 48036 19610 48092 19612
rect 48116 19610 48172 19612
rect 48196 19610 48252 19612
rect 47956 19558 48002 19610
rect 48002 19558 48012 19610
rect 48036 19558 48066 19610
rect 48066 19558 48078 19610
rect 48078 19558 48092 19610
rect 48116 19558 48130 19610
rect 48130 19558 48142 19610
rect 48142 19558 48172 19610
rect 48196 19558 48206 19610
rect 48206 19558 48252 19610
rect 47956 19556 48012 19558
rect 48036 19556 48092 19558
rect 48116 19556 48172 19558
rect 48196 19556 48252 19558
rect 49146 21392 49202 21448
rect 49054 20984 49110 21040
rect 49054 20576 49110 20632
rect 49054 19760 49110 19816
rect 48686 19352 48742 19408
rect 49330 19352 49386 19408
rect 47306 18808 47362 18864
rect 49146 18944 49202 19000
rect 47956 18522 48012 18524
rect 48036 18522 48092 18524
rect 48116 18522 48172 18524
rect 48196 18522 48252 18524
rect 47956 18470 48002 18522
rect 48002 18470 48012 18522
rect 48036 18470 48066 18522
rect 48066 18470 48078 18522
rect 48078 18470 48092 18522
rect 48116 18470 48130 18522
rect 48130 18470 48142 18522
rect 48142 18470 48172 18522
rect 48196 18470 48206 18522
rect 48206 18470 48252 18522
rect 47956 18468 48012 18470
rect 48036 18468 48092 18470
rect 48116 18468 48172 18470
rect 48196 18468 48252 18470
rect 41234 18264 41290 18320
rect 48594 18536 48650 18592
rect 42956 17978 43012 17980
rect 43036 17978 43092 17980
rect 43116 17978 43172 17980
rect 43196 17978 43252 17980
rect 42956 17926 43002 17978
rect 43002 17926 43012 17978
rect 43036 17926 43066 17978
rect 43066 17926 43078 17978
rect 43078 17926 43092 17978
rect 43116 17926 43130 17978
rect 43130 17926 43142 17978
rect 43142 17926 43172 17978
rect 43196 17926 43206 17978
rect 43206 17926 43252 17978
rect 42956 17924 43012 17926
rect 43036 17924 43092 17926
rect 43116 17924 43172 17926
rect 43196 17924 43252 17926
rect 41418 17176 41474 17232
rect 42956 16890 43012 16892
rect 43036 16890 43092 16892
rect 43116 16890 43172 16892
rect 43196 16890 43252 16892
rect 42956 16838 43002 16890
rect 43002 16838 43012 16890
rect 43036 16838 43066 16890
rect 43066 16838 43078 16890
rect 43078 16838 43092 16890
rect 43116 16838 43130 16890
rect 43130 16838 43142 16890
rect 43142 16838 43172 16890
rect 43196 16838 43206 16890
rect 43206 16838 43252 16890
rect 42956 16836 43012 16838
rect 43036 16836 43092 16838
rect 43116 16836 43172 16838
rect 43196 16836 43252 16838
rect 42956 15802 43012 15804
rect 43036 15802 43092 15804
rect 43116 15802 43172 15804
rect 43196 15802 43252 15804
rect 42956 15750 43002 15802
rect 43002 15750 43012 15802
rect 43036 15750 43066 15802
rect 43066 15750 43078 15802
rect 43078 15750 43092 15802
rect 43116 15750 43130 15802
rect 43130 15750 43142 15802
rect 43142 15750 43172 15802
rect 43196 15750 43206 15802
rect 43206 15750 43252 15802
rect 42956 15748 43012 15750
rect 43036 15748 43092 15750
rect 43116 15748 43172 15750
rect 43196 15748 43252 15750
rect 49146 18128 49202 18184
rect 49054 17720 49110 17776
rect 47956 17434 48012 17436
rect 48036 17434 48092 17436
rect 48116 17434 48172 17436
rect 48196 17434 48252 17436
rect 47956 17382 48002 17434
rect 48002 17382 48012 17434
rect 48036 17382 48066 17434
rect 48066 17382 48078 17434
rect 48078 17382 48092 17434
rect 48116 17382 48130 17434
rect 48130 17382 48142 17434
rect 48142 17382 48172 17434
rect 48196 17382 48206 17434
rect 48206 17382 48252 17434
rect 47956 17380 48012 17382
rect 48036 17380 48092 17382
rect 48116 17380 48172 17382
rect 48196 17380 48252 17382
rect 49054 17312 49110 17368
rect 48594 16904 48650 16960
rect 48226 16496 48282 16552
rect 47956 16346 48012 16348
rect 48036 16346 48092 16348
rect 48116 16346 48172 16348
rect 48196 16346 48252 16348
rect 47956 16294 48002 16346
rect 48002 16294 48012 16346
rect 48036 16294 48066 16346
rect 48066 16294 48078 16346
rect 48078 16294 48092 16346
rect 48116 16294 48130 16346
rect 48130 16294 48142 16346
rect 48142 16294 48172 16346
rect 48196 16294 48206 16346
rect 48206 16294 48252 16346
rect 47956 16292 48012 16294
rect 48036 16292 48092 16294
rect 48116 16292 48172 16294
rect 48196 16292 48252 16294
rect 49146 16088 49202 16144
rect 45558 15544 45614 15600
rect 47956 15258 48012 15260
rect 48036 15258 48092 15260
rect 48116 15258 48172 15260
rect 48196 15258 48252 15260
rect 47956 15206 48002 15258
rect 48002 15206 48012 15258
rect 48036 15206 48066 15258
rect 48066 15206 48078 15258
rect 48078 15206 48092 15258
rect 48116 15206 48130 15258
rect 48130 15206 48142 15258
rect 48142 15206 48172 15258
rect 48196 15206 48206 15258
rect 48206 15206 48252 15258
rect 47956 15204 48012 15206
rect 48036 15204 48092 15206
rect 48116 15204 48172 15206
rect 48196 15204 48252 15206
rect 48502 15000 48558 15056
rect 48318 14884 48374 14920
rect 48318 14864 48320 14884
rect 48320 14864 48372 14884
rect 48372 14864 48374 14884
rect 42956 14714 43012 14716
rect 43036 14714 43092 14716
rect 43116 14714 43172 14716
rect 43196 14714 43252 14716
rect 42956 14662 43002 14714
rect 43002 14662 43012 14714
rect 43036 14662 43066 14714
rect 43066 14662 43078 14714
rect 43078 14662 43092 14714
rect 43116 14662 43130 14714
rect 43130 14662 43142 14714
rect 43142 14662 43172 14714
rect 43196 14662 43206 14714
rect 43206 14662 43252 14714
rect 42956 14660 43012 14662
rect 43036 14660 43092 14662
rect 43116 14660 43172 14662
rect 43196 14660 43252 14662
rect 38474 13912 38530 13968
rect 36450 11056 36506 11112
rect 36542 10920 36598 10976
rect 47956 14170 48012 14172
rect 48036 14170 48092 14172
rect 48116 14170 48172 14172
rect 48196 14170 48252 14172
rect 47956 14118 48002 14170
rect 48002 14118 48012 14170
rect 48036 14118 48066 14170
rect 48066 14118 48078 14170
rect 48078 14118 48092 14170
rect 48116 14118 48130 14170
rect 48130 14118 48142 14170
rect 48142 14118 48172 14170
rect 48196 14118 48206 14170
rect 48206 14118 48252 14170
rect 47956 14116 48012 14118
rect 48036 14116 48092 14118
rect 48116 14116 48172 14118
rect 48196 14116 48252 14118
rect 42956 13626 43012 13628
rect 43036 13626 43092 13628
rect 43116 13626 43172 13628
rect 43196 13626 43252 13628
rect 42956 13574 43002 13626
rect 43002 13574 43012 13626
rect 43036 13574 43066 13626
rect 43066 13574 43078 13626
rect 43078 13574 43092 13626
rect 43116 13574 43130 13626
rect 43130 13574 43142 13626
rect 43142 13574 43172 13626
rect 43196 13574 43206 13626
rect 43206 13574 43252 13626
rect 42956 13572 43012 13574
rect 43036 13572 43092 13574
rect 43116 13572 43172 13574
rect 43196 13572 43252 13574
rect 37956 13082 38012 13084
rect 38036 13082 38092 13084
rect 38116 13082 38172 13084
rect 38196 13082 38252 13084
rect 37956 13030 38002 13082
rect 38002 13030 38012 13082
rect 38036 13030 38066 13082
rect 38066 13030 38078 13082
rect 38078 13030 38092 13082
rect 38116 13030 38130 13082
rect 38130 13030 38142 13082
rect 38142 13030 38172 13082
rect 38196 13030 38206 13082
rect 38206 13030 38252 13082
rect 37956 13028 38012 13030
rect 38036 13028 38092 13030
rect 38116 13028 38172 13030
rect 38196 13028 38252 13030
rect 37956 11994 38012 11996
rect 38036 11994 38092 11996
rect 38116 11994 38172 11996
rect 38196 11994 38252 11996
rect 37956 11942 38002 11994
rect 38002 11942 38012 11994
rect 38036 11942 38066 11994
rect 38066 11942 38078 11994
rect 38078 11942 38092 11994
rect 38116 11942 38130 11994
rect 38130 11942 38142 11994
rect 38142 11942 38172 11994
rect 38196 11942 38206 11994
rect 38206 11942 38252 11994
rect 37956 11940 38012 11942
rect 38036 11940 38092 11942
rect 38116 11940 38172 11942
rect 38196 11940 38252 11942
rect 49054 15680 49110 15736
rect 49238 15408 49294 15464
rect 49330 15272 49386 15328
rect 49054 14864 49110 14920
rect 49054 14456 49110 14512
rect 49238 14320 49294 14376
rect 49146 14048 49202 14104
rect 48226 13640 48282 13696
rect 49146 13268 49148 13288
rect 49148 13268 49200 13288
rect 49200 13268 49202 13288
rect 49146 13232 49202 13268
rect 47956 13082 48012 13084
rect 48036 13082 48092 13084
rect 48116 13082 48172 13084
rect 48196 13082 48252 13084
rect 47956 13030 48002 13082
rect 48002 13030 48012 13082
rect 48036 13030 48066 13082
rect 48066 13030 48078 13082
rect 48078 13030 48092 13082
rect 48116 13030 48130 13082
rect 48130 13030 48142 13082
rect 48142 13030 48172 13082
rect 48196 13030 48206 13082
rect 48206 13030 48252 13082
rect 47956 13028 48012 13030
rect 48036 13028 48092 13030
rect 48116 13028 48172 13030
rect 48196 13028 48252 13030
rect 49146 12844 49202 12880
rect 49146 12824 49148 12844
rect 49148 12824 49200 12844
rect 49200 12824 49202 12844
rect 46846 12688 46902 12744
rect 37956 10906 38012 10908
rect 38036 10906 38092 10908
rect 38116 10906 38172 10908
rect 38196 10906 38252 10908
rect 37956 10854 38002 10906
rect 38002 10854 38012 10906
rect 38036 10854 38066 10906
rect 38066 10854 38078 10906
rect 38078 10854 38092 10906
rect 38116 10854 38130 10906
rect 38130 10854 38142 10906
rect 38142 10854 38172 10906
rect 38196 10854 38206 10906
rect 38206 10854 38252 10906
rect 37956 10852 38012 10854
rect 38036 10852 38092 10854
rect 38116 10852 38172 10854
rect 38196 10852 38252 10854
rect 37956 9818 38012 9820
rect 38036 9818 38092 9820
rect 38116 9818 38172 9820
rect 38196 9818 38252 9820
rect 37956 9766 38002 9818
rect 38002 9766 38012 9818
rect 38036 9766 38066 9818
rect 38066 9766 38078 9818
rect 38078 9766 38092 9818
rect 38116 9766 38130 9818
rect 38130 9766 38142 9818
rect 38142 9766 38172 9818
rect 38196 9766 38206 9818
rect 38206 9766 38252 9818
rect 37956 9764 38012 9766
rect 38036 9764 38092 9766
rect 38116 9764 38172 9766
rect 38196 9764 38252 9766
rect 37956 8730 38012 8732
rect 38036 8730 38092 8732
rect 38116 8730 38172 8732
rect 38196 8730 38252 8732
rect 37956 8678 38002 8730
rect 38002 8678 38012 8730
rect 38036 8678 38066 8730
rect 38066 8678 38078 8730
rect 38078 8678 38092 8730
rect 38116 8678 38130 8730
rect 38130 8678 38142 8730
rect 38142 8678 38172 8730
rect 38196 8678 38206 8730
rect 38206 8678 38252 8730
rect 37956 8676 38012 8678
rect 38036 8676 38092 8678
rect 38116 8676 38172 8678
rect 38196 8676 38252 8678
rect 40130 11328 40186 11384
rect 39762 10104 39818 10160
rect 42956 12538 43012 12540
rect 43036 12538 43092 12540
rect 43116 12538 43172 12540
rect 43196 12538 43252 12540
rect 42956 12486 43002 12538
rect 43002 12486 43012 12538
rect 43036 12486 43066 12538
rect 43066 12486 43078 12538
rect 43078 12486 43092 12538
rect 43116 12486 43130 12538
rect 43130 12486 43142 12538
rect 43142 12486 43172 12538
rect 43196 12486 43206 12538
rect 43206 12486 43252 12538
rect 42956 12484 43012 12486
rect 43036 12484 43092 12486
rect 43116 12484 43172 12486
rect 43196 12484 43252 12486
rect 49146 12416 49202 12472
rect 42956 11450 43012 11452
rect 43036 11450 43092 11452
rect 43116 11450 43172 11452
rect 43196 11450 43252 11452
rect 42956 11398 43002 11450
rect 43002 11398 43012 11450
rect 43036 11398 43066 11450
rect 43066 11398 43078 11450
rect 43078 11398 43092 11450
rect 43116 11398 43130 11450
rect 43130 11398 43142 11450
rect 43142 11398 43172 11450
rect 43196 11398 43206 11450
rect 43206 11398 43252 11450
rect 42956 11396 43012 11398
rect 43036 11396 43092 11398
rect 43116 11396 43172 11398
rect 43196 11396 43252 11398
rect 42956 10362 43012 10364
rect 43036 10362 43092 10364
rect 43116 10362 43172 10364
rect 43196 10362 43252 10364
rect 42956 10310 43002 10362
rect 43002 10310 43012 10362
rect 43036 10310 43066 10362
rect 43066 10310 43078 10362
rect 43078 10310 43092 10362
rect 43116 10310 43130 10362
rect 43130 10310 43142 10362
rect 43142 10310 43172 10362
rect 43196 10310 43206 10362
rect 43206 10310 43252 10362
rect 42956 10308 43012 10310
rect 43036 10308 43092 10310
rect 43116 10308 43172 10310
rect 43196 10308 43252 10310
rect 38750 8880 38806 8936
rect 37956 7642 38012 7644
rect 38036 7642 38092 7644
rect 38116 7642 38172 7644
rect 38196 7642 38252 7644
rect 37956 7590 38002 7642
rect 38002 7590 38012 7642
rect 38036 7590 38066 7642
rect 38066 7590 38078 7642
rect 38078 7590 38092 7642
rect 38116 7590 38130 7642
rect 38130 7590 38142 7642
rect 38142 7590 38172 7642
rect 38196 7590 38206 7642
rect 38206 7590 38252 7642
rect 37956 7588 38012 7590
rect 38036 7588 38092 7590
rect 38116 7588 38172 7590
rect 38196 7588 38252 7590
rect 37956 6554 38012 6556
rect 38036 6554 38092 6556
rect 38116 6554 38172 6556
rect 38196 6554 38252 6556
rect 37956 6502 38002 6554
rect 38002 6502 38012 6554
rect 38036 6502 38066 6554
rect 38066 6502 38078 6554
rect 38078 6502 38092 6554
rect 38116 6502 38130 6554
rect 38130 6502 38142 6554
rect 38142 6502 38172 6554
rect 38196 6502 38206 6554
rect 38206 6502 38252 6554
rect 37956 6500 38012 6502
rect 38036 6500 38092 6502
rect 38116 6500 38172 6502
rect 38196 6500 38252 6502
rect 37956 5466 38012 5468
rect 38036 5466 38092 5468
rect 38116 5466 38172 5468
rect 38196 5466 38252 5468
rect 37956 5414 38002 5466
rect 38002 5414 38012 5466
rect 38036 5414 38066 5466
rect 38066 5414 38078 5466
rect 38078 5414 38092 5466
rect 38116 5414 38130 5466
rect 38130 5414 38142 5466
rect 38142 5414 38172 5466
rect 38196 5414 38206 5466
rect 38206 5414 38252 5466
rect 37956 5412 38012 5414
rect 38036 5412 38092 5414
rect 38116 5412 38172 5414
rect 38196 5412 38252 5414
rect 42956 9274 43012 9276
rect 43036 9274 43092 9276
rect 43116 9274 43172 9276
rect 43196 9274 43252 9276
rect 42956 9222 43002 9274
rect 43002 9222 43012 9274
rect 43036 9222 43066 9274
rect 43066 9222 43078 9274
rect 43078 9222 43092 9274
rect 43116 9222 43130 9274
rect 43130 9222 43142 9274
rect 43142 9222 43172 9274
rect 43196 9222 43206 9274
rect 43206 9222 43252 9274
rect 42956 9220 43012 9222
rect 43036 9220 43092 9222
rect 43116 9220 43172 9222
rect 43196 9220 43252 9222
rect 42956 8186 43012 8188
rect 43036 8186 43092 8188
rect 43116 8186 43172 8188
rect 43196 8186 43252 8188
rect 42956 8134 43002 8186
rect 43002 8134 43012 8186
rect 43036 8134 43066 8186
rect 43066 8134 43078 8186
rect 43078 8134 43092 8186
rect 43116 8134 43130 8186
rect 43130 8134 43142 8186
rect 43142 8134 43172 8186
rect 43196 8134 43206 8186
rect 43206 8134 43252 8186
rect 42956 8132 43012 8134
rect 43036 8132 43092 8134
rect 43116 8132 43172 8134
rect 43196 8132 43252 8134
rect 42956 7098 43012 7100
rect 43036 7098 43092 7100
rect 43116 7098 43172 7100
rect 43196 7098 43252 7100
rect 42956 7046 43002 7098
rect 43002 7046 43012 7098
rect 43036 7046 43066 7098
rect 43066 7046 43078 7098
rect 43078 7046 43092 7098
rect 43116 7046 43130 7098
rect 43130 7046 43142 7098
rect 43142 7046 43172 7098
rect 43196 7046 43206 7098
rect 43206 7046 43252 7098
rect 42956 7044 43012 7046
rect 43036 7044 43092 7046
rect 43116 7044 43172 7046
rect 43196 7044 43252 7046
rect 42956 6010 43012 6012
rect 43036 6010 43092 6012
rect 43116 6010 43172 6012
rect 43196 6010 43252 6012
rect 42956 5958 43002 6010
rect 43002 5958 43012 6010
rect 43036 5958 43066 6010
rect 43066 5958 43078 6010
rect 43078 5958 43092 6010
rect 43116 5958 43130 6010
rect 43130 5958 43142 6010
rect 43142 5958 43172 6010
rect 43196 5958 43206 6010
rect 43206 5958 43252 6010
rect 42956 5956 43012 5958
rect 43036 5956 43092 5958
rect 43116 5956 43172 5958
rect 43196 5956 43252 5958
rect 37956 4378 38012 4380
rect 38036 4378 38092 4380
rect 38116 4378 38172 4380
rect 38196 4378 38252 4380
rect 37956 4326 38002 4378
rect 38002 4326 38012 4378
rect 38036 4326 38066 4378
rect 38066 4326 38078 4378
rect 38078 4326 38092 4378
rect 38116 4326 38130 4378
rect 38130 4326 38142 4378
rect 38142 4326 38172 4378
rect 38196 4326 38206 4378
rect 38206 4326 38252 4378
rect 37956 4324 38012 4326
rect 38036 4324 38092 4326
rect 38116 4324 38172 4326
rect 38196 4324 38252 4326
rect 32956 2746 33012 2748
rect 33036 2746 33092 2748
rect 33116 2746 33172 2748
rect 33196 2746 33252 2748
rect 32956 2694 33002 2746
rect 33002 2694 33012 2746
rect 33036 2694 33066 2746
rect 33066 2694 33078 2746
rect 33078 2694 33092 2746
rect 33116 2694 33130 2746
rect 33130 2694 33142 2746
rect 33142 2694 33172 2746
rect 33196 2694 33206 2746
rect 33206 2694 33252 2746
rect 32956 2692 33012 2694
rect 33036 2692 33092 2694
rect 33116 2692 33172 2694
rect 33196 2692 33252 2694
rect 37956 3290 38012 3292
rect 38036 3290 38092 3292
rect 38116 3290 38172 3292
rect 38196 3290 38252 3292
rect 37956 3238 38002 3290
rect 38002 3238 38012 3290
rect 38036 3238 38066 3290
rect 38066 3238 38078 3290
rect 38078 3238 38092 3290
rect 38116 3238 38130 3290
rect 38130 3238 38142 3290
rect 38142 3238 38172 3290
rect 38196 3238 38206 3290
rect 38206 3238 38252 3290
rect 37956 3236 38012 3238
rect 38036 3236 38092 3238
rect 38116 3236 38172 3238
rect 38196 3236 38252 3238
rect 37956 2202 38012 2204
rect 38036 2202 38092 2204
rect 38116 2202 38172 2204
rect 38196 2202 38252 2204
rect 37956 2150 38002 2202
rect 38002 2150 38012 2202
rect 38036 2150 38066 2202
rect 38066 2150 38078 2202
rect 38078 2150 38092 2202
rect 38116 2150 38130 2202
rect 38130 2150 38142 2202
rect 38142 2150 38172 2202
rect 38196 2150 38206 2202
rect 38206 2150 38252 2202
rect 37956 2148 38012 2150
rect 38036 2148 38092 2150
rect 38116 2148 38172 2150
rect 38196 2148 38252 2150
rect 42956 4922 43012 4924
rect 43036 4922 43092 4924
rect 43116 4922 43172 4924
rect 43196 4922 43252 4924
rect 42956 4870 43002 4922
rect 43002 4870 43012 4922
rect 43036 4870 43066 4922
rect 43066 4870 43078 4922
rect 43078 4870 43092 4922
rect 43116 4870 43130 4922
rect 43130 4870 43142 4922
rect 43142 4870 43172 4922
rect 43196 4870 43206 4922
rect 43206 4870 43252 4922
rect 42956 4868 43012 4870
rect 43036 4868 43092 4870
rect 43116 4868 43172 4870
rect 43196 4868 43252 4870
rect 42956 3834 43012 3836
rect 43036 3834 43092 3836
rect 43116 3834 43172 3836
rect 43196 3834 43252 3836
rect 42956 3782 43002 3834
rect 43002 3782 43012 3834
rect 43036 3782 43066 3834
rect 43066 3782 43078 3834
rect 43078 3782 43092 3834
rect 43116 3782 43130 3834
rect 43130 3782 43142 3834
rect 43142 3782 43172 3834
rect 43196 3782 43206 3834
rect 43206 3782 43252 3834
rect 42956 3780 43012 3782
rect 43036 3780 43092 3782
rect 43116 3780 43172 3782
rect 43196 3780 43252 3782
rect 42956 2746 43012 2748
rect 43036 2746 43092 2748
rect 43116 2746 43172 2748
rect 43196 2746 43252 2748
rect 42956 2694 43002 2746
rect 43002 2694 43012 2746
rect 43036 2694 43066 2746
rect 43066 2694 43078 2746
rect 43078 2694 43092 2746
rect 43116 2694 43130 2746
rect 43130 2694 43142 2746
rect 43142 2694 43172 2746
rect 43196 2694 43206 2746
rect 43206 2694 43252 2746
rect 42956 2692 43012 2694
rect 43036 2692 43092 2694
rect 43116 2692 43172 2694
rect 43196 2692 43252 2694
rect 49146 12008 49202 12064
rect 47956 11994 48012 11996
rect 48036 11994 48092 11996
rect 48116 11994 48172 11996
rect 48196 11994 48252 11996
rect 47956 11942 48002 11994
rect 48002 11942 48012 11994
rect 48036 11942 48066 11994
rect 48066 11942 48078 11994
rect 48078 11942 48092 11994
rect 48116 11942 48130 11994
rect 48130 11942 48142 11994
rect 48142 11942 48172 11994
rect 48196 11942 48206 11994
rect 48206 11942 48252 11994
rect 47956 11940 48012 11942
rect 48036 11940 48092 11942
rect 48116 11940 48172 11942
rect 48196 11940 48252 11942
rect 49146 11600 49202 11656
rect 49238 11192 49294 11248
rect 47956 10906 48012 10908
rect 48036 10906 48092 10908
rect 48116 10906 48172 10908
rect 48196 10906 48252 10908
rect 47956 10854 48002 10906
rect 48002 10854 48012 10906
rect 48036 10854 48066 10906
rect 48066 10854 48078 10906
rect 48078 10854 48092 10906
rect 48116 10854 48130 10906
rect 48130 10854 48142 10906
rect 48142 10854 48172 10906
rect 48196 10854 48206 10906
rect 48206 10854 48252 10906
rect 47956 10852 48012 10854
rect 48036 10852 48092 10854
rect 48116 10852 48172 10854
rect 48196 10852 48252 10854
rect 49146 10784 49202 10840
rect 49330 10376 49386 10432
rect 49238 9968 49294 10024
rect 47956 9818 48012 9820
rect 48036 9818 48092 9820
rect 48116 9818 48172 9820
rect 48196 9818 48252 9820
rect 47956 9766 48002 9818
rect 48002 9766 48012 9818
rect 48036 9766 48066 9818
rect 48066 9766 48078 9818
rect 48078 9766 48092 9818
rect 48116 9766 48130 9818
rect 48130 9766 48142 9818
rect 48142 9766 48172 9818
rect 48196 9766 48206 9818
rect 48206 9766 48252 9818
rect 47956 9764 48012 9766
rect 48036 9764 48092 9766
rect 48116 9764 48172 9766
rect 48196 9764 48252 9766
rect 47306 9560 47362 9616
rect 49146 9152 49202 9208
rect 47956 8730 48012 8732
rect 48036 8730 48092 8732
rect 48116 8730 48172 8732
rect 48196 8730 48252 8732
rect 47956 8678 48002 8730
rect 48002 8678 48012 8730
rect 48036 8678 48066 8730
rect 48066 8678 48078 8730
rect 48078 8678 48092 8730
rect 48116 8678 48130 8730
rect 48130 8678 48142 8730
rect 48142 8678 48172 8730
rect 48196 8678 48206 8730
rect 48206 8678 48252 8730
rect 47956 8676 48012 8678
rect 48036 8676 48092 8678
rect 48116 8676 48172 8678
rect 48196 8676 48252 8678
rect 46846 7928 46902 7984
rect 46846 2624 46902 2680
rect 49238 8744 49294 8800
rect 49330 8336 49386 8392
rect 47956 7642 48012 7644
rect 48036 7642 48092 7644
rect 48116 7642 48172 7644
rect 48196 7642 48252 7644
rect 47956 7590 48002 7642
rect 48002 7590 48012 7642
rect 48036 7590 48066 7642
rect 48066 7590 48078 7642
rect 48078 7590 48092 7642
rect 48116 7590 48130 7642
rect 48130 7590 48142 7642
rect 48142 7590 48172 7642
rect 48196 7590 48206 7642
rect 48206 7590 48252 7642
rect 47956 7588 48012 7590
rect 48036 7588 48092 7590
rect 48116 7588 48172 7590
rect 48196 7588 48252 7590
rect 49146 7520 49202 7576
rect 49238 7112 49294 7168
rect 47956 6554 48012 6556
rect 48036 6554 48092 6556
rect 48116 6554 48172 6556
rect 48196 6554 48252 6556
rect 47956 6502 48002 6554
rect 48002 6502 48012 6554
rect 48036 6502 48066 6554
rect 48066 6502 48078 6554
rect 48078 6502 48092 6554
rect 48116 6502 48130 6554
rect 48130 6502 48142 6554
rect 48142 6502 48172 6554
rect 48196 6502 48206 6554
rect 48206 6502 48252 6554
rect 47956 6500 48012 6502
rect 48036 6500 48092 6502
rect 48116 6500 48172 6502
rect 48196 6500 48252 6502
rect 49422 6704 49478 6760
rect 48870 6296 48926 6352
rect 49146 5888 49202 5944
rect 47956 5466 48012 5468
rect 48036 5466 48092 5468
rect 48116 5466 48172 5468
rect 48196 5466 48252 5468
rect 47956 5414 48002 5466
rect 48002 5414 48012 5466
rect 48036 5414 48066 5466
rect 48066 5414 48078 5466
rect 48078 5414 48092 5466
rect 48116 5414 48130 5466
rect 48130 5414 48142 5466
rect 48142 5414 48172 5466
rect 48196 5414 48206 5466
rect 48206 5414 48252 5466
rect 47956 5412 48012 5414
rect 48036 5412 48092 5414
rect 48116 5412 48172 5414
rect 48196 5412 48252 5414
rect 49422 5480 49478 5536
rect 49330 5072 49386 5128
rect 48318 4664 48374 4720
rect 46754 1808 46810 1864
rect 46662 1400 46718 1456
rect 47956 4378 48012 4380
rect 48036 4378 48092 4380
rect 48116 4378 48172 4380
rect 48196 4378 48252 4380
rect 47956 4326 48002 4378
rect 48002 4326 48012 4378
rect 48036 4326 48066 4378
rect 48066 4326 48078 4378
rect 48078 4326 48092 4378
rect 48116 4326 48130 4378
rect 48130 4326 48142 4378
rect 48142 4326 48172 4378
rect 48196 4326 48206 4378
rect 48206 4326 48252 4378
rect 47956 4324 48012 4326
rect 48036 4324 48092 4326
rect 48116 4324 48172 4326
rect 48196 4324 48252 4326
rect 49146 4256 49202 4312
rect 49238 3848 49294 3904
rect 49146 3440 49202 3496
rect 47956 3290 48012 3292
rect 48036 3290 48092 3292
rect 48116 3290 48172 3292
rect 48196 3290 48252 3292
rect 47956 3238 48002 3290
rect 48002 3238 48012 3290
rect 48036 3238 48066 3290
rect 48066 3238 48078 3290
rect 48078 3238 48092 3290
rect 48116 3238 48130 3290
rect 48130 3238 48142 3290
rect 48142 3238 48172 3290
rect 48196 3238 48206 3290
rect 48206 3238 48252 3290
rect 47956 3236 48012 3238
rect 48036 3236 48092 3238
rect 48116 3236 48172 3238
rect 48196 3236 48252 3238
rect 48686 3032 48742 3088
rect 48502 2216 48558 2272
rect 47956 2202 48012 2204
rect 48036 2202 48092 2204
rect 48116 2202 48172 2204
rect 48196 2202 48252 2204
rect 47956 2150 48002 2202
rect 48002 2150 48012 2202
rect 48036 2150 48066 2202
rect 48066 2150 48078 2202
rect 48078 2150 48092 2202
rect 48116 2150 48130 2202
rect 48130 2150 48142 2202
rect 48142 2150 48172 2202
rect 48196 2150 48206 2202
rect 48206 2150 48252 2202
rect 47956 2148 48012 2150
rect 48036 2148 48092 2150
rect 48116 2148 48172 2150
rect 48196 2148 48252 2150
<< metal3 >>
rect 34513 26346 34579 26349
rect 43345 26346 43411 26349
rect 34513 26344 43411 26346
rect 34513 26288 34518 26344
rect 34574 26288 43350 26344
rect 43406 26288 43411 26344
rect 34513 26286 43411 26288
rect 34513 26283 34579 26286
rect 43345 26283 43411 26286
rect 0 25666 800 25696
rect 3417 25666 3483 25669
rect 0 25664 3483 25666
rect 0 25608 3422 25664
rect 3478 25608 3483 25664
rect 0 25606 3483 25608
rect 0 25576 800 25606
rect 3417 25603 3483 25606
rect 48221 25530 48287 25533
rect 50200 25530 51000 25560
rect 48221 25528 51000 25530
rect 48221 25472 48226 25528
rect 48282 25472 51000 25528
rect 48221 25470 51000 25472
rect 48221 25467 48287 25470
rect 50200 25440 51000 25470
rect 0 25258 800 25288
rect 3325 25258 3391 25261
rect 0 25256 3391 25258
rect 0 25200 3330 25256
rect 3386 25200 3391 25256
rect 0 25198 3391 25200
rect 0 25168 800 25198
rect 3325 25195 3391 25198
rect 46749 25122 46815 25125
rect 50200 25122 51000 25152
rect 46749 25120 51000 25122
rect 46749 25064 46754 25120
rect 46810 25064 51000 25120
rect 46749 25062 51000 25064
rect 46749 25059 46815 25062
rect 50200 25032 51000 25062
rect 35382 24924 35388 24988
rect 35452 24986 35458 24988
rect 48313 24986 48379 24989
rect 35452 24984 48379 24986
rect 35452 24928 48318 24984
rect 48374 24928 48379 24984
rect 35452 24926 48379 24928
rect 35452 24924 35458 24926
rect 48313 24923 48379 24926
rect 0 24850 800 24880
rect 3141 24850 3207 24853
rect 0 24848 3207 24850
rect 0 24792 3146 24848
rect 3202 24792 3207 24848
rect 0 24790 3207 24792
rect 0 24760 800 24790
rect 3141 24787 3207 24790
rect 26049 24850 26115 24853
rect 37917 24850 37983 24853
rect 39941 24850 40007 24853
rect 26049 24848 40007 24850
rect 26049 24792 26054 24848
rect 26110 24792 37922 24848
rect 37978 24792 39946 24848
rect 40002 24792 40007 24848
rect 26049 24790 40007 24792
rect 26049 24787 26115 24790
rect 37917 24787 37983 24790
rect 39941 24787 40007 24790
rect 7465 24714 7531 24717
rect 26325 24714 26391 24717
rect 7465 24712 26391 24714
rect 7465 24656 7470 24712
rect 7526 24656 26330 24712
rect 26386 24656 26391 24712
rect 7465 24654 26391 24656
rect 7465 24651 7531 24654
rect 26325 24651 26391 24654
rect 33133 24714 33199 24717
rect 38653 24714 38719 24717
rect 33133 24712 38719 24714
rect 33133 24656 33138 24712
rect 33194 24656 38658 24712
rect 38714 24656 38719 24712
rect 33133 24654 38719 24656
rect 33133 24651 33199 24654
rect 38653 24651 38719 24654
rect 46657 24714 46723 24717
rect 50200 24714 51000 24744
rect 46657 24712 51000 24714
rect 46657 24656 46662 24712
rect 46718 24656 51000 24712
rect 46657 24654 51000 24656
rect 46657 24651 46723 24654
rect 50200 24624 51000 24654
rect 2946 24512 3262 24513
rect 0 24442 800 24472
rect 2946 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3262 24512
rect 2946 24447 3262 24448
rect 12946 24512 13262 24513
rect 12946 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13262 24512
rect 12946 24447 13262 24448
rect 22946 24512 23262 24513
rect 22946 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23262 24512
rect 22946 24447 23262 24448
rect 32946 24512 33262 24513
rect 32946 24448 32952 24512
rect 33016 24448 33032 24512
rect 33096 24448 33112 24512
rect 33176 24448 33192 24512
rect 33256 24448 33262 24512
rect 32946 24447 33262 24448
rect 42946 24512 43262 24513
rect 42946 24448 42952 24512
rect 43016 24448 43032 24512
rect 43096 24448 43112 24512
rect 43176 24448 43192 24512
rect 43256 24448 43262 24512
rect 42946 24447 43262 24448
rect 2773 24442 2839 24445
rect 0 24440 2839 24442
rect 0 24384 2778 24440
rect 2834 24384 2839 24440
rect 0 24382 2839 24384
rect 0 24352 800 24382
rect 2773 24379 2839 24382
rect 32305 24306 32371 24309
rect 41229 24306 41295 24309
rect 32305 24304 41295 24306
rect 32305 24248 32310 24304
rect 32366 24248 41234 24304
rect 41290 24248 41295 24304
rect 32305 24246 41295 24248
rect 32305 24243 32371 24246
rect 41229 24243 41295 24246
rect 48405 24306 48471 24309
rect 50200 24306 51000 24336
rect 48405 24304 51000 24306
rect 48405 24248 48410 24304
rect 48466 24248 51000 24304
rect 48405 24246 51000 24248
rect 48405 24243 48471 24246
rect 50200 24216 51000 24246
rect 24945 24170 25011 24173
rect 48589 24170 48655 24173
rect 24945 24168 48655 24170
rect 24945 24112 24950 24168
rect 25006 24112 48594 24168
rect 48650 24112 48655 24168
rect 24945 24110 48655 24112
rect 24945 24107 25011 24110
rect 48589 24107 48655 24110
rect 0 24034 800 24064
rect 3693 24034 3759 24037
rect 0 24032 3759 24034
rect 0 23976 3698 24032
rect 3754 23976 3759 24032
rect 0 23974 3759 23976
rect 0 23944 800 23974
rect 3693 23971 3759 23974
rect 7946 23968 8262 23969
rect 7946 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8262 23968
rect 7946 23903 8262 23904
rect 17946 23968 18262 23969
rect 17946 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18262 23968
rect 17946 23903 18262 23904
rect 27946 23968 28262 23969
rect 27946 23904 27952 23968
rect 28016 23904 28032 23968
rect 28096 23904 28112 23968
rect 28176 23904 28192 23968
rect 28256 23904 28262 23968
rect 27946 23903 28262 23904
rect 37946 23968 38262 23969
rect 37946 23904 37952 23968
rect 38016 23904 38032 23968
rect 38096 23904 38112 23968
rect 38176 23904 38192 23968
rect 38256 23904 38262 23968
rect 37946 23903 38262 23904
rect 47946 23968 48262 23969
rect 47946 23904 47952 23968
rect 48016 23904 48032 23968
rect 48096 23904 48112 23968
rect 48176 23904 48192 23968
rect 48256 23904 48262 23968
rect 47946 23903 48262 23904
rect 50200 23898 51000 23928
rect 48454 23838 51000 23898
rect 28942 23700 28948 23764
rect 29012 23762 29018 23764
rect 45461 23762 45527 23765
rect 29012 23760 45527 23762
rect 29012 23704 45466 23760
rect 45522 23704 45527 23760
rect 29012 23702 45527 23704
rect 29012 23700 29018 23702
rect 45461 23699 45527 23702
rect 46289 23762 46355 23765
rect 48454 23762 48514 23838
rect 50200 23808 51000 23838
rect 46289 23760 48514 23762
rect 46289 23704 46294 23760
rect 46350 23704 48514 23760
rect 46289 23702 48514 23704
rect 46289 23699 46355 23702
rect 0 23626 800 23656
rect 3417 23626 3483 23629
rect 0 23624 3483 23626
rect 0 23568 3422 23624
rect 3478 23568 3483 23624
rect 0 23566 3483 23568
rect 0 23536 800 23566
rect 3417 23563 3483 23566
rect 16573 23626 16639 23629
rect 26233 23626 26299 23629
rect 16573 23624 26299 23626
rect 16573 23568 16578 23624
rect 16634 23568 26238 23624
rect 26294 23568 26299 23624
rect 16573 23566 26299 23568
rect 16573 23563 16639 23566
rect 26233 23563 26299 23566
rect 32765 23626 32831 23629
rect 36537 23626 36603 23629
rect 32765 23624 36603 23626
rect 32765 23568 32770 23624
rect 32826 23568 36542 23624
rect 36598 23568 36603 23624
rect 32765 23566 36603 23568
rect 32765 23563 32831 23566
rect 36537 23563 36603 23566
rect 37089 23626 37155 23629
rect 40769 23626 40835 23629
rect 37089 23624 40835 23626
rect 37089 23568 37094 23624
rect 37150 23568 40774 23624
rect 40830 23568 40835 23624
rect 37089 23566 40835 23568
rect 37089 23563 37155 23566
rect 40769 23563 40835 23566
rect 36629 23490 36695 23493
rect 41321 23490 41387 23493
rect 36629 23488 41387 23490
rect 36629 23432 36634 23488
rect 36690 23432 41326 23488
rect 41382 23432 41387 23488
rect 36629 23430 41387 23432
rect 36629 23427 36695 23430
rect 41321 23427 41387 23430
rect 47853 23490 47919 23493
rect 50200 23490 51000 23520
rect 47853 23488 51000 23490
rect 47853 23432 47858 23488
rect 47914 23432 51000 23488
rect 47853 23430 51000 23432
rect 47853 23427 47919 23430
rect 2946 23424 3262 23425
rect 2946 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3262 23424
rect 2946 23359 3262 23360
rect 12946 23424 13262 23425
rect 12946 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13262 23424
rect 12946 23359 13262 23360
rect 22946 23424 23262 23425
rect 22946 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23262 23424
rect 22946 23359 23262 23360
rect 32946 23424 33262 23425
rect 32946 23360 32952 23424
rect 33016 23360 33032 23424
rect 33096 23360 33112 23424
rect 33176 23360 33192 23424
rect 33256 23360 33262 23424
rect 32946 23359 33262 23360
rect 42946 23424 43262 23425
rect 42946 23360 42952 23424
rect 43016 23360 43032 23424
rect 43096 23360 43112 23424
rect 43176 23360 43192 23424
rect 43256 23360 43262 23424
rect 50200 23400 51000 23430
rect 42946 23359 43262 23360
rect 24761 23354 24827 23357
rect 27889 23354 27955 23357
rect 24761 23352 27955 23354
rect 24761 23296 24766 23352
rect 24822 23296 27894 23352
rect 27950 23296 27955 23352
rect 24761 23294 27955 23296
rect 24761 23291 24827 23294
rect 27889 23291 27955 23294
rect 34697 23354 34763 23357
rect 38377 23354 38443 23357
rect 40585 23354 40651 23357
rect 34697 23352 40651 23354
rect 34697 23296 34702 23352
rect 34758 23296 38382 23352
rect 38438 23296 40590 23352
rect 40646 23296 40651 23352
rect 34697 23294 40651 23296
rect 34697 23291 34763 23294
rect 38377 23291 38443 23294
rect 40585 23291 40651 23294
rect 0 23218 800 23248
rect 3325 23218 3391 23221
rect 0 23216 3391 23218
rect 0 23160 3330 23216
rect 3386 23160 3391 23216
rect 0 23158 3391 23160
rect 0 23128 800 23158
rect 3325 23155 3391 23158
rect 24945 23218 25011 23221
rect 28993 23218 29059 23221
rect 36169 23218 36235 23221
rect 24945 23216 29059 23218
rect 24945 23160 24950 23216
rect 25006 23160 28998 23216
rect 29054 23160 29059 23216
rect 24945 23158 29059 23160
rect 24945 23155 25011 23158
rect 28993 23155 29059 23158
rect 31710 23216 36235 23218
rect 31710 23160 36174 23216
rect 36230 23160 36235 23216
rect 31710 23158 36235 23160
rect 26693 23082 26759 23085
rect 31710 23082 31770 23158
rect 36169 23155 36235 23158
rect 26693 23080 31770 23082
rect 26693 23024 26698 23080
rect 26754 23024 31770 23080
rect 26693 23022 31770 23024
rect 32121 23082 32187 23085
rect 33685 23082 33751 23085
rect 34329 23082 34395 23085
rect 35801 23082 35867 23085
rect 32121 23080 35867 23082
rect 32121 23024 32126 23080
rect 32182 23024 33690 23080
rect 33746 23024 34334 23080
rect 34390 23024 35806 23080
rect 35862 23024 35867 23080
rect 32121 23022 35867 23024
rect 26693 23019 26759 23022
rect 32121 23019 32187 23022
rect 33685 23019 33751 23022
rect 34329 23019 34395 23022
rect 35801 23019 35867 23022
rect 48313 23082 48379 23085
rect 50200 23082 51000 23112
rect 48313 23080 51000 23082
rect 48313 23024 48318 23080
rect 48374 23024 51000 23080
rect 48313 23022 51000 23024
rect 48313 23019 48379 23022
rect 50200 22992 51000 23022
rect 32581 22946 32647 22949
rect 36261 22946 36327 22949
rect 32581 22944 36327 22946
rect 32581 22888 32586 22944
rect 32642 22888 36266 22944
rect 36322 22888 36327 22944
rect 32581 22886 36327 22888
rect 32581 22883 32647 22886
rect 36261 22883 36327 22886
rect 7946 22880 8262 22881
rect 0 22810 800 22840
rect 7946 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8262 22880
rect 7946 22815 8262 22816
rect 17946 22880 18262 22881
rect 17946 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18262 22880
rect 17946 22815 18262 22816
rect 27946 22880 28262 22881
rect 27946 22816 27952 22880
rect 28016 22816 28032 22880
rect 28096 22816 28112 22880
rect 28176 22816 28192 22880
rect 28256 22816 28262 22880
rect 27946 22815 28262 22816
rect 37946 22880 38262 22881
rect 37946 22816 37952 22880
rect 38016 22816 38032 22880
rect 38096 22816 38112 22880
rect 38176 22816 38192 22880
rect 38256 22816 38262 22880
rect 37946 22815 38262 22816
rect 47946 22880 48262 22881
rect 47946 22816 47952 22880
rect 48016 22816 48032 22880
rect 48096 22816 48112 22880
rect 48176 22816 48192 22880
rect 48256 22816 48262 22880
rect 47946 22815 48262 22816
rect 3417 22810 3483 22813
rect 0 22808 3483 22810
rect 0 22752 3422 22808
rect 3478 22752 3483 22808
rect 0 22750 3483 22752
rect 0 22720 800 22750
rect 3417 22747 3483 22750
rect 20529 22810 20595 22813
rect 22277 22810 22343 22813
rect 20529 22808 22343 22810
rect 20529 22752 20534 22808
rect 20590 22752 22282 22808
rect 22338 22752 22343 22808
rect 20529 22750 22343 22752
rect 20529 22747 20595 22750
rect 22277 22747 22343 22750
rect 31661 22810 31727 22813
rect 35433 22810 35499 22813
rect 31661 22808 35499 22810
rect 31661 22752 31666 22808
rect 31722 22752 35438 22808
rect 35494 22752 35499 22808
rect 31661 22750 35499 22752
rect 31661 22747 31727 22750
rect 35433 22747 35499 22750
rect 39021 22810 39087 22813
rect 41873 22810 41939 22813
rect 39021 22808 41939 22810
rect 39021 22752 39026 22808
rect 39082 22752 41878 22808
rect 41934 22752 41939 22808
rect 39021 22750 41939 22752
rect 39021 22747 39087 22750
rect 41873 22747 41939 22750
rect 12065 22674 12131 22677
rect 25589 22674 25655 22677
rect 12065 22672 25655 22674
rect 12065 22616 12070 22672
rect 12126 22616 25594 22672
rect 25650 22616 25655 22672
rect 12065 22614 25655 22616
rect 12065 22611 12131 22614
rect 25589 22611 25655 22614
rect 31109 22674 31175 22677
rect 36445 22674 36511 22677
rect 41045 22674 41111 22677
rect 43621 22674 43687 22677
rect 31109 22672 43687 22674
rect 31109 22616 31114 22672
rect 31170 22616 36450 22672
rect 36506 22616 41050 22672
rect 41106 22616 43626 22672
rect 43682 22616 43687 22672
rect 31109 22614 43687 22616
rect 31109 22611 31175 22614
rect 36445 22611 36511 22614
rect 41045 22611 41111 22614
rect 43621 22611 43687 22614
rect 49141 22674 49207 22677
rect 50200 22674 51000 22704
rect 49141 22672 51000 22674
rect 49141 22616 49146 22672
rect 49202 22616 51000 22672
rect 49141 22614 51000 22616
rect 49141 22611 49207 22614
rect 50200 22584 51000 22614
rect 4245 22538 4311 22541
rect 2454 22536 4311 22538
rect 2454 22480 4250 22536
rect 4306 22480 4311 22536
rect 2454 22478 4311 22480
rect 0 22402 800 22432
rect 2454 22402 2514 22478
rect 4245 22475 4311 22478
rect 29085 22538 29151 22541
rect 34789 22538 34855 22541
rect 29085 22536 34855 22538
rect 29085 22480 29090 22536
rect 29146 22480 34794 22536
rect 34850 22480 34855 22536
rect 29085 22478 34855 22480
rect 29085 22475 29151 22478
rect 34789 22475 34855 22478
rect 36169 22538 36235 22541
rect 40677 22538 40743 22541
rect 45185 22538 45251 22541
rect 36169 22536 45251 22538
rect 36169 22480 36174 22536
rect 36230 22480 40682 22536
rect 40738 22480 45190 22536
rect 45246 22480 45251 22536
rect 36169 22478 45251 22480
rect 36169 22475 36235 22478
rect 40677 22475 40743 22478
rect 45185 22475 45251 22478
rect 0 22342 2514 22402
rect 24669 22402 24735 22405
rect 31477 22402 31543 22405
rect 24669 22400 31543 22402
rect 24669 22344 24674 22400
rect 24730 22344 31482 22400
rect 31538 22344 31543 22400
rect 24669 22342 31543 22344
rect 0 22312 800 22342
rect 24669 22339 24735 22342
rect 31477 22339 31543 22342
rect 35249 22402 35315 22405
rect 41597 22402 41663 22405
rect 35249 22400 41663 22402
rect 35249 22344 35254 22400
rect 35310 22344 41602 22400
rect 41658 22344 41663 22400
rect 35249 22342 41663 22344
rect 35249 22339 35315 22342
rect 41597 22339 41663 22342
rect 2946 22336 3262 22337
rect 2946 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3262 22336
rect 2946 22271 3262 22272
rect 12946 22336 13262 22337
rect 12946 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13262 22336
rect 12946 22271 13262 22272
rect 22946 22336 23262 22337
rect 22946 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23262 22336
rect 22946 22271 23262 22272
rect 32946 22336 33262 22337
rect 32946 22272 32952 22336
rect 33016 22272 33032 22336
rect 33096 22272 33112 22336
rect 33176 22272 33192 22336
rect 33256 22272 33262 22336
rect 32946 22271 33262 22272
rect 42946 22336 43262 22337
rect 42946 22272 42952 22336
rect 43016 22272 43032 22336
rect 43096 22272 43112 22336
rect 43176 22272 43192 22336
rect 43256 22272 43262 22336
rect 42946 22271 43262 22272
rect 26417 22266 26483 22269
rect 30281 22266 30347 22269
rect 36169 22266 36235 22269
rect 49049 22266 49115 22269
rect 50200 22266 51000 22296
rect 26417 22264 30347 22266
rect 26417 22208 26422 22264
rect 26478 22208 30286 22264
rect 30342 22208 30347 22264
rect 26417 22206 30347 22208
rect 26417 22203 26483 22206
rect 30281 22203 30347 22206
rect 36126 22264 41430 22266
rect 36126 22208 36174 22264
rect 36230 22208 41430 22264
rect 36126 22206 41430 22208
rect 36126 22203 36235 22206
rect 27613 22130 27679 22133
rect 27797 22130 27863 22133
rect 27613 22128 27863 22130
rect 27613 22072 27618 22128
rect 27674 22072 27802 22128
rect 27858 22072 27863 22128
rect 27613 22070 27863 22072
rect 27613 22067 27679 22070
rect 27797 22067 27863 22070
rect 30741 22130 30807 22133
rect 36126 22130 36186 22203
rect 30741 22128 36186 22130
rect 30741 22072 30746 22128
rect 30802 22072 36186 22128
rect 30741 22070 36186 22072
rect 37733 22130 37799 22133
rect 40769 22130 40835 22133
rect 37733 22128 40835 22130
rect 37733 22072 37738 22128
rect 37794 22072 40774 22128
rect 40830 22072 40835 22128
rect 37733 22070 40835 22072
rect 41370 22130 41430 22206
rect 49049 22264 51000 22266
rect 49049 22208 49054 22264
rect 49110 22208 51000 22264
rect 49049 22206 51000 22208
rect 49049 22203 49115 22206
rect 50200 22176 51000 22206
rect 44725 22130 44791 22133
rect 41370 22128 44791 22130
rect 41370 22072 44730 22128
rect 44786 22072 44791 22128
rect 41370 22070 44791 22072
rect 30741 22067 30807 22070
rect 37733 22067 37799 22070
rect 40769 22067 40835 22070
rect 44725 22067 44791 22070
rect 0 21994 800 22024
rect 3785 21994 3851 21997
rect 0 21992 3851 21994
rect 0 21936 3790 21992
rect 3846 21936 3851 21992
rect 0 21934 3851 21936
rect 0 21904 800 21934
rect 3785 21931 3851 21934
rect 12065 21994 12131 21997
rect 23381 21994 23447 21997
rect 12065 21992 23447 21994
rect 12065 21936 12070 21992
rect 12126 21936 23386 21992
rect 23442 21936 23447 21992
rect 12065 21934 23447 21936
rect 12065 21931 12131 21934
rect 23381 21931 23447 21934
rect 29913 21994 29979 21997
rect 34145 21994 34211 21997
rect 38469 21994 38535 21997
rect 43805 21994 43871 21997
rect 29913 21992 34211 21994
rect 29913 21936 29918 21992
rect 29974 21936 34150 21992
rect 34206 21936 34211 21992
rect 29913 21934 34211 21936
rect 29913 21931 29979 21934
rect 34145 21931 34211 21934
rect 34286 21934 38394 21994
rect 22277 21858 22343 21861
rect 26601 21858 26667 21861
rect 22277 21856 26667 21858
rect 22277 21800 22282 21856
rect 22338 21800 26606 21856
rect 26662 21800 26667 21856
rect 22277 21798 26667 21800
rect 22277 21795 22343 21798
rect 26601 21795 26667 21798
rect 28441 21858 28507 21861
rect 28809 21858 28875 21861
rect 28441 21856 28875 21858
rect 28441 21800 28446 21856
rect 28502 21800 28814 21856
rect 28870 21800 28875 21856
rect 28441 21798 28875 21800
rect 28441 21795 28507 21798
rect 28809 21795 28875 21798
rect 32489 21858 32555 21861
rect 34286 21858 34346 21934
rect 32489 21856 34346 21858
rect 32489 21800 32494 21856
rect 32550 21800 34346 21856
rect 32489 21798 34346 21800
rect 36077 21858 36143 21861
rect 37457 21858 37523 21861
rect 36077 21856 37523 21858
rect 36077 21800 36082 21856
rect 36138 21800 37462 21856
rect 37518 21800 37523 21856
rect 36077 21798 37523 21800
rect 38334 21858 38394 21934
rect 38469 21992 43871 21994
rect 38469 21936 38474 21992
rect 38530 21936 43810 21992
rect 43866 21936 43871 21992
rect 38469 21934 43871 21936
rect 38469 21931 38535 21934
rect 43805 21931 43871 21934
rect 41321 21858 41387 21861
rect 38334 21856 41387 21858
rect 38334 21800 41326 21856
rect 41382 21800 41387 21856
rect 38334 21798 41387 21800
rect 32489 21795 32555 21798
rect 36077 21795 36143 21798
rect 37457 21795 37523 21798
rect 41321 21795 41387 21798
rect 48589 21858 48655 21861
rect 50200 21858 51000 21888
rect 48589 21856 51000 21858
rect 48589 21800 48594 21856
rect 48650 21800 51000 21856
rect 48589 21798 51000 21800
rect 48589 21795 48655 21798
rect 7946 21792 8262 21793
rect 7946 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8262 21792
rect 7946 21727 8262 21728
rect 17946 21792 18262 21793
rect 17946 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18262 21792
rect 17946 21727 18262 21728
rect 27946 21792 28262 21793
rect 27946 21728 27952 21792
rect 28016 21728 28032 21792
rect 28096 21728 28112 21792
rect 28176 21728 28192 21792
rect 28256 21728 28262 21792
rect 27946 21727 28262 21728
rect 37946 21792 38262 21793
rect 37946 21728 37952 21792
rect 38016 21728 38032 21792
rect 38096 21728 38112 21792
rect 38176 21728 38192 21792
rect 38256 21728 38262 21792
rect 37946 21727 38262 21728
rect 47946 21792 48262 21793
rect 47946 21728 47952 21792
rect 48016 21728 48032 21792
rect 48096 21728 48112 21792
rect 48176 21728 48192 21792
rect 48256 21728 48262 21792
rect 50200 21768 51000 21798
rect 47946 21727 48262 21728
rect 0 21586 800 21616
rect 2681 21586 2747 21589
rect 0 21584 2747 21586
rect 0 21528 2686 21584
rect 2742 21528 2747 21584
rect 0 21526 2747 21528
rect 0 21496 800 21526
rect 2681 21523 2747 21526
rect 27705 21586 27771 21589
rect 28942 21586 28948 21588
rect 27705 21584 28948 21586
rect 27705 21528 27710 21584
rect 27766 21528 28948 21584
rect 27705 21526 28948 21528
rect 27705 21523 27771 21526
rect 28942 21524 28948 21526
rect 29012 21524 29018 21588
rect 41597 21586 41663 21589
rect 31710 21584 41663 21586
rect 31710 21528 41602 21584
rect 41658 21528 41663 21584
rect 31710 21526 41663 21528
rect 25129 21450 25195 21453
rect 31710 21450 31770 21526
rect 41597 21523 41663 21526
rect 25129 21448 31770 21450
rect 25129 21392 25134 21448
rect 25190 21392 31770 21448
rect 25129 21390 31770 21392
rect 33777 21450 33843 21453
rect 42793 21450 42859 21453
rect 33777 21448 42859 21450
rect 33777 21392 33782 21448
rect 33838 21392 42798 21448
rect 42854 21392 42859 21448
rect 33777 21390 42859 21392
rect 25129 21387 25195 21390
rect 33777 21387 33843 21390
rect 42793 21387 42859 21390
rect 49141 21450 49207 21453
rect 50200 21450 51000 21480
rect 49141 21448 51000 21450
rect 49141 21392 49146 21448
rect 49202 21392 51000 21448
rect 49141 21390 51000 21392
rect 49141 21387 49207 21390
rect 50200 21360 51000 21390
rect 28533 21314 28599 21317
rect 29913 21314 29979 21317
rect 28533 21312 29979 21314
rect 28533 21256 28538 21312
rect 28594 21256 29918 21312
rect 29974 21256 29979 21312
rect 28533 21254 29979 21256
rect 28533 21251 28599 21254
rect 29913 21251 29979 21254
rect 37457 21314 37523 21317
rect 39665 21314 39731 21317
rect 37457 21312 39731 21314
rect 37457 21256 37462 21312
rect 37518 21256 39670 21312
rect 39726 21256 39731 21312
rect 37457 21254 39731 21256
rect 37457 21251 37523 21254
rect 39665 21251 39731 21254
rect 2946 21248 3262 21249
rect 0 21178 800 21208
rect 2946 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3262 21248
rect 2946 21183 3262 21184
rect 12946 21248 13262 21249
rect 12946 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13262 21248
rect 12946 21183 13262 21184
rect 22946 21248 23262 21249
rect 22946 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23262 21248
rect 22946 21183 23262 21184
rect 32946 21248 33262 21249
rect 32946 21184 32952 21248
rect 33016 21184 33032 21248
rect 33096 21184 33112 21248
rect 33176 21184 33192 21248
rect 33256 21184 33262 21248
rect 32946 21183 33262 21184
rect 42946 21248 43262 21249
rect 42946 21184 42952 21248
rect 43016 21184 43032 21248
rect 43096 21184 43112 21248
rect 43176 21184 43192 21248
rect 43256 21184 43262 21248
rect 42946 21183 43262 21184
rect 2773 21178 2839 21181
rect 0 21176 2839 21178
rect 0 21120 2778 21176
rect 2834 21120 2839 21176
rect 0 21118 2839 21120
rect 0 21088 800 21118
rect 2773 21115 2839 21118
rect 27337 21178 27403 21181
rect 30281 21178 30347 21181
rect 27337 21176 30347 21178
rect 27337 21120 27342 21176
rect 27398 21120 30286 21176
rect 30342 21120 30347 21176
rect 27337 21118 30347 21120
rect 27337 21115 27403 21118
rect 30281 21115 30347 21118
rect 11145 21042 11211 21045
rect 22185 21042 22251 21045
rect 11145 21040 22251 21042
rect 11145 20984 11150 21040
rect 11206 20984 22190 21040
rect 22246 20984 22251 21040
rect 11145 20982 22251 20984
rect 11145 20979 11211 20982
rect 22185 20979 22251 20982
rect 26417 21042 26483 21045
rect 29453 21042 29519 21045
rect 26417 21040 29519 21042
rect 26417 20984 26422 21040
rect 26478 20984 29458 21040
rect 29514 20984 29519 21040
rect 26417 20982 29519 20984
rect 26417 20979 26483 20982
rect 29453 20979 29519 20982
rect 29913 21042 29979 21045
rect 43989 21042 44055 21045
rect 29913 21040 44055 21042
rect 29913 20984 29918 21040
rect 29974 20984 43994 21040
rect 44050 20984 44055 21040
rect 29913 20982 44055 20984
rect 29913 20979 29979 20982
rect 43989 20979 44055 20982
rect 49049 21042 49115 21045
rect 50200 21042 51000 21072
rect 49049 21040 51000 21042
rect 49049 20984 49054 21040
rect 49110 20984 51000 21040
rect 49049 20982 51000 20984
rect 49049 20979 49115 20982
rect 50200 20952 51000 20982
rect 12433 20906 12499 20909
rect 25037 20906 25103 20909
rect 27613 20906 27679 20909
rect 12433 20904 27679 20906
rect 12433 20848 12438 20904
rect 12494 20848 25042 20904
rect 25098 20848 27618 20904
rect 27674 20848 27679 20904
rect 12433 20846 27679 20848
rect 12433 20843 12499 20846
rect 25037 20843 25103 20846
rect 27613 20843 27679 20846
rect 28349 20906 28415 20909
rect 31109 20906 31175 20909
rect 43529 20906 43595 20909
rect 28349 20904 31175 20906
rect 28349 20848 28354 20904
rect 28410 20848 31114 20904
rect 31170 20848 31175 20904
rect 28349 20846 31175 20848
rect 28349 20843 28415 20846
rect 31109 20843 31175 20846
rect 31710 20904 43595 20906
rect 31710 20848 43534 20904
rect 43590 20848 43595 20904
rect 31710 20846 43595 20848
rect 0 20770 800 20800
rect 1301 20770 1367 20773
rect 0 20768 1367 20770
rect 0 20712 1306 20768
rect 1362 20712 1367 20768
rect 0 20710 1367 20712
rect 0 20680 800 20710
rect 1301 20707 1367 20710
rect 11697 20770 11763 20773
rect 16481 20770 16547 20773
rect 11697 20768 16547 20770
rect 11697 20712 11702 20768
rect 11758 20712 16486 20768
rect 16542 20712 16547 20768
rect 11697 20710 16547 20712
rect 11697 20707 11763 20710
rect 16481 20707 16547 20710
rect 24209 20770 24275 20773
rect 27705 20770 27771 20773
rect 24209 20768 27771 20770
rect 24209 20712 24214 20768
rect 24270 20712 27710 20768
rect 27766 20712 27771 20768
rect 24209 20710 27771 20712
rect 24209 20707 24275 20710
rect 27705 20707 27771 20710
rect 29453 20770 29519 20773
rect 31710 20770 31770 20846
rect 43529 20843 43595 20846
rect 29453 20768 31770 20770
rect 29453 20712 29458 20768
rect 29514 20712 31770 20768
rect 29453 20710 31770 20712
rect 29453 20707 29519 20710
rect 7946 20704 8262 20705
rect 7946 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8262 20704
rect 7946 20639 8262 20640
rect 17946 20704 18262 20705
rect 17946 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18262 20704
rect 17946 20639 18262 20640
rect 27946 20704 28262 20705
rect 27946 20640 27952 20704
rect 28016 20640 28032 20704
rect 28096 20640 28112 20704
rect 28176 20640 28192 20704
rect 28256 20640 28262 20704
rect 27946 20639 28262 20640
rect 37946 20704 38262 20705
rect 37946 20640 37952 20704
rect 38016 20640 38032 20704
rect 38096 20640 38112 20704
rect 38176 20640 38192 20704
rect 38256 20640 38262 20704
rect 37946 20639 38262 20640
rect 47946 20704 48262 20705
rect 47946 20640 47952 20704
rect 48016 20640 48032 20704
rect 48096 20640 48112 20704
rect 48176 20640 48192 20704
rect 48256 20640 48262 20704
rect 47946 20639 48262 20640
rect 19149 20634 19215 20637
rect 31109 20634 31175 20637
rect 34513 20634 34579 20637
rect 35382 20634 35388 20636
rect 19149 20632 25882 20634
rect 19149 20576 19154 20632
rect 19210 20576 25882 20632
rect 19149 20574 25882 20576
rect 19149 20571 19215 20574
rect 25822 20501 25882 20574
rect 31109 20632 32138 20634
rect 31109 20576 31114 20632
rect 31170 20576 32138 20632
rect 31109 20574 32138 20576
rect 31109 20571 31175 20574
rect 13629 20498 13695 20501
rect 21173 20498 21239 20501
rect 25129 20498 25195 20501
rect 13629 20496 25195 20498
rect 13629 20440 13634 20496
rect 13690 20440 21178 20496
rect 21234 20440 25134 20496
rect 25190 20440 25195 20496
rect 13629 20438 25195 20440
rect 25822 20498 25931 20501
rect 32078 20498 32138 20574
rect 34513 20632 35388 20634
rect 34513 20576 34518 20632
rect 34574 20576 35388 20632
rect 34513 20574 35388 20576
rect 34513 20571 34579 20574
rect 35382 20572 35388 20574
rect 35452 20572 35458 20636
rect 49049 20634 49115 20637
rect 50200 20634 51000 20664
rect 49049 20632 51000 20634
rect 49049 20576 49054 20632
rect 49110 20576 51000 20632
rect 49049 20574 51000 20576
rect 49049 20571 49115 20574
rect 50200 20544 51000 20574
rect 25822 20496 31954 20498
rect 25822 20440 25870 20496
rect 25926 20440 31954 20496
rect 25822 20438 31954 20440
rect 32078 20438 41430 20498
rect 13629 20435 13695 20438
rect 21173 20435 21239 20438
rect 25129 20435 25195 20438
rect 25865 20435 25931 20438
rect 0 20362 800 20392
rect 3877 20362 3943 20365
rect 0 20360 3943 20362
rect 0 20304 3882 20360
rect 3938 20304 3943 20360
rect 0 20302 3943 20304
rect 0 20272 800 20302
rect 3877 20299 3943 20302
rect 15377 20362 15443 20365
rect 26141 20362 26207 20365
rect 15377 20360 26207 20362
rect 15377 20304 15382 20360
rect 15438 20304 26146 20360
rect 26202 20304 26207 20360
rect 15377 20302 26207 20304
rect 15377 20299 15443 20302
rect 26141 20299 26207 20302
rect 28533 20364 28599 20365
rect 28533 20360 28580 20364
rect 28644 20362 28650 20364
rect 29637 20362 29703 20365
rect 30097 20362 30163 20365
rect 28533 20304 28538 20360
rect 28533 20300 28580 20304
rect 28644 20302 28690 20362
rect 29637 20360 30163 20362
rect 29637 20304 29642 20360
rect 29698 20304 30102 20360
rect 30158 20304 30163 20360
rect 29637 20302 30163 20304
rect 31894 20362 31954 20438
rect 40309 20362 40375 20365
rect 31894 20360 40375 20362
rect 31894 20304 40314 20360
rect 40370 20304 40375 20360
rect 31894 20302 40375 20304
rect 41370 20362 41430 20438
rect 41689 20362 41755 20365
rect 41370 20360 41755 20362
rect 41370 20304 41694 20360
rect 41750 20304 41755 20360
rect 41370 20302 41755 20304
rect 28644 20300 28650 20302
rect 28533 20299 28599 20300
rect 29637 20299 29703 20302
rect 30097 20299 30163 20302
rect 40309 20299 40375 20302
rect 41689 20299 41755 20302
rect 25957 20226 26023 20229
rect 28441 20226 28507 20229
rect 32581 20226 32647 20229
rect 25957 20224 32647 20226
rect 25957 20168 25962 20224
rect 26018 20168 28446 20224
rect 28502 20168 32586 20224
rect 32642 20168 32647 20224
rect 25957 20166 32647 20168
rect 25957 20163 26023 20166
rect 28441 20163 28507 20166
rect 32581 20163 32647 20166
rect 33593 20226 33659 20229
rect 39941 20226 40007 20229
rect 33593 20224 40007 20226
rect 33593 20168 33598 20224
rect 33654 20168 39946 20224
rect 40002 20168 40007 20224
rect 33593 20166 40007 20168
rect 33593 20163 33659 20166
rect 39941 20163 40007 20166
rect 48589 20226 48655 20229
rect 50200 20226 51000 20256
rect 48589 20224 51000 20226
rect 48589 20168 48594 20224
rect 48650 20168 51000 20224
rect 48589 20166 51000 20168
rect 48589 20163 48655 20166
rect 2946 20160 3262 20161
rect 2946 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3262 20160
rect 2946 20095 3262 20096
rect 12946 20160 13262 20161
rect 12946 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13262 20160
rect 12946 20095 13262 20096
rect 22946 20160 23262 20161
rect 22946 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23262 20160
rect 22946 20095 23262 20096
rect 32946 20160 33262 20161
rect 32946 20096 32952 20160
rect 33016 20096 33032 20160
rect 33096 20096 33112 20160
rect 33176 20096 33192 20160
rect 33256 20096 33262 20160
rect 32946 20095 33262 20096
rect 42946 20160 43262 20161
rect 42946 20096 42952 20160
rect 43016 20096 43032 20160
rect 43096 20096 43112 20160
rect 43176 20096 43192 20160
rect 43256 20096 43262 20160
rect 50200 20136 51000 20166
rect 42946 20095 43262 20096
rect 28533 20090 28599 20093
rect 32213 20090 32279 20093
rect 28533 20088 32279 20090
rect 28533 20032 28538 20088
rect 28594 20032 32218 20088
rect 32274 20032 32279 20088
rect 28533 20030 32279 20032
rect 28533 20027 28599 20030
rect 32213 20027 32279 20030
rect 39113 20090 39179 20093
rect 41873 20090 41939 20093
rect 39113 20088 41939 20090
rect 39113 20032 39118 20088
rect 39174 20032 41878 20088
rect 41934 20032 41939 20088
rect 39113 20030 41939 20032
rect 39113 20027 39179 20030
rect 41873 20027 41939 20030
rect 0 19954 800 19984
rect 3325 19954 3391 19957
rect 0 19952 3391 19954
rect 0 19896 3330 19952
rect 3386 19896 3391 19952
rect 0 19894 3391 19896
rect 0 19864 800 19894
rect 3325 19891 3391 19894
rect 14641 19954 14707 19957
rect 19333 19954 19399 19957
rect 28257 19954 28323 19957
rect 14641 19952 19399 19954
rect 14641 19896 14646 19952
rect 14702 19896 19338 19952
rect 19394 19896 19399 19952
rect 14641 19894 19399 19896
rect 14641 19891 14707 19894
rect 19333 19891 19399 19894
rect 26558 19952 28323 19954
rect 26558 19896 28262 19952
rect 28318 19896 28323 19952
rect 26558 19894 28323 19896
rect 16665 19818 16731 19821
rect 26558 19818 26618 19894
rect 28257 19891 28323 19894
rect 30833 19954 30899 19957
rect 48497 19954 48563 19957
rect 30833 19952 48563 19954
rect 30833 19896 30838 19952
rect 30894 19896 48502 19952
rect 48558 19896 48563 19952
rect 30833 19894 48563 19896
rect 30833 19891 30899 19894
rect 48497 19891 48563 19894
rect 26785 19818 26851 19821
rect 40401 19818 40467 19821
rect 16665 19816 26618 19818
rect 16665 19760 16670 19816
rect 16726 19760 26618 19816
rect 16665 19758 26618 19760
rect 26742 19816 40467 19818
rect 26742 19760 26790 19816
rect 26846 19760 40406 19816
rect 40462 19760 40467 19816
rect 26742 19758 40467 19760
rect 16665 19755 16731 19758
rect 26742 19755 26851 19758
rect 40401 19755 40467 19758
rect 49049 19818 49115 19821
rect 50200 19818 51000 19848
rect 49049 19816 51000 19818
rect 49049 19760 49054 19816
rect 49110 19760 51000 19816
rect 49049 19758 51000 19760
rect 49049 19755 49115 19758
rect 18413 19682 18479 19685
rect 18873 19682 18939 19685
rect 26742 19682 26802 19755
rect 50200 19728 51000 19758
rect 28533 19684 28599 19685
rect 28533 19682 28580 19684
rect 18413 19680 26802 19682
rect 18413 19624 18418 19680
rect 18474 19624 18878 19680
rect 18934 19624 26802 19680
rect 18413 19622 26802 19624
rect 28488 19680 28580 19682
rect 28488 19624 28538 19680
rect 28488 19622 28580 19624
rect 18413 19619 18479 19622
rect 18873 19619 18939 19622
rect 28533 19620 28580 19622
rect 28644 19620 28650 19684
rect 30005 19682 30071 19685
rect 37365 19682 37431 19685
rect 30005 19680 37431 19682
rect 30005 19624 30010 19680
rect 30066 19624 37370 19680
rect 37426 19624 37431 19680
rect 30005 19622 37431 19624
rect 28533 19619 28599 19620
rect 30005 19619 30071 19622
rect 37365 19619 37431 19622
rect 38377 19682 38443 19685
rect 46105 19682 46171 19685
rect 38377 19680 46171 19682
rect 38377 19624 38382 19680
rect 38438 19624 46110 19680
rect 46166 19624 46171 19680
rect 38377 19622 46171 19624
rect 38377 19619 38443 19622
rect 46105 19619 46171 19622
rect 7946 19616 8262 19617
rect 0 19546 800 19576
rect 7946 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8262 19616
rect 7946 19551 8262 19552
rect 17946 19616 18262 19617
rect 17946 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18262 19616
rect 17946 19551 18262 19552
rect 27946 19616 28262 19617
rect 27946 19552 27952 19616
rect 28016 19552 28032 19616
rect 28096 19552 28112 19616
rect 28176 19552 28192 19616
rect 28256 19552 28262 19616
rect 27946 19551 28262 19552
rect 37946 19616 38262 19617
rect 37946 19552 37952 19616
rect 38016 19552 38032 19616
rect 38096 19552 38112 19616
rect 38176 19552 38192 19616
rect 38256 19552 38262 19616
rect 37946 19551 38262 19552
rect 47946 19616 48262 19617
rect 47946 19552 47952 19616
rect 48016 19552 48032 19616
rect 48096 19552 48112 19616
rect 48176 19552 48192 19616
rect 48256 19552 48262 19616
rect 47946 19551 48262 19552
rect 2681 19546 2747 19549
rect 0 19544 2747 19546
rect 0 19488 2686 19544
rect 2742 19488 2747 19544
rect 0 19486 2747 19488
rect 0 19456 800 19486
rect 2681 19483 2747 19486
rect 35709 19546 35775 19549
rect 37733 19546 37799 19549
rect 35709 19544 37799 19546
rect 35709 19488 35714 19544
rect 35770 19488 37738 19544
rect 37794 19488 37799 19544
rect 35709 19486 37799 19488
rect 35709 19483 35775 19486
rect 37733 19483 37799 19486
rect 17401 19410 17467 19413
rect 25957 19410 26023 19413
rect 17401 19408 26023 19410
rect 17401 19352 17406 19408
rect 17462 19352 25962 19408
rect 26018 19352 26023 19408
rect 17401 19350 26023 19352
rect 17401 19347 17467 19350
rect 25957 19347 26023 19350
rect 26141 19410 26207 19413
rect 33961 19410 34027 19413
rect 48681 19410 48747 19413
rect 26141 19408 48747 19410
rect 26141 19352 26146 19408
rect 26202 19352 33966 19408
rect 34022 19352 48686 19408
rect 48742 19352 48747 19408
rect 26141 19350 48747 19352
rect 26141 19347 26207 19350
rect 33961 19347 34027 19350
rect 48681 19347 48747 19350
rect 49325 19410 49391 19413
rect 50200 19410 51000 19440
rect 49325 19408 51000 19410
rect 49325 19352 49330 19408
rect 49386 19352 51000 19408
rect 49325 19350 51000 19352
rect 49325 19347 49391 19350
rect 50200 19320 51000 19350
rect 2957 19274 3023 19277
rect 1304 19272 3023 19274
rect 1304 19216 2962 19272
rect 3018 19216 3023 19272
rect 1304 19214 3023 19216
rect 0 19138 800 19168
rect 1304 19138 1364 19214
rect 2957 19211 3023 19214
rect 12709 19274 12775 19277
rect 13721 19274 13787 19277
rect 12709 19272 13787 19274
rect 12709 19216 12714 19272
rect 12770 19216 13726 19272
rect 13782 19216 13787 19272
rect 12709 19214 13787 19216
rect 12709 19211 12775 19214
rect 13721 19211 13787 19214
rect 21449 19274 21515 19277
rect 24669 19274 24735 19277
rect 21449 19272 24735 19274
rect 21449 19216 21454 19272
rect 21510 19216 24674 19272
rect 24730 19216 24735 19272
rect 21449 19214 24735 19216
rect 21449 19211 21515 19214
rect 24669 19211 24735 19214
rect 28942 19212 28948 19276
rect 29012 19274 29018 19276
rect 30189 19274 30255 19277
rect 38377 19274 38443 19277
rect 29012 19272 30255 19274
rect 29012 19216 30194 19272
rect 30250 19216 30255 19272
rect 29012 19214 30255 19216
rect 29012 19212 29018 19214
rect 30189 19211 30255 19214
rect 31710 19272 38443 19274
rect 31710 19216 38382 19272
rect 38438 19216 38443 19272
rect 31710 19214 38443 19216
rect 0 19078 1364 19138
rect 25037 19138 25103 19141
rect 30741 19138 30807 19141
rect 25037 19136 30807 19138
rect 25037 19080 25042 19136
rect 25098 19080 30746 19136
rect 30802 19080 30807 19136
rect 25037 19078 30807 19080
rect 0 19048 800 19078
rect 25037 19075 25103 19078
rect 30741 19075 30807 19078
rect 2946 19072 3262 19073
rect 2946 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3262 19072
rect 2946 19007 3262 19008
rect 12946 19072 13262 19073
rect 12946 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13262 19072
rect 12946 19007 13262 19008
rect 22946 19072 23262 19073
rect 22946 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23262 19072
rect 22946 19007 23262 19008
rect 20529 19002 20595 19005
rect 22277 19002 22343 19005
rect 20529 19000 22343 19002
rect 20529 18944 20534 19000
rect 20590 18944 22282 19000
rect 22338 18944 22343 19000
rect 20529 18942 22343 18944
rect 20529 18939 20595 18942
rect 22277 18939 22343 18942
rect 28349 19002 28415 19005
rect 31710 19002 31770 19214
rect 38377 19211 38443 19214
rect 32946 19072 33262 19073
rect 32946 19008 32952 19072
rect 33016 19008 33032 19072
rect 33096 19008 33112 19072
rect 33176 19008 33192 19072
rect 33256 19008 33262 19072
rect 32946 19007 33262 19008
rect 42946 19072 43262 19073
rect 42946 19008 42952 19072
rect 43016 19008 43032 19072
rect 43096 19008 43112 19072
rect 43176 19008 43192 19072
rect 43256 19008 43262 19072
rect 42946 19007 43262 19008
rect 28349 19000 31770 19002
rect 28349 18944 28354 19000
rect 28410 18944 31770 19000
rect 28349 18942 31770 18944
rect 49141 19002 49207 19005
rect 50200 19002 51000 19032
rect 49141 19000 51000 19002
rect 49141 18944 49146 19000
rect 49202 18944 51000 19000
rect 49141 18942 51000 18944
rect 28349 18939 28415 18942
rect 49141 18939 49207 18942
rect 50200 18912 51000 18942
rect 2773 18866 2839 18869
rect 1304 18864 2839 18866
rect 1304 18808 2778 18864
rect 2834 18808 2839 18864
rect 1304 18806 2839 18808
rect 0 18730 800 18760
rect 1304 18730 1364 18806
rect 2773 18803 2839 18806
rect 15653 18866 15719 18869
rect 22737 18866 22803 18869
rect 15653 18864 22803 18866
rect 15653 18808 15658 18864
rect 15714 18808 22742 18864
rect 22798 18808 22803 18864
rect 15653 18806 22803 18808
rect 15653 18803 15719 18806
rect 22737 18803 22803 18806
rect 33041 18866 33107 18869
rect 47301 18866 47367 18869
rect 33041 18864 47367 18866
rect 33041 18808 33046 18864
rect 33102 18808 47306 18864
rect 47362 18808 47367 18864
rect 33041 18806 47367 18808
rect 33041 18803 33107 18806
rect 47301 18803 47367 18806
rect 0 18670 1364 18730
rect 1761 18730 1827 18733
rect 16205 18730 16271 18733
rect 1761 18728 16271 18730
rect 1761 18672 1766 18728
rect 1822 18672 16210 18728
rect 16266 18672 16271 18728
rect 1761 18670 16271 18672
rect 0 18640 800 18670
rect 1761 18667 1827 18670
rect 16205 18667 16271 18670
rect 18413 18730 18479 18733
rect 37457 18730 37523 18733
rect 18413 18728 37523 18730
rect 18413 18672 18418 18728
rect 18474 18672 37462 18728
rect 37518 18672 37523 18728
rect 18413 18670 37523 18672
rect 18413 18667 18479 18670
rect 37457 18667 37523 18670
rect 19333 18594 19399 18597
rect 19701 18594 19767 18597
rect 25037 18594 25103 18597
rect 19333 18592 25103 18594
rect 19333 18536 19338 18592
rect 19394 18536 19706 18592
rect 19762 18536 25042 18592
rect 25098 18536 25103 18592
rect 19333 18534 25103 18536
rect 19333 18531 19399 18534
rect 19701 18531 19767 18534
rect 25037 18531 25103 18534
rect 30649 18594 30715 18597
rect 33041 18594 33107 18597
rect 30649 18592 33107 18594
rect 30649 18536 30654 18592
rect 30710 18536 33046 18592
rect 33102 18536 33107 18592
rect 30649 18534 33107 18536
rect 30649 18531 30715 18534
rect 33041 18531 33107 18534
rect 48589 18594 48655 18597
rect 50200 18594 51000 18624
rect 48589 18592 51000 18594
rect 48589 18536 48594 18592
rect 48650 18536 51000 18592
rect 48589 18534 51000 18536
rect 48589 18531 48655 18534
rect 7946 18528 8262 18529
rect 7946 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8262 18528
rect 7946 18463 8262 18464
rect 17946 18528 18262 18529
rect 17946 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18262 18528
rect 17946 18463 18262 18464
rect 27946 18528 28262 18529
rect 27946 18464 27952 18528
rect 28016 18464 28032 18528
rect 28096 18464 28112 18528
rect 28176 18464 28192 18528
rect 28256 18464 28262 18528
rect 27946 18463 28262 18464
rect 37946 18528 38262 18529
rect 37946 18464 37952 18528
rect 38016 18464 38032 18528
rect 38096 18464 38112 18528
rect 38176 18464 38192 18528
rect 38256 18464 38262 18528
rect 37946 18463 38262 18464
rect 47946 18528 48262 18529
rect 47946 18464 47952 18528
rect 48016 18464 48032 18528
rect 48096 18464 48112 18528
rect 48176 18464 48192 18528
rect 48256 18464 48262 18528
rect 50200 18504 51000 18534
rect 47946 18463 48262 18464
rect 19241 18458 19307 18461
rect 21265 18458 21331 18461
rect 22369 18458 22435 18461
rect 19241 18456 22435 18458
rect 19241 18400 19246 18456
rect 19302 18400 21270 18456
rect 21326 18400 22374 18456
rect 22430 18400 22435 18456
rect 19241 18398 22435 18400
rect 19241 18395 19307 18398
rect 21265 18395 21331 18398
rect 22369 18395 22435 18398
rect 34421 18458 34487 18461
rect 35249 18458 35315 18461
rect 36537 18458 36603 18461
rect 34421 18456 36603 18458
rect 34421 18400 34426 18456
rect 34482 18400 35254 18456
rect 35310 18400 36542 18456
rect 36598 18400 36603 18456
rect 34421 18398 36603 18400
rect 34421 18395 34487 18398
rect 35249 18395 35315 18398
rect 36537 18395 36603 18398
rect 0 18322 800 18352
rect 2865 18322 2931 18325
rect 0 18320 2931 18322
rect 0 18264 2870 18320
rect 2926 18264 2931 18320
rect 0 18262 2931 18264
rect 0 18232 800 18262
rect 2865 18259 2931 18262
rect 16481 18322 16547 18325
rect 30005 18322 30071 18325
rect 16481 18320 30071 18322
rect 16481 18264 16486 18320
rect 16542 18264 30010 18320
rect 30066 18264 30071 18320
rect 16481 18262 30071 18264
rect 16481 18259 16547 18262
rect 30005 18259 30071 18262
rect 30189 18322 30255 18325
rect 41229 18322 41295 18325
rect 30189 18320 41295 18322
rect 30189 18264 30194 18320
rect 30250 18264 41234 18320
rect 41290 18264 41295 18320
rect 30189 18262 41295 18264
rect 30189 18259 30255 18262
rect 41229 18259 41295 18262
rect 14825 18186 14891 18189
rect 24945 18186 25011 18189
rect 14825 18184 25011 18186
rect 14825 18128 14830 18184
rect 14886 18128 24950 18184
rect 25006 18128 25011 18184
rect 14825 18126 25011 18128
rect 14825 18123 14891 18126
rect 24945 18123 25011 18126
rect 49141 18186 49207 18189
rect 50200 18186 51000 18216
rect 49141 18184 51000 18186
rect 49141 18128 49146 18184
rect 49202 18128 51000 18184
rect 49141 18126 51000 18128
rect 49141 18123 49207 18126
rect 50200 18096 51000 18126
rect 14181 18050 14247 18053
rect 18781 18050 18847 18053
rect 14181 18048 18847 18050
rect 14181 17992 14186 18048
rect 14242 17992 18786 18048
rect 18842 17992 18847 18048
rect 14181 17990 18847 17992
rect 14181 17987 14247 17990
rect 18781 17987 18847 17990
rect 24669 18050 24735 18053
rect 26049 18050 26115 18053
rect 24669 18048 26115 18050
rect 24669 17992 24674 18048
rect 24730 17992 26054 18048
rect 26110 17992 26115 18048
rect 24669 17990 26115 17992
rect 24669 17987 24735 17990
rect 26049 17987 26115 17990
rect 2946 17984 3262 17985
rect 0 17914 800 17944
rect 2946 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3262 17984
rect 2946 17919 3262 17920
rect 12946 17984 13262 17985
rect 12946 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13262 17984
rect 12946 17919 13262 17920
rect 22946 17984 23262 17985
rect 22946 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23262 17984
rect 22946 17919 23262 17920
rect 32946 17984 33262 17985
rect 32946 17920 32952 17984
rect 33016 17920 33032 17984
rect 33096 17920 33112 17984
rect 33176 17920 33192 17984
rect 33256 17920 33262 17984
rect 32946 17919 33262 17920
rect 42946 17984 43262 17985
rect 42946 17920 42952 17984
rect 43016 17920 43032 17984
rect 43096 17920 43112 17984
rect 43176 17920 43192 17984
rect 43256 17920 43262 17984
rect 42946 17919 43262 17920
rect 2681 17914 2747 17917
rect 0 17912 2747 17914
rect 0 17856 2686 17912
rect 2742 17856 2747 17912
rect 0 17854 2747 17856
rect 0 17824 800 17854
rect 2681 17851 2747 17854
rect 12065 17778 12131 17781
rect 19241 17778 19307 17781
rect 22185 17778 22251 17781
rect 24301 17778 24367 17781
rect 12065 17776 24367 17778
rect 12065 17720 12070 17776
rect 12126 17720 19246 17776
rect 19302 17720 22190 17776
rect 22246 17720 24306 17776
rect 24362 17720 24367 17776
rect 12065 17718 24367 17720
rect 12065 17715 12131 17718
rect 19241 17715 19307 17718
rect 22185 17715 22251 17718
rect 24301 17715 24367 17718
rect 29729 17778 29795 17781
rect 35065 17778 35131 17781
rect 29729 17776 35131 17778
rect 29729 17720 29734 17776
rect 29790 17720 35070 17776
rect 35126 17720 35131 17776
rect 29729 17718 35131 17720
rect 29729 17715 29795 17718
rect 35065 17715 35131 17718
rect 49049 17778 49115 17781
rect 50200 17778 51000 17808
rect 49049 17776 51000 17778
rect 49049 17720 49054 17776
rect 49110 17720 51000 17776
rect 49049 17718 51000 17720
rect 49049 17715 49115 17718
rect 50200 17688 51000 17718
rect 25681 17642 25747 17645
rect 40585 17642 40651 17645
rect 25681 17640 40651 17642
rect 25681 17584 25686 17640
rect 25742 17584 40590 17640
rect 40646 17584 40651 17640
rect 25681 17582 40651 17584
rect 25681 17579 25747 17582
rect 40585 17579 40651 17582
rect 0 17506 800 17536
rect 2773 17506 2839 17509
rect 0 17504 2839 17506
rect 0 17448 2778 17504
rect 2834 17448 2839 17504
rect 0 17446 2839 17448
rect 0 17416 800 17446
rect 2773 17443 2839 17446
rect 20621 17506 20687 17509
rect 26325 17506 26391 17509
rect 20621 17504 26391 17506
rect 20621 17448 20626 17504
rect 20682 17448 26330 17504
rect 26386 17448 26391 17504
rect 20621 17446 26391 17448
rect 20621 17443 20687 17446
rect 26325 17443 26391 17446
rect 26601 17506 26667 17509
rect 27797 17506 27863 17509
rect 26601 17504 27863 17506
rect 26601 17448 26606 17504
rect 26662 17448 27802 17504
rect 27858 17448 27863 17504
rect 26601 17446 27863 17448
rect 26601 17443 26667 17446
rect 27797 17443 27863 17446
rect 7946 17440 8262 17441
rect 7946 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8262 17440
rect 7946 17375 8262 17376
rect 17946 17440 18262 17441
rect 17946 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18262 17440
rect 17946 17375 18262 17376
rect 27946 17440 28262 17441
rect 27946 17376 27952 17440
rect 28016 17376 28032 17440
rect 28096 17376 28112 17440
rect 28176 17376 28192 17440
rect 28256 17376 28262 17440
rect 27946 17375 28262 17376
rect 37946 17440 38262 17441
rect 37946 17376 37952 17440
rect 38016 17376 38032 17440
rect 38096 17376 38112 17440
rect 38176 17376 38192 17440
rect 38256 17376 38262 17440
rect 37946 17375 38262 17376
rect 47946 17440 48262 17441
rect 47946 17376 47952 17440
rect 48016 17376 48032 17440
rect 48096 17376 48112 17440
rect 48176 17376 48192 17440
rect 48256 17376 48262 17440
rect 47946 17375 48262 17376
rect 19977 17370 20043 17373
rect 20989 17370 21055 17373
rect 19977 17368 21055 17370
rect 19977 17312 19982 17368
rect 20038 17312 20994 17368
rect 21050 17312 21055 17368
rect 19977 17310 21055 17312
rect 19977 17307 20043 17310
rect 20989 17307 21055 17310
rect 49049 17370 49115 17373
rect 50200 17370 51000 17400
rect 49049 17368 51000 17370
rect 49049 17312 49054 17368
rect 49110 17312 51000 17368
rect 49049 17310 51000 17312
rect 49049 17307 49115 17310
rect 50200 17280 51000 17310
rect 14181 17234 14247 17237
rect 25589 17234 25655 17237
rect 14181 17232 25655 17234
rect 14181 17176 14186 17232
rect 14242 17176 25594 17232
rect 25650 17176 25655 17232
rect 14181 17174 25655 17176
rect 14181 17171 14247 17174
rect 25589 17171 25655 17174
rect 27705 17234 27771 17237
rect 41413 17234 41479 17237
rect 27705 17232 41479 17234
rect 27705 17176 27710 17232
rect 27766 17176 41418 17232
rect 41474 17176 41479 17232
rect 27705 17174 41479 17176
rect 27705 17171 27771 17174
rect 41413 17171 41479 17174
rect 0 17098 800 17128
rect 1209 17098 1275 17101
rect 0 17096 1275 17098
rect 0 17040 1214 17096
rect 1270 17040 1275 17096
rect 0 17038 1275 17040
rect 0 17008 800 17038
rect 1209 17035 1275 17038
rect 16573 17098 16639 17101
rect 27797 17098 27863 17101
rect 16573 17096 27863 17098
rect 16573 17040 16578 17096
rect 16634 17040 27802 17096
rect 27858 17040 27863 17096
rect 16573 17038 27863 17040
rect 16573 17035 16639 17038
rect 27797 17035 27863 17038
rect 48589 16962 48655 16965
rect 50200 16962 51000 16992
rect 48589 16960 51000 16962
rect 48589 16904 48594 16960
rect 48650 16904 51000 16960
rect 48589 16902 51000 16904
rect 48589 16899 48655 16902
rect 2946 16896 3262 16897
rect 2946 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3262 16896
rect 2946 16831 3262 16832
rect 12946 16896 13262 16897
rect 12946 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13262 16896
rect 12946 16831 13262 16832
rect 22946 16896 23262 16897
rect 22946 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23262 16896
rect 22946 16831 23262 16832
rect 32946 16896 33262 16897
rect 32946 16832 32952 16896
rect 33016 16832 33032 16896
rect 33096 16832 33112 16896
rect 33176 16832 33192 16896
rect 33256 16832 33262 16896
rect 32946 16831 33262 16832
rect 42946 16896 43262 16897
rect 42946 16832 42952 16896
rect 43016 16832 43032 16896
rect 43096 16832 43112 16896
rect 43176 16832 43192 16896
rect 43256 16832 43262 16896
rect 50200 16872 51000 16902
rect 42946 16831 43262 16832
rect 0 16690 800 16720
rect 1301 16690 1367 16693
rect 0 16688 1367 16690
rect 0 16632 1306 16688
rect 1362 16632 1367 16688
rect 0 16630 1367 16632
rect 0 16600 800 16630
rect 1301 16627 1367 16630
rect 16021 16554 16087 16557
rect 26049 16554 26115 16557
rect 16021 16552 26115 16554
rect 16021 16496 16026 16552
rect 16082 16496 26054 16552
rect 26110 16496 26115 16552
rect 16021 16494 26115 16496
rect 16021 16491 16087 16494
rect 26049 16491 26115 16494
rect 48221 16554 48287 16557
rect 50200 16554 51000 16584
rect 48221 16552 51000 16554
rect 48221 16496 48226 16552
rect 48282 16496 51000 16552
rect 48221 16494 51000 16496
rect 48221 16491 48287 16494
rect 50200 16464 51000 16494
rect 14917 16418 14983 16421
rect 16481 16418 16547 16421
rect 14917 16416 16547 16418
rect 14917 16360 14922 16416
rect 14978 16360 16486 16416
rect 16542 16360 16547 16416
rect 14917 16358 16547 16360
rect 14917 16355 14983 16358
rect 16481 16355 16547 16358
rect 7946 16352 8262 16353
rect 0 16282 800 16312
rect 7946 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8262 16352
rect 7946 16287 8262 16288
rect 17946 16352 18262 16353
rect 17946 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18262 16352
rect 17946 16287 18262 16288
rect 27946 16352 28262 16353
rect 27946 16288 27952 16352
rect 28016 16288 28032 16352
rect 28096 16288 28112 16352
rect 28176 16288 28192 16352
rect 28256 16288 28262 16352
rect 27946 16287 28262 16288
rect 37946 16352 38262 16353
rect 37946 16288 37952 16352
rect 38016 16288 38032 16352
rect 38096 16288 38112 16352
rect 38176 16288 38192 16352
rect 38256 16288 38262 16352
rect 37946 16287 38262 16288
rect 47946 16352 48262 16353
rect 47946 16288 47952 16352
rect 48016 16288 48032 16352
rect 48096 16288 48112 16352
rect 48176 16288 48192 16352
rect 48256 16288 48262 16352
rect 47946 16287 48262 16288
rect 1301 16282 1367 16285
rect 0 16280 1367 16282
rect 0 16224 1306 16280
rect 1362 16224 1367 16280
rect 0 16222 1367 16224
rect 0 16192 800 16222
rect 1301 16219 1367 16222
rect 21173 16282 21239 16285
rect 26325 16282 26391 16285
rect 21173 16280 26391 16282
rect 21173 16224 21178 16280
rect 21234 16224 26330 16280
rect 26386 16224 26391 16280
rect 21173 16222 26391 16224
rect 21173 16219 21239 16222
rect 26325 16219 26391 16222
rect 11881 16146 11947 16149
rect 14365 16146 14431 16149
rect 11881 16144 14431 16146
rect 11881 16088 11886 16144
rect 11942 16088 14370 16144
rect 14426 16088 14431 16144
rect 11881 16086 14431 16088
rect 11881 16083 11947 16086
rect 14365 16083 14431 16086
rect 24485 16146 24551 16149
rect 27705 16146 27771 16149
rect 24485 16144 27771 16146
rect 24485 16088 24490 16144
rect 24546 16088 27710 16144
rect 27766 16088 27771 16144
rect 24485 16086 27771 16088
rect 24485 16083 24551 16086
rect 27705 16083 27771 16086
rect 49141 16146 49207 16149
rect 50200 16146 51000 16176
rect 49141 16144 51000 16146
rect 49141 16088 49146 16144
rect 49202 16088 51000 16144
rect 49141 16086 51000 16088
rect 49141 16083 49207 16086
rect 50200 16056 51000 16086
rect 11329 16010 11395 16013
rect 24853 16010 24919 16013
rect 26141 16010 26207 16013
rect 11329 16008 26207 16010
rect 11329 15952 11334 16008
rect 11390 15952 24858 16008
rect 24914 15952 26146 16008
rect 26202 15952 26207 16008
rect 11329 15950 26207 15952
rect 11329 15947 11395 15950
rect 24853 15947 24919 15950
rect 26141 15947 26207 15950
rect 0 15874 800 15904
rect 1301 15874 1367 15877
rect 0 15872 1367 15874
rect 0 15816 1306 15872
rect 1362 15816 1367 15872
rect 0 15814 1367 15816
rect 0 15784 800 15814
rect 1301 15811 1367 15814
rect 2946 15808 3262 15809
rect 2946 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3262 15808
rect 2946 15743 3262 15744
rect 12946 15808 13262 15809
rect 12946 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13262 15808
rect 12946 15743 13262 15744
rect 22946 15808 23262 15809
rect 22946 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23262 15808
rect 22946 15743 23262 15744
rect 32946 15808 33262 15809
rect 32946 15744 32952 15808
rect 33016 15744 33032 15808
rect 33096 15744 33112 15808
rect 33176 15744 33192 15808
rect 33256 15744 33262 15808
rect 32946 15743 33262 15744
rect 42946 15808 43262 15809
rect 42946 15744 42952 15808
rect 43016 15744 43032 15808
rect 43096 15744 43112 15808
rect 43176 15744 43192 15808
rect 43256 15744 43262 15808
rect 42946 15743 43262 15744
rect 49049 15738 49115 15741
rect 50200 15738 51000 15768
rect 49049 15736 51000 15738
rect 49049 15680 49054 15736
rect 49110 15680 51000 15736
rect 49049 15678 51000 15680
rect 49049 15675 49115 15678
rect 50200 15648 51000 15678
rect 20897 15602 20963 15605
rect 22277 15602 22343 15605
rect 24853 15602 24919 15605
rect 20897 15600 24919 15602
rect 20897 15544 20902 15600
rect 20958 15544 22282 15600
rect 22338 15544 24858 15600
rect 24914 15544 24919 15600
rect 20897 15542 24919 15544
rect 20897 15539 20963 15542
rect 22277 15539 22343 15542
rect 24853 15539 24919 15542
rect 26233 15602 26299 15605
rect 45553 15602 45619 15605
rect 26233 15600 45619 15602
rect 26233 15544 26238 15600
rect 26294 15544 45558 15600
rect 45614 15544 45619 15600
rect 26233 15542 45619 15544
rect 26233 15539 26299 15542
rect 45553 15539 45619 15542
rect 0 15466 800 15496
rect 1301 15466 1367 15469
rect 0 15464 1367 15466
rect 0 15408 1306 15464
rect 1362 15408 1367 15464
rect 0 15406 1367 15408
rect 0 15376 800 15406
rect 1301 15403 1367 15406
rect 16297 15466 16363 15469
rect 18873 15466 18939 15469
rect 16297 15464 18939 15466
rect 16297 15408 16302 15464
rect 16358 15408 18878 15464
rect 18934 15408 18939 15464
rect 16297 15406 18939 15408
rect 16297 15403 16363 15406
rect 18873 15403 18939 15406
rect 25405 15466 25471 15469
rect 49233 15466 49299 15469
rect 25405 15464 49299 15466
rect 25405 15408 25410 15464
rect 25466 15408 49238 15464
rect 49294 15408 49299 15464
rect 25405 15406 49299 15408
rect 25405 15403 25471 15406
rect 49233 15403 49299 15406
rect 49325 15330 49391 15333
rect 50200 15330 51000 15360
rect 49325 15328 51000 15330
rect 49325 15272 49330 15328
rect 49386 15272 51000 15328
rect 49325 15270 51000 15272
rect 49325 15267 49391 15270
rect 7946 15264 8262 15265
rect 7946 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8262 15264
rect 7946 15199 8262 15200
rect 17946 15264 18262 15265
rect 17946 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18262 15264
rect 17946 15199 18262 15200
rect 27946 15264 28262 15265
rect 27946 15200 27952 15264
rect 28016 15200 28032 15264
rect 28096 15200 28112 15264
rect 28176 15200 28192 15264
rect 28256 15200 28262 15264
rect 27946 15199 28262 15200
rect 37946 15264 38262 15265
rect 37946 15200 37952 15264
rect 38016 15200 38032 15264
rect 38096 15200 38112 15264
rect 38176 15200 38192 15264
rect 38256 15200 38262 15264
rect 37946 15199 38262 15200
rect 47946 15264 48262 15265
rect 47946 15200 47952 15264
rect 48016 15200 48032 15264
rect 48096 15200 48112 15264
rect 48176 15200 48192 15264
rect 48256 15200 48262 15264
rect 50200 15240 51000 15270
rect 47946 15199 48262 15200
rect 14733 15194 14799 15197
rect 15101 15194 15167 15197
rect 17401 15194 17467 15197
rect 14733 15192 17467 15194
rect 14733 15136 14738 15192
rect 14794 15136 15106 15192
rect 15162 15136 17406 15192
rect 17462 15136 17467 15192
rect 14733 15134 17467 15136
rect 14733 15131 14799 15134
rect 15101 15131 15167 15134
rect 17401 15131 17467 15134
rect 21725 15194 21791 15197
rect 21725 15192 26986 15194
rect 21725 15136 21730 15192
rect 21786 15136 26986 15192
rect 21725 15134 26986 15136
rect 21725 15131 21791 15134
rect 0 15058 800 15088
rect 1301 15058 1367 15061
rect 0 15056 1367 15058
rect 0 15000 1306 15056
rect 1362 15000 1367 15056
rect 0 14998 1367 15000
rect 0 14968 800 14998
rect 1301 14995 1367 14998
rect 13169 15058 13235 15061
rect 26141 15058 26207 15061
rect 13169 15056 26207 15058
rect 13169 15000 13174 15056
rect 13230 15000 26146 15056
rect 26202 15000 26207 15056
rect 13169 14998 26207 15000
rect 13169 14995 13235 14998
rect 26141 14995 26207 14998
rect 13997 14922 14063 14925
rect 16849 14922 16915 14925
rect 26141 14922 26207 14925
rect 13997 14920 26207 14922
rect 13997 14864 14002 14920
rect 14058 14864 16854 14920
rect 16910 14864 26146 14920
rect 26202 14864 26207 14920
rect 13997 14862 26207 14864
rect 26926 14922 26986 15134
rect 27521 15058 27587 15061
rect 48497 15058 48563 15061
rect 27521 15056 48563 15058
rect 27521 15000 27526 15056
rect 27582 15000 48502 15056
rect 48558 15000 48563 15056
rect 27521 14998 48563 15000
rect 27521 14995 27587 14998
rect 48497 14995 48563 14998
rect 48313 14922 48379 14925
rect 26926 14920 48379 14922
rect 26926 14864 48318 14920
rect 48374 14864 48379 14920
rect 26926 14862 48379 14864
rect 13997 14859 14063 14862
rect 16849 14859 16915 14862
rect 26141 14859 26207 14862
rect 48313 14859 48379 14862
rect 49049 14922 49115 14925
rect 50200 14922 51000 14952
rect 49049 14920 51000 14922
rect 49049 14864 49054 14920
rect 49110 14864 51000 14920
rect 49049 14862 51000 14864
rect 49049 14859 49115 14862
rect 50200 14832 51000 14862
rect 29453 14786 29519 14789
rect 32213 14786 32279 14789
rect 29453 14784 32279 14786
rect 29453 14728 29458 14784
rect 29514 14728 32218 14784
rect 32274 14728 32279 14784
rect 29453 14726 32279 14728
rect 29453 14723 29519 14726
rect 32213 14723 32279 14726
rect 2946 14720 3262 14721
rect 0 14650 800 14680
rect 2946 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3262 14720
rect 2946 14655 3262 14656
rect 12946 14720 13262 14721
rect 12946 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13262 14720
rect 12946 14655 13262 14656
rect 22946 14720 23262 14721
rect 22946 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23262 14720
rect 22946 14655 23262 14656
rect 32946 14720 33262 14721
rect 32946 14656 32952 14720
rect 33016 14656 33032 14720
rect 33096 14656 33112 14720
rect 33176 14656 33192 14720
rect 33256 14656 33262 14720
rect 32946 14655 33262 14656
rect 42946 14720 43262 14721
rect 42946 14656 42952 14720
rect 43016 14656 43032 14720
rect 43096 14656 43112 14720
rect 43176 14656 43192 14720
rect 43256 14656 43262 14720
rect 42946 14655 43262 14656
rect 1301 14650 1367 14653
rect 0 14648 1367 14650
rect 0 14592 1306 14648
rect 1362 14592 1367 14648
rect 0 14590 1367 14592
rect 0 14560 800 14590
rect 1301 14587 1367 14590
rect 16205 14514 16271 14517
rect 17217 14514 17283 14517
rect 17953 14514 18019 14517
rect 16205 14512 18019 14514
rect 16205 14456 16210 14512
rect 16266 14456 17222 14512
rect 17278 14456 17958 14512
rect 18014 14456 18019 14512
rect 16205 14454 18019 14456
rect 16205 14451 16271 14454
rect 17217 14451 17283 14454
rect 17953 14451 18019 14454
rect 18597 14514 18663 14517
rect 32070 14514 32076 14516
rect 18597 14512 32076 14514
rect 18597 14456 18602 14512
rect 18658 14456 32076 14512
rect 18597 14454 32076 14456
rect 18597 14451 18663 14454
rect 32070 14452 32076 14454
rect 32140 14514 32146 14516
rect 32489 14514 32555 14517
rect 32140 14512 32555 14514
rect 32140 14456 32494 14512
rect 32550 14456 32555 14512
rect 32140 14454 32555 14456
rect 32140 14452 32146 14454
rect 32489 14451 32555 14454
rect 49049 14514 49115 14517
rect 50200 14514 51000 14544
rect 49049 14512 51000 14514
rect 49049 14456 49054 14512
rect 49110 14456 51000 14512
rect 49049 14454 51000 14456
rect 49049 14451 49115 14454
rect 50200 14424 51000 14454
rect 11145 14378 11211 14381
rect 22369 14378 22435 14381
rect 22553 14378 22619 14381
rect 49233 14378 49299 14381
rect 11145 14376 49299 14378
rect 11145 14320 11150 14376
rect 11206 14320 22374 14376
rect 22430 14320 22558 14376
rect 22614 14320 49238 14376
rect 49294 14320 49299 14376
rect 11145 14318 49299 14320
rect 11145 14315 11211 14318
rect 22369 14315 22435 14318
rect 22553 14315 22619 14318
rect 49233 14315 49299 14318
rect 0 14242 800 14272
rect 1301 14242 1367 14245
rect 0 14240 1367 14242
rect 0 14184 1306 14240
rect 1362 14184 1367 14240
rect 0 14182 1367 14184
rect 0 14152 800 14182
rect 1301 14179 1367 14182
rect 10133 14242 10199 14245
rect 16757 14242 16823 14245
rect 10133 14240 16823 14242
rect 10133 14184 10138 14240
rect 10194 14184 16762 14240
rect 16818 14184 16823 14240
rect 10133 14182 16823 14184
rect 10133 14179 10199 14182
rect 16757 14179 16823 14182
rect 29545 14242 29611 14245
rect 34881 14242 34947 14245
rect 29545 14240 34947 14242
rect 29545 14184 29550 14240
rect 29606 14184 34886 14240
rect 34942 14184 34947 14240
rect 29545 14182 34947 14184
rect 29545 14179 29611 14182
rect 34881 14179 34947 14182
rect 7946 14176 8262 14177
rect 7946 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8262 14176
rect 7946 14111 8262 14112
rect 17946 14176 18262 14177
rect 17946 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18262 14176
rect 17946 14111 18262 14112
rect 27946 14176 28262 14177
rect 27946 14112 27952 14176
rect 28016 14112 28032 14176
rect 28096 14112 28112 14176
rect 28176 14112 28192 14176
rect 28256 14112 28262 14176
rect 27946 14111 28262 14112
rect 37946 14176 38262 14177
rect 37946 14112 37952 14176
rect 38016 14112 38032 14176
rect 38096 14112 38112 14176
rect 38176 14112 38192 14176
rect 38256 14112 38262 14176
rect 37946 14111 38262 14112
rect 47946 14176 48262 14177
rect 47946 14112 47952 14176
rect 48016 14112 48032 14176
rect 48096 14112 48112 14176
rect 48176 14112 48192 14176
rect 48256 14112 48262 14176
rect 47946 14111 48262 14112
rect 20069 14106 20135 14109
rect 23657 14106 23723 14109
rect 20069 14104 23723 14106
rect 20069 14048 20074 14104
rect 20130 14048 23662 14104
rect 23718 14048 23723 14104
rect 20069 14046 23723 14048
rect 20069 14043 20135 14046
rect 23657 14043 23723 14046
rect 49141 14106 49207 14109
rect 50200 14106 51000 14136
rect 49141 14104 51000 14106
rect 49141 14048 49146 14104
rect 49202 14048 51000 14104
rect 49141 14046 51000 14048
rect 49141 14043 49207 14046
rect 50200 14016 51000 14046
rect 24669 13970 24735 13973
rect 25773 13970 25839 13973
rect 24669 13968 25839 13970
rect 24669 13912 24674 13968
rect 24730 13912 25778 13968
rect 25834 13912 25839 13968
rect 24669 13910 25839 13912
rect 24669 13907 24735 13910
rect 25773 13907 25839 13910
rect 32581 13970 32647 13973
rect 38469 13970 38535 13973
rect 32581 13968 38535 13970
rect 32581 13912 32586 13968
rect 32642 13912 38474 13968
rect 38530 13912 38535 13968
rect 32581 13910 38535 13912
rect 32581 13907 32647 13910
rect 38469 13907 38535 13910
rect 0 13834 800 13864
rect 2773 13834 2839 13837
rect 0 13832 2839 13834
rect 0 13776 2778 13832
rect 2834 13776 2839 13832
rect 0 13774 2839 13776
rect 0 13744 800 13774
rect 2773 13771 2839 13774
rect 15653 13836 15719 13837
rect 15653 13832 15700 13836
rect 15764 13834 15770 13836
rect 15653 13776 15658 13832
rect 15653 13772 15700 13776
rect 15764 13774 15810 13834
rect 15764 13772 15770 13774
rect 15653 13771 15719 13772
rect 15101 13698 15167 13701
rect 21173 13698 21239 13701
rect 15101 13696 21239 13698
rect 15101 13640 15106 13696
rect 15162 13640 21178 13696
rect 21234 13640 21239 13696
rect 15101 13638 21239 13640
rect 15101 13635 15167 13638
rect 21173 13635 21239 13638
rect 48221 13698 48287 13701
rect 50200 13698 51000 13728
rect 48221 13696 51000 13698
rect 48221 13640 48226 13696
rect 48282 13640 51000 13696
rect 48221 13638 51000 13640
rect 48221 13635 48287 13638
rect 2946 13632 3262 13633
rect 2946 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3262 13632
rect 2946 13567 3262 13568
rect 12946 13632 13262 13633
rect 12946 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13262 13632
rect 12946 13567 13262 13568
rect 22946 13632 23262 13633
rect 22946 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23262 13632
rect 22946 13567 23262 13568
rect 32946 13632 33262 13633
rect 32946 13568 32952 13632
rect 33016 13568 33032 13632
rect 33096 13568 33112 13632
rect 33176 13568 33192 13632
rect 33256 13568 33262 13632
rect 32946 13567 33262 13568
rect 42946 13632 43262 13633
rect 42946 13568 42952 13632
rect 43016 13568 43032 13632
rect 43096 13568 43112 13632
rect 43176 13568 43192 13632
rect 43256 13568 43262 13632
rect 50200 13608 51000 13638
rect 42946 13567 43262 13568
rect 0 13426 800 13456
rect 3509 13426 3575 13429
rect 0 13424 3575 13426
rect 0 13368 3514 13424
rect 3570 13368 3575 13424
rect 0 13366 3575 13368
rect 0 13336 800 13366
rect 3509 13363 3575 13366
rect 28809 13426 28875 13429
rect 33869 13426 33935 13429
rect 28809 13424 33935 13426
rect 28809 13368 28814 13424
rect 28870 13368 33874 13424
rect 33930 13368 33935 13424
rect 28809 13366 33935 13368
rect 28809 13363 28875 13366
rect 33869 13363 33935 13366
rect 10317 13290 10383 13293
rect 17953 13290 18019 13293
rect 10317 13288 18019 13290
rect 10317 13232 10322 13288
rect 10378 13232 17958 13288
rect 18014 13232 18019 13288
rect 10317 13230 18019 13232
rect 10317 13227 10383 13230
rect 17953 13227 18019 13230
rect 18781 13290 18847 13293
rect 34697 13290 34763 13293
rect 18781 13288 34763 13290
rect 18781 13232 18786 13288
rect 18842 13232 34702 13288
rect 34758 13232 34763 13288
rect 18781 13230 34763 13232
rect 18781 13227 18847 13230
rect 34697 13227 34763 13230
rect 49141 13290 49207 13293
rect 50200 13290 51000 13320
rect 49141 13288 51000 13290
rect 49141 13232 49146 13288
rect 49202 13232 51000 13288
rect 49141 13230 51000 13232
rect 49141 13227 49207 13230
rect 50200 13200 51000 13230
rect 7946 13088 8262 13089
rect 0 13018 800 13048
rect 7946 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8262 13088
rect 7946 13023 8262 13024
rect 17946 13088 18262 13089
rect 17946 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18262 13088
rect 17946 13023 18262 13024
rect 27946 13088 28262 13089
rect 27946 13024 27952 13088
rect 28016 13024 28032 13088
rect 28096 13024 28112 13088
rect 28176 13024 28192 13088
rect 28256 13024 28262 13088
rect 27946 13023 28262 13024
rect 37946 13088 38262 13089
rect 37946 13024 37952 13088
rect 38016 13024 38032 13088
rect 38096 13024 38112 13088
rect 38176 13024 38192 13088
rect 38256 13024 38262 13088
rect 37946 13023 38262 13024
rect 47946 13088 48262 13089
rect 47946 13024 47952 13088
rect 48016 13024 48032 13088
rect 48096 13024 48112 13088
rect 48176 13024 48192 13088
rect 48256 13024 48262 13088
rect 47946 13023 48262 13024
rect 933 13018 999 13021
rect 0 13016 999 13018
rect 0 12960 938 13016
rect 994 12960 999 13016
rect 0 12958 999 12960
rect 0 12928 800 12958
rect 933 12955 999 12958
rect 16297 13018 16363 13021
rect 16481 13018 16547 13021
rect 16297 13016 16547 13018
rect 16297 12960 16302 13016
rect 16358 12960 16486 13016
rect 16542 12960 16547 13016
rect 16297 12958 16547 12960
rect 16297 12955 16363 12958
rect 16481 12955 16547 12958
rect 15837 12882 15903 12885
rect 16297 12882 16363 12885
rect 25313 12882 25379 12885
rect 26233 12882 26299 12885
rect 15837 12880 26299 12882
rect 15837 12824 15842 12880
rect 15898 12824 16302 12880
rect 16358 12824 25318 12880
rect 25374 12824 26238 12880
rect 26294 12824 26299 12880
rect 15837 12822 26299 12824
rect 15837 12819 15903 12822
rect 16297 12819 16363 12822
rect 25313 12819 25379 12822
rect 26233 12819 26299 12822
rect 49141 12882 49207 12885
rect 50200 12882 51000 12912
rect 49141 12880 51000 12882
rect 49141 12824 49146 12880
rect 49202 12824 51000 12880
rect 49141 12822 51000 12824
rect 49141 12819 49207 12822
rect 50200 12792 51000 12822
rect 22369 12746 22435 12749
rect 46841 12746 46907 12749
rect 22369 12744 46907 12746
rect 22369 12688 22374 12744
rect 22430 12688 46846 12744
rect 46902 12688 46907 12744
rect 22369 12686 46907 12688
rect 22369 12683 22435 12686
rect 46841 12683 46907 12686
rect 0 12610 800 12640
rect 1301 12610 1367 12613
rect 0 12608 1367 12610
rect 0 12552 1306 12608
rect 1362 12552 1367 12608
rect 0 12550 1367 12552
rect 0 12520 800 12550
rect 1301 12547 1367 12550
rect 13537 12610 13603 12613
rect 15561 12610 15627 12613
rect 13537 12608 15627 12610
rect 13537 12552 13542 12608
rect 13598 12552 15566 12608
rect 15622 12552 15627 12608
rect 13537 12550 15627 12552
rect 13537 12547 13603 12550
rect 15561 12547 15627 12550
rect 2946 12544 3262 12545
rect 2946 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3262 12544
rect 2946 12479 3262 12480
rect 12946 12544 13262 12545
rect 12946 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13262 12544
rect 12946 12479 13262 12480
rect 22946 12544 23262 12545
rect 22946 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23262 12544
rect 22946 12479 23262 12480
rect 32946 12544 33262 12545
rect 32946 12480 32952 12544
rect 33016 12480 33032 12544
rect 33096 12480 33112 12544
rect 33176 12480 33192 12544
rect 33256 12480 33262 12544
rect 32946 12479 33262 12480
rect 42946 12544 43262 12545
rect 42946 12480 42952 12544
rect 43016 12480 43032 12544
rect 43096 12480 43112 12544
rect 43176 12480 43192 12544
rect 43256 12480 43262 12544
rect 42946 12479 43262 12480
rect 31937 12474 32003 12477
rect 32305 12474 32371 12477
rect 31937 12472 32371 12474
rect 31937 12416 31942 12472
rect 31998 12416 32310 12472
rect 32366 12416 32371 12472
rect 31937 12414 32371 12416
rect 31937 12411 32003 12414
rect 32305 12411 32371 12414
rect 49141 12474 49207 12477
rect 50200 12474 51000 12504
rect 49141 12472 51000 12474
rect 49141 12416 49146 12472
rect 49202 12416 51000 12472
rect 49141 12414 51000 12416
rect 49141 12411 49207 12414
rect 50200 12384 51000 12414
rect 11329 12338 11395 12341
rect 15469 12338 15535 12341
rect 11329 12336 15535 12338
rect 11329 12280 11334 12336
rect 11390 12280 15474 12336
rect 15530 12280 15535 12336
rect 11329 12278 15535 12280
rect 11329 12275 11395 12278
rect 15469 12275 15535 12278
rect 32489 12338 32555 12341
rect 32949 12338 33015 12341
rect 32489 12336 33015 12338
rect 32489 12280 32494 12336
rect 32550 12280 32954 12336
rect 33010 12280 33015 12336
rect 32489 12278 33015 12280
rect 32489 12275 32555 12278
rect 32949 12275 33015 12278
rect 0 12202 800 12232
rect 1025 12202 1091 12205
rect 0 12200 1091 12202
rect 0 12144 1030 12200
rect 1086 12144 1091 12200
rect 0 12142 1091 12144
rect 0 12112 800 12142
rect 1025 12139 1091 12142
rect 11053 12202 11119 12205
rect 15009 12202 15075 12205
rect 17217 12202 17283 12205
rect 11053 12200 17283 12202
rect 11053 12144 11058 12200
rect 11114 12144 15014 12200
rect 15070 12144 17222 12200
rect 17278 12144 17283 12200
rect 11053 12142 17283 12144
rect 11053 12139 11119 12142
rect 15009 12139 15075 12142
rect 17217 12139 17283 12142
rect 17769 12202 17835 12205
rect 32489 12202 32555 12205
rect 32765 12202 32831 12205
rect 17769 12200 22110 12202
rect 17769 12144 17774 12200
rect 17830 12144 22110 12200
rect 17769 12142 22110 12144
rect 17769 12139 17835 12142
rect 22050 12066 22110 12142
rect 32489 12200 32831 12202
rect 32489 12144 32494 12200
rect 32550 12144 32770 12200
rect 32826 12144 32831 12200
rect 32489 12142 32831 12144
rect 32489 12139 32555 12142
rect 32765 12139 32831 12142
rect 33317 12202 33383 12205
rect 33685 12202 33751 12205
rect 33317 12200 33751 12202
rect 33317 12144 33322 12200
rect 33378 12144 33690 12200
rect 33746 12144 33751 12200
rect 33317 12142 33751 12144
rect 33317 12139 33383 12142
rect 33685 12139 33751 12142
rect 22461 12066 22527 12069
rect 22050 12064 22527 12066
rect 22050 12008 22466 12064
rect 22522 12008 22527 12064
rect 22050 12006 22527 12008
rect 22461 12003 22527 12006
rect 23749 12066 23815 12069
rect 27705 12066 27771 12069
rect 23749 12064 27771 12066
rect 23749 12008 23754 12064
rect 23810 12008 27710 12064
rect 27766 12008 27771 12064
rect 23749 12006 27771 12008
rect 23749 12003 23815 12006
rect 27705 12003 27771 12006
rect 49141 12066 49207 12069
rect 50200 12066 51000 12096
rect 49141 12064 51000 12066
rect 49141 12008 49146 12064
rect 49202 12008 51000 12064
rect 49141 12006 51000 12008
rect 49141 12003 49207 12006
rect 7946 12000 8262 12001
rect 7946 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8262 12000
rect 7946 11935 8262 11936
rect 17946 12000 18262 12001
rect 17946 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18262 12000
rect 17946 11935 18262 11936
rect 27946 12000 28262 12001
rect 27946 11936 27952 12000
rect 28016 11936 28032 12000
rect 28096 11936 28112 12000
rect 28176 11936 28192 12000
rect 28256 11936 28262 12000
rect 27946 11935 28262 11936
rect 37946 12000 38262 12001
rect 37946 11936 37952 12000
rect 38016 11936 38032 12000
rect 38096 11936 38112 12000
rect 38176 11936 38192 12000
rect 38256 11936 38262 12000
rect 37946 11935 38262 11936
rect 47946 12000 48262 12001
rect 47946 11936 47952 12000
rect 48016 11936 48032 12000
rect 48096 11936 48112 12000
rect 48176 11936 48192 12000
rect 48256 11936 48262 12000
rect 50200 11976 51000 12006
rect 47946 11935 48262 11936
rect 32029 11930 32095 11933
rect 32305 11930 32371 11933
rect 32029 11928 32371 11930
rect 32029 11872 32034 11928
rect 32090 11872 32310 11928
rect 32366 11872 32371 11928
rect 32029 11870 32371 11872
rect 32029 11867 32095 11870
rect 32305 11867 32371 11870
rect 0 11794 800 11824
rect 933 11794 999 11797
rect 0 11792 999 11794
rect 0 11736 938 11792
rect 994 11736 999 11792
rect 0 11734 999 11736
rect 0 11704 800 11734
rect 933 11731 999 11734
rect 20989 11794 21055 11797
rect 27429 11794 27495 11797
rect 36169 11794 36235 11797
rect 20989 11792 36235 11794
rect 20989 11736 20994 11792
rect 21050 11736 27434 11792
rect 27490 11736 36174 11792
rect 36230 11736 36235 11792
rect 20989 11734 36235 11736
rect 20989 11731 21055 11734
rect 27429 11731 27495 11734
rect 36169 11731 36235 11734
rect 49141 11658 49207 11661
rect 50200 11658 51000 11688
rect 49141 11656 51000 11658
rect 49141 11600 49146 11656
rect 49202 11600 51000 11656
rect 49141 11598 51000 11600
rect 49141 11595 49207 11598
rect 50200 11568 51000 11598
rect 2946 11456 3262 11457
rect 0 11386 800 11416
rect 2946 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3262 11456
rect 2946 11391 3262 11392
rect 12946 11456 13262 11457
rect 12946 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13262 11456
rect 12946 11391 13262 11392
rect 22946 11456 23262 11457
rect 22946 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23262 11456
rect 22946 11391 23262 11392
rect 32946 11456 33262 11457
rect 32946 11392 32952 11456
rect 33016 11392 33032 11456
rect 33096 11392 33112 11456
rect 33176 11392 33192 11456
rect 33256 11392 33262 11456
rect 32946 11391 33262 11392
rect 42946 11456 43262 11457
rect 42946 11392 42952 11456
rect 43016 11392 43032 11456
rect 43096 11392 43112 11456
rect 43176 11392 43192 11456
rect 43256 11392 43262 11456
rect 42946 11391 43262 11392
rect 933 11386 999 11389
rect 0 11384 999 11386
rect 0 11328 938 11384
rect 994 11328 999 11384
rect 0 11326 999 11328
rect 0 11296 800 11326
rect 933 11323 999 11326
rect 36169 11386 36235 11389
rect 40125 11386 40191 11389
rect 36169 11384 40191 11386
rect 36169 11328 36174 11384
rect 36230 11328 40130 11384
rect 40186 11328 40191 11384
rect 36169 11326 40191 11328
rect 36169 11323 36235 11326
rect 40125 11323 40191 11326
rect 17217 11250 17283 11253
rect 23289 11250 23355 11253
rect 17217 11248 23355 11250
rect 17217 11192 17222 11248
rect 17278 11192 23294 11248
rect 23350 11192 23355 11248
rect 17217 11190 23355 11192
rect 17217 11187 17283 11190
rect 23289 11187 23355 11190
rect 49233 11250 49299 11253
rect 50200 11250 51000 11280
rect 49233 11248 51000 11250
rect 49233 11192 49238 11248
rect 49294 11192 51000 11248
rect 49233 11190 51000 11192
rect 49233 11187 49299 11190
rect 50200 11160 51000 11190
rect 32070 11052 32076 11116
rect 32140 11114 32146 11116
rect 36445 11114 36511 11117
rect 32140 11112 36511 11114
rect 32140 11056 36450 11112
rect 36506 11056 36511 11112
rect 32140 11054 36511 11056
rect 32140 11052 32146 11054
rect 36445 11051 36511 11054
rect 0 10978 800 11008
rect 1577 10978 1643 10981
rect 0 10976 1643 10978
rect 0 10920 1582 10976
rect 1638 10920 1643 10976
rect 0 10918 1643 10920
rect 0 10888 800 10918
rect 1577 10915 1643 10918
rect 31477 10978 31543 10981
rect 33777 10978 33843 10981
rect 31477 10976 33843 10978
rect 31477 10920 31482 10976
rect 31538 10920 33782 10976
rect 33838 10920 33843 10976
rect 31477 10918 33843 10920
rect 31477 10915 31543 10918
rect 33777 10915 33843 10918
rect 34237 10978 34303 10981
rect 36537 10978 36603 10981
rect 34237 10976 36603 10978
rect 34237 10920 34242 10976
rect 34298 10920 36542 10976
rect 36598 10920 36603 10976
rect 34237 10918 36603 10920
rect 34237 10915 34303 10918
rect 36537 10915 36603 10918
rect 7946 10912 8262 10913
rect 7946 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8262 10912
rect 7946 10847 8262 10848
rect 17946 10912 18262 10913
rect 17946 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18262 10912
rect 17946 10847 18262 10848
rect 27946 10912 28262 10913
rect 27946 10848 27952 10912
rect 28016 10848 28032 10912
rect 28096 10848 28112 10912
rect 28176 10848 28192 10912
rect 28256 10848 28262 10912
rect 27946 10847 28262 10848
rect 37946 10912 38262 10913
rect 37946 10848 37952 10912
rect 38016 10848 38032 10912
rect 38096 10848 38112 10912
rect 38176 10848 38192 10912
rect 38256 10848 38262 10912
rect 37946 10847 38262 10848
rect 47946 10912 48262 10913
rect 47946 10848 47952 10912
rect 48016 10848 48032 10912
rect 48096 10848 48112 10912
rect 48176 10848 48192 10912
rect 48256 10848 48262 10912
rect 47946 10847 48262 10848
rect 49141 10842 49207 10845
rect 50200 10842 51000 10872
rect 49141 10840 51000 10842
rect 49141 10784 49146 10840
rect 49202 10784 51000 10840
rect 49141 10782 51000 10784
rect 49141 10779 49207 10782
rect 50200 10752 51000 10782
rect 14457 10706 14523 10709
rect 19333 10706 19399 10709
rect 20621 10706 20687 10709
rect 14457 10704 20687 10706
rect 14457 10648 14462 10704
rect 14518 10648 19338 10704
rect 19394 10648 20626 10704
rect 20682 10648 20687 10704
rect 14457 10646 20687 10648
rect 14457 10643 14523 10646
rect 19333 10643 19399 10646
rect 20621 10643 20687 10646
rect 0 10570 800 10600
rect 933 10570 999 10573
rect 0 10568 999 10570
rect 0 10512 938 10568
rect 994 10512 999 10568
rect 0 10510 999 10512
rect 0 10480 800 10510
rect 933 10507 999 10510
rect 49325 10434 49391 10437
rect 50200 10434 51000 10464
rect 49325 10432 51000 10434
rect 49325 10376 49330 10432
rect 49386 10376 51000 10432
rect 49325 10374 51000 10376
rect 49325 10371 49391 10374
rect 2946 10368 3262 10369
rect 2946 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3262 10368
rect 2946 10303 3262 10304
rect 12946 10368 13262 10369
rect 12946 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13262 10368
rect 12946 10303 13262 10304
rect 22946 10368 23262 10369
rect 22946 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23262 10368
rect 22946 10303 23262 10304
rect 32946 10368 33262 10369
rect 32946 10304 32952 10368
rect 33016 10304 33032 10368
rect 33096 10304 33112 10368
rect 33176 10304 33192 10368
rect 33256 10304 33262 10368
rect 32946 10303 33262 10304
rect 42946 10368 43262 10369
rect 42946 10304 42952 10368
rect 43016 10304 43032 10368
rect 43096 10304 43112 10368
rect 43176 10304 43192 10368
rect 43256 10304 43262 10368
rect 50200 10344 51000 10374
rect 42946 10303 43262 10304
rect 0 10162 800 10192
rect 1209 10162 1275 10165
rect 0 10160 1275 10162
rect 0 10104 1214 10160
rect 1270 10104 1275 10160
rect 0 10102 1275 10104
rect 0 10072 800 10102
rect 1209 10099 1275 10102
rect 33593 10162 33659 10165
rect 34329 10162 34395 10165
rect 39757 10162 39823 10165
rect 33593 10160 39823 10162
rect 33593 10104 33598 10160
rect 33654 10104 34334 10160
rect 34390 10104 39762 10160
rect 39818 10104 39823 10160
rect 33593 10102 39823 10104
rect 33593 10099 33659 10102
rect 34329 10099 34395 10102
rect 39757 10099 39823 10102
rect 13261 10026 13327 10029
rect 33961 10026 34027 10029
rect 13261 10024 34027 10026
rect 13261 9968 13266 10024
rect 13322 9968 33966 10024
rect 34022 9968 34027 10024
rect 13261 9966 34027 9968
rect 13261 9963 13327 9966
rect 33961 9963 34027 9966
rect 49233 10026 49299 10029
rect 50200 10026 51000 10056
rect 49233 10024 51000 10026
rect 49233 9968 49238 10024
rect 49294 9968 51000 10024
rect 49233 9966 51000 9968
rect 49233 9963 49299 9966
rect 50200 9936 51000 9966
rect 7946 9824 8262 9825
rect 0 9754 800 9784
rect 7946 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8262 9824
rect 7946 9759 8262 9760
rect 17946 9824 18262 9825
rect 17946 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18262 9824
rect 17946 9759 18262 9760
rect 27946 9824 28262 9825
rect 27946 9760 27952 9824
rect 28016 9760 28032 9824
rect 28096 9760 28112 9824
rect 28176 9760 28192 9824
rect 28256 9760 28262 9824
rect 27946 9759 28262 9760
rect 37946 9824 38262 9825
rect 37946 9760 37952 9824
rect 38016 9760 38032 9824
rect 38096 9760 38112 9824
rect 38176 9760 38192 9824
rect 38256 9760 38262 9824
rect 37946 9759 38262 9760
rect 47946 9824 48262 9825
rect 47946 9760 47952 9824
rect 48016 9760 48032 9824
rect 48096 9760 48112 9824
rect 48176 9760 48192 9824
rect 48256 9760 48262 9824
rect 47946 9759 48262 9760
rect 933 9754 999 9757
rect 0 9752 999 9754
rect 0 9696 938 9752
rect 994 9696 999 9752
rect 0 9694 999 9696
rect 0 9664 800 9694
rect 933 9691 999 9694
rect 15469 9618 15535 9621
rect 15694 9618 15700 9620
rect 15469 9616 15700 9618
rect 15469 9560 15474 9616
rect 15530 9560 15700 9616
rect 15469 9558 15700 9560
rect 15469 9555 15535 9558
rect 15694 9556 15700 9558
rect 15764 9618 15770 9620
rect 26141 9618 26207 9621
rect 15764 9616 26207 9618
rect 15764 9560 26146 9616
rect 26202 9560 26207 9616
rect 15764 9558 26207 9560
rect 15764 9556 15770 9558
rect 26141 9555 26207 9558
rect 47301 9618 47367 9621
rect 50200 9618 51000 9648
rect 47301 9616 51000 9618
rect 47301 9560 47306 9616
rect 47362 9560 51000 9616
rect 47301 9558 51000 9560
rect 47301 9555 47367 9558
rect 50200 9528 51000 9558
rect 1761 9482 1827 9485
rect 33593 9482 33659 9485
rect 1761 9480 33659 9482
rect 1761 9424 1766 9480
rect 1822 9424 33598 9480
rect 33654 9424 33659 9480
rect 1761 9422 33659 9424
rect 1761 9419 1827 9422
rect 33593 9419 33659 9422
rect 0 9346 800 9376
rect 933 9346 999 9349
rect 0 9344 999 9346
rect 0 9288 938 9344
rect 994 9288 999 9344
rect 0 9286 999 9288
rect 0 9256 800 9286
rect 933 9283 999 9286
rect 2946 9280 3262 9281
rect 2946 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3262 9280
rect 2946 9215 3262 9216
rect 12946 9280 13262 9281
rect 12946 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13262 9280
rect 12946 9215 13262 9216
rect 22946 9280 23262 9281
rect 22946 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23262 9280
rect 22946 9215 23262 9216
rect 32946 9280 33262 9281
rect 32946 9216 32952 9280
rect 33016 9216 33032 9280
rect 33096 9216 33112 9280
rect 33176 9216 33192 9280
rect 33256 9216 33262 9280
rect 32946 9215 33262 9216
rect 42946 9280 43262 9281
rect 42946 9216 42952 9280
rect 43016 9216 43032 9280
rect 43096 9216 43112 9280
rect 43176 9216 43192 9280
rect 43256 9216 43262 9280
rect 42946 9215 43262 9216
rect 49141 9210 49207 9213
rect 50200 9210 51000 9240
rect 49141 9208 51000 9210
rect 49141 9152 49146 9208
rect 49202 9152 51000 9208
rect 49141 9150 51000 9152
rect 49141 9147 49207 9150
rect 50200 9120 51000 9150
rect 14825 9074 14891 9077
rect 18413 9074 18479 9077
rect 14825 9072 18479 9074
rect 14825 9016 14830 9072
rect 14886 9016 18418 9072
rect 18474 9016 18479 9072
rect 14825 9014 18479 9016
rect 14825 9011 14891 9014
rect 18413 9011 18479 9014
rect 0 8938 800 8968
rect 933 8938 999 8941
rect 0 8936 999 8938
rect 0 8880 938 8936
rect 994 8880 999 8936
rect 0 8878 999 8880
rect 0 8848 800 8878
rect 933 8875 999 8878
rect 28625 8938 28691 8941
rect 31845 8938 31911 8941
rect 38745 8938 38811 8941
rect 28625 8936 38811 8938
rect 28625 8880 28630 8936
rect 28686 8880 31850 8936
rect 31906 8880 38750 8936
rect 38806 8880 38811 8936
rect 28625 8878 38811 8880
rect 28625 8875 28691 8878
rect 31845 8875 31911 8878
rect 38745 8875 38811 8878
rect 49233 8802 49299 8805
rect 50200 8802 51000 8832
rect 49233 8800 51000 8802
rect 49233 8744 49238 8800
rect 49294 8744 51000 8800
rect 49233 8742 51000 8744
rect 49233 8739 49299 8742
rect 7946 8736 8262 8737
rect 7946 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8262 8736
rect 7946 8671 8262 8672
rect 17946 8736 18262 8737
rect 17946 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18262 8736
rect 17946 8671 18262 8672
rect 27946 8736 28262 8737
rect 27946 8672 27952 8736
rect 28016 8672 28032 8736
rect 28096 8672 28112 8736
rect 28176 8672 28192 8736
rect 28256 8672 28262 8736
rect 27946 8671 28262 8672
rect 37946 8736 38262 8737
rect 37946 8672 37952 8736
rect 38016 8672 38032 8736
rect 38096 8672 38112 8736
rect 38176 8672 38192 8736
rect 38256 8672 38262 8736
rect 37946 8671 38262 8672
rect 47946 8736 48262 8737
rect 47946 8672 47952 8736
rect 48016 8672 48032 8736
rect 48096 8672 48112 8736
rect 48176 8672 48192 8736
rect 48256 8672 48262 8736
rect 50200 8712 51000 8742
rect 47946 8671 48262 8672
rect 0 8530 800 8560
rect 1209 8530 1275 8533
rect 0 8528 1275 8530
rect 0 8472 1214 8528
rect 1270 8472 1275 8528
rect 0 8470 1275 8472
rect 0 8440 800 8470
rect 1209 8467 1275 8470
rect 49325 8394 49391 8397
rect 50200 8394 51000 8424
rect 49325 8392 51000 8394
rect 49325 8336 49330 8392
rect 49386 8336 51000 8392
rect 49325 8334 51000 8336
rect 49325 8331 49391 8334
rect 50200 8304 51000 8334
rect 2946 8192 3262 8193
rect 0 8122 800 8152
rect 2946 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3262 8192
rect 2946 8127 3262 8128
rect 12946 8192 13262 8193
rect 12946 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13262 8192
rect 12946 8127 13262 8128
rect 22946 8192 23262 8193
rect 22946 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23262 8192
rect 22946 8127 23262 8128
rect 32946 8192 33262 8193
rect 32946 8128 32952 8192
rect 33016 8128 33032 8192
rect 33096 8128 33112 8192
rect 33176 8128 33192 8192
rect 33256 8128 33262 8192
rect 32946 8127 33262 8128
rect 42946 8192 43262 8193
rect 42946 8128 42952 8192
rect 43016 8128 43032 8192
rect 43096 8128 43112 8192
rect 43176 8128 43192 8192
rect 43256 8128 43262 8192
rect 42946 8127 43262 8128
rect 1577 8122 1643 8125
rect 0 8120 1643 8122
rect 0 8064 1582 8120
rect 1638 8064 1643 8120
rect 0 8062 1643 8064
rect 0 8032 800 8062
rect 1577 8059 1643 8062
rect 46841 7986 46907 7989
rect 50200 7986 51000 8016
rect 46841 7984 51000 7986
rect 46841 7928 46846 7984
rect 46902 7928 51000 7984
rect 46841 7926 51000 7928
rect 46841 7923 46907 7926
rect 50200 7896 51000 7926
rect 0 7714 800 7744
rect 933 7714 999 7717
rect 0 7712 999 7714
rect 0 7656 938 7712
rect 994 7656 999 7712
rect 0 7654 999 7656
rect 0 7624 800 7654
rect 933 7651 999 7654
rect 7946 7648 8262 7649
rect 7946 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8262 7648
rect 7946 7583 8262 7584
rect 17946 7648 18262 7649
rect 17946 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18262 7648
rect 17946 7583 18262 7584
rect 27946 7648 28262 7649
rect 27946 7584 27952 7648
rect 28016 7584 28032 7648
rect 28096 7584 28112 7648
rect 28176 7584 28192 7648
rect 28256 7584 28262 7648
rect 27946 7583 28262 7584
rect 37946 7648 38262 7649
rect 37946 7584 37952 7648
rect 38016 7584 38032 7648
rect 38096 7584 38112 7648
rect 38176 7584 38192 7648
rect 38256 7584 38262 7648
rect 37946 7583 38262 7584
rect 47946 7648 48262 7649
rect 47946 7584 47952 7648
rect 48016 7584 48032 7648
rect 48096 7584 48112 7648
rect 48176 7584 48192 7648
rect 48256 7584 48262 7648
rect 47946 7583 48262 7584
rect 49141 7578 49207 7581
rect 50200 7578 51000 7608
rect 49141 7576 51000 7578
rect 49141 7520 49146 7576
rect 49202 7520 51000 7576
rect 49141 7518 51000 7520
rect 49141 7515 49207 7518
rect 50200 7488 51000 7518
rect 0 7306 800 7336
rect 933 7306 999 7309
rect 0 7304 999 7306
rect 0 7248 938 7304
rect 994 7248 999 7304
rect 0 7246 999 7248
rect 0 7216 800 7246
rect 933 7243 999 7246
rect 49233 7170 49299 7173
rect 50200 7170 51000 7200
rect 49233 7168 51000 7170
rect 49233 7112 49238 7168
rect 49294 7112 51000 7168
rect 49233 7110 51000 7112
rect 49233 7107 49299 7110
rect 2946 7104 3262 7105
rect 2946 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3262 7104
rect 2946 7039 3262 7040
rect 12946 7104 13262 7105
rect 12946 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13262 7104
rect 12946 7039 13262 7040
rect 22946 7104 23262 7105
rect 22946 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23262 7104
rect 22946 7039 23262 7040
rect 32946 7104 33262 7105
rect 32946 7040 32952 7104
rect 33016 7040 33032 7104
rect 33096 7040 33112 7104
rect 33176 7040 33192 7104
rect 33256 7040 33262 7104
rect 32946 7039 33262 7040
rect 42946 7104 43262 7105
rect 42946 7040 42952 7104
rect 43016 7040 43032 7104
rect 43096 7040 43112 7104
rect 43176 7040 43192 7104
rect 43256 7040 43262 7104
rect 50200 7080 51000 7110
rect 42946 7039 43262 7040
rect 0 6898 800 6928
rect 933 6898 999 6901
rect 0 6896 999 6898
rect 0 6840 938 6896
rect 994 6840 999 6896
rect 0 6838 999 6840
rect 0 6808 800 6838
rect 933 6835 999 6838
rect 49417 6762 49483 6765
rect 50200 6762 51000 6792
rect 49417 6760 51000 6762
rect 49417 6704 49422 6760
rect 49478 6704 51000 6760
rect 49417 6702 51000 6704
rect 49417 6699 49483 6702
rect 50200 6672 51000 6702
rect 7946 6560 8262 6561
rect 0 6490 800 6520
rect 7946 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8262 6560
rect 7946 6495 8262 6496
rect 17946 6560 18262 6561
rect 17946 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18262 6560
rect 17946 6495 18262 6496
rect 27946 6560 28262 6561
rect 27946 6496 27952 6560
rect 28016 6496 28032 6560
rect 28096 6496 28112 6560
rect 28176 6496 28192 6560
rect 28256 6496 28262 6560
rect 27946 6495 28262 6496
rect 37946 6560 38262 6561
rect 37946 6496 37952 6560
rect 38016 6496 38032 6560
rect 38096 6496 38112 6560
rect 38176 6496 38192 6560
rect 38256 6496 38262 6560
rect 37946 6495 38262 6496
rect 47946 6560 48262 6561
rect 47946 6496 47952 6560
rect 48016 6496 48032 6560
rect 48096 6496 48112 6560
rect 48176 6496 48192 6560
rect 48256 6496 48262 6560
rect 47946 6495 48262 6496
rect 1301 6490 1367 6493
rect 0 6488 1367 6490
rect 0 6432 1306 6488
rect 1362 6432 1367 6488
rect 0 6430 1367 6432
rect 0 6400 800 6430
rect 1301 6427 1367 6430
rect 48865 6354 48931 6357
rect 50200 6354 51000 6384
rect 48865 6352 51000 6354
rect 48865 6296 48870 6352
rect 48926 6296 51000 6352
rect 48865 6294 51000 6296
rect 48865 6291 48931 6294
rect 50200 6264 51000 6294
rect 0 6082 800 6112
rect 933 6082 999 6085
rect 0 6080 999 6082
rect 0 6024 938 6080
rect 994 6024 999 6080
rect 0 6022 999 6024
rect 0 5992 800 6022
rect 933 6019 999 6022
rect 2946 6016 3262 6017
rect 2946 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3262 6016
rect 2946 5951 3262 5952
rect 12946 6016 13262 6017
rect 12946 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13262 6016
rect 12946 5951 13262 5952
rect 22946 6016 23262 6017
rect 22946 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23262 6016
rect 22946 5951 23262 5952
rect 32946 6016 33262 6017
rect 32946 5952 32952 6016
rect 33016 5952 33032 6016
rect 33096 5952 33112 6016
rect 33176 5952 33192 6016
rect 33256 5952 33262 6016
rect 32946 5951 33262 5952
rect 42946 6016 43262 6017
rect 42946 5952 42952 6016
rect 43016 5952 43032 6016
rect 43096 5952 43112 6016
rect 43176 5952 43192 6016
rect 43256 5952 43262 6016
rect 42946 5951 43262 5952
rect 49141 5946 49207 5949
rect 50200 5946 51000 5976
rect 49141 5944 51000 5946
rect 49141 5888 49146 5944
rect 49202 5888 51000 5944
rect 49141 5886 51000 5888
rect 49141 5883 49207 5886
rect 50200 5856 51000 5886
rect 0 5674 800 5704
rect 933 5674 999 5677
rect 0 5672 999 5674
rect 0 5616 938 5672
rect 994 5616 999 5672
rect 0 5614 999 5616
rect 0 5584 800 5614
rect 933 5611 999 5614
rect 49417 5538 49483 5541
rect 50200 5538 51000 5568
rect 49417 5536 51000 5538
rect 49417 5480 49422 5536
rect 49478 5480 51000 5536
rect 49417 5478 51000 5480
rect 49417 5475 49483 5478
rect 7946 5472 8262 5473
rect 7946 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8262 5472
rect 7946 5407 8262 5408
rect 17946 5472 18262 5473
rect 17946 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18262 5472
rect 17946 5407 18262 5408
rect 27946 5472 28262 5473
rect 27946 5408 27952 5472
rect 28016 5408 28032 5472
rect 28096 5408 28112 5472
rect 28176 5408 28192 5472
rect 28256 5408 28262 5472
rect 27946 5407 28262 5408
rect 37946 5472 38262 5473
rect 37946 5408 37952 5472
rect 38016 5408 38032 5472
rect 38096 5408 38112 5472
rect 38176 5408 38192 5472
rect 38256 5408 38262 5472
rect 37946 5407 38262 5408
rect 47946 5472 48262 5473
rect 47946 5408 47952 5472
rect 48016 5408 48032 5472
rect 48096 5408 48112 5472
rect 48176 5408 48192 5472
rect 48256 5408 48262 5472
rect 50200 5448 51000 5478
rect 47946 5407 48262 5408
rect 0 5266 800 5296
rect 2313 5266 2379 5269
rect 0 5264 2379 5266
rect 0 5208 2318 5264
rect 2374 5208 2379 5264
rect 0 5206 2379 5208
rect 0 5176 800 5206
rect 2313 5203 2379 5206
rect 49325 5130 49391 5133
rect 50200 5130 51000 5160
rect 49325 5128 51000 5130
rect 49325 5072 49330 5128
rect 49386 5072 51000 5128
rect 49325 5070 51000 5072
rect 49325 5067 49391 5070
rect 50200 5040 51000 5070
rect 2946 4928 3262 4929
rect 0 4858 800 4888
rect 2946 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3262 4928
rect 2946 4863 3262 4864
rect 12946 4928 13262 4929
rect 12946 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13262 4928
rect 12946 4863 13262 4864
rect 22946 4928 23262 4929
rect 22946 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23262 4928
rect 22946 4863 23262 4864
rect 32946 4928 33262 4929
rect 32946 4864 32952 4928
rect 33016 4864 33032 4928
rect 33096 4864 33112 4928
rect 33176 4864 33192 4928
rect 33256 4864 33262 4928
rect 32946 4863 33262 4864
rect 42946 4928 43262 4929
rect 42946 4864 42952 4928
rect 43016 4864 43032 4928
rect 43096 4864 43112 4928
rect 43176 4864 43192 4928
rect 43256 4864 43262 4928
rect 42946 4863 43262 4864
rect 933 4858 999 4861
rect 0 4856 999 4858
rect 0 4800 938 4856
rect 994 4800 999 4856
rect 0 4798 999 4800
rect 0 4768 800 4798
rect 933 4795 999 4798
rect 48313 4722 48379 4725
rect 50200 4722 51000 4752
rect 48313 4720 51000 4722
rect 48313 4664 48318 4720
rect 48374 4664 51000 4720
rect 48313 4662 51000 4664
rect 48313 4659 48379 4662
rect 50200 4632 51000 4662
rect 0 4450 800 4480
rect 933 4450 999 4453
rect 0 4448 999 4450
rect 0 4392 938 4448
rect 994 4392 999 4448
rect 0 4390 999 4392
rect 0 4360 800 4390
rect 933 4387 999 4390
rect 7946 4384 8262 4385
rect 7946 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8262 4384
rect 7946 4319 8262 4320
rect 17946 4384 18262 4385
rect 17946 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18262 4384
rect 17946 4319 18262 4320
rect 27946 4384 28262 4385
rect 27946 4320 27952 4384
rect 28016 4320 28032 4384
rect 28096 4320 28112 4384
rect 28176 4320 28192 4384
rect 28256 4320 28262 4384
rect 27946 4319 28262 4320
rect 37946 4384 38262 4385
rect 37946 4320 37952 4384
rect 38016 4320 38032 4384
rect 38096 4320 38112 4384
rect 38176 4320 38192 4384
rect 38256 4320 38262 4384
rect 37946 4319 38262 4320
rect 47946 4384 48262 4385
rect 47946 4320 47952 4384
rect 48016 4320 48032 4384
rect 48096 4320 48112 4384
rect 48176 4320 48192 4384
rect 48256 4320 48262 4384
rect 47946 4319 48262 4320
rect 49141 4314 49207 4317
rect 50200 4314 51000 4344
rect 49141 4312 51000 4314
rect 49141 4256 49146 4312
rect 49202 4256 51000 4312
rect 49141 4254 51000 4256
rect 49141 4251 49207 4254
rect 50200 4224 51000 4254
rect 0 4042 800 4072
rect 1669 4042 1735 4045
rect 0 4040 1735 4042
rect 0 3984 1674 4040
rect 1730 3984 1735 4040
rect 0 3982 1735 3984
rect 0 3952 800 3982
rect 1669 3979 1735 3982
rect 49233 3906 49299 3909
rect 50200 3906 51000 3936
rect 49233 3904 51000 3906
rect 49233 3848 49238 3904
rect 49294 3848 51000 3904
rect 49233 3846 51000 3848
rect 49233 3843 49299 3846
rect 2946 3840 3262 3841
rect 2946 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3262 3840
rect 2946 3775 3262 3776
rect 12946 3840 13262 3841
rect 12946 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13262 3840
rect 12946 3775 13262 3776
rect 22946 3840 23262 3841
rect 22946 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23262 3840
rect 22946 3775 23262 3776
rect 32946 3840 33262 3841
rect 32946 3776 32952 3840
rect 33016 3776 33032 3840
rect 33096 3776 33112 3840
rect 33176 3776 33192 3840
rect 33256 3776 33262 3840
rect 32946 3775 33262 3776
rect 42946 3840 43262 3841
rect 42946 3776 42952 3840
rect 43016 3776 43032 3840
rect 43096 3776 43112 3840
rect 43176 3776 43192 3840
rect 43256 3776 43262 3840
rect 50200 3816 51000 3846
rect 42946 3775 43262 3776
rect 0 3634 800 3664
rect 933 3634 999 3637
rect 0 3632 999 3634
rect 0 3576 938 3632
rect 994 3576 999 3632
rect 0 3574 999 3576
rect 0 3544 800 3574
rect 933 3571 999 3574
rect 5349 3634 5415 3637
rect 24393 3634 24459 3637
rect 5349 3632 24459 3634
rect 5349 3576 5354 3632
rect 5410 3576 24398 3632
rect 24454 3576 24459 3632
rect 5349 3574 24459 3576
rect 5349 3571 5415 3574
rect 24393 3571 24459 3574
rect 1117 3498 1183 3501
rect 22185 3498 22251 3501
rect 27613 3498 27679 3501
rect 1117 3496 27679 3498
rect 1117 3440 1122 3496
rect 1178 3440 22190 3496
rect 22246 3440 27618 3496
rect 27674 3440 27679 3496
rect 1117 3438 27679 3440
rect 1117 3435 1183 3438
rect 22185 3435 22251 3438
rect 27613 3435 27679 3438
rect 49141 3498 49207 3501
rect 50200 3498 51000 3528
rect 49141 3496 51000 3498
rect 49141 3440 49146 3496
rect 49202 3440 51000 3496
rect 49141 3438 51000 3440
rect 49141 3435 49207 3438
rect 50200 3408 51000 3438
rect 7946 3296 8262 3297
rect 0 3226 800 3256
rect 7946 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8262 3296
rect 7946 3231 8262 3232
rect 17946 3296 18262 3297
rect 17946 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18262 3296
rect 17946 3231 18262 3232
rect 27946 3296 28262 3297
rect 27946 3232 27952 3296
rect 28016 3232 28032 3296
rect 28096 3232 28112 3296
rect 28176 3232 28192 3296
rect 28256 3232 28262 3296
rect 27946 3231 28262 3232
rect 37946 3296 38262 3297
rect 37946 3232 37952 3296
rect 38016 3232 38032 3296
rect 38096 3232 38112 3296
rect 38176 3232 38192 3296
rect 38256 3232 38262 3296
rect 37946 3231 38262 3232
rect 47946 3296 48262 3297
rect 47946 3232 47952 3296
rect 48016 3232 48032 3296
rect 48096 3232 48112 3296
rect 48176 3232 48192 3296
rect 48256 3232 48262 3296
rect 47946 3231 48262 3232
rect 933 3226 999 3229
rect 0 3224 999 3226
rect 0 3168 938 3224
rect 994 3168 999 3224
rect 0 3166 999 3168
rect 0 3136 800 3166
rect 933 3163 999 3166
rect 48681 3090 48747 3093
rect 50200 3090 51000 3120
rect 48681 3088 51000 3090
rect 48681 3032 48686 3088
rect 48742 3032 51000 3088
rect 48681 3030 51000 3032
rect 48681 3027 48747 3030
rect 50200 3000 51000 3030
rect 0 2818 800 2848
rect 933 2818 999 2821
rect 0 2816 999 2818
rect 0 2760 938 2816
rect 994 2760 999 2816
rect 0 2758 999 2760
rect 0 2728 800 2758
rect 933 2755 999 2758
rect 2946 2752 3262 2753
rect 2946 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3262 2752
rect 2946 2687 3262 2688
rect 12946 2752 13262 2753
rect 12946 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13262 2752
rect 12946 2687 13262 2688
rect 22946 2752 23262 2753
rect 22946 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23262 2752
rect 22946 2687 23262 2688
rect 32946 2752 33262 2753
rect 32946 2688 32952 2752
rect 33016 2688 33032 2752
rect 33096 2688 33112 2752
rect 33176 2688 33192 2752
rect 33256 2688 33262 2752
rect 32946 2687 33262 2688
rect 42946 2752 43262 2753
rect 42946 2688 42952 2752
rect 43016 2688 43032 2752
rect 43096 2688 43112 2752
rect 43176 2688 43192 2752
rect 43256 2688 43262 2752
rect 42946 2687 43262 2688
rect 46841 2682 46907 2685
rect 50200 2682 51000 2712
rect 46841 2680 51000 2682
rect 46841 2624 46846 2680
rect 46902 2624 51000 2680
rect 46841 2622 51000 2624
rect 46841 2619 46907 2622
rect 50200 2592 51000 2622
rect 0 2410 800 2440
rect 933 2410 999 2413
rect 0 2408 999 2410
rect 0 2352 938 2408
rect 994 2352 999 2408
rect 0 2350 999 2352
rect 0 2320 800 2350
rect 933 2347 999 2350
rect 48497 2274 48563 2277
rect 50200 2274 51000 2304
rect 48497 2272 51000 2274
rect 48497 2216 48502 2272
rect 48558 2216 51000 2272
rect 48497 2214 51000 2216
rect 48497 2211 48563 2214
rect 7946 2208 8262 2209
rect 7946 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8262 2208
rect 7946 2143 8262 2144
rect 17946 2208 18262 2209
rect 17946 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18262 2208
rect 17946 2143 18262 2144
rect 27946 2208 28262 2209
rect 27946 2144 27952 2208
rect 28016 2144 28032 2208
rect 28096 2144 28112 2208
rect 28176 2144 28192 2208
rect 28256 2144 28262 2208
rect 27946 2143 28262 2144
rect 37946 2208 38262 2209
rect 37946 2144 37952 2208
rect 38016 2144 38032 2208
rect 38096 2144 38112 2208
rect 38176 2144 38192 2208
rect 38256 2144 38262 2208
rect 37946 2143 38262 2144
rect 47946 2208 48262 2209
rect 47946 2144 47952 2208
rect 48016 2144 48032 2208
rect 48096 2144 48112 2208
rect 48176 2144 48192 2208
rect 48256 2144 48262 2208
rect 50200 2184 51000 2214
rect 47946 2143 48262 2144
rect 0 2002 800 2032
rect 1209 2002 1275 2005
rect 0 2000 1275 2002
rect 0 1944 1214 2000
rect 1270 1944 1275 2000
rect 0 1942 1275 1944
rect 0 1912 800 1942
rect 1209 1939 1275 1942
rect 46749 1866 46815 1869
rect 50200 1866 51000 1896
rect 46749 1864 51000 1866
rect 46749 1808 46754 1864
rect 46810 1808 51000 1864
rect 46749 1806 51000 1808
rect 46749 1803 46815 1806
rect 50200 1776 51000 1806
rect 0 1594 800 1624
rect 1301 1594 1367 1597
rect 0 1592 1367 1594
rect 0 1536 1306 1592
rect 1362 1536 1367 1592
rect 0 1534 1367 1536
rect 0 1504 800 1534
rect 1301 1531 1367 1534
rect 46657 1458 46723 1461
rect 50200 1458 51000 1488
rect 46657 1456 51000 1458
rect 46657 1400 46662 1456
rect 46718 1400 51000 1456
rect 46657 1398 51000 1400
rect 46657 1395 46723 1398
rect 50200 1368 51000 1398
<< via3 >>
rect 35388 24924 35452 24988
rect 2952 24508 3016 24512
rect 2952 24452 2956 24508
rect 2956 24452 3012 24508
rect 3012 24452 3016 24508
rect 2952 24448 3016 24452
rect 3032 24508 3096 24512
rect 3032 24452 3036 24508
rect 3036 24452 3092 24508
rect 3092 24452 3096 24508
rect 3032 24448 3096 24452
rect 3112 24508 3176 24512
rect 3112 24452 3116 24508
rect 3116 24452 3172 24508
rect 3172 24452 3176 24508
rect 3112 24448 3176 24452
rect 3192 24508 3256 24512
rect 3192 24452 3196 24508
rect 3196 24452 3252 24508
rect 3252 24452 3256 24508
rect 3192 24448 3256 24452
rect 12952 24508 13016 24512
rect 12952 24452 12956 24508
rect 12956 24452 13012 24508
rect 13012 24452 13016 24508
rect 12952 24448 13016 24452
rect 13032 24508 13096 24512
rect 13032 24452 13036 24508
rect 13036 24452 13092 24508
rect 13092 24452 13096 24508
rect 13032 24448 13096 24452
rect 13112 24508 13176 24512
rect 13112 24452 13116 24508
rect 13116 24452 13172 24508
rect 13172 24452 13176 24508
rect 13112 24448 13176 24452
rect 13192 24508 13256 24512
rect 13192 24452 13196 24508
rect 13196 24452 13252 24508
rect 13252 24452 13256 24508
rect 13192 24448 13256 24452
rect 22952 24508 23016 24512
rect 22952 24452 22956 24508
rect 22956 24452 23012 24508
rect 23012 24452 23016 24508
rect 22952 24448 23016 24452
rect 23032 24508 23096 24512
rect 23032 24452 23036 24508
rect 23036 24452 23092 24508
rect 23092 24452 23096 24508
rect 23032 24448 23096 24452
rect 23112 24508 23176 24512
rect 23112 24452 23116 24508
rect 23116 24452 23172 24508
rect 23172 24452 23176 24508
rect 23112 24448 23176 24452
rect 23192 24508 23256 24512
rect 23192 24452 23196 24508
rect 23196 24452 23252 24508
rect 23252 24452 23256 24508
rect 23192 24448 23256 24452
rect 32952 24508 33016 24512
rect 32952 24452 32956 24508
rect 32956 24452 33012 24508
rect 33012 24452 33016 24508
rect 32952 24448 33016 24452
rect 33032 24508 33096 24512
rect 33032 24452 33036 24508
rect 33036 24452 33092 24508
rect 33092 24452 33096 24508
rect 33032 24448 33096 24452
rect 33112 24508 33176 24512
rect 33112 24452 33116 24508
rect 33116 24452 33172 24508
rect 33172 24452 33176 24508
rect 33112 24448 33176 24452
rect 33192 24508 33256 24512
rect 33192 24452 33196 24508
rect 33196 24452 33252 24508
rect 33252 24452 33256 24508
rect 33192 24448 33256 24452
rect 42952 24508 43016 24512
rect 42952 24452 42956 24508
rect 42956 24452 43012 24508
rect 43012 24452 43016 24508
rect 42952 24448 43016 24452
rect 43032 24508 43096 24512
rect 43032 24452 43036 24508
rect 43036 24452 43092 24508
rect 43092 24452 43096 24508
rect 43032 24448 43096 24452
rect 43112 24508 43176 24512
rect 43112 24452 43116 24508
rect 43116 24452 43172 24508
rect 43172 24452 43176 24508
rect 43112 24448 43176 24452
rect 43192 24508 43256 24512
rect 43192 24452 43196 24508
rect 43196 24452 43252 24508
rect 43252 24452 43256 24508
rect 43192 24448 43256 24452
rect 7952 23964 8016 23968
rect 7952 23908 7956 23964
rect 7956 23908 8012 23964
rect 8012 23908 8016 23964
rect 7952 23904 8016 23908
rect 8032 23964 8096 23968
rect 8032 23908 8036 23964
rect 8036 23908 8092 23964
rect 8092 23908 8096 23964
rect 8032 23904 8096 23908
rect 8112 23964 8176 23968
rect 8112 23908 8116 23964
rect 8116 23908 8172 23964
rect 8172 23908 8176 23964
rect 8112 23904 8176 23908
rect 8192 23964 8256 23968
rect 8192 23908 8196 23964
rect 8196 23908 8252 23964
rect 8252 23908 8256 23964
rect 8192 23904 8256 23908
rect 17952 23964 18016 23968
rect 17952 23908 17956 23964
rect 17956 23908 18012 23964
rect 18012 23908 18016 23964
rect 17952 23904 18016 23908
rect 18032 23964 18096 23968
rect 18032 23908 18036 23964
rect 18036 23908 18092 23964
rect 18092 23908 18096 23964
rect 18032 23904 18096 23908
rect 18112 23964 18176 23968
rect 18112 23908 18116 23964
rect 18116 23908 18172 23964
rect 18172 23908 18176 23964
rect 18112 23904 18176 23908
rect 18192 23964 18256 23968
rect 18192 23908 18196 23964
rect 18196 23908 18252 23964
rect 18252 23908 18256 23964
rect 18192 23904 18256 23908
rect 27952 23964 28016 23968
rect 27952 23908 27956 23964
rect 27956 23908 28012 23964
rect 28012 23908 28016 23964
rect 27952 23904 28016 23908
rect 28032 23964 28096 23968
rect 28032 23908 28036 23964
rect 28036 23908 28092 23964
rect 28092 23908 28096 23964
rect 28032 23904 28096 23908
rect 28112 23964 28176 23968
rect 28112 23908 28116 23964
rect 28116 23908 28172 23964
rect 28172 23908 28176 23964
rect 28112 23904 28176 23908
rect 28192 23964 28256 23968
rect 28192 23908 28196 23964
rect 28196 23908 28252 23964
rect 28252 23908 28256 23964
rect 28192 23904 28256 23908
rect 37952 23964 38016 23968
rect 37952 23908 37956 23964
rect 37956 23908 38012 23964
rect 38012 23908 38016 23964
rect 37952 23904 38016 23908
rect 38032 23964 38096 23968
rect 38032 23908 38036 23964
rect 38036 23908 38092 23964
rect 38092 23908 38096 23964
rect 38032 23904 38096 23908
rect 38112 23964 38176 23968
rect 38112 23908 38116 23964
rect 38116 23908 38172 23964
rect 38172 23908 38176 23964
rect 38112 23904 38176 23908
rect 38192 23964 38256 23968
rect 38192 23908 38196 23964
rect 38196 23908 38252 23964
rect 38252 23908 38256 23964
rect 38192 23904 38256 23908
rect 47952 23964 48016 23968
rect 47952 23908 47956 23964
rect 47956 23908 48012 23964
rect 48012 23908 48016 23964
rect 47952 23904 48016 23908
rect 48032 23964 48096 23968
rect 48032 23908 48036 23964
rect 48036 23908 48092 23964
rect 48092 23908 48096 23964
rect 48032 23904 48096 23908
rect 48112 23964 48176 23968
rect 48112 23908 48116 23964
rect 48116 23908 48172 23964
rect 48172 23908 48176 23964
rect 48112 23904 48176 23908
rect 48192 23964 48256 23968
rect 48192 23908 48196 23964
rect 48196 23908 48252 23964
rect 48252 23908 48256 23964
rect 48192 23904 48256 23908
rect 28948 23700 29012 23764
rect 2952 23420 3016 23424
rect 2952 23364 2956 23420
rect 2956 23364 3012 23420
rect 3012 23364 3016 23420
rect 2952 23360 3016 23364
rect 3032 23420 3096 23424
rect 3032 23364 3036 23420
rect 3036 23364 3092 23420
rect 3092 23364 3096 23420
rect 3032 23360 3096 23364
rect 3112 23420 3176 23424
rect 3112 23364 3116 23420
rect 3116 23364 3172 23420
rect 3172 23364 3176 23420
rect 3112 23360 3176 23364
rect 3192 23420 3256 23424
rect 3192 23364 3196 23420
rect 3196 23364 3252 23420
rect 3252 23364 3256 23420
rect 3192 23360 3256 23364
rect 12952 23420 13016 23424
rect 12952 23364 12956 23420
rect 12956 23364 13012 23420
rect 13012 23364 13016 23420
rect 12952 23360 13016 23364
rect 13032 23420 13096 23424
rect 13032 23364 13036 23420
rect 13036 23364 13092 23420
rect 13092 23364 13096 23420
rect 13032 23360 13096 23364
rect 13112 23420 13176 23424
rect 13112 23364 13116 23420
rect 13116 23364 13172 23420
rect 13172 23364 13176 23420
rect 13112 23360 13176 23364
rect 13192 23420 13256 23424
rect 13192 23364 13196 23420
rect 13196 23364 13252 23420
rect 13252 23364 13256 23420
rect 13192 23360 13256 23364
rect 22952 23420 23016 23424
rect 22952 23364 22956 23420
rect 22956 23364 23012 23420
rect 23012 23364 23016 23420
rect 22952 23360 23016 23364
rect 23032 23420 23096 23424
rect 23032 23364 23036 23420
rect 23036 23364 23092 23420
rect 23092 23364 23096 23420
rect 23032 23360 23096 23364
rect 23112 23420 23176 23424
rect 23112 23364 23116 23420
rect 23116 23364 23172 23420
rect 23172 23364 23176 23420
rect 23112 23360 23176 23364
rect 23192 23420 23256 23424
rect 23192 23364 23196 23420
rect 23196 23364 23252 23420
rect 23252 23364 23256 23420
rect 23192 23360 23256 23364
rect 32952 23420 33016 23424
rect 32952 23364 32956 23420
rect 32956 23364 33012 23420
rect 33012 23364 33016 23420
rect 32952 23360 33016 23364
rect 33032 23420 33096 23424
rect 33032 23364 33036 23420
rect 33036 23364 33092 23420
rect 33092 23364 33096 23420
rect 33032 23360 33096 23364
rect 33112 23420 33176 23424
rect 33112 23364 33116 23420
rect 33116 23364 33172 23420
rect 33172 23364 33176 23420
rect 33112 23360 33176 23364
rect 33192 23420 33256 23424
rect 33192 23364 33196 23420
rect 33196 23364 33252 23420
rect 33252 23364 33256 23420
rect 33192 23360 33256 23364
rect 42952 23420 43016 23424
rect 42952 23364 42956 23420
rect 42956 23364 43012 23420
rect 43012 23364 43016 23420
rect 42952 23360 43016 23364
rect 43032 23420 43096 23424
rect 43032 23364 43036 23420
rect 43036 23364 43092 23420
rect 43092 23364 43096 23420
rect 43032 23360 43096 23364
rect 43112 23420 43176 23424
rect 43112 23364 43116 23420
rect 43116 23364 43172 23420
rect 43172 23364 43176 23420
rect 43112 23360 43176 23364
rect 43192 23420 43256 23424
rect 43192 23364 43196 23420
rect 43196 23364 43252 23420
rect 43252 23364 43256 23420
rect 43192 23360 43256 23364
rect 7952 22876 8016 22880
rect 7952 22820 7956 22876
rect 7956 22820 8012 22876
rect 8012 22820 8016 22876
rect 7952 22816 8016 22820
rect 8032 22876 8096 22880
rect 8032 22820 8036 22876
rect 8036 22820 8092 22876
rect 8092 22820 8096 22876
rect 8032 22816 8096 22820
rect 8112 22876 8176 22880
rect 8112 22820 8116 22876
rect 8116 22820 8172 22876
rect 8172 22820 8176 22876
rect 8112 22816 8176 22820
rect 8192 22876 8256 22880
rect 8192 22820 8196 22876
rect 8196 22820 8252 22876
rect 8252 22820 8256 22876
rect 8192 22816 8256 22820
rect 17952 22876 18016 22880
rect 17952 22820 17956 22876
rect 17956 22820 18012 22876
rect 18012 22820 18016 22876
rect 17952 22816 18016 22820
rect 18032 22876 18096 22880
rect 18032 22820 18036 22876
rect 18036 22820 18092 22876
rect 18092 22820 18096 22876
rect 18032 22816 18096 22820
rect 18112 22876 18176 22880
rect 18112 22820 18116 22876
rect 18116 22820 18172 22876
rect 18172 22820 18176 22876
rect 18112 22816 18176 22820
rect 18192 22876 18256 22880
rect 18192 22820 18196 22876
rect 18196 22820 18252 22876
rect 18252 22820 18256 22876
rect 18192 22816 18256 22820
rect 27952 22876 28016 22880
rect 27952 22820 27956 22876
rect 27956 22820 28012 22876
rect 28012 22820 28016 22876
rect 27952 22816 28016 22820
rect 28032 22876 28096 22880
rect 28032 22820 28036 22876
rect 28036 22820 28092 22876
rect 28092 22820 28096 22876
rect 28032 22816 28096 22820
rect 28112 22876 28176 22880
rect 28112 22820 28116 22876
rect 28116 22820 28172 22876
rect 28172 22820 28176 22876
rect 28112 22816 28176 22820
rect 28192 22876 28256 22880
rect 28192 22820 28196 22876
rect 28196 22820 28252 22876
rect 28252 22820 28256 22876
rect 28192 22816 28256 22820
rect 37952 22876 38016 22880
rect 37952 22820 37956 22876
rect 37956 22820 38012 22876
rect 38012 22820 38016 22876
rect 37952 22816 38016 22820
rect 38032 22876 38096 22880
rect 38032 22820 38036 22876
rect 38036 22820 38092 22876
rect 38092 22820 38096 22876
rect 38032 22816 38096 22820
rect 38112 22876 38176 22880
rect 38112 22820 38116 22876
rect 38116 22820 38172 22876
rect 38172 22820 38176 22876
rect 38112 22816 38176 22820
rect 38192 22876 38256 22880
rect 38192 22820 38196 22876
rect 38196 22820 38252 22876
rect 38252 22820 38256 22876
rect 38192 22816 38256 22820
rect 47952 22876 48016 22880
rect 47952 22820 47956 22876
rect 47956 22820 48012 22876
rect 48012 22820 48016 22876
rect 47952 22816 48016 22820
rect 48032 22876 48096 22880
rect 48032 22820 48036 22876
rect 48036 22820 48092 22876
rect 48092 22820 48096 22876
rect 48032 22816 48096 22820
rect 48112 22876 48176 22880
rect 48112 22820 48116 22876
rect 48116 22820 48172 22876
rect 48172 22820 48176 22876
rect 48112 22816 48176 22820
rect 48192 22876 48256 22880
rect 48192 22820 48196 22876
rect 48196 22820 48252 22876
rect 48252 22820 48256 22876
rect 48192 22816 48256 22820
rect 2952 22332 3016 22336
rect 2952 22276 2956 22332
rect 2956 22276 3012 22332
rect 3012 22276 3016 22332
rect 2952 22272 3016 22276
rect 3032 22332 3096 22336
rect 3032 22276 3036 22332
rect 3036 22276 3092 22332
rect 3092 22276 3096 22332
rect 3032 22272 3096 22276
rect 3112 22332 3176 22336
rect 3112 22276 3116 22332
rect 3116 22276 3172 22332
rect 3172 22276 3176 22332
rect 3112 22272 3176 22276
rect 3192 22332 3256 22336
rect 3192 22276 3196 22332
rect 3196 22276 3252 22332
rect 3252 22276 3256 22332
rect 3192 22272 3256 22276
rect 12952 22332 13016 22336
rect 12952 22276 12956 22332
rect 12956 22276 13012 22332
rect 13012 22276 13016 22332
rect 12952 22272 13016 22276
rect 13032 22332 13096 22336
rect 13032 22276 13036 22332
rect 13036 22276 13092 22332
rect 13092 22276 13096 22332
rect 13032 22272 13096 22276
rect 13112 22332 13176 22336
rect 13112 22276 13116 22332
rect 13116 22276 13172 22332
rect 13172 22276 13176 22332
rect 13112 22272 13176 22276
rect 13192 22332 13256 22336
rect 13192 22276 13196 22332
rect 13196 22276 13252 22332
rect 13252 22276 13256 22332
rect 13192 22272 13256 22276
rect 22952 22332 23016 22336
rect 22952 22276 22956 22332
rect 22956 22276 23012 22332
rect 23012 22276 23016 22332
rect 22952 22272 23016 22276
rect 23032 22332 23096 22336
rect 23032 22276 23036 22332
rect 23036 22276 23092 22332
rect 23092 22276 23096 22332
rect 23032 22272 23096 22276
rect 23112 22332 23176 22336
rect 23112 22276 23116 22332
rect 23116 22276 23172 22332
rect 23172 22276 23176 22332
rect 23112 22272 23176 22276
rect 23192 22332 23256 22336
rect 23192 22276 23196 22332
rect 23196 22276 23252 22332
rect 23252 22276 23256 22332
rect 23192 22272 23256 22276
rect 32952 22332 33016 22336
rect 32952 22276 32956 22332
rect 32956 22276 33012 22332
rect 33012 22276 33016 22332
rect 32952 22272 33016 22276
rect 33032 22332 33096 22336
rect 33032 22276 33036 22332
rect 33036 22276 33092 22332
rect 33092 22276 33096 22332
rect 33032 22272 33096 22276
rect 33112 22332 33176 22336
rect 33112 22276 33116 22332
rect 33116 22276 33172 22332
rect 33172 22276 33176 22332
rect 33112 22272 33176 22276
rect 33192 22332 33256 22336
rect 33192 22276 33196 22332
rect 33196 22276 33252 22332
rect 33252 22276 33256 22332
rect 33192 22272 33256 22276
rect 42952 22332 43016 22336
rect 42952 22276 42956 22332
rect 42956 22276 43012 22332
rect 43012 22276 43016 22332
rect 42952 22272 43016 22276
rect 43032 22332 43096 22336
rect 43032 22276 43036 22332
rect 43036 22276 43092 22332
rect 43092 22276 43096 22332
rect 43032 22272 43096 22276
rect 43112 22332 43176 22336
rect 43112 22276 43116 22332
rect 43116 22276 43172 22332
rect 43172 22276 43176 22332
rect 43112 22272 43176 22276
rect 43192 22332 43256 22336
rect 43192 22276 43196 22332
rect 43196 22276 43252 22332
rect 43252 22276 43256 22332
rect 43192 22272 43256 22276
rect 7952 21788 8016 21792
rect 7952 21732 7956 21788
rect 7956 21732 8012 21788
rect 8012 21732 8016 21788
rect 7952 21728 8016 21732
rect 8032 21788 8096 21792
rect 8032 21732 8036 21788
rect 8036 21732 8092 21788
rect 8092 21732 8096 21788
rect 8032 21728 8096 21732
rect 8112 21788 8176 21792
rect 8112 21732 8116 21788
rect 8116 21732 8172 21788
rect 8172 21732 8176 21788
rect 8112 21728 8176 21732
rect 8192 21788 8256 21792
rect 8192 21732 8196 21788
rect 8196 21732 8252 21788
rect 8252 21732 8256 21788
rect 8192 21728 8256 21732
rect 17952 21788 18016 21792
rect 17952 21732 17956 21788
rect 17956 21732 18012 21788
rect 18012 21732 18016 21788
rect 17952 21728 18016 21732
rect 18032 21788 18096 21792
rect 18032 21732 18036 21788
rect 18036 21732 18092 21788
rect 18092 21732 18096 21788
rect 18032 21728 18096 21732
rect 18112 21788 18176 21792
rect 18112 21732 18116 21788
rect 18116 21732 18172 21788
rect 18172 21732 18176 21788
rect 18112 21728 18176 21732
rect 18192 21788 18256 21792
rect 18192 21732 18196 21788
rect 18196 21732 18252 21788
rect 18252 21732 18256 21788
rect 18192 21728 18256 21732
rect 27952 21788 28016 21792
rect 27952 21732 27956 21788
rect 27956 21732 28012 21788
rect 28012 21732 28016 21788
rect 27952 21728 28016 21732
rect 28032 21788 28096 21792
rect 28032 21732 28036 21788
rect 28036 21732 28092 21788
rect 28092 21732 28096 21788
rect 28032 21728 28096 21732
rect 28112 21788 28176 21792
rect 28112 21732 28116 21788
rect 28116 21732 28172 21788
rect 28172 21732 28176 21788
rect 28112 21728 28176 21732
rect 28192 21788 28256 21792
rect 28192 21732 28196 21788
rect 28196 21732 28252 21788
rect 28252 21732 28256 21788
rect 28192 21728 28256 21732
rect 37952 21788 38016 21792
rect 37952 21732 37956 21788
rect 37956 21732 38012 21788
rect 38012 21732 38016 21788
rect 37952 21728 38016 21732
rect 38032 21788 38096 21792
rect 38032 21732 38036 21788
rect 38036 21732 38092 21788
rect 38092 21732 38096 21788
rect 38032 21728 38096 21732
rect 38112 21788 38176 21792
rect 38112 21732 38116 21788
rect 38116 21732 38172 21788
rect 38172 21732 38176 21788
rect 38112 21728 38176 21732
rect 38192 21788 38256 21792
rect 38192 21732 38196 21788
rect 38196 21732 38252 21788
rect 38252 21732 38256 21788
rect 38192 21728 38256 21732
rect 47952 21788 48016 21792
rect 47952 21732 47956 21788
rect 47956 21732 48012 21788
rect 48012 21732 48016 21788
rect 47952 21728 48016 21732
rect 48032 21788 48096 21792
rect 48032 21732 48036 21788
rect 48036 21732 48092 21788
rect 48092 21732 48096 21788
rect 48032 21728 48096 21732
rect 48112 21788 48176 21792
rect 48112 21732 48116 21788
rect 48116 21732 48172 21788
rect 48172 21732 48176 21788
rect 48112 21728 48176 21732
rect 48192 21788 48256 21792
rect 48192 21732 48196 21788
rect 48196 21732 48252 21788
rect 48252 21732 48256 21788
rect 48192 21728 48256 21732
rect 28948 21524 29012 21588
rect 2952 21244 3016 21248
rect 2952 21188 2956 21244
rect 2956 21188 3012 21244
rect 3012 21188 3016 21244
rect 2952 21184 3016 21188
rect 3032 21244 3096 21248
rect 3032 21188 3036 21244
rect 3036 21188 3092 21244
rect 3092 21188 3096 21244
rect 3032 21184 3096 21188
rect 3112 21244 3176 21248
rect 3112 21188 3116 21244
rect 3116 21188 3172 21244
rect 3172 21188 3176 21244
rect 3112 21184 3176 21188
rect 3192 21244 3256 21248
rect 3192 21188 3196 21244
rect 3196 21188 3252 21244
rect 3252 21188 3256 21244
rect 3192 21184 3256 21188
rect 12952 21244 13016 21248
rect 12952 21188 12956 21244
rect 12956 21188 13012 21244
rect 13012 21188 13016 21244
rect 12952 21184 13016 21188
rect 13032 21244 13096 21248
rect 13032 21188 13036 21244
rect 13036 21188 13092 21244
rect 13092 21188 13096 21244
rect 13032 21184 13096 21188
rect 13112 21244 13176 21248
rect 13112 21188 13116 21244
rect 13116 21188 13172 21244
rect 13172 21188 13176 21244
rect 13112 21184 13176 21188
rect 13192 21244 13256 21248
rect 13192 21188 13196 21244
rect 13196 21188 13252 21244
rect 13252 21188 13256 21244
rect 13192 21184 13256 21188
rect 22952 21244 23016 21248
rect 22952 21188 22956 21244
rect 22956 21188 23012 21244
rect 23012 21188 23016 21244
rect 22952 21184 23016 21188
rect 23032 21244 23096 21248
rect 23032 21188 23036 21244
rect 23036 21188 23092 21244
rect 23092 21188 23096 21244
rect 23032 21184 23096 21188
rect 23112 21244 23176 21248
rect 23112 21188 23116 21244
rect 23116 21188 23172 21244
rect 23172 21188 23176 21244
rect 23112 21184 23176 21188
rect 23192 21244 23256 21248
rect 23192 21188 23196 21244
rect 23196 21188 23252 21244
rect 23252 21188 23256 21244
rect 23192 21184 23256 21188
rect 32952 21244 33016 21248
rect 32952 21188 32956 21244
rect 32956 21188 33012 21244
rect 33012 21188 33016 21244
rect 32952 21184 33016 21188
rect 33032 21244 33096 21248
rect 33032 21188 33036 21244
rect 33036 21188 33092 21244
rect 33092 21188 33096 21244
rect 33032 21184 33096 21188
rect 33112 21244 33176 21248
rect 33112 21188 33116 21244
rect 33116 21188 33172 21244
rect 33172 21188 33176 21244
rect 33112 21184 33176 21188
rect 33192 21244 33256 21248
rect 33192 21188 33196 21244
rect 33196 21188 33252 21244
rect 33252 21188 33256 21244
rect 33192 21184 33256 21188
rect 42952 21244 43016 21248
rect 42952 21188 42956 21244
rect 42956 21188 43012 21244
rect 43012 21188 43016 21244
rect 42952 21184 43016 21188
rect 43032 21244 43096 21248
rect 43032 21188 43036 21244
rect 43036 21188 43092 21244
rect 43092 21188 43096 21244
rect 43032 21184 43096 21188
rect 43112 21244 43176 21248
rect 43112 21188 43116 21244
rect 43116 21188 43172 21244
rect 43172 21188 43176 21244
rect 43112 21184 43176 21188
rect 43192 21244 43256 21248
rect 43192 21188 43196 21244
rect 43196 21188 43252 21244
rect 43252 21188 43256 21244
rect 43192 21184 43256 21188
rect 7952 20700 8016 20704
rect 7952 20644 7956 20700
rect 7956 20644 8012 20700
rect 8012 20644 8016 20700
rect 7952 20640 8016 20644
rect 8032 20700 8096 20704
rect 8032 20644 8036 20700
rect 8036 20644 8092 20700
rect 8092 20644 8096 20700
rect 8032 20640 8096 20644
rect 8112 20700 8176 20704
rect 8112 20644 8116 20700
rect 8116 20644 8172 20700
rect 8172 20644 8176 20700
rect 8112 20640 8176 20644
rect 8192 20700 8256 20704
rect 8192 20644 8196 20700
rect 8196 20644 8252 20700
rect 8252 20644 8256 20700
rect 8192 20640 8256 20644
rect 17952 20700 18016 20704
rect 17952 20644 17956 20700
rect 17956 20644 18012 20700
rect 18012 20644 18016 20700
rect 17952 20640 18016 20644
rect 18032 20700 18096 20704
rect 18032 20644 18036 20700
rect 18036 20644 18092 20700
rect 18092 20644 18096 20700
rect 18032 20640 18096 20644
rect 18112 20700 18176 20704
rect 18112 20644 18116 20700
rect 18116 20644 18172 20700
rect 18172 20644 18176 20700
rect 18112 20640 18176 20644
rect 18192 20700 18256 20704
rect 18192 20644 18196 20700
rect 18196 20644 18252 20700
rect 18252 20644 18256 20700
rect 18192 20640 18256 20644
rect 27952 20700 28016 20704
rect 27952 20644 27956 20700
rect 27956 20644 28012 20700
rect 28012 20644 28016 20700
rect 27952 20640 28016 20644
rect 28032 20700 28096 20704
rect 28032 20644 28036 20700
rect 28036 20644 28092 20700
rect 28092 20644 28096 20700
rect 28032 20640 28096 20644
rect 28112 20700 28176 20704
rect 28112 20644 28116 20700
rect 28116 20644 28172 20700
rect 28172 20644 28176 20700
rect 28112 20640 28176 20644
rect 28192 20700 28256 20704
rect 28192 20644 28196 20700
rect 28196 20644 28252 20700
rect 28252 20644 28256 20700
rect 28192 20640 28256 20644
rect 37952 20700 38016 20704
rect 37952 20644 37956 20700
rect 37956 20644 38012 20700
rect 38012 20644 38016 20700
rect 37952 20640 38016 20644
rect 38032 20700 38096 20704
rect 38032 20644 38036 20700
rect 38036 20644 38092 20700
rect 38092 20644 38096 20700
rect 38032 20640 38096 20644
rect 38112 20700 38176 20704
rect 38112 20644 38116 20700
rect 38116 20644 38172 20700
rect 38172 20644 38176 20700
rect 38112 20640 38176 20644
rect 38192 20700 38256 20704
rect 38192 20644 38196 20700
rect 38196 20644 38252 20700
rect 38252 20644 38256 20700
rect 38192 20640 38256 20644
rect 47952 20700 48016 20704
rect 47952 20644 47956 20700
rect 47956 20644 48012 20700
rect 48012 20644 48016 20700
rect 47952 20640 48016 20644
rect 48032 20700 48096 20704
rect 48032 20644 48036 20700
rect 48036 20644 48092 20700
rect 48092 20644 48096 20700
rect 48032 20640 48096 20644
rect 48112 20700 48176 20704
rect 48112 20644 48116 20700
rect 48116 20644 48172 20700
rect 48172 20644 48176 20700
rect 48112 20640 48176 20644
rect 48192 20700 48256 20704
rect 48192 20644 48196 20700
rect 48196 20644 48252 20700
rect 48252 20644 48256 20700
rect 48192 20640 48256 20644
rect 35388 20572 35452 20636
rect 28580 20360 28644 20364
rect 28580 20304 28594 20360
rect 28594 20304 28644 20360
rect 28580 20300 28644 20304
rect 2952 20156 3016 20160
rect 2952 20100 2956 20156
rect 2956 20100 3012 20156
rect 3012 20100 3016 20156
rect 2952 20096 3016 20100
rect 3032 20156 3096 20160
rect 3032 20100 3036 20156
rect 3036 20100 3092 20156
rect 3092 20100 3096 20156
rect 3032 20096 3096 20100
rect 3112 20156 3176 20160
rect 3112 20100 3116 20156
rect 3116 20100 3172 20156
rect 3172 20100 3176 20156
rect 3112 20096 3176 20100
rect 3192 20156 3256 20160
rect 3192 20100 3196 20156
rect 3196 20100 3252 20156
rect 3252 20100 3256 20156
rect 3192 20096 3256 20100
rect 12952 20156 13016 20160
rect 12952 20100 12956 20156
rect 12956 20100 13012 20156
rect 13012 20100 13016 20156
rect 12952 20096 13016 20100
rect 13032 20156 13096 20160
rect 13032 20100 13036 20156
rect 13036 20100 13092 20156
rect 13092 20100 13096 20156
rect 13032 20096 13096 20100
rect 13112 20156 13176 20160
rect 13112 20100 13116 20156
rect 13116 20100 13172 20156
rect 13172 20100 13176 20156
rect 13112 20096 13176 20100
rect 13192 20156 13256 20160
rect 13192 20100 13196 20156
rect 13196 20100 13252 20156
rect 13252 20100 13256 20156
rect 13192 20096 13256 20100
rect 22952 20156 23016 20160
rect 22952 20100 22956 20156
rect 22956 20100 23012 20156
rect 23012 20100 23016 20156
rect 22952 20096 23016 20100
rect 23032 20156 23096 20160
rect 23032 20100 23036 20156
rect 23036 20100 23092 20156
rect 23092 20100 23096 20156
rect 23032 20096 23096 20100
rect 23112 20156 23176 20160
rect 23112 20100 23116 20156
rect 23116 20100 23172 20156
rect 23172 20100 23176 20156
rect 23112 20096 23176 20100
rect 23192 20156 23256 20160
rect 23192 20100 23196 20156
rect 23196 20100 23252 20156
rect 23252 20100 23256 20156
rect 23192 20096 23256 20100
rect 32952 20156 33016 20160
rect 32952 20100 32956 20156
rect 32956 20100 33012 20156
rect 33012 20100 33016 20156
rect 32952 20096 33016 20100
rect 33032 20156 33096 20160
rect 33032 20100 33036 20156
rect 33036 20100 33092 20156
rect 33092 20100 33096 20156
rect 33032 20096 33096 20100
rect 33112 20156 33176 20160
rect 33112 20100 33116 20156
rect 33116 20100 33172 20156
rect 33172 20100 33176 20156
rect 33112 20096 33176 20100
rect 33192 20156 33256 20160
rect 33192 20100 33196 20156
rect 33196 20100 33252 20156
rect 33252 20100 33256 20156
rect 33192 20096 33256 20100
rect 42952 20156 43016 20160
rect 42952 20100 42956 20156
rect 42956 20100 43012 20156
rect 43012 20100 43016 20156
rect 42952 20096 43016 20100
rect 43032 20156 43096 20160
rect 43032 20100 43036 20156
rect 43036 20100 43092 20156
rect 43092 20100 43096 20156
rect 43032 20096 43096 20100
rect 43112 20156 43176 20160
rect 43112 20100 43116 20156
rect 43116 20100 43172 20156
rect 43172 20100 43176 20156
rect 43112 20096 43176 20100
rect 43192 20156 43256 20160
rect 43192 20100 43196 20156
rect 43196 20100 43252 20156
rect 43252 20100 43256 20156
rect 43192 20096 43256 20100
rect 28580 19680 28644 19684
rect 28580 19624 28594 19680
rect 28594 19624 28644 19680
rect 28580 19620 28644 19624
rect 7952 19612 8016 19616
rect 7952 19556 7956 19612
rect 7956 19556 8012 19612
rect 8012 19556 8016 19612
rect 7952 19552 8016 19556
rect 8032 19612 8096 19616
rect 8032 19556 8036 19612
rect 8036 19556 8092 19612
rect 8092 19556 8096 19612
rect 8032 19552 8096 19556
rect 8112 19612 8176 19616
rect 8112 19556 8116 19612
rect 8116 19556 8172 19612
rect 8172 19556 8176 19612
rect 8112 19552 8176 19556
rect 8192 19612 8256 19616
rect 8192 19556 8196 19612
rect 8196 19556 8252 19612
rect 8252 19556 8256 19612
rect 8192 19552 8256 19556
rect 17952 19612 18016 19616
rect 17952 19556 17956 19612
rect 17956 19556 18012 19612
rect 18012 19556 18016 19612
rect 17952 19552 18016 19556
rect 18032 19612 18096 19616
rect 18032 19556 18036 19612
rect 18036 19556 18092 19612
rect 18092 19556 18096 19612
rect 18032 19552 18096 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 27952 19612 28016 19616
rect 27952 19556 27956 19612
rect 27956 19556 28012 19612
rect 28012 19556 28016 19612
rect 27952 19552 28016 19556
rect 28032 19612 28096 19616
rect 28032 19556 28036 19612
rect 28036 19556 28092 19612
rect 28092 19556 28096 19612
rect 28032 19552 28096 19556
rect 28112 19612 28176 19616
rect 28112 19556 28116 19612
rect 28116 19556 28172 19612
rect 28172 19556 28176 19612
rect 28112 19552 28176 19556
rect 28192 19612 28256 19616
rect 28192 19556 28196 19612
rect 28196 19556 28252 19612
rect 28252 19556 28256 19612
rect 28192 19552 28256 19556
rect 37952 19612 38016 19616
rect 37952 19556 37956 19612
rect 37956 19556 38012 19612
rect 38012 19556 38016 19612
rect 37952 19552 38016 19556
rect 38032 19612 38096 19616
rect 38032 19556 38036 19612
rect 38036 19556 38092 19612
rect 38092 19556 38096 19612
rect 38032 19552 38096 19556
rect 38112 19612 38176 19616
rect 38112 19556 38116 19612
rect 38116 19556 38172 19612
rect 38172 19556 38176 19612
rect 38112 19552 38176 19556
rect 38192 19612 38256 19616
rect 38192 19556 38196 19612
rect 38196 19556 38252 19612
rect 38252 19556 38256 19612
rect 38192 19552 38256 19556
rect 47952 19612 48016 19616
rect 47952 19556 47956 19612
rect 47956 19556 48012 19612
rect 48012 19556 48016 19612
rect 47952 19552 48016 19556
rect 48032 19612 48096 19616
rect 48032 19556 48036 19612
rect 48036 19556 48092 19612
rect 48092 19556 48096 19612
rect 48032 19552 48096 19556
rect 48112 19612 48176 19616
rect 48112 19556 48116 19612
rect 48116 19556 48172 19612
rect 48172 19556 48176 19612
rect 48112 19552 48176 19556
rect 48192 19612 48256 19616
rect 48192 19556 48196 19612
rect 48196 19556 48252 19612
rect 48252 19556 48256 19612
rect 48192 19552 48256 19556
rect 28948 19212 29012 19276
rect 2952 19068 3016 19072
rect 2952 19012 2956 19068
rect 2956 19012 3012 19068
rect 3012 19012 3016 19068
rect 2952 19008 3016 19012
rect 3032 19068 3096 19072
rect 3032 19012 3036 19068
rect 3036 19012 3092 19068
rect 3092 19012 3096 19068
rect 3032 19008 3096 19012
rect 3112 19068 3176 19072
rect 3112 19012 3116 19068
rect 3116 19012 3172 19068
rect 3172 19012 3176 19068
rect 3112 19008 3176 19012
rect 3192 19068 3256 19072
rect 3192 19012 3196 19068
rect 3196 19012 3252 19068
rect 3252 19012 3256 19068
rect 3192 19008 3256 19012
rect 12952 19068 13016 19072
rect 12952 19012 12956 19068
rect 12956 19012 13012 19068
rect 13012 19012 13016 19068
rect 12952 19008 13016 19012
rect 13032 19068 13096 19072
rect 13032 19012 13036 19068
rect 13036 19012 13092 19068
rect 13092 19012 13096 19068
rect 13032 19008 13096 19012
rect 13112 19068 13176 19072
rect 13112 19012 13116 19068
rect 13116 19012 13172 19068
rect 13172 19012 13176 19068
rect 13112 19008 13176 19012
rect 13192 19068 13256 19072
rect 13192 19012 13196 19068
rect 13196 19012 13252 19068
rect 13252 19012 13256 19068
rect 13192 19008 13256 19012
rect 22952 19068 23016 19072
rect 22952 19012 22956 19068
rect 22956 19012 23012 19068
rect 23012 19012 23016 19068
rect 22952 19008 23016 19012
rect 23032 19068 23096 19072
rect 23032 19012 23036 19068
rect 23036 19012 23092 19068
rect 23092 19012 23096 19068
rect 23032 19008 23096 19012
rect 23112 19068 23176 19072
rect 23112 19012 23116 19068
rect 23116 19012 23172 19068
rect 23172 19012 23176 19068
rect 23112 19008 23176 19012
rect 23192 19068 23256 19072
rect 23192 19012 23196 19068
rect 23196 19012 23252 19068
rect 23252 19012 23256 19068
rect 23192 19008 23256 19012
rect 32952 19068 33016 19072
rect 32952 19012 32956 19068
rect 32956 19012 33012 19068
rect 33012 19012 33016 19068
rect 32952 19008 33016 19012
rect 33032 19068 33096 19072
rect 33032 19012 33036 19068
rect 33036 19012 33092 19068
rect 33092 19012 33096 19068
rect 33032 19008 33096 19012
rect 33112 19068 33176 19072
rect 33112 19012 33116 19068
rect 33116 19012 33172 19068
rect 33172 19012 33176 19068
rect 33112 19008 33176 19012
rect 33192 19068 33256 19072
rect 33192 19012 33196 19068
rect 33196 19012 33252 19068
rect 33252 19012 33256 19068
rect 33192 19008 33256 19012
rect 42952 19068 43016 19072
rect 42952 19012 42956 19068
rect 42956 19012 43012 19068
rect 43012 19012 43016 19068
rect 42952 19008 43016 19012
rect 43032 19068 43096 19072
rect 43032 19012 43036 19068
rect 43036 19012 43092 19068
rect 43092 19012 43096 19068
rect 43032 19008 43096 19012
rect 43112 19068 43176 19072
rect 43112 19012 43116 19068
rect 43116 19012 43172 19068
rect 43172 19012 43176 19068
rect 43112 19008 43176 19012
rect 43192 19068 43256 19072
rect 43192 19012 43196 19068
rect 43196 19012 43252 19068
rect 43252 19012 43256 19068
rect 43192 19008 43256 19012
rect 7952 18524 8016 18528
rect 7952 18468 7956 18524
rect 7956 18468 8012 18524
rect 8012 18468 8016 18524
rect 7952 18464 8016 18468
rect 8032 18524 8096 18528
rect 8032 18468 8036 18524
rect 8036 18468 8092 18524
rect 8092 18468 8096 18524
rect 8032 18464 8096 18468
rect 8112 18524 8176 18528
rect 8112 18468 8116 18524
rect 8116 18468 8172 18524
rect 8172 18468 8176 18524
rect 8112 18464 8176 18468
rect 8192 18524 8256 18528
rect 8192 18468 8196 18524
rect 8196 18468 8252 18524
rect 8252 18468 8256 18524
rect 8192 18464 8256 18468
rect 17952 18524 18016 18528
rect 17952 18468 17956 18524
rect 17956 18468 18012 18524
rect 18012 18468 18016 18524
rect 17952 18464 18016 18468
rect 18032 18524 18096 18528
rect 18032 18468 18036 18524
rect 18036 18468 18092 18524
rect 18092 18468 18096 18524
rect 18032 18464 18096 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 27952 18524 28016 18528
rect 27952 18468 27956 18524
rect 27956 18468 28012 18524
rect 28012 18468 28016 18524
rect 27952 18464 28016 18468
rect 28032 18524 28096 18528
rect 28032 18468 28036 18524
rect 28036 18468 28092 18524
rect 28092 18468 28096 18524
rect 28032 18464 28096 18468
rect 28112 18524 28176 18528
rect 28112 18468 28116 18524
rect 28116 18468 28172 18524
rect 28172 18468 28176 18524
rect 28112 18464 28176 18468
rect 28192 18524 28256 18528
rect 28192 18468 28196 18524
rect 28196 18468 28252 18524
rect 28252 18468 28256 18524
rect 28192 18464 28256 18468
rect 37952 18524 38016 18528
rect 37952 18468 37956 18524
rect 37956 18468 38012 18524
rect 38012 18468 38016 18524
rect 37952 18464 38016 18468
rect 38032 18524 38096 18528
rect 38032 18468 38036 18524
rect 38036 18468 38092 18524
rect 38092 18468 38096 18524
rect 38032 18464 38096 18468
rect 38112 18524 38176 18528
rect 38112 18468 38116 18524
rect 38116 18468 38172 18524
rect 38172 18468 38176 18524
rect 38112 18464 38176 18468
rect 38192 18524 38256 18528
rect 38192 18468 38196 18524
rect 38196 18468 38252 18524
rect 38252 18468 38256 18524
rect 38192 18464 38256 18468
rect 47952 18524 48016 18528
rect 47952 18468 47956 18524
rect 47956 18468 48012 18524
rect 48012 18468 48016 18524
rect 47952 18464 48016 18468
rect 48032 18524 48096 18528
rect 48032 18468 48036 18524
rect 48036 18468 48092 18524
rect 48092 18468 48096 18524
rect 48032 18464 48096 18468
rect 48112 18524 48176 18528
rect 48112 18468 48116 18524
rect 48116 18468 48172 18524
rect 48172 18468 48176 18524
rect 48112 18464 48176 18468
rect 48192 18524 48256 18528
rect 48192 18468 48196 18524
rect 48196 18468 48252 18524
rect 48252 18468 48256 18524
rect 48192 18464 48256 18468
rect 2952 17980 3016 17984
rect 2952 17924 2956 17980
rect 2956 17924 3012 17980
rect 3012 17924 3016 17980
rect 2952 17920 3016 17924
rect 3032 17980 3096 17984
rect 3032 17924 3036 17980
rect 3036 17924 3092 17980
rect 3092 17924 3096 17980
rect 3032 17920 3096 17924
rect 3112 17980 3176 17984
rect 3112 17924 3116 17980
rect 3116 17924 3172 17980
rect 3172 17924 3176 17980
rect 3112 17920 3176 17924
rect 3192 17980 3256 17984
rect 3192 17924 3196 17980
rect 3196 17924 3252 17980
rect 3252 17924 3256 17980
rect 3192 17920 3256 17924
rect 12952 17980 13016 17984
rect 12952 17924 12956 17980
rect 12956 17924 13012 17980
rect 13012 17924 13016 17980
rect 12952 17920 13016 17924
rect 13032 17980 13096 17984
rect 13032 17924 13036 17980
rect 13036 17924 13092 17980
rect 13092 17924 13096 17980
rect 13032 17920 13096 17924
rect 13112 17980 13176 17984
rect 13112 17924 13116 17980
rect 13116 17924 13172 17980
rect 13172 17924 13176 17980
rect 13112 17920 13176 17924
rect 13192 17980 13256 17984
rect 13192 17924 13196 17980
rect 13196 17924 13252 17980
rect 13252 17924 13256 17980
rect 13192 17920 13256 17924
rect 22952 17980 23016 17984
rect 22952 17924 22956 17980
rect 22956 17924 23012 17980
rect 23012 17924 23016 17980
rect 22952 17920 23016 17924
rect 23032 17980 23096 17984
rect 23032 17924 23036 17980
rect 23036 17924 23092 17980
rect 23092 17924 23096 17980
rect 23032 17920 23096 17924
rect 23112 17980 23176 17984
rect 23112 17924 23116 17980
rect 23116 17924 23172 17980
rect 23172 17924 23176 17980
rect 23112 17920 23176 17924
rect 23192 17980 23256 17984
rect 23192 17924 23196 17980
rect 23196 17924 23252 17980
rect 23252 17924 23256 17980
rect 23192 17920 23256 17924
rect 32952 17980 33016 17984
rect 32952 17924 32956 17980
rect 32956 17924 33012 17980
rect 33012 17924 33016 17980
rect 32952 17920 33016 17924
rect 33032 17980 33096 17984
rect 33032 17924 33036 17980
rect 33036 17924 33092 17980
rect 33092 17924 33096 17980
rect 33032 17920 33096 17924
rect 33112 17980 33176 17984
rect 33112 17924 33116 17980
rect 33116 17924 33172 17980
rect 33172 17924 33176 17980
rect 33112 17920 33176 17924
rect 33192 17980 33256 17984
rect 33192 17924 33196 17980
rect 33196 17924 33252 17980
rect 33252 17924 33256 17980
rect 33192 17920 33256 17924
rect 42952 17980 43016 17984
rect 42952 17924 42956 17980
rect 42956 17924 43012 17980
rect 43012 17924 43016 17980
rect 42952 17920 43016 17924
rect 43032 17980 43096 17984
rect 43032 17924 43036 17980
rect 43036 17924 43092 17980
rect 43092 17924 43096 17980
rect 43032 17920 43096 17924
rect 43112 17980 43176 17984
rect 43112 17924 43116 17980
rect 43116 17924 43172 17980
rect 43172 17924 43176 17980
rect 43112 17920 43176 17924
rect 43192 17980 43256 17984
rect 43192 17924 43196 17980
rect 43196 17924 43252 17980
rect 43252 17924 43256 17980
rect 43192 17920 43256 17924
rect 7952 17436 8016 17440
rect 7952 17380 7956 17436
rect 7956 17380 8012 17436
rect 8012 17380 8016 17436
rect 7952 17376 8016 17380
rect 8032 17436 8096 17440
rect 8032 17380 8036 17436
rect 8036 17380 8092 17436
rect 8092 17380 8096 17436
rect 8032 17376 8096 17380
rect 8112 17436 8176 17440
rect 8112 17380 8116 17436
rect 8116 17380 8172 17436
rect 8172 17380 8176 17436
rect 8112 17376 8176 17380
rect 8192 17436 8256 17440
rect 8192 17380 8196 17436
rect 8196 17380 8252 17436
rect 8252 17380 8256 17436
rect 8192 17376 8256 17380
rect 17952 17436 18016 17440
rect 17952 17380 17956 17436
rect 17956 17380 18012 17436
rect 18012 17380 18016 17436
rect 17952 17376 18016 17380
rect 18032 17436 18096 17440
rect 18032 17380 18036 17436
rect 18036 17380 18092 17436
rect 18092 17380 18096 17436
rect 18032 17376 18096 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 27952 17436 28016 17440
rect 27952 17380 27956 17436
rect 27956 17380 28012 17436
rect 28012 17380 28016 17436
rect 27952 17376 28016 17380
rect 28032 17436 28096 17440
rect 28032 17380 28036 17436
rect 28036 17380 28092 17436
rect 28092 17380 28096 17436
rect 28032 17376 28096 17380
rect 28112 17436 28176 17440
rect 28112 17380 28116 17436
rect 28116 17380 28172 17436
rect 28172 17380 28176 17436
rect 28112 17376 28176 17380
rect 28192 17436 28256 17440
rect 28192 17380 28196 17436
rect 28196 17380 28252 17436
rect 28252 17380 28256 17436
rect 28192 17376 28256 17380
rect 37952 17436 38016 17440
rect 37952 17380 37956 17436
rect 37956 17380 38012 17436
rect 38012 17380 38016 17436
rect 37952 17376 38016 17380
rect 38032 17436 38096 17440
rect 38032 17380 38036 17436
rect 38036 17380 38092 17436
rect 38092 17380 38096 17436
rect 38032 17376 38096 17380
rect 38112 17436 38176 17440
rect 38112 17380 38116 17436
rect 38116 17380 38172 17436
rect 38172 17380 38176 17436
rect 38112 17376 38176 17380
rect 38192 17436 38256 17440
rect 38192 17380 38196 17436
rect 38196 17380 38252 17436
rect 38252 17380 38256 17436
rect 38192 17376 38256 17380
rect 47952 17436 48016 17440
rect 47952 17380 47956 17436
rect 47956 17380 48012 17436
rect 48012 17380 48016 17436
rect 47952 17376 48016 17380
rect 48032 17436 48096 17440
rect 48032 17380 48036 17436
rect 48036 17380 48092 17436
rect 48092 17380 48096 17436
rect 48032 17376 48096 17380
rect 48112 17436 48176 17440
rect 48112 17380 48116 17436
rect 48116 17380 48172 17436
rect 48172 17380 48176 17436
rect 48112 17376 48176 17380
rect 48192 17436 48256 17440
rect 48192 17380 48196 17436
rect 48196 17380 48252 17436
rect 48252 17380 48256 17436
rect 48192 17376 48256 17380
rect 2952 16892 3016 16896
rect 2952 16836 2956 16892
rect 2956 16836 3012 16892
rect 3012 16836 3016 16892
rect 2952 16832 3016 16836
rect 3032 16892 3096 16896
rect 3032 16836 3036 16892
rect 3036 16836 3092 16892
rect 3092 16836 3096 16892
rect 3032 16832 3096 16836
rect 3112 16892 3176 16896
rect 3112 16836 3116 16892
rect 3116 16836 3172 16892
rect 3172 16836 3176 16892
rect 3112 16832 3176 16836
rect 3192 16892 3256 16896
rect 3192 16836 3196 16892
rect 3196 16836 3252 16892
rect 3252 16836 3256 16892
rect 3192 16832 3256 16836
rect 12952 16892 13016 16896
rect 12952 16836 12956 16892
rect 12956 16836 13012 16892
rect 13012 16836 13016 16892
rect 12952 16832 13016 16836
rect 13032 16892 13096 16896
rect 13032 16836 13036 16892
rect 13036 16836 13092 16892
rect 13092 16836 13096 16892
rect 13032 16832 13096 16836
rect 13112 16892 13176 16896
rect 13112 16836 13116 16892
rect 13116 16836 13172 16892
rect 13172 16836 13176 16892
rect 13112 16832 13176 16836
rect 13192 16892 13256 16896
rect 13192 16836 13196 16892
rect 13196 16836 13252 16892
rect 13252 16836 13256 16892
rect 13192 16832 13256 16836
rect 22952 16892 23016 16896
rect 22952 16836 22956 16892
rect 22956 16836 23012 16892
rect 23012 16836 23016 16892
rect 22952 16832 23016 16836
rect 23032 16892 23096 16896
rect 23032 16836 23036 16892
rect 23036 16836 23092 16892
rect 23092 16836 23096 16892
rect 23032 16832 23096 16836
rect 23112 16892 23176 16896
rect 23112 16836 23116 16892
rect 23116 16836 23172 16892
rect 23172 16836 23176 16892
rect 23112 16832 23176 16836
rect 23192 16892 23256 16896
rect 23192 16836 23196 16892
rect 23196 16836 23252 16892
rect 23252 16836 23256 16892
rect 23192 16832 23256 16836
rect 32952 16892 33016 16896
rect 32952 16836 32956 16892
rect 32956 16836 33012 16892
rect 33012 16836 33016 16892
rect 32952 16832 33016 16836
rect 33032 16892 33096 16896
rect 33032 16836 33036 16892
rect 33036 16836 33092 16892
rect 33092 16836 33096 16892
rect 33032 16832 33096 16836
rect 33112 16892 33176 16896
rect 33112 16836 33116 16892
rect 33116 16836 33172 16892
rect 33172 16836 33176 16892
rect 33112 16832 33176 16836
rect 33192 16892 33256 16896
rect 33192 16836 33196 16892
rect 33196 16836 33252 16892
rect 33252 16836 33256 16892
rect 33192 16832 33256 16836
rect 42952 16892 43016 16896
rect 42952 16836 42956 16892
rect 42956 16836 43012 16892
rect 43012 16836 43016 16892
rect 42952 16832 43016 16836
rect 43032 16892 43096 16896
rect 43032 16836 43036 16892
rect 43036 16836 43092 16892
rect 43092 16836 43096 16892
rect 43032 16832 43096 16836
rect 43112 16892 43176 16896
rect 43112 16836 43116 16892
rect 43116 16836 43172 16892
rect 43172 16836 43176 16892
rect 43112 16832 43176 16836
rect 43192 16892 43256 16896
rect 43192 16836 43196 16892
rect 43196 16836 43252 16892
rect 43252 16836 43256 16892
rect 43192 16832 43256 16836
rect 7952 16348 8016 16352
rect 7952 16292 7956 16348
rect 7956 16292 8012 16348
rect 8012 16292 8016 16348
rect 7952 16288 8016 16292
rect 8032 16348 8096 16352
rect 8032 16292 8036 16348
rect 8036 16292 8092 16348
rect 8092 16292 8096 16348
rect 8032 16288 8096 16292
rect 8112 16348 8176 16352
rect 8112 16292 8116 16348
rect 8116 16292 8172 16348
rect 8172 16292 8176 16348
rect 8112 16288 8176 16292
rect 8192 16348 8256 16352
rect 8192 16292 8196 16348
rect 8196 16292 8252 16348
rect 8252 16292 8256 16348
rect 8192 16288 8256 16292
rect 17952 16348 18016 16352
rect 17952 16292 17956 16348
rect 17956 16292 18012 16348
rect 18012 16292 18016 16348
rect 17952 16288 18016 16292
rect 18032 16348 18096 16352
rect 18032 16292 18036 16348
rect 18036 16292 18092 16348
rect 18092 16292 18096 16348
rect 18032 16288 18096 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 27952 16348 28016 16352
rect 27952 16292 27956 16348
rect 27956 16292 28012 16348
rect 28012 16292 28016 16348
rect 27952 16288 28016 16292
rect 28032 16348 28096 16352
rect 28032 16292 28036 16348
rect 28036 16292 28092 16348
rect 28092 16292 28096 16348
rect 28032 16288 28096 16292
rect 28112 16348 28176 16352
rect 28112 16292 28116 16348
rect 28116 16292 28172 16348
rect 28172 16292 28176 16348
rect 28112 16288 28176 16292
rect 28192 16348 28256 16352
rect 28192 16292 28196 16348
rect 28196 16292 28252 16348
rect 28252 16292 28256 16348
rect 28192 16288 28256 16292
rect 37952 16348 38016 16352
rect 37952 16292 37956 16348
rect 37956 16292 38012 16348
rect 38012 16292 38016 16348
rect 37952 16288 38016 16292
rect 38032 16348 38096 16352
rect 38032 16292 38036 16348
rect 38036 16292 38092 16348
rect 38092 16292 38096 16348
rect 38032 16288 38096 16292
rect 38112 16348 38176 16352
rect 38112 16292 38116 16348
rect 38116 16292 38172 16348
rect 38172 16292 38176 16348
rect 38112 16288 38176 16292
rect 38192 16348 38256 16352
rect 38192 16292 38196 16348
rect 38196 16292 38252 16348
rect 38252 16292 38256 16348
rect 38192 16288 38256 16292
rect 47952 16348 48016 16352
rect 47952 16292 47956 16348
rect 47956 16292 48012 16348
rect 48012 16292 48016 16348
rect 47952 16288 48016 16292
rect 48032 16348 48096 16352
rect 48032 16292 48036 16348
rect 48036 16292 48092 16348
rect 48092 16292 48096 16348
rect 48032 16288 48096 16292
rect 48112 16348 48176 16352
rect 48112 16292 48116 16348
rect 48116 16292 48172 16348
rect 48172 16292 48176 16348
rect 48112 16288 48176 16292
rect 48192 16348 48256 16352
rect 48192 16292 48196 16348
rect 48196 16292 48252 16348
rect 48252 16292 48256 16348
rect 48192 16288 48256 16292
rect 2952 15804 3016 15808
rect 2952 15748 2956 15804
rect 2956 15748 3012 15804
rect 3012 15748 3016 15804
rect 2952 15744 3016 15748
rect 3032 15804 3096 15808
rect 3032 15748 3036 15804
rect 3036 15748 3092 15804
rect 3092 15748 3096 15804
rect 3032 15744 3096 15748
rect 3112 15804 3176 15808
rect 3112 15748 3116 15804
rect 3116 15748 3172 15804
rect 3172 15748 3176 15804
rect 3112 15744 3176 15748
rect 3192 15804 3256 15808
rect 3192 15748 3196 15804
rect 3196 15748 3252 15804
rect 3252 15748 3256 15804
rect 3192 15744 3256 15748
rect 12952 15804 13016 15808
rect 12952 15748 12956 15804
rect 12956 15748 13012 15804
rect 13012 15748 13016 15804
rect 12952 15744 13016 15748
rect 13032 15804 13096 15808
rect 13032 15748 13036 15804
rect 13036 15748 13092 15804
rect 13092 15748 13096 15804
rect 13032 15744 13096 15748
rect 13112 15804 13176 15808
rect 13112 15748 13116 15804
rect 13116 15748 13172 15804
rect 13172 15748 13176 15804
rect 13112 15744 13176 15748
rect 13192 15804 13256 15808
rect 13192 15748 13196 15804
rect 13196 15748 13252 15804
rect 13252 15748 13256 15804
rect 13192 15744 13256 15748
rect 22952 15804 23016 15808
rect 22952 15748 22956 15804
rect 22956 15748 23012 15804
rect 23012 15748 23016 15804
rect 22952 15744 23016 15748
rect 23032 15804 23096 15808
rect 23032 15748 23036 15804
rect 23036 15748 23092 15804
rect 23092 15748 23096 15804
rect 23032 15744 23096 15748
rect 23112 15804 23176 15808
rect 23112 15748 23116 15804
rect 23116 15748 23172 15804
rect 23172 15748 23176 15804
rect 23112 15744 23176 15748
rect 23192 15804 23256 15808
rect 23192 15748 23196 15804
rect 23196 15748 23252 15804
rect 23252 15748 23256 15804
rect 23192 15744 23256 15748
rect 32952 15804 33016 15808
rect 32952 15748 32956 15804
rect 32956 15748 33012 15804
rect 33012 15748 33016 15804
rect 32952 15744 33016 15748
rect 33032 15804 33096 15808
rect 33032 15748 33036 15804
rect 33036 15748 33092 15804
rect 33092 15748 33096 15804
rect 33032 15744 33096 15748
rect 33112 15804 33176 15808
rect 33112 15748 33116 15804
rect 33116 15748 33172 15804
rect 33172 15748 33176 15804
rect 33112 15744 33176 15748
rect 33192 15804 33256 15808
rect 33192 15748 33196 15804
rect 33196 15748 33252 15804
rect 33252 15748 33256 15804
rect 33192 15744 33256 15748
rect 42952 15804 43016 15808
rect 42952 15748 42956 15804
rect 42956 15748 43012 15804
rect 43012 15748 43016 15804
rect 42952 15744 43016 15748
rect 43032 15804 43096 15808
rect 43032 15748 43036 15804
rect 43036 15748 43092 15804
rect 43092 15748 43096 15804
rect 43032 15744 43096 15748
rect 43112 15804 43176 15808
rect 43112 15748 43116 15804
rect 43116 15748 43172 15804
rect 43172 15748 43176 15804
rect 43112 15744 43176 15748
rect 43192 15804 43256 15808
rect 43192 15748 43196 15804
rect 43196 15748 43252 15804
rect 43252 15748 43256 15804
rect 43192 15744 43256 15748
rect 7952 15260 8016 15264
rect 7952 15204 7956 15260
rect 7956 15204 8012 15260
rect 8012 15204 8016 15260
rect 7952 15200 8016 15204
rect 8032 15260 8096 15264
rect 8032 15204 8036 15260
rect 8036 15204 8092 15260
rect 8092 15204 8096 15260
rect 8032 15200 8096 15204
rect 8112 15260 8176 15264
rect 8112 15204 8116 15260
rect 8116 15204 8172 15260
rect 8172 15204 8176 15260
rect 8112 15200 8176 15204
rect 8192 15260 8256 15264
rect 8192 15204 8196 15260
rect 8196 15204 8252 15260
rect 8252 15204 8256 15260
rect 8192 15200 8256 15204
rect 17952 15260 18016 15264
rect 17952 15204 17956 15260
rect 17956 15204 18012 15260
rect 18012 15204 18016 15260
rect 17952 15200 18016 15204
rect 18032 15260 18096 15264
rect 18032 15204 18036 15260
rect 18036 15204 18092 15260
rect 18092 15204 18096 15260
rect 18032 15200 18096 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 27952 15260 28016 15264
rect 27952 15204 27956 15260
rect 27956 15204 28012 15260
rect 28012 15204 28016 15260
rect 27952 15200 28016 15204
rect 28032 15260 28096 15264
rect 28032 15204 28036 15260
rect 28036 15204 28092 15260
rect 28092 15204 28096 15260
rect 28032 15200 28096 15204
rect 28112 15260 28176 15264
rect 28112 15204 28116 15260
rect 28116 15204 28172 15260
rect 28172 15204 28176 15260
rect 28112 15200 28176 15204
rect 28192 15260 28256 15264
rect 28192 15204 28196 15260
rect 28196 15204 28252 15260
rect 28252 15204 28256 15260
rect 28192 15200 28256 15204
rect 37952 15260 38016 15264
rect 37952 15204 37956 15260
rect 37956 15204 38012 15260
rect 38012 15204 38016 15260
rect 37952 15200 38016 15204
rect 38032 15260 38096 15264
rect 38032 15204 38036 15260
rect 38036 15204 38092 15260
rect 38092 15204 38096 15260
rect 38032 15200 38096 15204
rect 38112 15260 38176 15264
rect 38112 15204 38116 15260
rect 38116 15204 38172 15260
rect 38172 15204 38176 15260
rect 38112 15200 38176 15204
rect 38192 15260 38256 15264
rect 38192 15204 38196 15260
rect 38196 15204 38252 15260
rect 38252 15204 38256 15260
rect 38192 15200 38256 15204
rect 47952 15260 48016 15264
rect 47952 15204 47956 15260
rect 47956 15204 48012 15260
rect 48012 15204 48016 15260
rect 47952 15200 48016 15204
rect 48032 15260 48096 15264
rect 48032 15204 48036 15260
rect 48036 15204 48092 15260
rect 48092 15204 48096 15260
rect 48032 15200 48096 15204
rect 48112 15260 48176 15264
rect 48112 15204 48116 15260
rect 48116 15204 48172 15260
rect 48172 15204 48176 15260
rect 48112 15200 48176 15204
rect 48192 15260 48256 15264
rect 48192 15204 48196 15260
rect 48196 15204 48252 15260
rect 48252 15204 48256 15260
rect 48192 15200 48256 15204
rect 2952 14716 3016 14720
rect 2952 14660 2956 14716
rect 2956 14660 3012 14716
rect 3012 14660 3016 14716
rect 2952 14656 3016 14660
rect 3032 14716 3096 14720
rect 3032 14660 3036 14716
rect 3036 14660 3092 14716
rect 3092 14660 3096 14716
rect 3032 14656 3096 14660
rect 3112 14716 3176 14720
rect 3112 14660 3116 14716
rect 3116 14660 3172 14716
rect 3172 14660 3176 14716
rect 3112 14656 3176 14660
rect 3192 14716 3256 14720
rect 3192 14660 3196 14716
rect 3196 14660 3252 14716
rect 3252 14660 3256 14716
rect 3192 14656 3256 14660
rect 12952 14716 13016 14720
rect 12952 14660 12956 14716
rect 12956 14660 13012 14716
rect 13012 14660 13016 14716
rect 12952 14656 13016 14660
rect 13032 14716 13096 14720
rect 13032 14660 13036 14716
rect 13036 14660 13092 14716
rect 13092 14660 13096 14716
rect 13032 14656 13096 14660
rect 13112 14716 13176 14720
rect 13112 14660 13116 14716
rect 13116 14660 13172 14716
rect 13172 14660 13176 14716
rect 13112 14656 13176 14660
rect 13192 14716 13256 14720
rect 13192 14660 13196 14716
rect 13196 14660 13252 14716
rect 13252 14660 13256 14716
rect 13192 14656 13256 14660
rect 22952 14716 23016 14720
rect 22952 14660 22956 14716
rect 22956 14660 23012 14716
rect 23012 14660 23016 14716
rect 22952 14656 23016 14660
rect 23032 14716 23096 14720
rect 23032 14660 23036 14716
rect 23036 14660 23092 14716
rect 23092 14660 23096 14716
rect 23032 14656 23096 14660
rect 23112 14716 23176 14720
rect 23112 14660 23116 14716
rect 23116 14660 23172 14716
rect 23172 14660 23176 14716
rect 23112 14656 23176 14660
rect 23192 14716 23256 14720
rect 23192 14660 23196 14716
rect 23196 14660 23252 14716
rect 23252 14660 23256 14716
rect 23192 14656 23256 14660
rect 32952 14716 33016 14720
rect 32952 14660 32956 14716
rect 32956 14660 33012 14716
rect 33012 14660 33016 14716
rect 32952 14656 33016 14660
rect 33032 14716 33096 14720
rect 33032 14660 33036 14716
rect 33036 14660 33092 14716
rect 33092 14660 33096 14716
rect 33032 14656 33096 14660
rect 33112 14716 33176 14720
rect 33112 14660 33116 14716
rect 33116 14660 33172 14716
rect 33172 14660 33176 14716
rect 33112 14656 33176 14660
rect 33192 14716 33256 14720
rect 33192 14660 33196 14716
rect 33196 14660 33252 14716
rect 33252 14660 33256 14716
rect 33192 14656 33256 14660
rect 42952 14716 43016 14720
rect 42952 14660 42956 14716
rect 42956 14660 43012 14716
rect 43012 14660 43016 14716
rect 42952 14656 43016 14660
rect 43032 14716 43096 14720
rect 43032 14660 43036 14716
rect 43036 14660 43092 14716
rect 43092 14660 43096 14716
rect 43032 14656 43096 14660
rect 43112 14716 43176 14720
rect 43112 14660 43116 14716
rect 43116 14660 43172 14716
rect 43172 14660 43176 14716
rect 43112 14656 43176 14660
rect 43192 14716 43256 14720
rect 43192 14660 43196 14716
rect 43196 14660 43252 14716
rect 43252 14660 43256 14716
rect 43192 14656 43256 14660
rect 32076 14452 32140 14516
rect 7952 14172 8016 14176
rect 7952 14116 7956 14172
rect 7956 14116 8012 14172
rect 8012 14116 8016 14172
rect 7952 14112 8016 14116
rect 8032 14172 8096 14176
rect 8032 14116 8036 14172
rect 8036 14116 8092 14172
rect 8092 14116 8096 14172
rect 8032 14112 8096 14116
rect 8112 14172 8176 14176
rect 8112 14116 8116 14172
rect 8116 14116 8172 14172
rect 8172 14116 8176 14172
rect 8112 14112 8176 14116
rect 8192 14172 8256 14176
rect 8192 14116 8196 14172
rect 8196 14116 8252 14172
rect 8252 14116 8256 14172
rect 8192 14112 8256 14116
rect 17952 14172 18016 14176
rect 17952 14116 17956 14172
rect 17956 14116 18012 14172
rect 18012 14116 18016 14172
rect 17952 14112 18016 14116
rect 18032 14172 18096 14176
rect 18032 14116 18036 14172
rect 18036 14116 18092 14172
rect 18092 14116 18096 14172
rect 18032 14112 18096 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 27952 14172 28016 14176
rect 27952 14116 27956 14172
rect 27956 14116 28012 14172
rect 28012 14116 28016 14172
rect 27952 14112 28016 14116
rect 28032 14172 28096 14176
rect 28032 14116 28036 14172
rect 28036 14116 28092 14172
rect 28092 14116 28096 14172
rect 28032 14112 28096 14116
rect 28112 14172 28176 14176
rect 28112 14116 28116 14172
rect 28116 14116 28172 14172
rect 28172 14116 28176 14172
rect 28112 14112 28176 14116
rect 28192 14172 28256 14176
rect 28192 14116 28196 14172
rect 28196 14116 28252 14172
rect 28252 14116 28256 14172
rect 28192 14112 28256 14116
rect 37952 14172 38016 14176
rect 37952 14116 37956 14172
rect 37956 14116 38012 14172
rect 38012 14116 38016 14172
rect 37952 14112 38016 14116
rect 38032 14172 38096 14176
rect 38032 14116 38036 14172
rect 38036 14116 38092 14172
rect 38092 14116 38096 14172
rect 38032 14112 38096 14116
rect 38112 14172 38176 14176
rect 38112 14116 38116 14172
rect 38116 14116 38172 14172
rect 38172 14116 38176 14172
rect 38112 14112 38176 14116
rect 38192 14172 38256 14176
rect 38192 14116 38196 14172
rect 38196 14116 38252 14172
rect 38252 14116 38256 14172
rect 38192 14112 38256 14116
rect 47952 14172 48016 14176
rect 47952 14116 47956 14172
rect 47956 14116 48012 14172
rect 48012 14116 48016 14172
rect 47952 14112 48016 14116
rect 48032 14172 48096 14176
rect 48032 14116 48036 14172
rect 48036 14116 48092 14172
rect 48092 14116 48096 14172
rect 48032 14112 48096 14116
rect 48112 14172 48176 14176
rect 48112 14116 48116 14172
rect 48116 14116 48172 14172
rect 48172 14116 48176 14172
rect 48112 14112 48176 14116
rect 48192 14172 48256 14176
rect 48192 14116 48196 14172
rect 48196 14116 48252 14172
rect 48252 14116 48256 14172
rect 48192 14112 48256 14116
rect 15700 13832 15764 13836
rect 15700 13776 15714 13832
rect 15714 13776 15764 13832
rect 15700 13772 15764 13776
rect 2952 13628 3016 13632
rect 2952 13572 2956 13628
rect 2956 13572 3012 13628
rect 3012 13572 3016 13628
rect 2952 13568 3016 13572
rect 3032 13628 3096 13632
rect 3032 13572 3036 13628
rect 3036 13572 3092 13628
rect 3092 13572 3096 13628
rect 3032 13568 3096 13572
rect 3112 13628 3176 13632
rect 3112 13572 3116 13628
rect 3116 13572 3172 13628
rect 3172 13572 3176 13628
rect 3112 13568 3176 13572
rect 3192 13628 3256 13632
rect 3192 13572 3196 13628
rect 3196 13572 3252 13628
rect 3252 13572 3256 13628
rect 3192 13568 3256 13572
rect 12952 13628 13016 13632
rect 12952 13572 12956 13628
rect 12956 13572 13012 13628
rect 13012 13572 13016 13628
rect 12952 13568 13016 13572
rect 13032 13628 13096 13632
rect 13032 13572 13036 13628
rect 13036 13572 13092 13628
rect 13092 13572 13096 13628
rect 13032 13568 13096 13572
rect 13112 13628 13176 13632
rect 13112 13572 13116 13628
rect 13116 13572 13172 13628
rect 13172 13572 13176 13628
rect 13112 13568 13176 13572
rect 13192 13628 13256 13632
rect 13192 13572 13196 13628
rect 13196 13572 13252 13628
rect 13252 13572 13256 13628
rect 13192 13568 13256 13572
rect 22952 13628 23016 13632
rect 22952 13572 22956 13628
rect 22956 13572 23012 13628
rect 23012 13572 23016 13628
rect 22952 13568 23016 13572
rect 23032 13628 23096 13632
rect 23032 13572 23036 13628
rect 23036 13572 23092 13628
rect 23092 13572 23096 13628
rect 23032 13568 23096 13572
rect 23112 13628 23176 13632
rect 23112 13572 23116 13628
rect 23116 13572 23172 13628
rect 23172 13572 23176 13628
rect 23112 13568 23176 13572
rect 23192 13628 23256 13632
rect 23192 13572 23196 13628
rect 23196 13572 23252 13628
rect 23252 13572 23256 13628
rect 23192 13568 23256 13572
rect 32952 13628 33016 13632
rect 32952 13572 32956 13628
rect 32956 13572 33012 13628
rect 33012 13572 33016 13628
rect 32952 13568 33016 13572
rect 33032 13628 33096 13632
rect 33032 13572 33036 13628
rect 33036 13572 33092 13628
rect 33092 13572 33096 13628
rect 33032 13568 33096 13572
rect 33112 13628 33176 13632
rect 33112 13572 33116 13628
rect 33116 13572 33172 13628
rect 33172 13572 33176 13628
rect 33112 13568 33176 13572
rect 33192 13628 33256 13632
rect 33192 13572 33196 13628
rect 33196 13572 33252 13628
rect 33252 13572 33256 13628
rect 33192 13568 33256 13572
rect 42952 13628 43016 13632
rect 42952 13572 42956 13628
rect 42956 13572 43012 13628
rect 43012 13572 43016 13628
rect 42952 13568 43016 13572
rect 43032 13628 43096 13632
rect 43032 13572 43036 13628
rect 43036 13572 43092 13628
rect 43092 13572 43096 13628
rect 43032 13568 43096 13572
rect 43112 13628 43176 13632
rect 43112 13572 43116 13628
rect 43116 13572 43172 13628
rect 43172 13572 43176 13628
rect 43112 13568 43176 13572
rect 43192 13628 43256 13632
rect 43192 13572 43196 13628
rect 43196 13572 43252 13628
rect 43252 13572 43256 13628
rect 43192 13568 43256 13572
rect 7952 13084 8016 13088
rect 7952 13028 7956 13084
rect 7956 13028 8012 13084
rect 8012 13028 8016 13084
rect 7952 13024 8016 13028
rect 8032 13084 8096 13088
rect 8032 13028 8036 13084
rect 8036 13028 8092 13084
rect 8092 13028 8096 13084
rect 8032 13024 8096 13028
rect 8112 13084 8176 13088
rect 8112 13028 8116 13084
rect 8116 13028 8172 13084
rect 8172 13028 8176 13084
rect 8112 13024 8176 13028
rect 8192 13084 8256 13088
rect 8192 13028 8196 13084
rect 8196 13028 8252 13084
rect 8252 13028 8256 13084
rect 8192 13024 8256 13028
rect 17952 13084 18016 13088
rect 17952 13028 17956 13084
rect 17956 13028 18012 13084
rect 18012 13028 18016 13084
rect 17952 13024 18016 13028
rect 18032 13084 18096 13088
rect 18032 13028 18036 13084
rect 18036 13028 18092 13084
rect 18092 13028 18096 13084
rect 18032 13024 18096 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 27952 13084 28016 13088
rect 27952 13028 27956 13084
rect 27956 13028 28012 13084
rect 28012 13028 28016 13084
rect 27952 13024 28016 13028
rect 28032 13084 28096 13088
rect 28032 13028 28036 13084
rect 28036 13028 28092 13084
rect 28092 13028 28096 13084
rect 28032 13024 28096 13028
rect 28112 13084 28176 13088
rect 28112 13028 28116 13084
rect 28116 13028 28172 13084
rect 28172 13028 28176 13084
rect 28112 13024 28176 13028
rect 28192 13084 28256 13088
rect 28192 13028 28196 13084
rect 28196 13028 28252 13084
rect 28252 13028 28256 13084
rect 28192 13024 28256 13028
rect 37952 13084 38016 13088
rect 37952 13028 37956 13084
rect 37956 13028 38012 13084
rect 38012 13028 38016 13084
rect 37952 13024 38016 13028
rect 38032 13084 38096 13088
rect 38032 13028 38036 13084
rect 38036 13028 38092 13084
rect 38092 13028 38096 13084
rect 38032 13024 38096 13028
rect 38112 13084 38176 13088
rect 38112 13028 38116 13084
rect 38116 13028 38172 13084
rect 38172 13028 38176 13084
rect 38112 13024 38176 13028
rect 38192 13084 38256 13088
rect 38192 13028 38196 13084
rect 38196 13028 38252 13084
rect 38252 13028 38256 13084
rect 38192 13024 38256 13028
rect 47952 13084 48016 13088
rect 47952 13028 47956 13084
rect 47956 13028 48012 13084
rect 48012 13028 48016 13084
rect 47952 13024 48016 13028
rect 48032 13084 48096 13088
rect 48032 13028 48036 13084
rect 48036 13028 48092 13084
rect 48092 13028 48096 13084
rect 48032 13024 48096 13028
rect 48112 13084 48176 13088
rect 48112 13028 48116 13084
rect 48116 13028 48172 13084
rect 48172 13028 48176 13084
rect 48112 13024 48176 13028
rect 48192 13084 48256 13088
rect 48192 13028 48196 13084
rect 48196 13028 48252 13084
rect 48252 13028 48256 13084
rect 48192 13024 48256 13028
rect 2952 12540 3016 12544
rect 2952 12484 2956 12540
rect 2956 12484 3012 12540
rect 3012 12484 3016 12540
rect 2952 12480 3016 12484
rect 3032 12540 3096 12544
rect 3032 12484 3036 12540
rect 3036 12484 3092 12540
rect 3092 12484 3096 12540
rect 3032 12480 3096 12484
rect 3112 12540 3176 12544
rect 3112 12484 3116 12540
rect 3116 12484 3172 12540
rect 3172 12484 3176 12540
rect 3112 12480 3176 12484
rect 3192 12540 3256 12544
rect 3192 12484 3196 12540
rect 3196 12484 3252 12540
rect 3252 12484 3256 12540
rect 3192 12480 3256 12484
rect 12952 12540 13016 12544
rect 12952 12484 12956 12540
rect 12956 12484 13012 12540
rect 13012 12484 13016 12540
rect 12952 12480 13016 12484
rect 13032 12540 13096 12544
rect 13032 12484 13036 12540
rect 13036 12484 13092 12540
rect 13092 12484 13096 12540
rect 13032 12480 13096 12484
rect 13112 12540 13176 12544
rect 13112 12484 13116 12540
rect 13116 12484 13172 12540
rect 13172 12484 13176 12540
rect 13112 12480 13176 12484
rect 13192 12540 13256 12544
rect 13192 12484 13196 12540
rect 13196 12484 13252 12540
rect 13252 12484 13256 12540
rect 13192 12480 13256 12484
rect 22952 12540 23016 12544
rect 22952 12484 22956 12540
rect 22956 12484 23012 12540
rect 23012 12484 23016 12540
rect 22952 12480 23016 12484
rect 23032 12540 23096 12544
rect 23032 12484 23036 12540
rect 23036 12484 23092 12540
rect 23092 12484 23096 12540
rect 23032 12480 23096 12484
rect 23112 12540 23176 12544
rect 23112 12484 23116 12540
rect 23116 12484 23172 12540
rect 23172 12484 23176 12540
rect 23112 12480 23176 12484
rect 23192 12540 23256 12544
rect 23192 12484 23196 12540
rect 23196 12484 23252 12540
rect 23252 12484 23256 12540
rect 23192 12480 23256 12484
rect 32952 12540 33016 12544
rect 32952 12484 32956 12540
rect 32956 12484 33012 12540
rect 33012 12484 33016 12540
rect 32952 12480 33016 12484
rect 33032 12540 33096 12544
rect 33032 12484 33036 12540
rect 33036 12484 33092 12540
rect 33092 12484 33096 12540
rect 33032 12480 33096 12484
rect 33112 12540 33176 12544
rect 33112 12484 33116 12540
rect 33116 12484 33172 12540
rect 33172 12484 33176 12540
rect 33112 12480 33176 12484
rect 33192 12540 33256 12544
rect 33192 12484 33196 12540
rect 33196 12484 33252 12540
rect 33252 12484 33256 12540
rect 33192 12480 33256 12484
rect 42952 12540 43016 12544
rect 42952 12484 42956 12540
rect 42956 12484 43012 12540
rect 43012 12484 43016 12540
rect 42952 12480 43016 12484
rect 43032 12540 43096 12544
rect 43032 12484 43036 12540
rect 43036 12484 43092 12540
rect 43092 12484 43096 12540
rect 43032 12480 43096 12484
rect 43112 12540 43176 12544
rect 43112 12484 43116 12540
rect 43116 12484 43172 12540
rect 43172 12484 43176 12540
rect 43112 12480 43176 12484
rect 43192 12540 43256 12544
rect 43192 12484 43196 12540
rect 43196 12484 43252 12540
rect 43252 12484 43256 12540
rect 43192 12480 43256 12484
rect 7952 11996 8016 12000
rect 7952 11940 7956 11996
rect 7956 11940 8012 11996
rect 8012 11940 8016 11996
rect 7952 11936 8016 11940
rect 8032 11996 8096 12000
rect 8032 11940 8036 11996
rect 8036 11940 8092 11996
rect 8092 11940 8096 11996
rect 8032 11936 8096 11940
rect 8112 11996 8176 12000
rect 8112 11940 8116 11996
rect 8116 11940 8172 11996
rect 8172 11940 8176 11996
rect 8112 11936 8176 11940
rect 8192 11996 8256 12000
rect 8192 11940 8196 11996
rect 8196 11940 8252 11996
rect 8252 11940 8256 11996
rect 8192 11936 8256 11940
rect 17952 11996 18016 12000
rect 17952 11940 17956 11996
rect 17956 11940 18012 11996
rect 18012 11940 18016 11996
rect 17952 11936 18016 11940
rect 18032 11996 18096 12000
rect 18032 11940 18036 11996
rect 18036 11940 18092 11996
rect 18092 11940 18096 11996
rect 18032 11936 18096 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 27952 11996 28016 12000
rect 27952 11940 27956 11996
rect 27956 11940 28012 11996
rect 28012 11940 28016 11996
rect 27952 11936 28016 11940
rect 28032 11996 28096 12000
rect 28032 11940 28036 11996
rect 28036 11940 28092 11996
rect 28092 11940 28096 11996
rect 28032 11936 28096 11940
rect 28112 11996 28176 12000
rect 28112 11940 28116 11996
rect 28116 11940 28172 11996
rect 28172 11940 28176 11996
rect 28112 11936 28176 11940
rect 28192 11996 28256 12000
rect 28192 11940 28196 11996
rect 28196 11940 28252 11996
rect 28252 11940 28256 11996
rect 28192 11936 28256 11940
rect 37952 11996 38016 12000
rect 37952 11940 37956 11996
rect 37956 11940 38012 11996
rect 38012 11940 38016 11996
rect 37952 11936 38016 11940
rect 38032 11996 38096 12000
rect 38032 11940 38036 11996
rect 38036 11940 38092 11996
rect 38092 11940 38096 11996
rect 38032 11936 38096 11940
rect 38112 11996 38176 12000
rect 38112 11940 38116 11996
rect 38116 11940 38172 11996
rect 38172 11940 38176 11996
rect 38112 11936 38176 11940
rect 38192 11996 38256 12000
rect 38192 11940 38196 11996
rect 38196 11940 38252 11996
rect 38252 11940 38256 11996
rect 38192 11936 38256 11940
rect 47952 11996 48016 12000
rect 47952 11940 47956 11996
rect 47956 11940 48012 11996
rect 48012 11940 48016 11996
rect 47952 11936 48016 11940
rect 48032 11996 48096 12000
rect 48032 11940 48036 11996
rect 48036 11940 48092 11996
rect 48092 11940 48096 11996
rect 48032 11936 48096 11940
rect 48112 11996 48176 12000
rect 48112 11940 48116 11996
rect 48116 11940 48172 11996
rect 48172 11940 48176 11996
rect 48112 11936 48176 11940
rect 48192 11996 48256 12000
rect 48192 11940 48196 11996
rect 48196 11940 48252 11996
rect 48252 11940 48256 11996
rect 48192 11936 48256 11940
rect 2952 11452 3016 11456
rect 2952 11396 2956 11452
rect 2956 11396 3012 11452
rect 3012 11396 3016 11452
rect 2952 11392 3016 11396
rect 3032 11452 3096 11456
rect 3032 11396 3036 11452
rect 3036 11396 3092 11452
rect 3092 11396 3096 11452
rect 3032 11392 3096 11396
rect 3112 11452 3176 11456
rect 3112 11396 3116 11452
rect 3116 11396 3172 11452
rect 3172 11396 3176 11452
rect 3112 11392 3176 11396
rect 3192 11452 3256 11456
rect 3192 11396 3196 11452
rect 3196 11396 3252 11452
rect 3252 11396 3256 11452
rect 3192 11392 3256 11396
rect 12952 11452 13016 11456
rect 12952 11396 12956 11452
rect 12956 11396 13012 11452
rect 13012 11396 13016 11452
rect 12952 11392 13016 11396
rect 13032 11452 13096 11456
rect 13032 11396 13036 11452
rect 13036 11396 13092 11452
rect 13092 11396 13096 11452
rect 13032 11392 13096 11396
rect 13112 11452 13176 11456
rect 13112 11396 13116 11452
rect 13116 11396 13172 11452
rect 13172 11396 13176 11452
rect 13112 11392 13176 11396
rect 13192 11452 13256 11456
rect 13192 11396 13196 11452
rect 13196 11396 13252 11452
rect 13252 11396 13256 11452
rect 13192 11392 13256 11396
rect 22952 11452 23016 11456
rect 22952 11396 22956 11452
rect 22956 11396 23012 11452
rect 23012 11396 23016 11452
rect 22952 11392 23016 11396
rect 23032 11452 23096 11456
rect 23032 11396 23036 11452
rect 23036 11396 23092 11452
rect 23092 11396 23096 11452
rect 23032 11392 23096 11396
rect 23112 11452 23176 11456
rect 23112 11396 23116 11452
rect 23116 11396 23172 11452
rect 23172 11396 23176 11452
rect 23112 11392 23176 11396
rect 23192 11452 23256 11456
rect 23192 11396 23196 11452
rect 23196 11396 23252 11452
rect 23252 11396 23256 11452
rect 23192 11392 23256 11396
rect 32952 11452 33016 11456
rect 32952 11396 32956 11452
rect 32956 11396 33012 11452
rect 33012 11396 33016 11452
rect 32952 11392 33016 11396
rect 33032 11452 33096 11456
rect 33032 11396 33036 11452
rect 33036 11396 33092 11452
rect 33092 11396 33096 11452
rect 33032 11392 33096 11396
rect 33112 11452 33176 11456
rect 33112 11396 33116 11452
rect 33116 11396 33172 11452
rect 33172 11396 33176 11452
rect 33112 11392 33176 11396
rect 33192 11452 33256 11456
rect 33192 11396 33196 11452
rect 33196 11396 33252 11452
rect 33252 11396 33256 11452
rect 33192 11392 33256 11396
rect 42952 11452 43016 11456
rect 42952 11396 42956 11452
rect 42956 11396 43012 11452
rect 43012 11396 43016 11452
rect 42952 11392 43016 11396
rect 43032 11452 43096 11456
rect 43032 11396 43036 11452
rect 43036 11396 43092 11452
rect 43092 11396 43096 11452
rect 43032 11392 43096 11396
rect 43112 11452 43176 11456
rect 43112 11396 43116 11452
rect 43116 11396 43172 11452
rect 43172 11396 43176 11452
rect 43112 11392 43176 11396
rect 43192 11452 43256 11456
rect 43192 11396 43196 11452
rect 43196 11396 43252 11452
rect 43252 11396 43256 11452
rect 43192 11392 43256 11396
rect 32076 11052 32140 11116
rect 7952 10908 8016 10912
rect 7952 10852 7956 10908
rect 7956 10852 8012 10908
rect 8012 10852 8016 10908
rect 7952 10848 8016 10852
rect 8032 10908 8096 10912
rect 8032 10852 8036 10908
rect 8036 10852 8092 10908
rect 8092 10852 8096 10908
rect 8032 10848 8096 10852
rect 8112 10908 8176 10912
rect 8112 10852 8116 10908
rect 8116 10852 8172 10908
rect 8172 10852 8176 10908
rect 8112 10848 8176 10852
rect 8192 10908 8256 10912
rect 8192 10852 8196 10908
rect 8196 10852 8252 10908
rect 8252 10852 8256 10908
rect 8192 10848 8256 10852
rect 17952 10908 18016 10912
rect 17952 10852 17956 10908
rect 17956 10852 18012 10908
rect 18012 10852 18016 10908
rect 17952 10848 18016 10852
rect 18032 10908 18096 10912
rect 18032 10852 18036 10908
rect 18036 10852 18092 10908
rect 18092 10852 18096 10908
rect 18032 10848 18096 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 27952 10908 28016 10912
rect 27952 10852 27956 10908
rect 27956 10852 28012 10908
rect 28012 10852 28016 10908
rect 27952 10848 28016 10852
rect 28032 10908 28096 10912
rect 28032 10852 28036 10908
rect 28036 10852 28092 10908
rect 28092 10852 28096 10908
rect 28032 10848 28096 10852
rect 28112 10908 28176 10912
rect 28112 10852 28116 10908
rect 28116 10852 28172 10908
rect 28172 10852 28176 10908
rect 28112 10848 28176 10852
rect 28192 10908 28256 10912
rect 28192 10852 28196 10908
rect 28196 10852 28252 10908
rect 28252 10852 28256 10908
rect 28192 10848 28256 10852
rect 37952 10908 38016 10912
rect 37952 10852 37956 10908
rect 37956 10852 38012 10908
rect 38012 10852 38016 10908
rect 37952 10848 38016 10852
rect 38032 10908 38096 10912
rect 38032 10852 38036 10908
rect 38036 10852 38092 10908
rect 38092 10852 38096 10908
rect 38032 10848 38096 10852
rect 38112 10908 38176 10912
rect 38112 10852 38116 10908
rect 38116 10852 38172 10908
rect 38172 10852 38176 10908
rect 38112 10848 38176 10852
rect 38192 10908 38256 10912
rect 38192 10852 38196 10908
rect 38196 10852 38252 10908
rect 38252 10852 38256 10908
rect 38192 10848 38256 10852
rect 47952 10908 48016 10912
rect 47952 10852 47956 10908
rect 47956 10852 48012 10908
rect 48012 10852 48016 10908
rect 47952 10848 48016 10852
rect 48032 10908 48096 10912
rect 48032 10852 48036 10908
rect 48036 10852 48092 10908
rect 48092 10852 48096 10908
rect 48032 10848 48096 10852
rect 48112 10908 48176 10912
rect 48112 10852 48116 10908
rect 48116 10852 48172 10908
rect 48172 10852 48176 10908
rect 48112 10848 48176 10852
rect 48192 10908 48256 10912
rect 48192 10852 48196 10908
rect 48196 10852 48252 10908
rect 48252 10852 48256 10908
rect 48192 10848 48256 10852
rect 2952 10364 3016 10368
rect 2952 10308 2956 10364
rect 2956 10308 3012 10364
rect 3012 10308 3016 10364
rect 2952 10304 3016 10308
rect 3032 10364 3096 10368
rect 3032 10308 3036 10364
rect 3036 10308 3092 10364
rect 3092 10308 3096 10364
rect 3032 10304 3096 10308
rect 3112 10364 3176 10368
rect 3112 10308 3116 10364
rect 3116 10308 3172 10364
rect 3172 10308 3176 10364
rect 3112 10304 3176 10308
rect 3192 10364 3256 10368
rect 3192 10308 3196 10364
rect 3196 10308 3252 10364
rect 3252 10308 3256 10364
rect 3192 10304 3256 10308
rect 12952 10364 13016 10368
rect 12952 10308 12956 10364
rect 12956 10308 13012 10364
rect 13012 10308 13016 10364
rect 12952 10304 13016 10308
rect 13032 10364 13096 10368
rect 13032 10308 13036 10364
rect 13036 10308 13092 10364
rect 13092 10308 13096 10364
rect 13032 10304 13096 10308
rect 13112 10364 13176 10368
rect 13112 10308 13116 10364
rect 13116 10308 13172 10364
rect 13172 10308 13176 10364
rect 13112 10304 13176 10308
rect 13192 10364 13256 10368
rect 13192 10308 13196 10364
rect 13196 10308 13252 10364
rect 13252 10308 13256 10364
rect 13192 10304 13256 10308
rect 22952 10364 23016 10368
rect 22952 10308 22956 10364
rect 22956 10308 23012 10364
rect 23012 10308 23016 10364
rect 22952 10304 23016 10308
rect 23032 10364 23096 10368
rect 23032 10308 23036 10364
rect 23036 10308 23092 10364
rect 23092 10308 23096 10364
rect 23032 10304 23096 10308
rect 23112 10364 23176 10368
rect 23112 10308 23116 10364
rect 23116 10308 23172 10364
rect 23172 10308 23176 10364
rect 23112 10304 23176 10308
rect 23192 10364 23256 10368
rect 23192 10308 23196 10364
rect 23196 10308 23252 10364
rect 23252 10308 23256 10364
rect 23192 10304 23256 10308
rect 32952 10364 33016 10368
rect 32952 10308 32956 10364
rect 32956 10308 33012 10364
rect 33012 10308 33016 10364
rect 32952 10304 33016 10308
rect 33032 10364 33096 10368
rect 33032 10308 33036 10364
rect 33036 10308 33092 10364
rect 33092 10308 33096 10364
rect 33032 10304 33096 10308
rect 33112 10364 33176 10368
rect 33112 10308 33116 10364
rect 33116 10308 33172 10364
rect 33172 10308 33176 10364
rect 33112 10304 33176 10308
rect 33192 10364 33256 10368
rect 33192 10308 33196 10364
rect 33196 10308 33252 10364
rect 33252 10308 33256 10364
rect 33192 10304 33256 10308
rect 42952 10364 43016 10368
rect 42952 10308 42956 10364
rect 42956 10308 43012 10364
rect 43012 10308 43016 10364
rect 42952 10304 43016 10308
rect 43032 10364 43096 10368
rect 43032 10308 43036 10364
rect 43036 10308 43092 10364
rect 43092 10308 43096 10364
rect 43032 10304 43096 10308
rect 43112 10364 43176 10368
rect 43112 10308 43116 10364
rect 43116 10308 43172 10364
rect 43172 10308 43176 10364
rect 43112 10304 43176 10308
rect 43192 10364 43256 10368
rect 43192 10308 43196 10364
rect 43196 10308 43252 10364
rect 43252 10308 43256 10364
rect 43192 10304 43256 10308
rect 7952 9820 8016 9824
rect 7952 9764 7956 9820
rect 7956 9764 8012 9820
rect 8012 9764 8016 9820
rect 7952 9760 8016 9764
rect 8032 9820 8096 9824
rect 8032 9764 8036 9820
rect 8036 9764 8092 9820
rect 8092 9764 8096 9820
rect 8032 9760 8096 9764
rect 8112 9820 8176 9824
rect 8112 9764 8116 9820
rect 8116 9764 8172 9820
rect 8172 9764 8176 9820
rect 8112 9760 8176 9764
rect 8192 9820 8256 9824
rect 8192 9764 8196 9820
rect 8196 9764 8252 9820
rect 8252 9764 8256 9820
rect 8192 9760 8256 9764
rect 17952 9820 18016 9824
rect 17952 9764 17956 9820
rect 17956 9764 18012 9820
rect 18012 9764 18016 9820
rect 17952 9760 18016 9764
rect 18032 9820 18096 9824
rect 18032 9764 18036 9820
rect 18036 9764 18092 9820
rect 18092 9764 18096 9820
rect 18032 9760 18096 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 27952 9820 28016 9824
rect 27952 9764 27956 9820
rect 27956 9764 28012 9820
rect 28012 9764 28016 9820
rect 27952 9760 28016 9764
rect 28032 9820 28096 9824
rect 28032 9764 28036 9820
rect 28036 9764 28092 9820
rect 28092 9764 28096 9820
rect 28032 9760 28096 9764
rect 28112 9820 28176 9824
rect 28112 9764 28116 9820
rect 28116 9764 28172 9820
rect 28172 9764 28176 9820
rect 28112 9760 28176 9764
rect 28192 9820 28256 9824
rect 28192 9764 28196 9820
rect 28196 9764 28252 9820
rect 28252 9764 28256 9820
rect 28192 9760 28256 9764
rect 37952 9820 38016 9824
rect 37952 9764 37956 9820
rect 37956 9764 38012 9820
rect 38012 9764 38016 9820
rect 37952 9760 38016 9764
rect 38032 9820 38096 9824
rect 38032 9764 38036 9820
rect 38036 9764 38092 9820
rect 38092 9764 38096 9820
rect 38032 9760 38096 9764
rect 38112 9820 38176 9824
rect 38112 9764 38116 9820
rect 38116 9764 38172 9820
rect 38172 9764 38176 9820
rect 38112 9760 38176 9764
rect 38192 9820 38256 9824
rect 38192 9764 38196 9820
rect 38196 9764 38252 9820
rect 38252 9764 38256 9820
rect 38192 9760 38256 9764
rect 47952 9820 48016 9824
rect 47952 9764 47956 9820
rect 47956 9764 48012 9820
rect 48012 9764 48016 9820
rect 47952 9760 48016 9764
rect 48032 9820 48096 9824
rect 48032 9764 48036 9820
rect 48036 9764 48092 9820
rect 48092 9764 48096 9820
rect 48032 9760 48096 9764
rect 48112 9820 48176 9824
rect 48112 9764 48116 9820
rect 48116 9764 48172 9820
rect 48172 9764 48176 9820
rect 48112 9760 48176 9764
rect 48192 9820 48256 9824
rect 48192 9764 48196 9820
rect 48196 9764 48252 9820
rect 48252 9764 48256 9820
rect 48192 9760 48256 9764
rect 15700 9556 15764 9620
rect 2952 9276 3016 9280
rect 2952 9220 2956 9276
rect 2956 9220 3012 9276
rect 3012 9220 3016 9276
rect 2952 9216 3016 9220
rect 3032 9276 3096 9280
rect 3032 9220 3036 9276
rect 3036 9220 3092 9276
rect 3092 9220 3096 9276
rect 3032 9216 3096 9220
rect 3112 9276 3176 9280
rect 3112 9220 3116 9276
rect 3116 9220 3172 9276
rect 3172 9220 3176 9276
rect 3112 9216 3176 9220
rect 3192 9276 3256 9280
rect 3192 9220 3196 9276
rect 3196 9220 3252 9276
rect 3252 9220 3256 9276
rect 3192 9216 3256 9220
rect 12952 9276 13016 9280
rect 12952 9220 12956 9276
rect 12956 9220 13012 9276
rect 13012 9220 13016 9276
rect 12952 9216 13016 9220
rect 13032 9276 13096 9280
rect 13032 9220 13036 9276
rect 13036 9220 13092 9276
rect 13092 9220 13096 9276
rect 13032 9216 13096 9220
rect 13112 9276 13176 9280
rect 13112 9220 13116 9276
rect 13116 9220 13172 9276
rect 13172 9220 13176 9276
rect 13112 9216 13176 9220
rect 13192 9276 13256 9280
rect 13192 9220 13196 9276
rect 13196 9220 13252 9276
rect 13252 9220 13256 9276
rect 13192 9216 13256 9220
rect 22952 9276 23016 9280
rect 22952 9220 22956 9276
rect 22956 9220 23012 9276
rect 23012 9220 23016 9276
rect 22952 9216 23016 9220
rect 23032 9276 23096 9280
rect 23032 9220 23036 9276
rect 23036 9220 23092 9276
rect 23092 9220 23096 9276
rect 23032 9216 23096 9220
rect 23112 9276 23176 9280
rect 23112 9220 23116 9276
rect 23116 9220 23172 9276
rect 23172 9220 23176 9276
rect 23112 9216 23176 9220
rect 23192 9276 23256 9280
rect 23192 9220 23196 9276
rect 23196 9220 23252 9276
rect 23252 9220 23256 9276
rect 23192 9216 23256 9220
rect 32952 9276 33016 9280
rect 32952 9220 32956 9276
rect 32956 9220 33012 9276
rect 33012 9220 33016 9276
rect 32952 9216 33016 9220
rect 33032 9276 33096 9280
rect 33032 9220 33036 9276
rect 33036 9220 33092 9276
rect 33092 9220 33096 9276
rect 33032 9216 33096 9220
rect 33112 9276 33176 9280
rect 33112 9220 33116 9276
rect 33116 9220 33172 9276
rect 33172 9220 33176 9276
rect 33112 9216 33176 9220
rect 33192 9276 33256 9280
rect 33192 9220 33196 9276
rect 33196 9220 33252 9276
rect 33252 9220 33256 9276
rect 33192 9216 33256 9220
rect 42952 9276 43016 9280
rect 42952 9220 42956 9276
rect 42956 9220 43012 9276
rect 43012 9220 43016 9276
rect 42952 9216 43016 9220
rect 43032 9276 43096 9280
rect 43032 9220 43036 9276
rect 43036 9220 43092 9276
rect 43092 9220 43096 9276
rect 43032 9216 43096 9220
rect 43112 9276 43176 9280
rect 43112 9220 43116 9276
rect 43116 9220 43172 9276
rect 43172 9220 43176 9276
rect 43112 9216 43176 9220
rect 43192 9276 43256 9280
rect 43192 9220 43196 9276
rect 43196 9220 43252 9276
rect 43252 9220 43256 9276
rect 43192 9216 43256 9220
rect 7952 8732 8016 8736
rect 7952 8676 7956 8732
rect 7956 8676 8012 8732
rect 8012 8676 8016 8732
rect 7952 8672 8016 8676
rect 8032 8732 8096 8736
rect 8032 8676 8036 8732
rect 8036 8676 8092 8732
rect 8092 8676 8096 8732
rect 8032 8672 8096 8676
rect 8112 8732 8176 8736
rect 8112 8676 8116 8732
rect 8116 8676 8172 8732
rect 8172 8676 8176 8732
rect 8112 8672 8176 8676
rect 8192 8732 8256 8736
rect 8192 8676 8196 8732
rect 8196 8676 8252 8732
rect 8252 8676 8256 8732
rect 8192 8672 8256 8676
rect 17952 8732 18016 8736
rect 17952 8676 17956 8732
rect 17956 8676 18012 8732
rect 18012 8676 18016 8732
rect 17952 8672 18016 8676
rect 18032 8732 18096 8736
rect 18032 8676 18036 8732
rect 18036 8676 18092 8732
rect 18092 8676 18096 8732
rect 18032 8672 18096 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 27952 8732 28016 8736
rect 27952 8676 27956 8732
rect 27956 8676 28012 8732
rect 28012 8676 28016 8732
rect 27952 8672 28016 8676
rect 28032 8732 28096 8736
rect 28032 8676 28036 8732
rect 28036 8676 28092 8732
rect 28092 8676 28096 8732
rect 28032 8672 28096 8676
rect 28112 8732 28176 8736
rect 28112 8676 28116 8732
rect 28116 8676 28172 8732
rect 28172 8676 28176 8732
rect 28112 8672 28176 8676
rect 28192 8732 28256 8736
rect 28192 8676 28196 8732
rect 28196 8676 28252 8732
rect 28252 8676 28256 8732
rect 28192 8672 28256 8676
rect 37952 8732 38016 8736
rect 37952 8676 37956 8732
rect 37956 8676 38012 8732
rect 38012 8676 38016 8732
rect 37952 8672 38016 8676
rect 38032 8732 38096 8736
rect 38032 8676 38036 8732
rect 38036 8676 38092 8732
rect 38092 8676 38096 8732
rect 38032 8672 38096 8676
rect 38112 8732 38176 8736
rect 38112 8676 38116 8732
rect 38116 8676 38172 8732
rect 38172 8676 38176 8732
rect 38112 8672 38176 8676
rect 38192 8732 38256 8736
rect 38192 8676 38196 8732
rect 38196 8676 38252 8732
rect 38252 8676 38256 8732
rect 38192 8672 38256 8676
rect 47952 8732 48016 8736
rect 47952 8676 47956 8732
rect 47956 8676 48012 8732
rect 48012 8676 48016 8732
rect 47952 8672 48016 8676
rect 48032 8732 48096 8736
rect 48032 8676 48036 8732
rect 48036 8676 48092 8732
rect 48092 8676 48096 8732
rect 48032 8672 48096 8676
rect 48112 8732 48176 8736
rect 48112 8676 48116 8732
rect 48116 8676 48172 8732
rect 48172 8676 48176 8732
rect 48112 8672 48176 8676
rect 48192 8732 48256 8736
rect 48192 8676 48196 8732
rect 48196 8676 48252 8732
rect 48252 8676 48256 8732
rect 48192 8672 48256 8676
rect 2952 8188 3016 8192
rect 2952 8132 2956 8188
rect 2956 8132 3012 8188
rect 3012 8132 3016 8188
rect 2952 8128 3016 8132
rect 3032 8188 3096 8192
rect 3032 8132 3036 8188
rect 3036 8132 3092 8188
rect 3092 8132 3096 8188
rect 3032 8128 3096 8132
rect 3112 8188 3176 8192
rect 3112 8132 3116 8188
rect 3116 8132 3172 8188
rect 3172 8132 3176 8188
rect 3112 8128 3176 8132
rect 3192 8188 3256 8192
rect 3192 8132 3196 8188
rect 3196 8132 3252 8188
rect 3252 8132 3256 8188
rect 3192 8128 3256 8132
rect 12952 8188 13016 8192
rect 12952 8132 12956 8188
rect 12956 8132 13012 8188
rect 13012 8132 13016 8188
rect 12952 8128 13016 8132
rect 13032 8188 13096 8192
rect 13032 8132 13036 8188
rect 13036 8132 13092 8188
rect 13092 8132 13096 8188
rect 13032 8128 13096 8132
rect 13112 8188 13176 8192
rect 13112 8132 13116 8188
rect 13116 8132 13172 8188
rect 13172 8132 13176 8188
rect 13112 8128 13176 8132
rect 13192 8188 13256 8192
rect 13192 8132 13196 8188
rect 13196 8132 13252 8188
rect 13252 8132 13256 8188
rect 13192 8128 13256 8132
rect 22952 8188 23016 8192
rect 22952 8132 22956 8188
rect 22956 8132 23012 8188
rect 23012 8132 23016 8188
rect 22952 8128 23016 8132
rect 23032 8188 23096 8192
rect 23032 8132 23036 8188
rect 23036 8132 23092 8188
rect 23092 8132 23096 8188
rect 23032 8128 23096 8132
rect 23112 8188 23176 8192
rect 23112 8132 23116 8188
rect 23116 8132 23172 8188
rect 23172 8132 23176 8188
rect 23112 8128 23176 8132
rect 23192 8188 23256 8192
rect 23192 8132 23196 8188
rect 23196 8132 23252 8188
rect 23252 8132 23256 8188
rect 23192 8128 23256 8132
rect 32952 8188 33016 8192
rect 32952 8132 32956 8188
rect 32956 8132 33012 8188
rect 33012 8132 33016 8188
rect 32952 8128 33016 8132
rect 33032 8188 33096 8192
rect 33032 8132 33036 8188
rect 33036 8132 33092 8188
rect 33092 8132 33096 8188
rect 33032 8128 33096 8132
rect 33112 8188 33176 8192
rect 33112 8132 33116 8188
rect 33116 8132 33172 8188
rect 33172 8132 33176 8188
rect 33112 8128 33176 8132
rect 33192 8188 33256 8192
rect 33192 8132 33196 8188
rect 33196 8132 33252 8188
rect 33252 8132 33256 8188
rect 33192 8128 33256 8132
rect 42952 8188 43016 8192
rect 42952 8132 42956 8188
rect 42956 8132 43012 8188
rect 43012 8132 43016 8188
rect 42952 8128 43016 8132
rect 43032 8188 43096 8192
rect 43032 8132 43036 8188
rect 43036 8132 43092 8188
rect 43092 8132 43096 8188
rect 43032 8128 43096 8132
rect 43112 8188 43176 8192
rect 43112 8132 43116 8188
rect 43116 8132 43172 8188
rect 43172 8132 43176 8188
rect 43112 8128 43176 8132
rect 43192 8188 43256 8192
rect 43192 8132 43196 8188
rect 43196 8132 43252 8188
rect 43252 8132 43256 8188
rect 43192 8128 43256 8132
rect 7952 7644 8016 7648
rect 7952 7588 7956 7644
rect 7956 7588 8012 7644
rect 8012 7588 8016 7644
rect 7952 7584 8016 7588
rect 8032 7644 8096 7648
rect 8032 7588 8036 7644
rect 8036 7588 8092 7644
rect 8092 7588 8096 7644
rect 8032 7584 8096 7588
rect 8112 7644 8176 7648
rect 8112 7588 8116 7644
rect 8116 7588 8172 7644
rect 8172 7588 8176 7644
rect 8112 7584 8176 7588
rect 8192 7644 8256 7648
rect 8192 7588 8196 7644
rect 8196 7588 8252 7644
rect 8252 7588 8256 7644
rect 8192 7584 8256 7588
rect 17952 7644 18016 7648
rect 17952 7588 17956 7644
rect 17956 7588 18012 7644
rect 18012 7588 18016 7644
rect 17952 7584 18016 7588
rect 18032 7644 18096 7648
rect 18032 7588 18036 7644
rect 18036 7588 18092 7644
rect 18092 7588 18096 7644
rect 18032 7584 18096 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 27952 7644 28016 7648
rect 27952 7588 27956 7644
rect 27956 7588 28012 7644
rect 28012 7588 28016 7644
rect 27952 7584 28016 7588
rect 28032 7644 28096 7648
rect 28032 7588 28036 7644
rect 28036 7588 28092 7644
rect 28092 7588 28096 7644
rect 28032 7584 28096 7588
rect 28112 7644 28176 7648
rect 28112 7588 28116 7644
rect 28116 7588 28172 7644
rect 28172 7588 28176 7644
rect 28112 7584 28176 7588
rect 28192 7644 28256 7648
rect 28192 7588 28196 7644
rect 28196 7588 28252 7644
rect 28252 7588 28256 7644
rect 28192 7584 28256 7588
rect 37952 7644 38016 7648
rect 37952 7588 37956 7644
rect 37956 7588 38012 7644
rect 38012 7588 38016 7644
rect 37952 7584 38016 7588
rect 38032 7644 38096 7648
rect 38032 7588 38036 7644
rect 38036 7588 38092 7644
rect 38092 7588 38096 7644
rect 38032 7584 38096 7588
rect 38112 7644 38176 7648
rect 38112 7588 38116 7644
rect 38116 7588 38172 7644
rect 38172 7588 38176 7644
rect 38112 7584 38176 7588
rect 38192 7644 38256 7648
rect 38192 7588 38196 7644
rect 38196 7588 38252 7644
rect 38252 7588 38256 7644
rect 38192 7584 38256 7588
rect 47952 7644 48016 7648
rect 47952 7588 47956 7644
rect 47956 7588 48012 7644
rect 48012 7588 48016 7644
rect 47952 7584 48016 7588
rect 48032 7644 48096 7648
rect 48032 7588 48036 7644
rect 48036 7588 48092 7644
rect 48092 7588 48096 7644
rect 48032 7584 48096 7588
rect 48112 7644 48176 7648
rect 48112 7588 48116 7644
rect 48116 7588 48172 7644
rect 48172 7588 48176 7644
rect 48112 7584 48176 7588
rect 48192 7644 48256 7648
rect 48192 7588 48196 7644
rect 48196 7588 48252 7644
rect 48252 7588 48256 7644
rect 48192 7584 48256 7588
rect 2952 7100 3016 7104
rect 2952 7044 2956 7100
rect 2956 7044 3012 7100
rect 3012 7044 3016 7100
rect 2952 7040 3016 7044
rect 3032 7100 3096 7104
rect 3032 7044 3036 7100
rect 3036 7044 3092 7100
rect 3092 7044 3096 7100
rect 3032 7040 3096 7044
rect 3112 7100 3176 7104
rect 3112 7044 3116 7100
rect 3116 7044 3172 7100
rect 3172 7044 3176 7100
rect 3112 7040 3176 7044
rect 3192 7100 3256 7104
rect 3192 7044 3196 7100
rect 3196 7044 3252 7100
rect 3252 7044 3256 7100
rect 3192 7040 3256 7044
rect 12952 7100 13016 7104
rect 12952 7044 12956 7100
rect 12956 7044 13012 7100
rect 13012 7044 13016 7100
rect 12952 7040 13016 7044
rect 13032 7100 13096 7104
rect 13032 7044 13036 7100
rect 13036 7044 13092 7100
rect 13092 7044 13096 7100
rect 13032 7040 13096 7044
rect 13112 7100 13176 7104
rect 13112 7044 13116 7100
rect 13116 7044 13172 7100
rect 13172 7044 13176 7100
rect 13112 7040 13176 7044
rect 13192 7100 13256 7104
rect 13192 7044 13196 7100
rect 13196 7044 13252 7100
rect 13252 7044 13256 7100
rect 13192 7040 13256 7044
rect 22952 7100 23016 7104
rect 22952 7044 22956 7100
rect 22956 7044 23012 7100
rect 23012 7044 23016 7100
rect 22952 7040 23016 7044
rect 23032 7100 23096 7104
rect 23032 7044 23036 7100
rect 23036 7044 23092 7100
rect 23092 7044 23096 7100
rect 23032 7040 23096 7044
rect 23112 7100 23176 7104
rect 23112 7044 23116 7100
rect 23116 7044 23172 7100
rect 23172 7044 23176 7100
rect 23112 7040 23176 7044
rect 23192 7100 23256 7104
rect 23192 7044 23196 7100
rect 23196 7044 23252 7100
rect 23252 7044 23256 7100
rect 23192 7040 23256 7044
rect 32952 7100 33016 7104
rect 32952 7044 32956 7100
rect 32956 7044 33012 7100
rect 33012 7044 33016 7100
rect 32952 7040 33016 7044
rect 33032 7100 33096 7104
rect 33032 7044 33036 7100
rect 33036 7044 33092 7100
rect 33092 7044 33096 7100
rect 33032 7040 33096 7044
rect 33112 7100 33176 7104
rect 33112 7044 33116 7100
rect 33116 7044 33172 7100
rect 33172 7044 33176 7100
rect 33112 7040 33176 7044
rect 33192 7100 33256 7104
rect 33192 7044 33196 7100
rect 33196 7044 33252 7100
rect 33252 7044 33256 7100
rect 33192 7040 33256 7044
rect 42952 7100 43016 7104
rect 42952 7044 42956 7100
rect 42956 7044 43012 7100
rect 43012 7044 43016 7100
rect 42952 7040 43016 7044
rect 43032 7100 43096 7104
rect 43032 7044 43036 7100
rect 43036 7044 43092 7100
rect 43092 7044 43096 7100
rect 43032 7040 43096 7044
rect 43112 7100 43176 7104
rect 43112 7044 43116 7100
rect 43116 7044 43172 7100
rect 43172 7044 43176 7100
rect 43112 7040 43176 7044
rect 43192 7100 43256 7104
rect 43192 7044 43196 7100
rect 43196 7044 43252 7100
rect 43252 7044 43256 7100
rect 43192 7040 43256 7044
rect 7952 6556 8016 6560
rect 7952 6500 7956 6556
rect 7956 6500 8012 6556
rect 8012 6500 8016 6556
rect 7952 6496 8016 6500
rect 8032 6556 8096 6560
rect 8032 6500 8036 6556
rect 8036 6500 8092 6556
rect 8092 6500 8096 6556
rect 8032 6496 8096 6500
rect 8112 6556 8176 6560
rect 8112 6500 8116 6556
rect 8116 6500 8172 6556
rect 8172 6500 8176 6556
rect 8112 6496 8176 6500
rect 8192 6556 8256 6560
rect 8192 6500 8196 6556
rect 8196 6500 8252 6556
rect 8252 6500 8256 6556
rect 8192 6496 8256 6500
rect 17952 6556 18016 6560
rect 17952 6500 17956 6556
rect 17956 6500 18012 6556
rect 18012 6500 18016 6556
rect 17952 6496 18016 6500
rect 18032 6556 18096 6560
rect 18032 6500 18036 6556
rect 18036 6500 18092 6556
rect 18092 6500 18096 6556
rect 18032 6496 18096 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 27952 6556 28016 6560
rect 27952 6500 27956 6556
rect 27956 6500 28012 6556
rect 28012 6500 28016 6556
rect 27952 6496 28016 6500
rect 28032 6556 28096 6560
rect 28032 6500 28036 6556
rect 28036 6500 28092 6556
rect 28092 6500 28096 6556
rect 28032 6496 28096 6500
rect 28112 6556 28176 6560
rect 28112 6500 28116 6556
rect 28116 6500 28172 6556
rect 28172 6500 28176 6556
rect 28112 6496 28176 6500
rect 28192 6556 28256 6560
rect 28192 6500 28196 6556
rect 28196 6500 28252 6556
rect 28252 6500 28256 6556
rect 28192 6496 28256 6500
rect 37952 6556 38016 6560
rect 37952 6500 37956 6556
rect 37956 6500 38012 6556
rect 38012 6500 38016 6556
rect 37952 6496 38016 6500
rect 38032 6556 38096 6560
rect 38032 6500 38036 6556
rect 38036 6500 38092 6556
rect 38092 6500 38096 6556
rect 38032 6496 38096 6500
rect 38112 6556 38176 6560
rect 38112 6500 38116 6556
rect 38116 6500 38172 6556
rect 38172 6500 38176 6556
rect 38112 6496 38176 6500
rect 38192 6556 38256 6560
rect 38192 6500 38196 6556
rect 38196 6500 38252 6556
rect 38252 6500 38256 6556
rect 38192 6496 38256 6500
rect 47952 6556 48016 6560
rect 47952 6500 47956 6556
rect 47956 6500 48012 6556
rect 48012 6500 48016 6556
rect 47952 6496 48016 6500
rect 48032 6556 48096 6560
rect 48032 6500 48036 6556
rect 48036 6500 48092 6556
rect 48092 6500 48096 6556
rect 48032 6496 48096 6500
rect 48112 6556 48176 6560
rect 48112 6500 48116 6556
rect 48116 6500 48172 6556
rect 48172 6500 48176 6556
rect 48112 6496 48176 6500
rect 48192 6556 48256 6560
rect 48192 6500 48196 6556
rect 48196 6500 48252 6556
rect 48252 6500 48256 6556
rect 48192 6496 48256 6500
rect 2952 6012 3016 6016
rect 2952 5956 2956 6012
rect 2956 5956 3012 6012
rect 3012 5956 3016 6012
rect 2952 5952 3016 5956
rect 3032 6012 3096 6016
rect 3032 5956 3036 6012
rect 3036 5956 3092 6012
rect 3092 5956 3096 6012
rect 3032 5952 3096 5956
rect 3112 6012 3176 6016
rect 3112 5956 3116 6012
rect 3116 5956 3172 6012
rect 3172 5956 3176 6012
rect 3112 5952 3176 5956
rect 3192 6012 3256 6016
rect 3192 5956 3196 6012
rect 3196 5956 3252 6012
rect 3252 5956 3256 6012
rect 3192 5952 3256 5956
rect 12952 6012 13016 6016
rect 12952 5956 12956 6012
rect 12956 5956 13012 6012
rect 13012 5956 13016 6012
rect 12952 5952 13016 5956
rect 13032 6012 13096 6016
rect 13032 5956 13036 6012
rect 13036 5956 13092 6012
rect 13092 5956 13096 6012
rect 13032 5952 13096 5956
rect 13112 6012 13176 6016
rect 13112 5956 13116 6012
rect 13116 5956 13172 6012
rect 13172 5956 13176 6012
rect 13112 5952 13176 5956
rect 13192 6012 13256 6016
rect 13192 5956 13196 6012
rect 13196 5956 13252 6012
rect 13252 5956 13256 6012
rect 13192 5952 13256 5956
rect 22952 6012 23016 6016
rect 22952 5956 22956 6012
rect 22956 5956 23012 6012
rect 23012 5956 23016 6012
rect 22952 5952 23016 5956
rect 23032 6012 23096 6016
rect 23032 5956 23036 6012
rect 23036 5956 23092 6012
rect 23092 5956 23096 6012
rect 23032 5952 23096 5956
rect 23112 6012 23176 6016
rect 23112 5956 23116 6012
rect 23116 5956 23172 6012
rect 23172 5956 23176 6012
rect 23112 5952 23176 5956
rect 23192 6012 23256 6016
rect 23192 5956 23196 6012
rect 23196 5956 23252 6012
rect 23252 5956 23256 6012
rect 23192 5952 23256 5956
rect 32952 6012 33016 6016
rect 32952 5956 32956 6012
rect 32956 5956 33012 6012
rect 33012 5956 33016 6012
rect 32952 5952 33016 5956
rect 33032 6012 33096 6016
rect 33032 5956 33036 6012
rect 33036 5956 33092 6012
rect 33092 5956 33096 6012
rect 33032 5952 33096 5956
rect 33112 6012 33176 6016
rect 33112 5956 33116 6012
rect 33116 5956 33172 6012
rect 33172 5956 33176 6012
rect 33112 5952 33176 5956
rect 33192 6012 33256 6016
rect 33192 5956 33196 6012
rect 33196 5956 33252 6012
rect 33252 5956 33256 6012
rect 33192 5952 33256 5956
rect 42952 6012 43016 6016
rect 42952 5956 42956 6012
rect 42956 5956 43012 6012
rect 43012 5956 43016 6012
rect 42952 5952 43016 5956
rect 43032 6012 43096 6016
rect 43032 5956 43036 6012
rect 43036 5956 43092 6012
rect 43092 5956 43096 6012
rect 43032 5952 43096 5956
rect 43112 6012 43176 6016
rect 43112 5956 43116 6012
rect 43116 5956 43172 6012
rect 43172 5956 43176 6012
rect 43112 5952 43176 5956
rect 43192 6012 43256 6016
rect 43192 5956 43196 6012
rect 43196 5956 43252 6012
rect 43252 5956 43256 6012
rect 43192 5952 43256 5956
rect 7952 5468 8016 5472
rect 7952 5412 7956 5468
rect 7956 5412 8012 5468
rect 8012 5412 8016 5468
rect 7952 5408 8016 5412
rect 8032 5468 8096 5472
rect 8032 5412 8036 5468
rect 8036 5412 8092 5468
rect 8092 5412 8096 5468
rect 8032 5408 8096 5412
rect 8112 5468 8176 5472
rect 8112 5412 8116 5468
rect 8116 5412 8172 5468
rect 8172 5412 8176 5468
rect 8112 5408 8176 5412
rect 8192 5468 8256 5472
rect 8192 5412 8196 5468
rect 8196 5412 8252 5468
rect 8252 5412 8256 5468
rect 8192 5408 8256 5412
rect 17952 5468 18016 5472
rect 17952 5412 17956 5468
rect 17956 5412 18012 5468
rect 18012 5412 18016 5468
rect 17952 5408 18016 5412
rect 18032 5468 18096 5472
rect 18032 5412 18036 5468
rect 18036 5412 18092 5468
rect 18092 5412 18096 5468
rect 18032 5408 18096 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 27952 5468 28016 5472
rect 27952 5412 27956 5468
rect 27956 5412 28012 5468
rect 28012 5412 28016 5468
rect 27952 5408 28016 5412
rect 28032 5468 28096 5472
rect 28032 5412 28036 5468
rect 28036 5412 28092 5468
rect 28092 5412 28096 5468
rect 28032 5408 28096 5412
rect 28112 5468 28176 5472
rect 28112 5412 28116 5468
rect 28116 5412 28172 5468
rect 28172 5412 28176 5468
rect 28112 5408 28176 5412
rect 28192 5468 28256 5472
rect 28192 5412 28196 5468
rect 28196 5412 28252 5468
rect 28252 5412 28256 5468
rect 28192 5408 28256 5412
rect 37952 5468 38016 5472
rect 37952 5412 37956 5468
rect 37956 5412 38012 5468
rect 38012 5412 38016 5468
rect 37952 5408 38016 5412
rect 38032 5468 38096 5472
rect 38032 5412 38036 5468
rect 38036 5412 38092 5468
rect 38092 5412 38096 5468
rect 38032 5408 38096 5412
rect 38112 5468 38176 5472
rect 38112 5412 38116 5468
rect 38116 5412 38172 5468
rect 38172 5412 38176 5468
rect 38112 5408 38176 5412
rect 38192 5468 38256 5472
rect 38192 5412 38196 5468
rect 38196 5412 38252 5468
rect 38252 5412 38256 5468
rect 38192 5408 38256 5412
rect 47952 5468 48016 5472
rect 47952 5412 47956 5468
rect 47956 5412 48012 5468
rect 48012 5412 48016 5468
rect 47952 5408 48016 5412
rect 48032 5468 48096 5472
rect 48032 5412 48036 5468
rect 48036 5412 48092 5468
rect 48092 5412 48096 5468
rect 48032 5408 48096 5412
rect 48112 5468 48176 5472
rect 48112 5412 48116 5468
rect 48116 5412 48172 5468
rect 48172 5412 48176 5468
rect 48112 5408 48176 5412
rect 48192 5468 48256 5472
rect 48192 5412 48196 5468
rect 48196 5412 48252 5468
rect 48252 5412 48256 5468
rect 48192 5408 48256 5412
rect 2952 4924 3016 4928
rect 2952 4868 2956 4924
rect 2956 4868 3012 4924
rect 3012 4868 3016 4924
rect 2952 4864 3016 4868
rect 3032 4924 3096 4928
rect 3032 4868 3036 4924
rect 3036 4868 3092 4924
rect 3092 4868 3096 4924
rect 3032 4864 3096 4868
rect 3112 4924 3176 4928
rect 3112 4868 3116 4924
rect 3116 4868 3172 4924
rect 3172 4868 3176 4924
rect 3112 4864 3176 4868
rect 3192 4924 3256 4928
rect 3192 4868 3196 4924
rect 3196 4868 3252 4924
rect 3252 4868 3256 4924
rect 3192 4864 3256 4868
rect 12952 4924 13016 4928
rect 12952 4868 12956 4924
rect 12956 4868 13012 4924
rect 13012 4868 13016 4924
rect 12952 4864 13016 4868
rect 13032 4924 13096 4928
rect 13032 4868 13036 4924
rect 13036 4868 13092 4924
rect 13092 4868 13096 4924
rect 13032 4864 13096 4868
rect 13112 4924 13176 4928
rect 13112 4868 13116 4924
rect 13116 4868 13172 4924
rect 13172 4868 13176 4924
rect 13112 4864 13176 4868
rect 13192 4924 13256 4928
rect 13192 4868 13196 4924
rect 13196 4868 13252 4924
rect 13252 4868 13256 4924
rect 13192 4864 13256 4868
rect 22952 4924 23016 4928
rect 22952 4868 22956 4924
rect 22956 4868 23012 4924
rect 23012 4868 23016 4924
rect 22952 4864 23016 4868
rect 23032 4924 23096 4928
rect 23032 4868 23036 4924
rect 23036 4868 23092 4924
rect 23092 4868 23096 4924
rect 23032 4864 23096 4868
rect 23112 4924 23176 4928
rect 23112 4868 23116 4924
rect 23116 4868 23172 4924
rect 23172 4868 23176 4924
rect 23112 4864 23176 4868
rect 23192 4924 23256 4928
rect 23192 4868 23196 4924
rect 23196 4868 23252 4924
rect 23252 4868 23256 4924
rect 23192 4864 23256 4868
rect 32952 4924 33016 4928
rect 32952 4868 32956 4924
rect 32956 4868 33012 4924
rect 33012 4868 33016 4924
rect 32952 4864 33016 4868
rect 33032 4924 33096 4928
rect 33032 4868 33036 4924
rect 33036 4868 33092 4924
rect 33092 4868 33096 4924
rect 33032 4864 33096 4868
rect 33112 4924 33176 4928
rect 33112 4868 33116 4924
rect 33116 4868 33172 4924
rect 33172 4868 33176 4924
rect 33112 4864 33176 4868
rect 33192 4924 33256 4928
rect 33192 4868 33196 4924
rect 33196 4868 33252 4924
rect 33252 4868 33256 4924
rect 33192 4864 33256 4868
rect 42952 4924 43016 4928
rect 42952 4868 42956 4924
rect 42956 4868 43012 4924
rect 43012 4868 43016 4924
rect 42952 4864 43016 4868
rect 43032 4924 43096 4928
rect 43032 4868 43036 4924
rect 43036 4868 43092 4924
rect 43092 4868 43096 4924
rect 43032 4864 43096 4868
rect 43112 4924 43176 4928
rect 43112 4868 43116 4924
rect 43116 4868 43172 4924
rect 43172 4868 43176 4924
rect 43112 4864 43176 4868
rect 43192 4924 43256 4928
rect 43192 4868 43196 4924
rect 43196 4868 43252 4924
rect 43252 4868 43256 4924
rect 43192 4864 43256 4868
rect 7952 4380 8016 4384
rect 7952 4324 7956 4380
rect 7956 4324 8012 4380
rect 8012 4324 8016 4380
rect 7952 4320 8016 4324
rect 8032 4380 8096 4384
rect 8032 4324 8036 4380
rect 8036 4324 8092 4380
rect 8092 4324 8096 4380
rect 8032 4320 8096 4324
rect 8112 4380 8176 4384
rect 8112 4324 8116 4380
rect 8116 4324 8172 4380
rect 8172 4324 8176 4380
rect 8112 4320 8176 4324
rect 8192 4380 8256 4384
rect 8192 4324 8196 4380
rect 8196 4324 8252 4380
rect 8252 4324 8256 4380
rect 8192 4320 8256 4324
rect 17952 4380 18016 4384
rect 17952 4324 17956 4380
rect 17956 4324 18012 4380
rect 18012 4324 18016 4380
rect 17952 4320 18016 4324
rect 18032 4380 18096 4384
rect 18032 4324 18036 4380
rect 18036 4324 18092 4380
rect 18092 4324 18096 4380
rect 18032 4320 18096 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 27952 4380 28016 4384
rect 27952 4324 27956 4380
rect 27956 4324 28012 4380
rect 28012 4324 28016 4380
rect 27952 4320 28016 4324
rect 28032 4380 28096 4384
rect 28032 4324 28036 4380
rect 28036 4324 28092 4380
rect 28092 4324 28096 4380
rect 28032 4320 28096 4324
rect 28112 4380 28176 4384
rect 28112 4324 28116 4380
rect 28116 4324 28172 4380
rect 28172 4324 28176 4380
rect 28112 4320 28176 4324
rect 28192 4380 28256 4384
rect 28192 4324 28196 4380
rect 28196 4324 28252 4380
rect 28252 4324 28256 4380
rect 28192 4320 28256 4324
rect 37952 4380 38016 4384
rect 37952 4324 37956 4380
rect 37956 4324 38012 4380
rect 38012 4324 38016 4380
rect 37952 4320 38016 4324
rect 38032 4380 38096 4384
rect 38032 4324 38036 4380
rect 38036 4324 38092 4380
rect 38092 4324 38096 4380
rect 38032 4320 38096 4324
rect 38112 4380 38176 4384
rect 38112 4324 38116 4380
rect 38116 4324 38172 4380
rect 38172 4324 38176 4380
rect 38112 4320 38176 4324
rect 38192 4380 38256 4384
rect 38192 4324 38196 4380
rect 38196 4324 38252 4380
rect 38252 4324 38256 4380
rect 38192 4320 38256 4324
rect 47952 4380 48016 4384
rect 47952 4324 47956 4380
rect 47956 4324 48012 4380
rect 48012 4324 48016 4380
rect 47952 4320 48016 4324
rect 48032 4380 48096 4384
rect 48032 4324 48036 4380
rect 48036 4324 48092 4380
rect 48092 4324 48096 4380
rect 48032 4320 48096 4324
rect 48112 4380 48176 4384
rect 48112 4324 48116 4380
rect 48116 4324 48172 4380
rect 48172 4324 48176 4380
rect 48112 4320 48176 4324
rect 48192 4380 48256 4384
rect 48192 4324 48196 4380
rect 48196 4324 48252 4380
rect 48252 4324 48256 4380
rect 48192 4320 48256 4324
rect 2952 3836 3016 3840
rect 2952 3780 2956 3836
rect 2956 3780 3012 3836
rect 3012 3780 3016 3836
rect 2952 3776 3016 3780
rect 3032 3836 3096 3840
rect 3032 3780 3036 3836
rect 3036 3780 3092 3836
rect 3092 3780 3096 3836
rect 3032 3776 3096 3780
rect 3112 3836 3176 3840
rect 3112 3780 3116 3836
rect 3116 3780 3172 3836
rect 3172 3780 3176 3836
rect 3112 3776 3176 3780
rect 3192 3836 3256 3840
rect 3192 3780 3196 3836
rect 3196 3780 3252 3836
rect 3252 3780 3256 3836
rect 3192 3776 3256 3780
rect 12952 3836 13016 3840
rect 12952 3780 12956 3836
rect 12956 3780 13012 3836
rect 13012 3780 13016 3836
rect 12952 3776 13016 3780
rect 13032 3836 13096 3840
rect 13032 3780 13036 3836
rect 13036 3780 13092 3836
rect 13092 3780 13096 3836
rect 13032 3776 13096 3780
rect 13112 3836 13176 3840
rect 13112 3780 13116 3836
rect 13116 3780 13172 3836
rect 13172 3780 13176 3836
rect 13112 3776 13176 3780
rect 13192 3836 13256 3840
rect 13192 3780 13196 3836
rect 13196 3780 13252 3836
rect 13252 3780 13256 3836
rect 13192 3776 13256 3780
rect 22952 3836 23016 3840
rect 22952 3780 22956 3836
rect 22956 3780 23012 3836
rect 23012 3780 23016 3836
rect 22952 3776 23016 3780
rect 23032 3836 23096 3840
rect 23032 3780 23036 3836
rect 23036 3780 23092 3836
rect 23092 3780 23096 3836
rect 23032 3776 23096 3780
rect 23112 3836 23176 3840
rect 23112 3780 23116 3836
rect 23116 3780 23172 3836
rect 23172 3780 23176 3836
rect 23112 3776 23176 3780
rect 23192 3836 23256 3840
rect 23192 3780 23196 3836
rect 23196 3780 23252 3836
rect 23252 3780 23256 3836
rect 23192 3776 23256 3780
rect 32952 3836 33016 3840
rect 32952 3780 32956 3836
rect 32956 3780 33012 3836
rect 33012 3780 33016 3836
rect 32952 3776 33016 3780
rect 33032 3836 33096 3840
rect 33032 3780 33036 3836
rect 33036 3780 33092 3836
rect 33092 3780 33096 3836
rect 33032 3776 33096 3780
rect 33112 3836 33176 3840
rect 33112 3780 33116 3836
rect 33116 3780 33172 3836
rect 33172 3780 33176 3836
rect 33112 3776 33176 3780
rect 33192 3836 33256 3840
rect 33192 3780 33196 3836
rect 33196 3780 33252 3836
rect 33252 3780 33256 3836
rect 33192 3776 33256 3780
rect 42952 3836 43016 3840
rect 42952 3780 42956 3836
rect 42956 3780 43012 3836
rect 43012 3780 43016 3836
rect 42952 3776 43016 3780
rect 43032 3836 43096 3840
rect 43032 3780 43036 3836
rect 43036 3780 43092 3836
rect 43092 3780 43096 3836
rect 43032 3776 43096 3780
rect 43112 3836 43176 3840
rect 43112 3780 43116 3836
rect 43116 3780 43172 3836
rect 43172 3780 43176 3836
rect 43112 3776 43176 3780
rect 43192 3836 43256 3840
rect 43192 3780 43196 3836
rect 43196 3780 43252 3836
rect 43252 3780 43256 3836
rect 43192 3776 43256 3780
rect 7952 3292 8016 3296
rect 7952 3236 7956 3292
rect 7956 3236 8012 3292
rect 8012 3236 8016 3292
rect 7952 3232 8016 3236
rect 8032 3292 8096 3296
rect 8032 3236 8036 3292
rect 8036 3236 8092 3292
rect 8092 3236 8096 3292
rect 8032 3232 8096 3236
rect 8112 3292 8176 3296
rect 8112 3236 8116 3292
rect 8116 3236 8172 3292
rect 8172 3236 8176 3292
rect 8112 3232 8176 3236
rect 8192 3292 8256 3296
rect 8192 3236 8196 3292
rect 8196 3236 8252 3292
rect 8252 3236 8256 3292
rect 8192 3232 8256 3236
rect 17952 3292 18016 3296
rect 17952 3236 17956 3292
rect 17956 3236 18012 3292
rect 18012 3236 18016 3292
rect 17952 3232 18016 3236
rect 18032 3292 18096 3296
rect 18032 3236 18036 3292
rect 18036 3236 18092 3292
rect 18092 3236 18096 3292
rect 18032 3232 18096 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 27952 3292 28016 3296
rect 27952 3236 27956 3292
rect 27956 3236 28012 3292
rect 28012 3236 28016 3292
rect 27952 3232 28016 3236
rect 28032 3292 28096 3296
rect 28032 3236 28036 3292
rect 28036 3236 28092 3292
rect 28092 3236 28096 3292
rect 28032 3232 28096 3236
rect 28112 3292 28176 3296
rect 28112 3236 28116 3292
rect 28116 3236 28172 3292
rect 28172 3236 28176 3292
rect 28112 3232 28176 3236
rect 28192 3292 28256 3296
rect 28192 3236 28196 3292
rect 28196 3236 28252 3292
rect 28252 3236 28256 3292
rect 28192 3232 28256 3236
rect 37952 3292 38016 3296
rect 37952 3236 37956 3292
rect 37956 3236 38012 3292
rect 38012 3236 38016 3292
rect 37952 3232 38016 3236
rect 38032 3292 38096 3296
rect 38032 3236 38036 3292
rect 38036 3236 38092 3292
rect 38092 3236 38096 3292
rect 38032 3232 38096 3236
rect 38112 3292 38176 3296
rect 38112 3236 38116 3292
rect 38116 3236 38172 3292
rect 38172 3236 38176 3292
rect 38112 3232 38176 3236
rect 38192 3292 38256 3296
rect 38192 3236 38196 3292
rect 38196 3236 38252 3292
rect 38252 3236 38256 3292
rect 38192 3232 38256 3236
rect 47952 3292 48016 3296
rect 47952 3236 47956 3292
rect 47956 3236 48012 3292
rect 48012 3236 48016 3292
rect 47952 3232 48016 3236
rect 48032 3292 48096 3296
rect 48032 3236 48036 3292
rect 48036 3236 48092 3292
rect 48092 3236 48096 3292
rect 48032 3232 48096 3236
rect 48112 3292 48176 3296
rect 48112 3236 48116 3292
rect 48116 3236 48172 3292
rect 48172 3236 48176 3292
rect 48112 3232 48176 3236
rect 48192 3292 48256 3296
rect 48192 3236 48196 3292
rect 48196 3236 48252 3292
rect 48252 3236 48256 3292
rect 48192 3232 48256 3236
rect 2952 2748 3016 2752
rect 2952 2692 2956 2748
rect 2956 2692 3012 2748
rect 3012 2692 3016 2748
rect 2952 2688 3016 2692
rect 3032 2748 3096 2752
rect 3032 2692 3036 2748
rect 3036 2692 3092 2748
rect 3092 2692 3096 2748
rect 3032 2688 3096 2692
rect 3112 2748 3176 2752
rect 3112 2692 3116 2748
rect 3116 2692 3172 2748
rect 3172 2692 3176 2748
rect 3112 2688 3176 2692
rect 3192 2748 3256 2752
rect 3192 2692 3196 2748
rect 3196 2692 3252 2748
rect 3252 2692 3256 2748
rect 3192 2688 3256 2692
rect 12952 2748 13016 2752
rect 12952 2692 12956 2748
rect 12956 2692 13012 2748
rect 13012 2692 13016 2748
rect 12952 2688 13016 2692
rect 13032 2748 13096 2752
rect 13032 2692 13036 2748
rect 13036 2692 13092 2748
rect 13092 2692 13096 2748
rect 13032 2688 13096 2692
rect 13112 2748 13176 2752
rect 13112 2692 13116 2748
rect 13116 2692 13172 2748
rect 13172 2692 13176 2748
rect 13112 2688 13176 2692
rect 13192 2748 13256 2752
rect 13192 2692 13196 2748
rect 13196 2692 13252 2748
rect 13252 2692 13256 2748
rect 13192 2688 13256 2692
rect 22952 2748 23016 2752
rect 22952 2692 22956 2748
rect 22956 2692 23012 2748
rect 23012 2692 23016 2748
rect 22952 2688 23016 2692
rect 23032 2748 23096 2752
rect 23032 2692 23036 2748
rect 23036 2692 23092 2748
rect 23092 2692 23096 2748
rect 23032 2688 23096 2692
rect 23112 2748 23176 2752
rect 23112 2692 23116 2748
rect 23116 2692 23172 2748
rect 23172 2692 23176 2748
rect 23112 2688 23176 2692
rect 23192 2748 23256 2752
rect 23192 2692 23196 2748
rect 23196 2692 23252 2748
rect 23252 2692 23256 2748
rect 23192 2688 23256 2692
rect 32952 2748 33016 2752
rect 32952 2692 32956 2748
rect 32956 2692 33012 2748
rect 33012 2692 33016 2748
rect 32952 2688 33016 2692
rect 33032 2748 33096 2752
rect 33032 2692 33036 2748
rect 33036 2692 33092 2748
rect 33092 2692 33096 2748
rect 33032 2688 33096 2692
rect 33112 2748 33176 2752
rect 33112 2692 33116 2748
rect 33116 2692 33172 2748
rect 33172 2692 33176 2748
rect 33112 2688 33176 2692
rect 33192 2748 33256 2752
rect 33192 2692 33196 2748
rect 33196 2692 33252 2748
rect 33252 2692 33256 2748
rect 33192 2688 33256 2692
rect 42952 2748 43016 2752
rect 42952 2692 42956 2748
rect 42956 2692 43012 2748
rect 43012 2692 43016 2748
rect 42952 2688 43016 2692
rect 43032 2748 43096 2752
rect 43032 2692 43036 2748
rect 43036 2692 43092 2748
rect 43092 2692 43096 2748
rect 43032 2688 43096 2692
rect 43112 2748 43176 2752
rect 43112 2692 43116 2748
rect 43116 2692 43172 2748
rect 43172 2692 43176 2748
rect 43112 2688 43176 2692
rect 43192 2748 43256 2752
rect 43192 2692 43196 2748
rect 43196 2692 43252 2748
rect 43252 2692 43256 2748
rect 43192 2688 43256 2692
rect 7952 2204 8016 2208
rect 7952 2148 7956 2204
rect 7956 2148 8012 2204
rect 8012 2148 8016 2204
rect 7952 2144 8016 2148
rect 8032 2204 8096 2208
rect 8032 2148 8036 2204
rect 8036 2148 8092 2204
rect 8092 2148 8096 2204
rect 8032 2144 8096 2148
rect 8112 2204 8176 2208
rect 8112 2148 8116 2204
rect 8116 2148 8172 2204
rect 8172 2148 8176 2204
rect 8112 2144 8176 2148
rect 8192 2204 8256 2208
rect 8192 2148 8196 2204
rect 8196 2148 8252 2204
rect 8252 2148 8256 2204
rect 8192 2144 8256 2148
rect 17952 2204 18016 2208
rect 17952 2148 17956 2204
rect 17956 2148 18012 2204
rect 18012 2148 18016 2204
rect 17952 2144 18016 2148
rect 18032 2204 18096 2208
rect 18032 2148 18036 2204
rect 18036 2148 18092 2204
rect 18092 2148 18096 2204
rect 18032 2144 18096 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
rect 27952 2204 28016 2208
rect 27952 2148 27956 2204
rect 27956 2148 28012 2204
rect 28012 2148 28016 2204
rect 27952 2144 28016 2148
rect 28032 2204 28096 2208
rect 28032 2148 28036 2204
rect 28036 2148 28092 2204
rect 28092 2148 28096 2204
rect 28032 2144 28096 2148
rect 28112 2204 28176 2208
rect 28112 2148 28116 2204
rect 28116 2148 28172 2204
rect 28172 2148 28176 2204
rect 28112 2144 28176 2148
rect 28192 2204 28256 2208
rect 28192 2148 28196 2204
rect 28196 2148 28252 2204
rect 28252 2148 28256 2204
rect 28192 2144 28256 2148
rect 37952 2204 38016 2208
rect 37952 2148 37956 2204
rect 37956 2148 38012 2204
rect 38012 2148 38016 2204
rect 37952 2144 38016 2148
rect 38032 2204 38096 2208
rect 38032 2148 38036 2204
rect 38036 2148 38092 2204
rect 38092 2148 38096 2204
rect 38032 2144 38096 2148
rect 38112 2204 38176 2208
rect 38112 2148 38116 2204
rect 38116 2148 38172 2204
rect 38172 2148 38176 2204
rect 38112 2144 38176 2148
rect 38192 2204 38256 2208
rect 38192 2148 38196 2204
rect 38196 2148 38252 2204
rect 38252 2148 38256 2204
rect 38192 2144 38256 2148
rect 47952 2204 48016 2208
rect 47952 2148 47956 2204
rect 47956 2148 48012 2204
rect 48012 2148 48016 2204
rect 47952 2144 48016 2148
rect 48032 2204 48096 2208
rect 48032 2148 48036 2204
rect 48036 2148 48092 2204
rect 48092 2148 48096 2204
rect 48032 2144 48096 2148
rect 48112 2204 48176 2208
rect 48112 2148 48116 2204
rect 48116 2148 48172 2204
rect 48172 2148 48176 2204
rect 48112 2144 48176 2148
rect 48192 2204 48256 2208
rect 48192 2148 48196 2204
rect 48196 2148 48252 2204
rect 48252 2148 48256 2204
rect 48192 2144 48256 2148
<< metal4 >>
rect 35387 24988 35453 24989
rect 35387 24924 35388 24988
rect 35452 24924 35453 24988
rect 35387 24923 35453 24924
rect 2944 24512 3264 24528
rect 2944 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3264 24512
rect 2944 23424 3264 24448
rect 2944 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3264 23424
rect 2944 22336 3264 23360
rect 2944 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3264 22336
rect 2944 21248 3264 22272
rect 2944 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3264 21248
rect 2944 20160 3264 21184
rect 2944 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3264 20160
rect 2944 19072 3264 20096
rect 2944 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3264 19072
rect 2944 17984 3264 19008
rect 2944 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3264 17984
rect 2944 16896 3264 17920
rect 2944 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3264 16896
rect 2944 15808 3264 16832
rect 2944 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3264 15808
rect 2944 14720 3264 15744
rect 2944 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3264 14720
rect 2944 13632 3264 14656
rect 2944 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3264 13632
rect 2944 12544 3264 13568
rect 2944 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3264 12544
rect 2944 11456 3264 12480
rect 2944 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3264 11456
rect 2944 10368 3264 11392
rect 2944 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3264 10368
rect 2944 9280 3264 10304
rect 2944 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3264 9280
rect 2944 8192 3264 9216
rect 2944 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3264 8192
rect 2944 7104 3264 8128
rect 2944 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3264 7104
rect 2944 6016 3264 7040
rect 2944 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3264 6016
rect 2944 4928 3264 5952
rect 2944 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3264 4928
rect 2944 3840 3264 4864
rect 2944 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3264 3840
rect 2944 2752 3264 3776
rect 2944 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3264 2752
rect 2944 2128 3264 2688
rect 7944 23968 8264 24528
rect 7944 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8264 23968
rect 7944 22880 8264 23904
rect 7944 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8264 22880
rect 7944 21792 8264 22816
rect 7944 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8264 21792
rect 7944 20704 8264 21728
rect 7944 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8264 20704
rect 7944 19616 8264 20640
rect 7944 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8264 19616
rect 7944 18528 8264 19552
rect 7944 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8264 18528
rect 7944 17440 8264 18464
rect 7944 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8264 17440
rect 7944 16352 8264 17376
rect 7944 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8264 16352
rect 7944 15264 8264 16288
rect 7944 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8264 15264
rect 7944 14176 8264 15200
rect 7944 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8264 14176
rect 7944 13088 8264 14112
rect 7944 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8264 13088
rect 7944 12000 8264 13024
rect 7944 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8264 12000
rect 7944 10912 8264 11936
rect 7944 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8264 10912
rect 7944 9824 8264 10848
rect 7944 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8264 9824
rect 7944 8736 8264 9760
rect 7944 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8264 8736
rect 7944 7648 8264 8672
rect 7944 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8264 7648
rect 7944 6560 8264 7584
rect 7944 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8264 6560
rect 7944 5472 8264 6496
rect 7944 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8264 5472
rect 7944 4384 8264 5408
rect 7944 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8264 4384
rect 7944 3296 8264 4320
rect 7944 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8264 3296
rect 7944 2208 8264 3232
rect 7944 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8264 2208
rect 7944 2128 8264 2144
rect 12944 24512 13264 24528
rect 12944 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13264 24512
rect 12944 23424 13264 24448
rect 12944 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13264 23424
rect 12944 22336 13264 23360
rect 12944 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13264 22336
rect 12944 21248 13264 22272
rect 12944 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13264 21248
rect 12944 20160 13264 21184
rect 12944 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13264 20160
rect 12944 19072 13264 20096
rect 12944 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13264 19072
rect 12944 17984 13264 19008
rect 12944 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13264 17984
rect 12944 16896 13264 17920
rect 12944 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13264 16896
rect 12944 15808 13264 16832
rect 12944 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13264 15808
rect 12944 14720 13264 15744
rect 12944 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13264 14720
rect 12944 13632 13264 14656
rect 17944 23968 18264 24528
rect 17944 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18264 23968
rect 17944 22880 18264 23904
rect 17944 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18264 22880
rect 17944 21792 18264 22816
rect 17944 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18264 21792
rect 17944 20704 18264 21728
rect 17944 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18264 20704
rect 17944 19616 18264 20640
rect 17944 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18264 19616
rect 17944 18528 18264 19552
rect 17944 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18264 18528
rect 17944 17440 18264 18464
rect 17944 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18264 17440
rect 17944 16352 18264 17376
rect 17944 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18264 16352
rect 17944 15264 18264 16288
rect 17944 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18264 15264
rect 17944 14176 18264 15200
rect 17944 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18264 14176
rect 15699 13836 15765 13837
rect 15699 13772 15700 13836
rect 15764 13772 15765 13836
rect 15699 13771 15765 13772
rect 12944 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13264 13632
rect 12944 12544 13264 13568
rect 12944 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13264 12544
rect 12944 11456 13264 12480
rect 12944 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13264 11456
rect 12944 10368 13264 11392
rect 12944 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13264 10368
rect 12944 9280 13264 10304
rect 15702 9621 15762 13771
rect 17944 13088 18264 14112
rect 17944 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18264 13088
rect 17944 12000 18264 13024
rect 17944 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18264 12000
rect 17944 10912 18264 11936
rect 17944 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18264 10912
rect 17944 9824 18264 10848
rect 17944 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18264 9824
rect 15699 9620 15765 9621
rect 15699 9556 15700 9620
rect 15764 9556 15765 9620
rect 15699 9555 15765 9556
rect 12944 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13264 9280
rect 12944 8192 13264 9216
rect 12944 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13264 8192
rect 12944 7104 13264 8128
rect 12944 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13264 7104
rect 12944 6016 13264 7040
rect 12944 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13264 6016
rect 12944 4928 13264 5952
rect 12944 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13264 4928
rect 12944 3840 13264 4864
rect 12944 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13264 3840
rect 12944 2752 13264 3776
rect 12944 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13264 2752
rect 12944 2128 13264 2688
rect 17944 8736 18264 9760
rect 17944 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18264 8736
rect 17944 7648 18264 8672
rect 17944 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18264 7648
rect 17944 6560 18264 7584
rect 17944 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18264 6560
rect 17944 5472 18264 6496
rect 17944 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18264 5472
rect 17944 4384 18264 5408
rect 17944 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18264 4384
rect 17944 3296 18264 4320
rect 17944 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18264 3296
rect 17944 2208 18264 3232
rect 17944 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18264 2208
rect 17944 2128 18264 2144
rect 22944 24512 23264 24528
rect 22944 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23264 24512
rect 22944 23424 23264 24448
rect 22944 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23264 23424
rect 22944 22336 23264 23360
rect 22944 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23264 22336
rect 22944 21248 23264 22272
rect 22944 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23264 21248
rect 22944 20160 23264 21184
rect 22944 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23264 20160
rect 22944 19072 23264 20096
rect 22944 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23264 19072
rect 22944 17984 23264 19008
rect 22944 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23264 17984
rect 22944 16896 23264 17920
rect 22944 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23264 16896
rect 22944 15808 23264 16832
rect 22944 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23264 15808
rect 22944 14720 23264 15744
rect 22944 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23264 14720
rect 22944 13632 23264 14656
rect 22944 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23264 13632
rect 22944 12544 23264 13568
rect 22944 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23264 12544
rect 22944 11456 23264 12480
rect 22944 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23264 11456
rect 22944 10368 23264 11392
rect 22944 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23264 10368
rect 22944 9280 23264 10304
rect 22944 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23264 9280
rect 22944 8192 23264 9216
rect 22944 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23264 8192
rect 22944 7104 23264 8128
rect 22944 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23264 7104
rect 22944 6016 23264 7040
rect 22944 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23264 6016
rect 22944 4928 23264 5952
rect 22944 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23264 4928
rect 22944 3840 23264 4864
rect 22944 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23264 3840
rect 22944 2752 23264 3776
rect 22944 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23264 2752
rect 22944 2128 23264 2688
rect 27944 23968 28264 24528
rect 27944 23904 27952 23968
rect 28016 23904 28032 23968
rect 28096 23904 28112 23968
rect 28176 23904 28192 23968
rect 28256 23904 28264 23968
rect 27944 22880 28264 23904
rect 32944 24512 33264 24528
rect 32944 24448 32952 24512
rect 33016 24448 33032 24512
rect 33096 24448 33112 24512
rect 33176 24448 33192 24512
rect 33256 24448 33264 24512
rect 28947 23764 29013 23765
rect 28947 23700 28948 23764
rect 29012 23700 29013 23764
rect 28947 23699 29013 23700
rect 27944 22816 27952 22880
rect 28016 22816 28032 22880
rect 28096 22816 28112 22880
rect 28176 22816 28192 22880
rect 28256 22816 28264 22880
rect 27944 21792 28264 22816
rect 27944 21728 27952 21792
rect 28016 21728 28032 21792
rect 28096 21728 28112 21792
rect 28176 21728 28192 21792
rect 28256 21728 28264 21792
rect 27944 20704 28264 21728
rect 28950 21589 29010 23699
rect 32944 23424 33264 24448
rect 32944 23360 32952 23424
rect 33016 23360 33032 23424
rect 33096 23360 33112 23424
rect 33176 23360 33192 23424
rect 33256 23360 33264 23424
rect 32944 22336 33264 23360
rect 32944 22272 32952 22336
rect 33016 22272 33032 22336
rect 33096 22272 33112 22336
rect 33176 22272 33192 22336
rect 33256 22272 33264 22336
rect 28947 21588 29013 21589
rect 28947 21524 28948 21588
rect 29012 21524 29013 21588
rect 28947 21523 29013 21524
rect 27944 20640 27952 20704
rect 28016 20640 28032 20704
rect 28096 20640 28112 20704
rect 28176 20640 28192 20704
rect 28256 20640 28264 20704
rect 27944 19616 28264 20640
rect 28579 20364 28645 20365
rect 28579 20300 28580 20364
rect 28644 20300 28645 20364
rect 28579 20299 28645 20300
rect 28582 19685 28642 20299
rect 28579 19684 28645 19685
rect 28579 19620 28580 19684
rect 28644 19620 28645 19684
rect 28579 19619 28645 19620
rect 27944 19552 27952 19616
rect 28016 19552 28032 19616
rect 28096 19552 28112 19616
rect 28176 19552 28192 19616
rect 28256 19552 28264 19616
rect 27944 18528 28264 19552
rect 28950 19277 29010 21523
rect 32944 21248 33264 22272
rect 32944 21184 32952 21248
rect 33016 21184 33032 21248
rect 33096 21184 33112 21248
rect 33176 21184 33192 21248
rect 33256 21184 33264 21248
rect 32944 20160 33264 21184
rect 35390 20637 35450 24923
rect 37944 23968 38264 24528
rect 37944 23904 37952 23968
rect 38016 23904 38032 23968
rect 38096 23904 38112 23968
rect 38176 23904 38192 23968
rect 38256 23904 38264 23968
rect 37944 22880 38264 23904
rect 37944 22816 37952 22880
rect 38016 22816 38032 22880
rect 38096 22816 38112 22880
rect 38176 22816 38192 22880
rect 38256 22816 38264 22880
rect 37944 21792 38264 22816
rect 37944 21728 37952 21792
rect 38016 21728 38032 21792
rect 38096 21728 38112 21792
rect 38176 21728 38192 21792
rect 38256 21728 38264 21792
rect 37944 20704 38264 21728
rect 37944 20640 37952 20704
rect 38016 20640 38032 20704
rect 38096 20640 38112 20704
rect 38176 20640 38192 20704
rect 38256 20640 38264 20704
rect 35387 20636 35453 20637
rect 35387 20572 35388 20636
rect 35452 20572 35453 20636
rect 35387 20571 35453 20572
rect 32944 20096 32952 20160
rect 33016 20096 33032 20160
rect 33096 20096 33112 20160
rect 33176 20096 33192 20160
rect 33256 20096 33264 20160
rect 28947 19276 29013 19277
rect 28947 19212 28948 19276
rect 29012 19212 29013 19276
rect 28947 19211 29013 19212
rect 27944 18464 27952 18528
rect 28016 18464 28032 18528
rect 28096 18464 28112 18528
rect 28176 18464 28192 18528
rect 28256 18464 28264 18528
rect 27944 17440 28264 18464
rect 27944 17376 27952 17440
rect 28016 17376 28032 17440
rect 28096 17376 28112 17440
rect 28176 17376 28192 17440
rect 28256 17376 28264 17440
rect 27944 16352 28264 17376
rect 27944 16288 27952 16352
rect 28016 16288 28032 16352
rect 28096 16288 28112 16352
rect 28176 16288 28192 16352
rect 28256 16288 28264 16352
rect 27944 15264 28264 16288
rect 27944 15200 27952 15264
rect 28016 15200 28032 15264
rect 28096 15200 28112 15264
rect 28176 15200 28192 15264
rect 28256 15200 28264 15264
rect 27944 14176 28264 15200
rect 32944 19072 33264 20096
rect 32944 19008 32952 19072
rect 33016 19008 33032 19072
rect 33096 19008 33112 19072
rect 33176 19008 33192 19072
rect 33256 19008 33264 19072
rect 32944 17984 33264 19008
rect 32944 17920 32952 17984
rect 33016 17920 33032 17984
rect 33096 17920 33112 17984
rect 33176 17920 33192 17984
rect 33256 17920 33264 17984
rect 32944 16896 33264 17920
rect 32944 16832 32952 16896
rect 33016 16832 33032 16896
rect 33096 16832 33112 16896
rect 33176 16832 33192 16896
rect 33256 16832 33264 16896
rect 32944 15808 33264 16832
rect 32944 15744 32952 15808
rect 33016 15744 33032 15808
rect 33096 15744 33112 15808
rect 33176 15744 33192 15808
rect 33256 15744 33264 15808
rect 32944 14720 33264 15744
rect 32944 14656 32952 14720
rect 33016 14656 33032 14720
rect 33096 14656 33112 14720
rect 33176 14656 33192 14720
rect 33256 14656 33264 14720
rect 32075 14516 32141 14517
rect 32075 14452 32076 14516
rect 32140 14452 32141 14516
rect 32075 14451 32141 14452
rect 27944 14112 27952 14176
rect 28016 14112 28032 14176
rect 28096 14112 28112 14176
rect 28176 14112 28192 14176
rect 28256 14112 28264 14176
rect 27944 13088 28264 14112
rect 27944 13024 27952 13088
rect 28016 13024 28032 13088
rect 28096 13024 28112 13088
rect 28176 13024 28192 13088
rect 28256 13024 28264 13088
rect 27944 12000 28264 13024
rect 27944 11936 27952 12000
rect 28016 11936 28032 12000
rect 28096 11936 28112 12000
rect 28176 11936 28192 12000
rect 28256 11936 28264 12000
rect 27944 10912 28264 11936
rect 32078 11117 32138 14451
rect 32944 13632 33264 14656
rect 32944 13568 32952 13632
rect 33016 13568 33032 13632
rect 33096 13568 33112 13632
rect 33176 13568 33192 13632
rect 33256 13568 33264 13632
rect 32944 12544 33264 13568
rect 32944 12480 32952 12544
rect 33016 12480 33032 12544
rect 33096 12480 33112 12544
rect 33176 12480 33192 12544
rect 33256 12480 33264 12544
rect 32944 11456 33264 12480
rect 32944 11392 32952 11456
rect 33016 11392 33032 11456
rect 33096 11392 33112 11456
rect 33176 11392 33192 11456
rect 33256 11392 33264 11456
rect 32075 11116 32141 11117
rect 32075 11052 32076 11116
rect 32140 11052 32141 11116
rect 32075 11051 32141 11052
rect 27944 10848 27952 10912
rect 28016 10848 28032 10912
rect 28096 10848 28112 10912
rect 28176 10848 28192 10912
rect 28256 10848 28264 10912
rect 27944 9824 28264 10848
rect 27944 9760 27952 9824
rect 28016 9760 28032 9824
rect 28096 9760 28112 9824
rect 28176 9760 28192 9824
rect 28256 9760 28264 9824
rect 27944 8736 28264 9760
rect 27944 8672 27952 8736
rect 28016 8672 28032 8736
rect 28096 8672 28112 8736
rect 28176 8672 28192 8736
rect 28256 8672 28264 8736
rect 27944 7648 28264 8672
rect 27944 7584 27952 7648
rect 28016 7584 28032 7648
rect 28096 7584 28112 7648
rect 28176 7584 28192 7648
rect 28256 7584 28264 7648
rect 27944 6560 28264 7584
rect 27944 6496 27952 6560
rect 28016 6496 28032 6560
rect 28096 6496 28112 6560
rect 28176 6496 28192 6560
rect 28256 6496 28264 6560
rect 27944 5472 28264 6496
rect 27944 5408 27952 5472
rect 28016 5408 28032 5472
rect 28096 5408 28112 5472
rect 28176 5408 28192 5472
rect 28256 5408 28264 5472
rect 27944 4384 28264 5408
rect 27944 4320 27952 4384
rect 28016 4320 28032 4384
rect 28096 4320 28112 4384
rect 28176 4320 28192 4384
rect 28256 4320 28264 4384
rect 27944 3296 28264 4320
rect 27944 3232 27952 3296
rect 28016 3232 28032 3296
rect 28096 3232 28112 3296
rect 28176 3232 28192 3296
rect 28256 3232 28264 3296
rect 27944 2208 28264 3232
rect 27944 2144 27952 2208
rect 28016 2144 28032 2208
rect 28096 2144 28112 2208
rect 28176 2144 28192 2208
rect 28256 2144 28264 2208
rect 27944 2128 28264 2144
rect 32944 10368 33264 11392
rect 32944 10304 32952 10368
rect 33016 10304 33032 10368
rect 33096 10304 33112 10368
rect 33176 10304 33192 10368
rect 33256 10304 33264 10368
rect 32944 9280 33264 10304
rect 32944 9216 32952 9280
rect 33016 9216 33032 9280
rect 33096 9216 33112 9280
rect 33176 9216 33192 9280
rect 33256 9216 33264 9280
rect 32944 8192 33264 9216
rect 32944 8128 32952 8192
rect 33016 8128 33032 8192
rect 33096 8128 33112 8192
rect 33176 8128 33192 8192
rect 33256 8128 33264 8192
rect 32944 7104 33264 8128
rect 32944 7040 32952 7104
rect 33016 7040 33032 7104
rect 33096 7040 33112 7104
rect 33176 7040 33192 7104
rect 33256 7040 33264 7104
rect 32944 6016 33264 7040
rect 32944 5952 32952 6016
rect 33016 5952 33032 6016
rect 33096 5952 33112 6016
rect 33176 5952 33192 6016
rect 33256 5952 33264 6016
rect 32944 4928 33264 5952
rect 32944 4864 32952 4928
rect 33016 4864 33032 4928
rect 33096 4864 33112 4928
rect 33176 4864 33192 4928
rect 33256 4864 33264 4928
rect 32944 3840 33264 4864
rect 32944 3776 32952 3840
rect 33016 3776 33032 3840
rect 33096 3776 33112 3840
rect 33176 3776 33192 3840
rect 33256 3776 33264 3840
rect 32944 2752 33264 3776
rect 32944 2688 32952 2752
rect 33016 2688 33032 2752
rect 33096 2688 33112 2752
rect 33176 2688 33192 2752
rect 33256 2688 33264 2752
rect 32944 2128 33264 2688
rect 37944 19616 38264 20640
rect 37944 19552 37952 19616
rect 38016 19552 38032 19616
rect 38096 19552 38112 19616
rect 38176 19552 38192 19616
rect 38256 19552 38264 19616
rect 37944 18528 38264 19552
rect 37944 18464 37952 18528
rect 38016 18464 38032 18528
rect 38096 18464 38112 18528
rect 38176 18464 38192 18528
rect 38256 18464 38264 18528
rect 37944 17440 38264 18464
rect 37944 17376 37952 17440
rect 38016 17376 38032 17440
rect 38096 17376 38112 17440
rect 38176 17376 38192 17440
rect 38256 17376 38264 17440
rect 37944 16352 38264 17376
rect 37944 16288 37952 16352
rect 38016 16288 38032 16352
rect 38096 16288 38112 16352
rect 38176 16288 38192 16352
rect 38256 16288 38264 16352
rect 37944 15264 38264 16288
rect 37944 15200 37952 15264
rect 38016 15200 38032 15264
rect 38096 15200 38112 15264
rect 38176 15200 38192 15264
rect 38256 15200 38264 15264
rect 37944 14176 38264 15200
rect 37944 14112 37952 14176
rect 38016 14112 38032 14176
rect 38096 14112 38112 14176
rect 38176 14112 38192 14176
rect 38256 14112 38264 14176
rect 37944 13088 38264 14112
rect 37944 13024 37952 13088
rect 38016 13024 38032 13088
rect 38096 13024 38112 13088
rect 38176 13024 38192 13088
rect 38256 13024 38264 13088
rect 37944 12000 38264 13024
rect 37944 11936 37952 12000
rect 38016 11936 38032 12000
rect 38096 11936 38112 12000
rect 38176 11936 38192 12000
rect 38256 11936 38264 12000
rect 37944 10912 38264 11936
rect 37944 10848 37952 10912
rect 38016 10848 38032 10912
rect 38096 10848 38112 10912
rect 38176 10848 38192 10912
rect 38256 10848 38264 10912
rect 37944 9824 38264 10848
rect 37944 9760 37952 9824
rect 38016 9760 38032 9824
rect 38096 9760 38112 9824
rect 38176 9760 38192 9824
rect 38256 9760 38264 9824
rect 37944 8736 38264 9760
rect 37944 8672 37952 8736
rect 38016 8672 38032 8736
rect 38096 8672 38112 8736
rect 38176 8672 38192 8736
rect 38256 8672 38264 8736
rect 37944 7648 38264 8672
rect 37944 7584 37952 7648
rect 38016 7584 38032 7648
rect 38096 7584 38112 7648
rect 38176 7584 38192 7648
rect 38256 7584 38264 7648
rect 37944 6560 38264 7584
rect 37944 6496 37952 6560
rect 38016 6496 38032 6560
rect 38096 6496 38112 6560
rect 38176 6496 38192 6560
rect 38256 6496 38264 6560
rect 37944 5472 38264 6496
rect 37944 5408 37952 5472
rect 38016 5408 38032 5472
rect 38096 5408 38112 5472
rect 38176 5408 38192 5472
rect 38256 5408 38264 5472
rect 37944 4384 38264 5408
rect 37944 4320 37952 4384
rect 38016 4320 38032 4384
rect 38096 4320 38112 4384
rect 38176 4320 38192 4384
rect 38256 4320 38264 4384
rect 37944 3296 38264 4320
rect 37944 3232 37952 3296
rect 38016 3232 38032 3296
rect 38096 3232 38112 3296
rect 38176 3232 38192 3296
rect 38256 3232 38264 3296
rect 37944 2208 38264 3232
rect 37944 2144 37952 2208
rect 38016 2144 38032 2208
rect 38096 2144 38112 2208
rect 38176 2144 38192 2208
rect 38256 2144 38264 2208
rect 37944 2128 38264 2144
rect 42944 24512 43264 24528
rect 42944 24448 42952 24512
rect 43016 24448 43032 24512
rect 43096 24448 43112 24512
rect 43176 24448 43192 24512
rect 43256 24448 43264 24512
rect 42944 23424 43264 24448
rect 42944 23360 42952 23424
rect 43016 23360 43032 23424
rect 43096 23360 43112 23424
rect 43176 23360 43192 23424
rect 43256 23360 43264 23424
rect 42944 22336 43264 23360
rect 42944 22272 42952 22336
rect 43016 22272 43032 22336
rect 43096 22272 43112 22336
rect 43176 22272 43192 22336
rect 43256 22272 43264 22336
rect 42944 21248 43264 22272
rect 42944 21184 42952 21248
rect 43016 21184 43032 21248
rect 43096 21184 43112 21248
rect 43176 21184 43192 21248
rect 43256 21184 43264 21248
rect 42944 20160 43264 21184
rect 42944 20096 42952 20160
rect 43016 20096 43032 20160
rect 43096 20096 43112 20160
rect 43176 20096 43192 20160
rect 43256 20096 43264 20160
rect 42944 19072 43264 20096
rect 42944 19008 42952 19072
rect 43016 19008 43032 19072
rect 43096 19008 43112 19072
rect 43176 19008 43192 19072
rect 43256 19008 43264 19072
rect 42944 17984 43264 19008
rect 42944 17920 42952 17984
rect 43016 17920 43032 17984
rect 43096 17920 43112 17984
rect 43176 17920 43192 17984
rect 43256 17920 43264 17984
rect 42944 16896 43264 17920
rect 42944 16832 42952 16896
rect 43016 16832 43032 16896
rect 43096 16832 43112 16896
rect 43176 16832 43192 16896
rect 43256 16832 43264 16896
rect 42944 15808 43264 16832
rect 42944 15744 42952 15808
rect 43016 15744 43032 15808
rect 43096 15744 43112 15808
rect 43176 15744 43192 15808
rect 43256 15744 43264 15808
rect 42944 14720 43264 15744
rect 42944 14656 42952 14720
rect 43016 14656 43032 14720
rect 43096 14656 43112 14720
rect 43176 14656 43192 14720
rect 43256 14656 43264 14720
rect 42944 13632 43264 14656
rect 42944 13568 42952 13632
rect 43016 13568 43032 13632
rect 43096 13568 43112 13632
rect 43176 13568 43192 13632
rect 43256 13568 43264 13632
rect 42944 12544 43264 13568
rect 42944 12480 42952 12544
rect 43016 12480 43032 12544
rect 43096 12480 43112 12544
rect 43176 12480 43192 12544
rect 43256 12480 43264 12544
rect 42944 11456 43264 12480
rect 42944 11392 42952 11456
rect 43016 11392 43032 11456
rect 43096 11392 43112 11456
rect 43176 11392 43192 11456
rect 43256 11392 43264 11456
rect 42944 10368 43264 11392
rect 42944 10304 42952 10368
rect 43016 10304 43032 10368
rect 43096 10304 43112 10368
rect 43176 10304 43192 10368
rect 43256 10304 43264 10368
rect 42944 9280 43264 10304
rect 42944 9216 42952 9280
rect 43016 9216 43032 9280
rect 43096 9216 43112 9280
rect 43176 9216 43192 9280
rect 43256 9216 43264 9280
rect 42944 8192 43264 9216
rect 42944 8128 42952 8192
rect 43016 8128 43032 8192
rect 43096 8128 43112 8192
rect 43176 8128 43192 8192
rect 43256 8128 43264 8192
rect 42944 7104 43264 8128
rect 42944 7040 42952 7104
rect 43016 7040 43032 7104
rect 43096 7040 43112 7104
rect 43176 7040 43192 7104
rect 43256 7040 43264 7104
rect 42944 6016 43264 7040
rect 42944 5952 42952 6016
rect 43016 5952 43032 6016
rect 43096 5952 43112 6016
rect 43176 5952 43192 6016
rect 43256 5952 43264 6016
rect 42944 4928 43264 5952
rect 42944 4864 42952 4928
rect 43016 4864 43032 4928
rect 43096 4864 43112 4928
rect 43176 4864 43192 4928
rect 43256 4864 43264 4928
rect 42944 3840 43264 4864
rect 42944 3776 42952 3840
rect 43016 3776 43032 3840
rect 43096 3776 43112 3840
rect 43176 3776 43192 3840
rect 43256 3776 43264 3840
rect 42944 2752 43264 3776
rect 42944 2688 42952 2752
rect 43016 2688 43032 2752
rect 43096 2688 43112 2752
rect 43176 2688 43192 2752
rect 43256 2688 43264 2752
rect 42944 2128 43264 2688
rect 47944 23968 48264 24528
rect 47944 23904 47952 23968
rect 48016 23904 48032 23968
rect 48096 23904 48112 23968
rect 48176 23904 48192 23968
rect 48256 23904 48264 23968
rect 47944 22880 48264 23904
rect 47944 22816 47952 22880
rect 48016 22816 48032 22880
rect 48096 22816 48112 22880
rect 48176 22816 48192 22880
rect 48256 22816 48264 22880
rect 47944 21792 48264 22816
rect 47944 21728 47952 21792
rect 48016 21728 48032 21792
rect 48096 21728 48112 21792
rect 48176 21728 48192 21792
rect 48256 21728 48264 21792
rect 47944 20704 48264 21728
rect 47944 20640 47952 20704
rect 48016 20640 48032 20704
rect 48096 20640 48112 20704
rect 48176 20640 48192 20704
rect 48256 20640 48264 20704
rect 47944 19616 48264 20640
rect 47944 19552 47952 19616
rect 48016 19552 48032 19616
rect 48096 19552 48112 19616
rect 48176 19552 48192 19616
rect 48256 19552 48264 19616
rect 47944 18528 48264 19552
rect 47944 18464 47952 18528
rect 48016 18464 48032 18528
rect 48096 18464 48112 18528
rect 48176 18464 48192 18528
rect 48256 18464 48264 18528
rect 47944 17440 48264 18464
rect 47944 17376 47952 17440
rect 48016 17376 48032 17440
rect 48096 17376 48112 17440
rect 48176 17376 48192 17440
rect 48256 17376 48264 17440
rect 47944 16352 48264 17376
rect 47944 16288 47952 16352
rect 48016 16288 48032 16352
rect 48096 16288 48112 16352
rect 48176 16288 48192 16352
rect 48256 16288 48264 16352
rect 47944 15264 48264 16288
rect 47944 15200 47952 15264
rect 48016 15200 48032 15264
rect 48096 15200 48112 15264
rect 48176 15200 48192 15264
rect 48256 15200 48264 15264
rect 47944 14176 48264 15200
rect 47944 14112 47952 14176
rect 48016 14112 48032 14176
rect 48096 14112 48112 14176
rect 48176 14112 48192 14176
rect 48256 14112 48264 14176
rect 47944 13088 48264 14112
rect 47944 13024 47952 13088
rect 48016 13024 48032 13088
rect 48096 13024 48112 13088
rect 48176 13024 48192 13088
rect 48256 13024 48264 13088
rect 47944 12000 48264 13024
rect 47944 11936 47952 12000
rect 48016 11936 48032 12000
rect 48096 11936 48112 12000
rect 48176 11936 48192 12000
rect 48256 11936 48264 12000
rect 47944 10912 48264 11936
rect 47944 10848 47952 10912
rect 48016 10848 48032 10912
rect 48096 10848 48112 10912
rect 48176 10848 48192 10912
rect 48256 10848 48264 10912
rect 47944 9824 48264 10848
rect 47944 9760 47952 9824
rect 48016 9760 48032 9824
rect 48096 9760 48112 9824
rect 48176 9760 48192 9824
rect 48256 9760 48264 9824
rect 47944 8736 48264 9760
rect 47944 8672 47952 8736
rect 48016 8672 48032 8736
rect 48096 8672 48112 8736
rect 48176 8672 48192 8736
rect 48256 8672 48264 8736
rect 47944 7648 48264 8672
rect 47944 7584 47952 7648
rect 48016 7584 48032 7648
rect 48096 7584 48112 7648
rect 48176 7584 48192 7648
rect 48256 7584 48264 7648
rect 47944 6560 48264 7584
rect 47944 6496 47952 6560
rect 48016 6496 48032 6560
rect 48096 6496 48112 6560
rect 48176 6496 48192 6560
rect 48256 6496 48264 6560
rect 47944 5472 48264 6496
rect 47944 5408 47952 5472
rect 48016 5408 48032 5472
rect 48096 5408 48112 5472
rect 48176 5408 48192 5472
rect 48256 5408 48264 5472
rect 47944 4384 48264 5408
rect 47944 4320 47952 4384
rect 48016 4320 48032 4384
rect 48096 4320 48112 4384
rect 48176 4320 48192 4384
rect 48256 4320 48264 4384
rect 47944 3296 48264 4320
rect 47944 3232 47952 3296
rect 48016 3232 48032 3296
rect 48096 3232 48112 3296
rect 48176 3232 48192 3296
rect 48256 3232 48264 3296
rect 47944 2208 48264 3232
rect 47944 2144 47952 2208
rect 48016 2144 48032 2208
rect 48096 2144 48112 2208
rect 48176 2144 48192 2208
rect 48256 2144 48264 2208
rect 47944 2128 48264 2144
use sky130_fd_sc_hd__clkbuf_2  _104_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14260 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _105_
timestamp 1676037725
transform 1 0 11040 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _106_
timestamp 1676037725
transform 1 0 9476 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _107_
timestamp 1676037725
transform 1 0 6440 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _108_
timestamp 1676037725
transform 1 0 10212 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _109_
timestamp 1676037725
transform 1 0 10856 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _110_
timestamp 1676037725
transform 1 0 14076 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _111_
timestamp 1676037725
transform 1 0 8096 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _112_
timestamp 1676037725
transform 1 0 10304 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _113_
timestamp 1676037725
transform 1 0 10856 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _114_
timestamp 1676037725
transform 1 0 11684 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _115_
timestamp 1676037725
transform 1 0 9108 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _116_
timestamp 1676037725
transform 1 0 16560 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _117_
timestamp 1676037725
transform 1 0 16008 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _118_
timestamp 1676037725
transform 1 0 11960 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _119_
timestamp 1676037725
transform 1 0 7636 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _120_
timestamp 1676037725
transform 1 0 11224 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _121_
timestamp 1676037725
transform 1 0 12420 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _122_
timestamp 1676037725
transform 1 0 15272 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _123_
timestamp 1676037725
transform 1 0 7636 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _124_
timestamp 1676037725
transform 1 0 11684 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _125_
timestamp 1676037725
transform 1 0 12144 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _126_
timestamp 1676037725
transform 1 0 11776 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _127_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7820 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _128_
timestamp 1676037725
transform 1 0 5244 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _129_
timestamp 1676037725
transform 1 0 11408 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _130_
timestamp 1676037725
transform 1 0 7728 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _131_
timestamp 1676037725
transform 1 0 3864 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _132_
timestamp 1676037725
transform 1 0 5704 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _133_
timestamp 1676037725
transform 1 0 6624 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _134_
timestamp 1676037725
transform 1 0 36340 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _135_
timestamp 1676037725
transform 1 0 37168 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _136_
timestamp 1676037725
transform 1 0 37904 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _137_
timestamp 1676037725
transform 1 0 43608 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _138_
timestamp 1676037725
transform 1 0 38364 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _139_
timestamp 1676037725
transform 1 0 37628 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _140_
timestamp 1676037725
transform 1 0 37444 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _141_
timestamp 1676037725
transform 1 0 43884 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _142_
timestamp 1676037725
transform 1 0 38456 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _143_
timestamp 1676037725
transform 1 0 37720 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _144_
timestamp 1676037725
transform 1 0 37904 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _145_
timestamp 1676037725
transform 1 0 44804 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _146_
timestamp 1676037725
transform 1 0 38640 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _147_
timestamp 1676037725
transform 1 0 40204 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _148_
timestamp 1676037725
transform 1 0 39192 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _149_
timestamp 1676037725
transform 1 0 44160 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _150_
timestamp 1676037725
transform 1 0 40020 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _151_
timestamp 1676037725
transform 1 0 38640 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _152_
timestamp 1676037725
transform 1 0 39652 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _153_
timestamp 1676037725
transform 1 0 44252 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _154_
timestamp 1676037725
transform 1 0 40020 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _155_
timestamp 1676037725
transform 1 0 39284 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _156_
timestamp 1676037725
transform 1 0 39836 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _157_
timestamp 1676037725
transform 1 0 44988 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _158_
timestamp 1676037725
transform 1 0 45540 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _159_
timestamp 1676037725
transform 1 0 39928 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _160_
timestamp 1676037725
transform 1 0 45908 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _161_
timestamp 1676037725
transform 1 0 45908 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _162_
timestamp 1676037725
transform 1 0 45632 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _163_
timestamp 1676037725
transform 1 0 44896 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _164_
timestamp 1676037725
transform 1 0 9108 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _165_
timestamp 1676037725
transform 1 0 4048 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _166_
timestamp 1676037725
transform 1 0 5244 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _167_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4140 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _168_
timestamp 1676037725
transform 1 0 7268 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _169_
timestamp 1676037725
transform 1 0 3956 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _170_
timestamp 1676037725
transform 1 0 4692 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _171_
timestamp 1676037725
transform 1 0 6532 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _172_
timestamp 1676037725
transform 1 0 6532 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _173_
timestamp 1676037725
transform 1 0 8372 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _174_
timestamp 1676037725
transform 1 0 26036 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _175_
timestamp 1676037725
transform 1 0 12696 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _176_
timestamp 1676037725
transform 1 0 11960 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _177_
timestamp 1676037725
transform 1 0 13064 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _178_
timestamp 1676037725
transform 1 0 10948 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _179_
timestamp 1676037725
transform 1 0 13432 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _180_
timestamp 1676037725
transform 1 0 14628 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _181_
timestamp 1676037725
transform 1 0 16008 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _182_
timestamp 1676037725
transform 1 0 14444 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _183_
timestamp 1676037725
transform 1 0 14260 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _184_
timestamp 1676037725
transform 1 0 20792 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _185_
timestamp 1676037725
transform 1 0 19596 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _186_
timestamp 1676037725
transform 1 0 19596 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _187_
timestamp 1676037725
transform 1 0 23736 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _188_
timestamp 1676037725
transform 1 0 27140 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _189_
timestamp 1676037725
transform 1 0 24564 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _190_
timestamp 1676037725
transform 1 0 21252 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _191_
timestamp 1676037725
transform 1 0 27140 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _192_
timestamp 1676037725
transform 1 0 22632 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _193_
timestamp 1676037725
transform 1 0 19412 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _194_
timestamp 1676037725
transform 1 0 16376 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _195_
timestamp 1676037725
transform 1 0 17388 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _196_
timestamp 1676037725
transform 1 0 18676 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _197_
timestamp 1676037725
transform 1 0 19964 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _198_
timestamp 1676037725
transform 1 0 19412 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _199_
timestamp 1676037725
transform 1 0 20608 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _200_
timestamp 1676037725
transform 1 0 21252 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _201_
timestamp 1676037725
transform 1 0 26312 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 47932 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1676037725
transform 1 0 39192 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1676037725
transform 1 0 41308 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1676037725
transform 1 0 42964 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1676037725
transform 1 0 11224 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1676037725
transform 1 0 44528 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1676037725
transform 1 0 13064 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1676037725
transform 1 0 27600 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1676037725
transform 1 0 17572 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1676037725
transform 1 0 20700 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1676037725
transform 1 0 38548 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1676037725
transform 1 0 29532 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1676037725
transform 1 0 25760 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1676037725
transform 1 0 23460 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1676037725
transform 1 0 23184 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1676037725
transform 1 0 31740 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1676037725
transform 1 0 23828 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1676037725
transform 1 0 10672 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 1676037725
transform 1 0 18032 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 1676037725
transform 1 0 25760 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 1676037725
transform 1 0 28336 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp 1676037725
transform 1 0 28520 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp 1676037725
transform 1 0 14996 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp 1676037725
transform 1 0 16376 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp 1676037725
transform 1 0 26312 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp 1676037725
transform 1 0 43516 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp 1676037725
transform 1 0 28336 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_28
timestamp 1676037725
transform 1 0 39376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_29
timestamp 1676037725
transform 1 0 14996 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_30
timestamp 1676037725
transform 1 0 13800 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_31
timestamp 1676037725
transform 1 0 27232 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_32
timestamp 1676037725
transform 1 0 27876 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_33
timestamp 1676037725
transform 1 0 20332 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_34
timestamp 1676037725
transform 1 0 28336 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_35
timestamp 1676037725
transform 1 0 35328 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_36
timestamp 1676037725
transform 1 0 37444 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_37
timestamp 1676037725
transform 1 0 17940 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_38
timestamp 1676037725
transform 1 0 39652 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_39
timestamp 1676037725
transform 1 0 13064 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_40
timestamp 1676037725
transform 1 0 26312 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_41
timestamp 1676037725
transform 1 0 18032 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  cbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18032 0 -1 19584
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16376 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16284 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 16836 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 16836 0 -1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 14260 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 14260 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 13524 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 13248 0 -1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 10764 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 10488 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 10948 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 12052 0 -1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 13248 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 10764 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  cbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 9108 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14444 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_1_
timestamp 1676037725
transform 1 0 15548 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_2_
timestamp 1676037725
transform 1 0 15548 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_3_
timestamp 1676037725
transform 1 0 20700 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_4_
timestamp 1676037725
transform 1 0 15548 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_0_
timestamp 1676037725
transform 1 0 15180 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_1_
timestamp 1676037725
transform 1 0 17112 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_2_
timestamp 1676037725
transform 1 0 16560 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_3_
timestamp 1676037725
transform 1 0 20148 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_3__254 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18676 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l3_in_0_
timestamp 1676037725
transform 1 0 15548 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l3_in_1_
timestamp 1676037725
transform 1 0 17756 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l4_in_0_
timestamp 1676037725
transform 1 0 17664 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19688 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_0_
timestamp 1676037725
transform 1 0 10396 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_1_
timestamp 1676037725
transform 1 0 12696 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_2_
timestamp 1676037725
transform 1 0 19504 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_3_
timestamp 1676037725
transform 1 0 16836 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_4_
timestamp 1676037725
transform 1 0 17940 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12604 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_1_
timestamp 1676037725
transform 1 0 15548 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_2_
timestamp 1676037725
transform 1 0 14352 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_3_
timestamp 1676037725
transform 1 0 17756 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_3__255
timestamp 1676037725
transform 1 0 19044 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l3_in_0_
timestamp 1676037725
transform 1 0 12972 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l3_in_1_
timestamp 1676037725
transform 1 0 13156 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l4_in_0_
timestamp 1676037725
transform 1 0 15548 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 17664 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_0_
timestamp 1676037725
transform 1 0 7728 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_1_
timestamp 1676037725
transform 1 0 7912 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_2_
timestamp 1676037725
transform 1 0 18124 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_3_
timestamp 1676037725
transform 1 0 15088 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_4_
timestamp 1676037725
transform 1 0 16652 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_0_
timestamp 1676037725
transform 1 0 9384 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_1_
timestamp 1676037725
transform 1 0 14260 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_2_
timestamp 1676037725
transform 1 0 14352 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_3__256
timestamp 1676037725
transform 1 0 10948 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_3_
timestamp 1676037725
transform 1 0 11684 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l3_in_0_
timestamp 1676037725
transform 1 0 11684 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l3_in_1_
timestamp 1676037725
transform 1 0 11592 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l4_in_0_
timestamp 1676037725
transform 1 0 12052 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 15640 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_0_
timestamp 1676037725
transform 1 0 12972 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_1_
timestamp 1676037725
transform 1 0 14352 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_2_
timestamp 1676037725
transform 1 0 15640 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_3_
timestamp 1676037725
transform 1 0 18308 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_4_
timestamp 1676037725
transform 1 0 15088 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_0_
timestamp 1676037725
transform 1 0 13156 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_1_
timestamp 1676037725
transform 1 0 15548 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_2_
timestamp 1676037725
transform 1 0 14352 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_3__257
timestamp 1676037725
transform 1 0 15916 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_3_
timestamp 1676037725
transform 1 0 16376 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l3_in_0_
timestamp 1676037725
transform 1 0 11776 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l3_in_1_
timestamp 1676037725
transform 1 0 12972 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l4_in_0_
timestamp 1676037725
transform 1 0 11040 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 13524 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 27140 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23460 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 22172 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21896 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 14536 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1676037725
transform 1 0 25116 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1676037725
transform 1 0 23368 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1676037725
transform 1 0 23184 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1676037725
transform 1 0 20424 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 20884 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1676037725
transform 1 0 24104 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1676037725
transform 1 0 22632 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1676037725
transform 1 0 23552 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1676037725
transform 1 0 18952 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 24104 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1676037725
transform 1 0 24564 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1676037725
transform 1 0 22540 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1676037725
transform 1 0 27416 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1676037725
transform 1 0 18032 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_2  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 28888 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 27140 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17848 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_prog_clk
timestamp 1676037725
transform 1 0 17848 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_prog_clk
timestamp 1676037725
transform 1 0 22448 0 1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_prog_clk
timestamp 1676037725
transform 1 0 22540 0 -1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_prog_clk
timestamp 1676037725
transform 1 0 17848 0 -1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_prog_clk
timestamp 1676037725
transform 1 0 17940 0 1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_prog_clk
timestamp 1676037725
transform 1 0 23276 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_prog_clk
timestamp 1676037725
transform 1 0 21988 0 -1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_prog_clk
timestamp 1676037725
transform 1 0 28796 0 -1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_prog_clk
timestamp 1676037725
transform 1 0 28244 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_prog_clk
timestamp 1676037725
transform 1 0 33764 0 -1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_prog_clk
timestamp 1676037725
transform 1 0 34500 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_prog_clk
timestamp 1676037725
transform 1 0 30176 0 1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_prog_clk
timestamp 1676037725
transform 1 0 30820 0 -1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_prog_clk
timestamp 1676037725
transform 1 0 34592 0 -1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_prog_clk
timestamp 1676037725
transform 1 0 34868 0 1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17
timestamp 1676037725
transform 1 0 2668 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24
timestamp 1676037725
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1676037725
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1676037725
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1676037725
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1676037725
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_85 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8924 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96
timestamp 1676037725
transform 1 0 9936 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_108
timestamp 1676037725
transform 1 0 11040 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_113
timestamp 1676037725
transform 1 0 11500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_132
timestamp 1676037725
transform 1 0 13248 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1676037725
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_159
timestamp 1676037725
transform 1 0 15732 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1676037725
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_187
timestamp 1676037725
transform 1 0 18308 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1676037725
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1676037725
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_202
timestamp 1676037725
transform 1 0 19688 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1676037725
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_225 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21804 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_247
timestamp 1676037725
transform 1 0 23828 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251
timestamp 1676037725
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1676037725
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_271
timestamp 1676037725
transform 1 0 26036 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_279
timestamp 1676037725
transform 1 0 26772 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1676037725
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_299
timestamp 1676037725
transform 1 0 28612 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_306
timestamp 1676037725
transform 1 0 29256 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_309
timestamp 1676037725
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_321
timestamp 1676037725
transform 1 0 30636 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_326
timestamp 1676037725
transform 1 0 31096 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_334
timestamp 1676037725
transform 1 0 31832 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_337
timestamp 1676037725
transform 1 0 32108 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_345
timestamp 1676037725
transform 1 0 32844 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_349
timestamp 1676037725
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 1676037725
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_365
timestamp 1676037725
transform 1 0 34684 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_372
timestamp 1676037725
transform 1 0 35328 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_384
timestamp 1676037725
transform 1 0 36432 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_393
timestamp 1676037725
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_405
timestamp 1676037725
transform 1 0 38364 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_417
timestamp 1676037725
transform 1 0 39468 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_421
timestamp 1676037725
transform 1 0 39836 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_429
timestamp 1676037725
transform 1 0 40572 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_446
timestamp 1676037725
transform 1 0 42136 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_449
timestamp 1676037725
transform 1 0 42412 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_471
timestamp 1676037725
transform 1 0 44436 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_475
timestamp 1676037725
transform 1 0 44804 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_477
timestamp 1676037725
transform 1 0 44988 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_485
timestamp 1676037725
transform 1 0 45724 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_502
timestamp 1676037725
transform 1 0 47288 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_505
timestamp 1676037725
transform 1 0 47564 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_525
timestamp 1676037725
transform 1 0 49404 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_9
timestamp 1676037725
transform 1 0 1932 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_21
timestamp 1676037725
transform 1 0 3036 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_33
timestamp 1676037725
transform 1 0 4140 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_45
timestamp 1676037725
transform 1 0 5244 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_53
timestamp 1676037725
transform 1 0 5980 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1676037725
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1676037725
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1676037725
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1676037725
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1676037725
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1676037725
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1676037725
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_137
timestamp 1676037725
transform 1 0 13708 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_145
timestamp 1676037725
transform 1 0 14444 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp 1676037725
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_169
timestamp 1676037725
transform 1 0 16652 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_180
timestamp 1676037725
transform 1 0 17664 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_184
timestamp 1676037725
transform 1 0 18032 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_201
timestamp 1676037725
transform 1 0 19596 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_208
timestamp 1676037725
transform 1 0 20240 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_215
timestamp 1676037725
transform 1 0 20884 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp 1676037725
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_225
timestamp 1676037725
transform 1 0 21804 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_235
timestamp 1676037725
transform 1 0 22724 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_239
timestamp 1676037725
transform 1 0 23092 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_246
timestamp 1676037725
transform 1 0 23736 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_270
timestamp 1676037725
transform 1 0 25944 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_277
timestamp 1676037725
transform 1 0 26588 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_281
timestamp 1676037725
transform 1 0 26956 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_285
timestamp 1676037725
transform 1 0 27324 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_292
timestamp 1676037725
transform 1 0 27968 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_300
timestamp 1676037725
transform 1 0 28704 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_323
timestamp 1676037725
transform 1 0 30820 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1676037725
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1676037725
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1676037725
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1676037725
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1676037725
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 1676037725
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1676037725
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_393
timestamp 1676037725
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_405
timestamp 1676037725
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_417
timestamp 1676037725
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_429
timestamp 1676037725
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_441
timestamp 1676037725
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1676037725
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_449
timestamp 1676037725
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_461
timestamp 1676037725
transform 1 0 43516 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_465
timestamp 1676037725
transform 1 0 43884 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_482
timestamp 1676037725
transform 1 0 45448 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_502
timestamp 1676037725
transform 1 0 47288 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_505
timestamp 1676037725
transform 1 0 47564 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_525
timestamp 1676037725
transform 1 0 49404 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1676037725
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1676037725
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1676037725
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1676037725
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1676037725
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1676037725
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1676037725
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1676037725
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1676037725
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1676037725
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1676037725
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1676037725
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1676037725
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1676037725
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1676037725
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_165
timestamp 1676037725
transform 1 0 16284 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_170
timestamp 1676037725
transform 1 0 16744 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_182
timestamp 1676037725
transform 1 0 17848 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp 1676037725
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1676037725
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_209
timestamp 1676037725
transform 1 0 20332 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_235
timestamp 1676037725
transform 1 0 22724 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_243
timestamp 1676037725
transform 1 0 23460 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_250
timestamp 1676037725
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_253
timestamp 1676037725
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_276
timestamp 1676037725
transform 1 0 26496 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_288
timestamp 1676037725
transform 1 0 27600 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_300
timestamp 1676037725
transform 1 0 28704 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1676037725
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1676037725
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1676037725
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1676037725
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1676037725
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1676037725
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1676037725
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_377
timestamp 1676037725
transform 1 0 35788 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_387
timestamp 1676037725
transform 1 0 36708 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_399
timestamp 1676037725
transform 1 0 37812 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_411
timestamp 1676037725
transform 1 0 38916 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1676037725
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_421
timestamp 1676037725
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_433
timestamp 1676037725
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_445
timestamp 1676037725
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_457
timestamp 1676037725
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_469
timestamp 1676037725
transform 1 0 44252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 1676037725
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_477
timestamp 1676037725
transform 1 0 44988 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_485
timestamp 1676037725
transform 1 0 45724 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_505
timestamp 1676037725
transform 1 0 47564 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_525
timestamp 1676037725
transform 1 0 49404 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_9
timestamp 1676037725
transform 1 0 1932 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_17
timestamp 1676037725
transform 1 0 2668 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_29
timestamp 1676037725
transform 1 0 3772 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_41
timestamp 1676037725
transform 1 0 4876 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_53
timestamp 1676037725
transform 1 0 5980 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1676037725
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1676037725
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1676037725
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1676037725
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1676037725
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1676037725
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1676037725
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1676037725
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1676037725
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1676037725
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1676037725
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1676037725
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1676037725
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1676037725
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1676037725
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1676037725
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1676037725
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_225
timestamp 1676037725
transform 1 0 21804 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_3_236
timestamp 1676037725
transform 1 0 22816 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_242
timestamp 1676037725
transform 1 0 23368 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_246
timestamp 1676037725
transform 1 0 23736 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_271
timestamp 1676037725
transform 1 0 26036 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1676037725
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_281
timestamp 1676037725
transform 1 0 26956 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_304
timestamp 1676037725
transform 1 0 29072 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_316
timestamp 1676037725
transform 1 0 30176 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_328
timestamp 1676037725
transform 1 0 31280 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1676037725
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1676037725
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1676037725
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1676037725
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1676037725
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1676037725
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1676037725
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1676037725
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1676037725
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1676037725
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1676037725
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1676037725
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1676037725
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 1676037725
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_473
timestamp 1676037725
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_485
timestamp 1676037725
transform 1 0 45724 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_502
timestamp 1676037725
transform 1 0 47288 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_505
timestamp 1676037725
transform 1 0 47564 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_525
timestamp 1676037725
transform 1 0 49404 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_9
timestamp 1676037725
transform 1 0 1932 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_21
timestamp 1676037725
transform 1 0 3036 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1676037725
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1676037725
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1676037725
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1676037725
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1676037725
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1676037725
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1676037725
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1676037725
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1676037725
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1676037725
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1676037725
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1676037725
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1676037725
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1676037725
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1676037725
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1676037725
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1676037725
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1676037725
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_209
timestamp 1676037725
transform 1 0 20332 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_218
timestamp 1676037725
transform 1 0 21160 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_4_234
timestamp 1676037725
transform 1 0 22632 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1676037725
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1676037725
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_253
timestamp 1676037725
transform 1 0 24380 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_282
timestamp 1676037725
transform 1 0 27048 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_294
timestamp 1676037725
transform 1 0 28152 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_306
timestamp 1676037725
transform 1 0 29256 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1676037725
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1676037725
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1676037725
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1676037725
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1676037725
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1676037725
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1676037725
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1676037725
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_389
timestamp 1676037725
transform 1 0 36892 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_396
timestamp 1676037725
transform 1 0 37536 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_404
timestamp 1676037725
transform 1 0 38272 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_416
timestamp 1676037725
transform 1 0 39376 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1676037725
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1676037725
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1676037725
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_457
timestamp 1676037725
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1676037725
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1676037725
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1676037725
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_489
timestamp 1676037725
transform 1 0 46092 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_497
timestamp 1676037725
transform 1 0 46828 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_505
timestamp 1676037725
transform 1 0 47564 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_525
timestamp 1676037725
transform 1 0 49404 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1676037725
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1676037725
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1676037725
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1676037725
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1676037725
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1676037725
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1676037725
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1676037725
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1676037725
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1676037725
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1676037725
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1676037725
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1676037725
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1676037725
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1676037725
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1676037725
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1676037725
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1676037725
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_193
timestamp 1676037725
transform 1 0 18860 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_202
timestamp 1676037725
transform 1 0 19688 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_214
timestamp 1676037725
transform 1 0 20792 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_222
timestamp 1676037725
transform 1 0 21528 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_225
timestamp 1676037725
transform 1 0 21804 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_233
timestamp 1676037725
transform 1 0 22540 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1676037725
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1676037725
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1676037725
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1676037725
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1676037725
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1676037725
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1676037725
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1676037725
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1676037725
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1676037725
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1676037725
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1676037725
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1676037725
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1676037725
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1676037725
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1676037725
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1676037725
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_393
timestamp 1676037725
transform 1 0 37260 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_401
timestamp 1676037725
transform 1 0 37996 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_409
timestamp 1676037725
transform 1 0 38732 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_421
timestamp 1676037725
transform 1 0 39836 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_433
timestamp 1676037725
transform 1 0 40940 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_445
timestamp 1676037725
transform 1 0 42044 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1676037725
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1676037725
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_473
timestamp 1676037725
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_485
timestamp 1676037725
transform 1 0 45724 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_502
timestamp 1676037725
transform 1 0 47288 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_505
timestamp 1676037725
transform 1 0 47564 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_525
timestamp 1676037725
transform 1 0 49404 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_9
timestamp 1676037725
transform 1 0 1932 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_17
timestamp 1676037725
transform 1 0 2668 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_25
timestamp 1676037725
transform 1 0 3404 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1676037725
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1676037725
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1676037725
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1676037725
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1676037725
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1676037725
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1676037725
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1676037725
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1676037725
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1676037725
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1676037725
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1676037725
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1676037725
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1676037725
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1676037725
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1676037725
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1676037725
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1676037725
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1676037725
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1676037725
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1676037725
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1676037725
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1676037725
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1676037725
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1676037725
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1676037725
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1676037725
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1676037725
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1676037725
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1676037725
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1676037725
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1676037725
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1676037725
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1676037725
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1676037725
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1676037725
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1676037725
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_401
timestamp 1676037725
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1676037725
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1676037725
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1676037725
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1676037725
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1676037725
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_457
timestamp 1676037725
transform 1 0 43148 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_461
timestamp 1676037725
transform 1 0 43516 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_466
timestamp 1676037725
transform 1 0 43976 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_474
timestamp 1676037725
transform 1 0 44712 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1676037725
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1676037725
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_501
timestamp 1676037725
transform 1 0 47196 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_525
timestamp 1676037725
transform 1 0 49404 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_9
timestamp 1676037725
transform 1 0 1932 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_21
timestamp 1676037725
transform 1 0 3036 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_33
timestamp 1676037725
transform 1 0 4140 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_45
timestamp 1676037725
transform 1 0 5244 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_53
timestamp 1676037725
transform 1 0 5980 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1676037725
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1676037725
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1676037725
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1676037725
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1676037725
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1676037725
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1676037725
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1676037725
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1676037725
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1676037725
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1676037725
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1676037725
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_181
timestamp 1676037725
transform 1 0 17756 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_192
timestamp 1676037725
transform 1 0 18768 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_204
timestamp 1676037725
transform 1 0 19872 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_216
timestamp 1676037725
transform 1 0 20976 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1676037725
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1676037725
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1676037725
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1676037725
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1676037725
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1676037725
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1676037725
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1676037725
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1676037725
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1676037725
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1676037725
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1676037725
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1676037725
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1676037725
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1676037725
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1676037725
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1676037725
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1676037725
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_393
timestamp 1676037725
transform 1 0 37260 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_399
timestamp 1676037725
transform 1 0 37812 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_411
timestamp 1676037725
transform 1 0 38916 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_423
timestamp 1676037725
transform 1 0 40020 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_435
timestamp 1676037725
transform 1 0 41124 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1676037725
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1676037725
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_461
timestamp 1676037725
transform 1 0 43516 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_469
timestamp 1676037725
transform 1 0 44252 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_481
timestamp 1676037725
transform 1 0 45356 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_493
timestamp 1676037725
transform 1 0 46460 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_501
timestamp 1676037725
transform 1 0 47196 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_505
timestamp 1676037725
transform 1 0 47564 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_525
timestamp 1676037725
transform 1 0 49404 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_9
timestamp 1676037725
transform 1 0 1932 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_16
timestamp 1676037725
transform 1 0 2576 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1676037725
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1676037725
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1676037725
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1676037725
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1676037725
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1676037725
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1676037725
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1676037725
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1676037725
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1676037725
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1676037725
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1676037725
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1676037725
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1676037725
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1676037725
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1676037725
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_197
timestamp 1676037725
transform 1 0 19228 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_201
timestamp 1676037725
transform 1 0 19596 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_205
timestamp 1676037725
transform 1 0 19964 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_217
timestamp 1676037725
transform 1 0 21068 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_229
timestamp 1676037725
transform 1 0 22172 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_241
timestamp 1676037725
transform 1 0 23276 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_249
timestamp 1676037725
transform 1 0 24012 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1676037725
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1676037725
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1676037725
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1676037725
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1676037725
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1676037725
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1676037725
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1676037725
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1676037725
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1676037725
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1676037725
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1676037725
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1676037725
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1676037725
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1676037725
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_401
timestamp 1676037725
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1676037725
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1676037725
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1676037725
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1676037725
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1676037725
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 1676037725
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1676037725
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1676037725
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1676037725
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_505
timestamp 1676037725
transform 1 0 47564 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_525
timestamp 1676037725
transform 1 0 49404 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_9
timestamp 1676037725
transform 1 0 1932 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_21
timestamp 1676037725
transform 1 0 3036 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_33
timestamp 1676037725
transform 1 0 4140 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_45
timestamp 1676037725
transform 1 0 5244 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_53
timestamp 1676037725
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1676037725
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1676037725
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1676037725
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1676037725
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1676037725
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1676037725
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1676037725
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1676037725
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1676037725
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1676037725
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1676037725
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_169
timestamp 1676037725
transform 1 0 16652 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_177
timestamp 1676037725
transform 1 0 17388 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_183
timestamp 1676037725
transform 1 0 17940 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_195
timestamp 1676037725
transform 1 0 19044 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_207
timestamp 1676037725
transform 1 0 20148 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_219
timestamp 1676037725
transform 1 0 21252 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1676037725
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_225
timestamp 1676037725
transform 1 0 21804 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_236
timestamp 1676037725
transform 1 0 22816 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_242
timestamp 1676037725
transform 1 0 23368 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_254
timestamp 1676037725
transform 1 0 24472 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_266
timestamp 1676037725
transform 1 0 25576 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_278
timestamp 1676037725
transform 1 0 26680 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1676037725
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1676037725
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1676037725
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_317
timestamp 1676037725
transform 1 0 30268 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_323
timestamp 1676037725
transform 1 0 30820 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_327
timestamp 1676037725
transform 1 0 31188 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1676037725
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1676037725
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1676037725
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1676037725
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1676037725
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1676037725
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1676037725
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_393
timestamp 1676037725
transform 1 0 37260 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_397
timestamp 1676037725
transform 1 0 37628 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_402
timestamp 1676037725
transform 1 0 38088 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_410
timestamp 1676037725
transform 1 0 38824 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_422
timestamp 1676037725
transform 1 0 39928 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_434
timestamp 1676037725
transform 1 0 41032 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_446
timestamp 1676037725
transform 1 0 42136 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1676037725
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1676037725
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_473
timestamp 1676037725
transform 1 0 44620 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_479
timestamp 1676037725
transform 1 0 45172 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_491
timestamp 1676037725
transform 1 0 46276 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1676037725
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_505
timestamp 1676037725
transform 1 0 47564 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_525
timestamp 1676037725
transform 1 0 49404 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_9
timestamp 1676037725
transform 1 0 1932 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_21
timestamp 1676037725
transform 1 0 3036 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1676037725
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1676037725
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1676037725
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1676037725
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1676037725
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1676037725
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1676037725
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1676037725
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1676037725
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1676037725
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1676037725
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1676037725
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1676037725
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_153
timestamp 1676037725
transform 1 0 15180 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_157
timestamp 1676037725
transform 1 0 15548 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_161
timestamp 1676037725
transform 1 0 15916 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_173
timestamp 1676037725
transform 1 0 17020 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_179
timestamp 1676037725
transform 1 0 17572 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1676037725
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1676037725
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1676037725
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_219
timestamp 1676037725
transform 1 0 21252 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_10_236
timestamp 1676037725
transform 1 0 22816 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_248
timestamp 1676037725
transform 1 0 23920 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1676037725
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1676037725
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1676037725
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1676037725
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1676037725
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1676037725
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_309
timestamp 1676037725
transform 1 0 29532 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_314
timestamp 1676037725
transform 1 0 29992 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_329
timestamp 1676037725
transform 1 0 31372 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_335
timestamp 1676037725
transform 1 0 31924 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_348
timestamp 1676037725
transform 1 0 33120 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_360
timestamp 1676037725
transform 1 0 34224 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1676037725
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1676037725
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_389
timestamp 1676037725
transform 1 0 36892 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_397
timestamp 1676037725
transform 1 0 37628 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_404
timestamp 1676037725
transform 1 0 38272 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_412
timestamp 1676037725
transform 1 0 39008 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 1676037725
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_433
timestamp 1676037725
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_445
timestamp 1676037725
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_457
timestamp 1676037725
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1676037725
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1676037725
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_477
timestamp 1676037725
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_489
timestamp 1676037725
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_501
timestamp 1676037725
transform 1 0 47196 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_525
timestamp 1676037725
transform 1 0 49404 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1676037725
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1676037725
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1676037725
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1676037725
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1676037725
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1676037725
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1676037725
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1676037725
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1676037725
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1676037725
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1676037725
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1676037725
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1676037725
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_125
timestamp 1676037725
transform 1 0 12604 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_133
timestamp 1676037725
transform 1 0 13340 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_155
timestamp 1676037725
transform 1 0 15364 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1676037725
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp 1676037725
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_191
timestamp 1676037725
transform 1 0 18676 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_198
timestamp 1676037725
transform 1 0 19320 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_222
timestamp 1676037725
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_225
timestamp 1676037725
transform 1 0 21804 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_247
timestamp 1676037725
transform 1 0 23828 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_259
timestamp 1676037725
transform 1 0 24932 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_271
timestamp 1676037725
transform 1 0 26036 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1676037725
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1676037725
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_293
timestamp 1676037725
transform 1 0 28060 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_321
timestamp 1676037725
transform 1 0 30636 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_334
timestamp 1676037725
transform 1 0 31832 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_337
timestamp 1676037725
transform 1 0 32108 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_359
timestamp 1676037725
transform 1 0 34132 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_371
timestamp 1676037725
transform 1 0 35236 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_383
timestamp 1676037725
transform 1 0 36340 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1676037725
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_393
timestamp 1676037725
transform 1 0 37260 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_398
timestamp 1676037725
transform 1 0 37720 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_410
timestamp 1676037725
transform 1 0 38824 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_414
timestamp 1676037725
transform 1 0 39192 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_422
timestamp 1676037725
transform 1 0 39928 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_429
timestamp 1676037725
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1676037725
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1676037725
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_449
timestamp 1676037725
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_461
timestamp 1676037725
transform 1 0 43516 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_467
timestamp 1676037725
transform 1 0 44068 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_472
timestamp 1676037725
transform 1 0 44528 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_484
timestamp 1676037725
transform 1 0 45632 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_502
timestamp 1676037725
transform 1 0 47288 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_505
timestamp 1676037725
transform 1 0 47564 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_525
timestamp 1676037725
transform 1 0 49404 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1676037725
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_9
timestamp 1676037725
transform 1 0 1932 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_17
timestamp 1676037725
transform 1 0 2668 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_25
timestamp 1676037725
transform 1 0 3404 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1676037725
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1676037725
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1676037725
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1676037725
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1676037725
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1676037725
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1676037725
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1676037725
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1676037725
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1676037725
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_133
timestamp 1676037725
transform 1 0 13340 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1676037725
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_141
timestamp 1676037725
transform 1 0 14076 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1676037725
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_185
timestamp 1676037725
transform 1 0 18124 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1676037725
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_197
timestamp 1676037725
transform 1 0 19228 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_219
timestamp 1676037725
transform 1 0 21252 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_226
timestamp 1676037725
transform 1 0 21896 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_250
timestamp 1676037725
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_253
timestamp 1676037725
transform 1 0 24380 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_264
timestamp 1676037725
transform 1 0 25392 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_276
timestamp 1676037725
transform 1 0 26496 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_290
timestamp 1676037725
transform 1 0 27784 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_303
timestamp 1676037725
transform 1 0 28980 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1676037725
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_309
timestamp 1676037725
transform 1 0 29532 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_314
timestamp 1676037725
transform 1 0 29992 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_12_342
timestamp 1676037725
transform 1 0 32568 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_359
timestamp 1676037725
transform 1 0 34132 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1676037725
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_365
timestamp 1676037725
transform 1 0 34684 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_376
timestamp 1676037725
transform 1 0 35696 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_384
timestamp 1676037725
transform 1 0 36432 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_389
timestamp 1676037725
transform 1 0 36892 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_12_400
timestamp 1676037725
transform 1 0 37904 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_412
timestamp 1676037725
transform 1 0 39008 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_418
timestamp 1676037725
transform 1 0 39560 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_421
timestamp 1676037725
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_433
timestamp 1676037725
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_445
timestamp 1676037725
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_457
timestamp 1676037725
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1676037725
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1676037725
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_477
timestamp 1676037725
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_489
timestamp 1676037725
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_501
timestamp 1676037725
transform 1 0 47196 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_525
timestamp 1676037725
transform 1 0 49404 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1676037725
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_9
timestamp 1676037725
transform 1 0 1932 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_21
timestamp 1676037725
transform 1 0 3036 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_33
timestamp 1676037725
transform 1 0 4140 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_45
timestamp 1676037725
transform 1 0 5244 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_53
timestamp 1676037725
transform 1 0 5980 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1676037725
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1676037725
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1676037725
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1676037725
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1676037725
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1676037725
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_113
timestamp 1676037725
transform 1 0 11500 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_128
timestamp 1676037725
transform 1 0 12880 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_155
timestamp 1676037725
transform 1 0 15364 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1676037725
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1676037725
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_194
timestamp 1676037725
transform 1 0 18952 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_218
timestamp 1676037725
transform 1 0 21160 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_225
timestamp 1676037725
transform 1 0 21804 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_229
timestamp 1676037725
transform 1 0 22172 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_239
timestamp 1676037725
transform 1 0 23092 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_265
timestamp 1676037725
transform 1 0 25484 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_276
timestamp 1676037725
transform 1 0 26496 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_281
timestamp 1676037725
transform 1 0 26956 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_307
timestamp 1676037725
transform 1 0 29348 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_331
timestamp 1676037725
transform 1 0 31556 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1676037725
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_337
timestamp 1676037725
transform 1 0 32108 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_341
timestamp 1676037725
transform 1 0 32476 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_351
timestamp 1676037725
transform 1 0 33396 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_355
timestamp 1676037725
transform 1 0 33764 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_376
timestamp 1676037725
transform 1 0 35696 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_388
timestamp 1676037725
transform 1 0 36800 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1676037725
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_405
timestamp 1676037725
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_417
timestamp 1676037725
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_429
timestamp 1676037725
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1676037725
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1676037725
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_449
timestamp 1676037725
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_461
timestamp 1676037725
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_473
timestamp 1676037725
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_485
timestamp 1676037725
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1676037725
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1676037725
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_505
timestamp 1676037725
transform 1 0 47564 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_525
timestamp 1676037725
transform 1 0 49404 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1676037725
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1676037725
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1676037725
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1676037725
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1676037725
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1676037725
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1676037725
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1676037725
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1676037725
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1676037725
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1676037725
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_109
timestamp 1676037725
transform 1 0 11132 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_113
timestamp 1676037725
transform 1 0 11500 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_123
timestamp 1676037725
transform 1 0 12420 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_136
timestamp 1676037725
transform 1 0 13616 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_141
timestamp 1676037725
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_163
timestamp 1676037725
transform 1 0 16100 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_167
timestamp 1676037725
transform 1 0 16468 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_177
timestamp 1676037725
transform 1 0 17388 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_190
timestamp 1676037725
transform 1 0 18584 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_14_197
timestamp 1676037725
transform 1 0 19228 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_203
timestamp 1676037725
transform 1 0 19780 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_207
timestamp 1676037725
transform 1 0 20148 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_228
timestamp 1676037725
transform 1 0 22080 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_243
timestamp 1676037725
transform 1 0 23460 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_250
timestamp 1676037725
transform 1 0 24104 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1676037725
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_275
timestamp 1676037725
transform 1 0 26404 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1676037725
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1676037725
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_309
timestamp 1676037725
transform 1 0 29532 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_314
timestamp 1676037725
transform 1 0 29992 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_338
timestamp 1676037725
transform 1 0 32200 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_351
timestamp 1676037725
transform 1 0 33396 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_358
timestamp 1676037725
transform 1 0 34040 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_365
timestamp 1676037725
transform 1 0 34684 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_387
timestamp 1676037725
transform 1 0 36708 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_404
timestamp 1676037725
transform 1 0 38272 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_412
timestamp 1676037725
transform 1 0 39008 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_421
timestamp 1676037725
transform 1 0 39836 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_427
timestamp 1676037725
transform 1 0 40388 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_439
timestamp 1676037725
transform 1 0 41492 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_451
timestamp 1676037725
transform 1 0 42596 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_463
timestamp 1676037725
transform 1 0 43700 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_14_473
timestamp 1676037725
transform 1 0 44620 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_477
timestamp 1676037725
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_505
timestamp 1676037725
transform 1 0 47564 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_525
timestamp 1676037725
transform 1 0 49404 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1676037725
transform 1 0 1380 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_9
timestamp 1676037725
transform 1 0 1932 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_17
timestamp 1676037725
transform 1 0 2668 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_29
timestamp 1676037725
transform 1 0 3772 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_41
timestamp 1676037725
transform 1 0 4876 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_53
timestamp 1676037725
transform 1 0 5980 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1676037725
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1676037725
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1676037725
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1676037725
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1676037725
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1676037725
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1676037725
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_125
timestamp 1676037725
transform 1 0 12604 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_140
timestamp 1676037725
transform 1 0 13984 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_153
timestamp 1676037725
transform 1 0 15180 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1676037725
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_169
timestamp 1676037725
transform 1 0 16652 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_173
timestamp 1676037725
transform 1 0 17020 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_177
timestamp 1676037725
transform 1 0 17388 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_190
timestamp 1676037725
transform 1 0 18584 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_203
timestamp 1676037725
transform 1 0 19780 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_216
timestamp 1676037725
transform 1 0 20976 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_225
timestamp 1676037725
transform 1 0 21804 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_247
timestamp 1676037725
transform 1 0 23828 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_260
timestamp 1676037725
transform 1 0 25024 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_267
timestamp 1676037725
transform 1 0 25668 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1676037725
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_281
timestamp 1676037725
transform 1 0 26956 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_292
timestamp 1676037725
transform 1 0 27968 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_298
timestamp 1676037725
transform 1 0 28520 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_312
timestamp 1676037725
transform 1 0 29808 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_325
timestamp 1676037725
transform 1 0 31004 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_332
timestamp 1676037725
transform 1 0 31648 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_337
timestamp 1676037725
transform 1 0 32108 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_348
timestamp 1676037725
transform 1 0 33120 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_354
timestamp 1676037725
transform 1 0 33672 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_376
timestamp 1676037725
transform 1 0 35696 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_389
timestamp 1676037725
transform 1 0 36892 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_393
timestamp 1676037725
transform 1 0 37260 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_404
timestamp 1676037725
transform 1 0 38272 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_416
timestamp 1676037725
transform 1 0 39376 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_423
timestamp 1676037725
transform 1 0 40020 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_435
timestamp 1676037725
transform 1 0 41124 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1676037725
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_449
timestamp 1676037725
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_461
timestamp 1676037725
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_473
timestamp 1676037725
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_485
timestamp 1676037725
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1676037725
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1676037725
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_505
timestamp 1676037725
transform 1 0 47564 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_525
timestamp 1676037725
transform 1 0 49404 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1676037725
transform 1 0 1380 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_9
timestamp 1676037725
transform 1 0 1932 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_21
timestamp 1676037725
transform 1 0 3036 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1676037725
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1676037725
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1676037725
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1676037725
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1676037725
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1676037725
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1676037725
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1676037725
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_97
timestamp 1676037725
transform 1 0 10028 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_105
timestamp 1676037725
transform 1 0 10764 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_127
timestamp 1676037725
transform 1 0 12788 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1676037725
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_141
timestamp 1676037725
transform 1 0 14076 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_153
timestamp 1676037725
transform 1 0 15180 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_166
timestamp 1676037725
transform 1 0 16376 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_179
timestamp 1676037725
transform 1 0 17572 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_192
timestamp 1676037725
transform 1 0 18768 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_197
timestamp 1676037725
transform 1 0 19228 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_206
timestamp 1676037725
transform 1 0 20056 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_230
timestamp 1676037725
transform 1 0 22264 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_234
timestamp 1676037725
transform 1 0 22632 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_244
timestamp 1676037725
transform 1 0 23552 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_253
timestamp 1676037725
transform 1 0 24380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_275
timestamp 1676037725
transform 1 0 26404 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_279
timestamp 1676037725
transform 1 0 26772 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_300
timestamp 1676037725
transform 1 0 28704 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_309
timestamp 1676037725
transform 1 0 29532 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_320
timestamp 1676037725
transform 1 0 30544 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_346
timestamp 1676037725
transform 1 0 32936 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_359
timestamp 1676037725
transform 1 0 34132 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1676037725
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1676037725
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_400
timestamp 1676037725
transform 1 0 37904 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_407
timestamp 1676037725
transform 1 0 38548 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1676037725
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_421
timestamp 1676037725
transform 1 0 39836 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_427
timestamp 1676037725
transform 1 0 40388 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_434
timestamp 1676037725
transform 1 0 41032 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_446
timestamp 1676037725
transform 1 0 42136 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_458
timestamp 1676037725
transform 1 0 43240 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_470
timestamp 1676037725
transform 1 0 44344 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_16_477
timestamp 1676037725
transform 1 0 44988 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_487
timestamp 1676037725
transform 1 0 45908 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_499
timestamp 1676037725
transform 1 0 47012 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_507
timestamp 1676037725
transform 1 0 47748 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_525
timestamp 1676037725
transform 1 0 49404 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1676037725
transform 1 0 1380 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_9
timestamp 1676037725
transform 1 0 1932 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_16
timestamp 1676037725
transform 1 0 2576 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_28
timestamp 1676037725
transform 1 0 3680 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_40
timestamp 1676037725
transform 1 0 4784 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_52
timestamp 1676037725
transform 1 0 5888 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1676037725
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1676037725
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1676037725
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1676037725
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1676037725
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1676037725
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_113
timestamp 1676037725
transform 1 0 11500 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_17_142
timestamp 1676037725
transform 1 0 14168 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_150
timestamp 1676037725
transform 1 0 14904 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1676037725
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1676037725
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1676037725
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_191
timestamp 1676037725
transform 1 0 18676 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_199
timestamp 1676037725
transform 1 0 19412 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_209
timestamp 1676037725
transform 1 0 20332 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_222
timestamp 1676037725
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_225
timestamp 1676037725
transform 1 0 21804 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_244
timestamp 1676037725
transform 1 0 23552 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_268
timestamp 1676037725
transform 1 0 25760 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_274
timestamp 1676037725
transform 1 0 26312 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_278
timestamp 1676037725
transform 1 0 26680 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_281
timestamp 1676037725
transform 1 0 26956 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_292
timestamp 1676037725
transform 1 0 27968 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_296
timestamp 1676037725
transform 1 0 28336 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_318
timestamp 1676037725
transform 1 0 30360 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_331
timestamp 1676037725
transform 1 0 31556 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1676037725
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_337
timestamp 1676037725
transform 1 0 32108 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_348
timestamp 1676037725
transform 1 0 33120 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_354
timestamp 1676037725
transform 1 0 33672 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_366
timestamp 1676037725
transform 1 0 34776 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_390
timestamp 1676037725
transform 1 0 36984 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_411
timestamp 1676037725
transform 1 0 38916 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_419
timestamp 1676037725
transform 1 0 39652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_431
timestamp 1676037725
transform 1 0 40756 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_443
timestamp 1676037725
transform 1 0 41860 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1676037725
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_449
timestamp 1676037725
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_461
timestamp 1676037725
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_473
timestamp 1676037725
transform 1 0 44620 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_481
timestamp 1676037725
transform 1 0 45356 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_493
timestamp 1676037725
transform 1 0 46460 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_501
timestamp 1676037725
transform 1 0 47196 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_505
timestamp 1676037725
transform 1 0 47564 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_525
timestamp 1676037725
transform 1 0 49404 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1676037725
transform 1 0 1380 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1676037725
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1676037725
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1676037725
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1676037725
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1676037725
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1676037725
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1676037725
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1676037725
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1676037725
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_97
timestamp 1676037725
transform 1 0 10028 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_101
timestamp 1676037725
transform 1 0 10396 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_122
timestamp 1676037725
transform 1 0 12328 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_128
timestamp 1676037725
transform 1 0 12880 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1676037725
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1676037725
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_164
timestamp 1676037725
transform 1 0 16192 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_168
timestamp 1676037725
transform 1 0 16560 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_178
timestamp 1676037725
transform 1 0 17480 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_193
timestamp 1676037725
transform 1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_197
timestamp 1676037725
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_208
timestamp 1676037725
transform 1 0 20240 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_223
timestamp 1676037725
transform 1 0 21620 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_227
timestamp 1676037725
transform 1 0 21988 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_237
timestamp 1676037725
transform 1 0 22908 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_250
timestamp 1676037725
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1676037725
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_275
timestamp 1676037725
transform 1 0 26404 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_290
timestamp 1676037725
transform 1 0 27784 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_294
timestamp 1676037725
transform 1 0 28152 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_306
timestamp 1676037725
transform 1 0 29256 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_309
timestamp 1676037725
transform 1 0 29532 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_331
timestamp 1676037725
transform 1 0 31556 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1676037725
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1676037725
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_365
timestamp 1676037725
transform 1 0 34684 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_387
timestamp 1676037725
transform 1 0 36708 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_418
timestamp 1676037725
transform 1 0 39560 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_428
timestamp 1676037725
transform 1 0 40480 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_18_439
timestamp 1676037725
transform 1 0 41492 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_451
timestamp 1676037725
transform 1 0 42596 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_463
timestamp 1676037725
transform 1 0 43700 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1676037725
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_477
timestamp 1676037725
transform 1 0 44988 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_485
timestamp 1676037725
transform 1 0 45724 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_490
timestamp 1676037725
transform 1 0 46184 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_502
timestamp 1676037725
transform 1 0 47288 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_508
timestamp 1676037725
transform 1 0 47840 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_525
timestamp 1676037725
transform 1 0 49404 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1676037725
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_9
timestamp 1676037725
transform 1 0 1932 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_17
timestamp 1676037725
transform 1 0 2668 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_22
timestamp 1676037725
transform 1 0 3128 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_34
timestamp 1676037725
transform 1 0 4232 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_46
timestamp 1676037725
transform 1 0 5336 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_54
timestamp 1676037725
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1676037725
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1676037725
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1676037725
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1676037725
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1676037725
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1676037725
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_113
timestamp 1676037725
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_124
timestamp 1676037725
transform 1 0 12512 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_128
timestamp 1676037725
transform 1 0 12880 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_149
timestamp 1676037725
transform 1 0 14812 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1676037725
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_169
timestamp 1676037725
transform 1 0 16652 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_178
timestamp 1676037725
transform 1 0 17480 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_211
timestamp 1676037725
transform 1 0 20516 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1676037725
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1676037725
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_230
timestamp 1676037725
transform 1 0 22264 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_243
timestamp 1676037725
transform 1 0 23460 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_269
timestamp 1676037725
transform 1 0 25852 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_277
timestamp 1676037725
transform 1 0 26588 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_281
timestamp 1676037725
transform 1 0 26956 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_288
timestamp 1676037725
transform 1 0 27600 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_312
timestamp 1676037725
transform 1 0 29808 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_325
timestamp 1676037725
transform 1 0 31004 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_332
timestamp 1676037725
transform 1 0 31648 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_337
timestamp 1676037725
transform 1 0 32108 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_359
timestamp 1676037725
transform 1 0 34132 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_374
timestamp 1676037725
transform 1 0 35512 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_387
timestamp 1676037725
transform 1 0 36708 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1676037725
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_393
timestamp 1676037725
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_405
timestamp 1676037725
transform 1 0 38364 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_409
timestamp 1676037725
transform 1 0 38732 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_415
timestamp 1676037725
transform 1 0 39284 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_418
timestamp 1676037725
transform 1 0 39560 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_426
timestamp 1676037725
transform 1 0 40296 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_438
timestamp 1676037725
transform 1 0 41400 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_446
timestamp 1676037725
transform 1 0 42136 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_449
timestamp 1676037725
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_461
timestamp 1676037725
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_473
timestamp 1676037725
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_485
timestamp 1676037725
transform 1 0 45724 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_490
timestamp 1676037725
transform 1 0 46184 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_502
timestamp 1676037725
transform 1 0 47288 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_505
timestamp 1676037725
transform 1 0 47564 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_525
timestamp 1676037725
transform 1 0 49404 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1676037725
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_21
timestamp 1676037725
transform 1 0 3036 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1676037725
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1676037725
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1676037725
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1676037725
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1676037725
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1676037725
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1676037725
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1676037725
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_97
timestamp 1676037725
transform 1 0 10028 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_126
timestamp 1676037725
transform 1 0 12696 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1676037725
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1676037725
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1676037725
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_147
timestamp 1676037725
transform 1 0 14628 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_162
timestamp 1676037725
transform 1 0 16008 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_187
timestamp 1676037725
transform 1 0 18308 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1676037725
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1676037725
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_211
timestamp 1676037725
transform 1 0 20516 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_224
timestamp 1676037725
transform 1 0 21712 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_237
timestamp 1676037725
transform 1 0 22908 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_250
timestamp 1676037725
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_253
timestamp 1676037725
transform 1 0 24380 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_257
timestamp 1676037725
transform 1 0 24748 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_267
timestamp 1676037725
transform 1 0 25668 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_274
timestamp 1676037725
transform 1 0 26312 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_278
timestamp 1676037725
transform 1 0 26680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_302
timestamp 1676037725
transform 1 0 28888 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_309
timestamp 1676037725
transform 1 0 29532 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_320
timestamp 1676037725
transform 1 0 30544 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_324
timestamp 1676037725
transform 1 0 30912 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_346
timestamp 1676037725
transform 1 0 32936 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_359
timestamp 1676037725
transform 1 0 34132 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1676037725
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_365
timestamp 1676037725
transform 1 0 34684 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_376
timestamp 1676037725
transform 1 0 35696 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_382
timestamp 1676037725
transform 1 0 36248 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_403
timestamp 1676037725
transform 1 0 38180 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_415
timestamp 1676037725
transform 1 0 39284 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1676037725
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_421
timestamp 1676037725
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_433
timestamp 1676037725
transform 1 0 40940 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_440
timestamp 1676037725
transform 1 0 41584 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_452
timestamp 1676037725
transform 1 0 42688 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_464
timestamp 1676037725
transform 1 0 43792 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_477
timestamp 1676037725
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_489
timestamp 1676037725
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_501
timestamp 1676037725
transform 1 0 47196 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_525
timestamp 1676037725
transform 1 0 49404 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1676037725
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_21
timestamp 1676037725
transform 1 0 3036 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_29
timestamp 1676037725
transform 1 0 3772 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_41
timestamp 1676037725
transform 1 0 4876 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_53
timestamp 1676037725
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1676037725
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1676037725
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1676037725
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1676037725
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_105
timestamp 1676037725
transform 1 0 10764 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1676037725
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_113
timestamp 1676037725
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_124
timestamp 1676037725
transform 1 0 12512 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_148
timestamp 1676037725
transform 1 0 14720 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_156
timestamp 1676037725
transform 1 0 15456 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1676037725
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_169
timestamp 1676037725
transform 1 0 16652 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_173
timestamp 1676037725
transform 1 0 17020 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_183
timestamp 1676037725
transform 1 0 17940 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_196
timestamp 1676037725
transform 1 0 19136 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1676037725
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_225
timestamp 1676037725
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_247
timestamp 1676037725
transform 1 0 23828 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_254
timestamp 1676037725
transform 1 0 24472 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_278
timestamp 1676037725
transform 1 0 26680 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_281
timestamp 1676037725
transform 1 0 26956 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_303
timestamp 1676037725
transform 1 0 28980 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_327
timestamp 1676037725
transform 1 0 31188 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_334
timestamp 1676037725
transform 1 0 31832 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_337
timestamp 1676037725
transform 1 0 32108 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_359
timestamp 1676037725
transform 1 0 34132 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_372
timestamp 1676037725
transform 1 0 35328 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1676037725
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1676037725
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_393
timestamp 1676037725
transform 1 0 37260 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_404
timestamp 1676037725
transform 1 0 38272 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_411
timestamp 1676037725
transform 1 0 38916 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_423
timestamp 1676037725
transform 1 0 40020 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_435
timestamp 1676037725
transform 1 0 41124 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1676037725
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_449
timestamp 1676037725
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_461
timestamp 1676037725
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_473
timestamp 1676037725
transform 1 0 44620 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_480
timestamp 1676037725
transform 1 0 45264 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_487
timestamp 1676037725
transform 1 0 45908 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_499
timestamp 1676037725
transform 1 0 47012 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1676037725
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_505
timestamp 1676037725
transform 1 0 47564 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_513
timestamp 1676037725
transform 1 0 48300 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_517
timestamp 1676037725
transform 1 0 48668 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_525
timestamp 1676037725
transform 1 0 49404 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1676037725
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_21
timestamp 1676037725
transform 1 0 3036 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1676037725
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1676037725
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1676037725
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1676037725
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1676037725
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1676037725
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1676037725
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_85
timestamp 1676037725
transform 1 0 8924 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_95
timestamp 1676037725
transform 1 0 9844 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_103
timestamp 1676037725
transform 1 0 10580 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_107
timestamp 1676037725
transform 1 0 10948 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_112
timestamp 1676037725
transform 1 0 11408 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_125
timestamp 1676037725
transform 1 0 12604 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1676037725
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1676037725
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_164
timestamp 1676037725
transform 1 0 16192 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_175
timestamp 1676037725
transform 1 0 17204 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_181
timestamp 1676037725
transform 1 0 17756 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1676037725
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_197
timestamp 1676037725
transform 1 0 19228 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_209
timestamp 1676037725
transform 1 0 20332 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_215
timestamp 1676037725
transform 1 0 20884 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_238
timestamp 1676037725
transform 1 0 23000 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_246
timestamp 1676037725
transform 1 0 23736 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_250
timestamp 1676037725
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_253
timestamp 1676037725
transform 1 0 24380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_280
timestamp 1676037725
transform 1 0 26864 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_286
timestamp 1676037725
transform 1 0 27416 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_299
timestamp 1676037725
transform 1 0 28612 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1676037725
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_309
timestamp 1676037725
transform 1 0 29532 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_320
timestamp 1676037725
transform 1 0 30544 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_324
timestamp 1676037725
transform 1 0 30912 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_334
timestamp 1676037725
transform 1 0 31832 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_347
timestamp 1676037725
transform 1 0 33028 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_360
timestamp 1676037725
transform 1 0 34224 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_365
timestamp 1676037725
transform 1 0 34684 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_387
timestamp 1676037725
transform 1 0 36708 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_411
timestamp 1676037725
transform 1 0 38916 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_418
timestamp 1676037725
transform 1 0 39560 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_421
timestamp 1676037725
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_433
timestamp 1676037725
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_445
timestamp 1676037725
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_457
timestamp 1676037725
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_469
timestamp 1676037725
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1676037725
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_477
timestamp 1676037725
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_489
timestamp 1676037725
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_501
timestamp 1676037725
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_513
timestamp 1676037725
transform 1 0 48300 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_525
timestamp 1676037725
transform 1 0 49404 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1676037725
transform 1 0 1380 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_21
timestamp 1676037725
transform 1 0 3036 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_33
timestamp 1676037725
transform 1 0 4140 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_45
timestamp 1676037725
transform 1 0 5244 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_53
timestamp 1676037725
transform 1 0 5980 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1676037725
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1676037725
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_81
timestamp 1676037725
transform 1 0 8556 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_89
timestamp 1676037725
transform 1 0 9292 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_99
timestamp 1676037725
transform 1 0 10212 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_105
timestamp 1676037725
transform 1 0 10764 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1676037725
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_113
timestamp 1676037725
transform 1 0 11500 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_126
timestamp 1676037725
transform 1 0 12696 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_153
timestamp 1676037725
transform 1 0 15180 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1676037725
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_169
timestamp 1676037725
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_180
timestamp 1676037725
transform 1 0 17664 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_186
timestamp 1676037725
transform 1 0 18216 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_196
timestamp 1676037725
transform 1 0 19136 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_209
timestamp 1676037725
transform 1 0 20332 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_222
timestamp 1676037725
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_225
timestamp 1676037725
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_246
timestamp 1676037725
transform 1 0 23736 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_259
timestamp 1676037725
transform 1 0 24932 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_270
timestamp 1676037725
transform 1 0 25944 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_276
timestamp 1676037725
transform 1 0 26496 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_281
timestamp 1676037725
transform 1 0 26956 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_292
timestamp 1676037725
transform 1 0 27968 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_305
timestamp 1676037725
transform 1 0 29164 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_320
timestamp 1676037725
transform 1 0 30544 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_324
timestamp 1676037725
transform 1 0 30912 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_334
timestamp 1676037725
transform 1 0 31832 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_337
timestamp 1676037725
transform 1 0 32108 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_348
timestamp 1676037725
transform 1 0 33120 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_361
timestamp 1676037725
transform 1 0 34316 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_374
timestamp 1676037725
transform 1 0 35512 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_387
timestamp 1676037725
transform 1 0 36708 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1676037725
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_393
timestamp 1676037725
transform 1 0 37260 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_415
timestamp 1676037725
transform 1 0 39284 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_428
timestamp 1676037725
transform 1 0 40480 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_435
timestamp 1676037725
transform 1 0 41124 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1676037725
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_449
timestamp 1676037725
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_461
timestamp 1676037725
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_473
timestamp 1676037725
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_485
timestamp 1676037725
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 1676037725
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1676037725
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_505
timestamp 1676037725
transform 1 0 47564 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_517
timestamp 1676037725
transform 1 0 48668 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_525
timestamp 1676037725
transform 1 0 49404 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1676037725
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_21
timestamp 1676037725
transform 1 0 3036 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1676037725
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1676037725
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1676037725
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_53
timestamp 1676037725
transform 1 0 5980 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_57
timestamp 1676037725
transform 1 0 6348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_62
timestamp 1676037725
transform 1 0 6808 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_74
timestamp 1676037725
transform 1 0 7912 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1676037725
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1676037725
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_97
timestamp 1676037725
transform 1 0 10028 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_24_125
timestamp 1676037725
transform 1 0 12604 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_24_141
timestamp 1676037725
transform 1 0 14076 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_149
timestamp 1676037725
transform 1 0 14812 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_153
timestamp 1676037725
transform 1 0 15180 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_166
timestamp 1676037725
transform 1 0 16376 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_179
timestamp 1676037725
transform 1 0 17572 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_185
timestamp 1676037725
transform 1 0 18124 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_191
timestamp 1676037725
transform 1 0 18676 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1676037725
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_197
timestamp 1676037725
transform 1 0 19228 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_203
timestamp 1676037725
transform 1 0 19780 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_213
timestamp 1676037725
transform 1 0 20700 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_217
timestamp 1676037725
transform 1 0 21068 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_227
timestamp 1676037725
transform 1 0 21988 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_248
timestamp 1676037725
transform 1 0 23920 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_253
timestamp 1676037725
transform 1 0 24380 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_265
timestamp 1676037725
transform 1 0 25484 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_278
timestamp 1676037725
transform 1 0 26680 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_24_295
timestamp 1676037725
transform 1 0 28244 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_306
timestamp 1676037725
transform 1 0 29256 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_309
timestamp 1676037725
transform 1 0 29532 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_315
timestamp 1676037725
transform 1 0 30084 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_339
timestamp 1676037725
transform 1 0 32292 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_352
timestamp 1676037725
transform 1 0 33488 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_359
timestamp 1676037725
transform 1 0 34132 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1676037725
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_365
timestamp 1676037725
transform 1 0 34684 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_387
timestamp 1676037725
transform 1 0 36708 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_394
timestamp 1676037725
transform 1 0 37352 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_418
timestamp 1676037725
transform 1 0 39560 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_421
timestamp 1676037725
transform 1 0 39836 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_443
timestamp 1676037725
transform 1 0 41860 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_455
timestamp 1676037725
transform 1 0 42964 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_467
timestamp 1676037725
transform 1 0 44068 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1676037725
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_477
timestamp 1676037725
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_489
timestamp 1676037725
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_501
timestamp 1676037725
transform 1 0 47196 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_513
timestamp 1676037725
transform 1 0 48300 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_521
timestamp 1676037725
transform 1 0 49036 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_525
timestamp 1676037725
transform 1 0 49404 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1676037725
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_21
timestamp 1676037725
transform 1 0 3036 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_33
timestamp 1676037725
transform 1 0 4140 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_45
timestamp 1676037725
transform 1 0 5244 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_53
timestamp 1676037725
transform 1 0 5980 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1676037725
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_69
timestamp 1676037725
transform 1 0 7452 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_73
timestamp 1676037725
transform 1 0 7820 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_83
timestamp 1676037725
transform 1 0 8740 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_91
timestamp 1676037725
transform 1 0 9476 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_103
timestamp 1676037725
transform 1 0 10580 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1676037725
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_113
timestamp 1676037725
transform 1 0 11500 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_134
timestamp 1676037725
transform 1 0 13432 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_140
timestamp 1676037725
transform 1 0 13984 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_153
timestamp 1676037725
transform 1 0 15180 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1676037725
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_169
timestamp 1676037725
transform 1 0 16652 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_25_186
timestamp 1676037725
transform 1 0 18216 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_194
timestamp 1676037725
transform 1 0 18952 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1676037725
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1676037725
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1676037725
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_237
timestamp 1676037725
transform 1 0 22908 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_247
timestamp 1676037725
transform 1 0 23828 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_270
timestamp 1676037725
transform 1 0 25944 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_276
timestamp 1676037725
transform 1 0 26496 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_281
timestamp 1676037725
transform 1 0 26956 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_292
timestamp 1676037725
transform 1 0 27968 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_318
timestamp 1676037725
transform 1 0 30360 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_25_330
timestamp 1676037725
transform 1 0 31464 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_337
timestamp 1676037725
transform 1 0 32108 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_348
timestamp 1676037725
transform 1 0 33120 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_361
timestamp 1676037725
transform 1 0 34316 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_390
timestamp 1676037725
transform 1 0 36984 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_393
timestamp 1676037725
transform 1 0 37260 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_401
timestamp 1676037725
transform 1 0 37996 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_423
timestamp 1676037725
transform 1 0 40020 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_427
timestamp 1676037725
transform 1 0 40388 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_437
timestamp 1676037725
transform 1 0 41308 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_445
timestamp 1676037725
transform 1 0 42044 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_449
timestamp 1676037725
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_461
timestamp 1676037725
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_473
timestamp 1676037725
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_485
timestamp 1676037725
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 1676037725
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1676037725
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_505
timestamp 1676037725
transform 1 0 47564 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_517
timestamp 1676037725
transform 1 0 48668 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_525
timestamp 1676037725
transform 1 0 49404 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1676037725
transform 1 0 1380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_21
timestamp 1676037725
transform 1 0 3036 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1676037725
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1676037725
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1676037725
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1676037725
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_65
timestamp 1676037725
transform 1 0 7084 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_71
timestamp 1676037725
transform 1 0 7636 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_81
timestamp 1676037725
transform 1 0 8556 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1676037725
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_97
timestamp 1676037725
transform 1 0 10028 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_104
timestamp 1676037725
transform 1 0 10672 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_117
timestamp 1676037725
transform 1 0 11868 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_121
timestamp 1676037725
transform 1 0 12236 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_125
timestamp 1676037725
transform 1 0 12604 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1676037725
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_141
timestamp 1676037725
transform 1 0 14076 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_154
timestamp 1676037725
transform 1 0 15272 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_167
timestamp 1676037725
transform 1 0 16468 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_173
timestamp 1676037725
transform 1 0 17020 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1676037725
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1676037725
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_202
timestamp 1676037725
transform 1 0 19688 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_209
timestamp 1676037725
transform 1 0 20332 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_215
timestamp 1676037725
transform 1 0 20884 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_236
timestamp 1676037725
transform 1 0 22816 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_240
timestamp 1676037725
transform 1 0 23184 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_250
timestamp 1676037725
transform 1 0 24104 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_253
timestamp 1676037725
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_258
timestamp 1676037725
transform 1 0 24840 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_26_286
timestamp 1676037725
transform 1 0 27416 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_298
timestamp 1676037725
transform 1 0 28520 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_306
timestamp 1676037725
transform 1 0 29256 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_309
timestamp 1676037725
transform 1 0 29532 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_320
timestamp 1676037725
transform 1 0 30544 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_333
timestamp 1676037725
transform 1 0 31740 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_359
timestamp 1676037725
transform 1 0 34132 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1676037725
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_365
timestamp 1676037725
transform 1 0 34684 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_378
timestamp 1676037725
transform 1 0 35880 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_391
timestamp 1676037725
transform 1 0 37076 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_397
timestamp 1676037725
transform 1 0 37628 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_418
timestamp 1676037725
transform 1 0 39560 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_421
timestamp 1676037725
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_433
timestamp 1676037725
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_445
timestamp 1676037725
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_457
timestamp 1676037725
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_469
timestamp 1676037725
transform 1 0 44252 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1676037725
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_477
timestamp 1676037725
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_489
timestamp 1676037725
transform 1 0 46092 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_501
timestamp 1676037725
transform 1 0 47196 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_513
timestamp 1676037725
transform 1 0 48300 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_525
timestamp 1676037725
transform 1 0 49404 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1676037725
transform 1 0 1380 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_21
timestamp 1676037725
transform 1 0 3036 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_33
timestamp 1676037725
transform 1 0 4140 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_45
timestamp 1676037725
transform 1 0 5244 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_53
timestamp 1676037725
transform 1 0 5980 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1676037725
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1676037725
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1676037725
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_93
timestamp 1676037725
transform 1 0 9660 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 1676037725
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 1676037725
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_119
timestamp 1676037725
transform 1 0 12052 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_125
timestamp 1676037725
transform 1 0 12604 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_135
timestamp 1676037725
transform 1 0 13524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_27_145
timestamp 1676037725
transform 1 0 14444 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_156
timestamp 1676037725
transform 1 0 15456 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1676037725
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1676037725
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_175
timestamp 1676037725
transform 1 0 17204 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_181
timestamp 1676037725
transform 1 0 17756 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_193
timestamp 1676037725
transform 1 0 18860 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1676037725
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1676037725
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_225
timestamp 1676037725
transform 1 0 21804 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_233
timestamp 1676037725
transform 1 0 22540 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_255
timestamp 1676037725
transform 1 0 24564 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_268
timestamp 1676037725
transform 1 0 25760 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_281
timestamp 1676037725
transform 1 0 26956 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_294
timestamp 1676037725
transform 1 0 28152 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_309
timestamp 1676037725
transform 1 0 29532 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_321
timestamp 1676037725
transform 1 0 30636 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_334
timestamp 1676037725
transform 1 0 31832 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_337
timestamp 1676037725
transform 1 0 32108 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_360
timestamp 1676037725
transform 1 0 34224 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_375
timestamp 1676037725
transform 1 0 35604 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_388
timestamp 1676037725
transform 1 0 36800 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_393
timestamp 1676037725
transform 1 0 37260 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_404
timestamp 1676037725
transform 1 0 38272 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_410
timestamp 1676037725
transform 1 0 38824 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_431
timestamp 1676037725
transform 1 0 40756 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_443
timestamp 1676037725
transform 1 0 41860 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1676037725
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_449
timestamp 1676037725
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_461
timestamp 1676037725
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_473
timestamp 1676037725
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_485
timestamp 1676037725
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_497
timestamp 1676037725
transform 1 0 46828 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1676037725
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_505
timestamp 1676037725
transform 1 0 47564 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_513
timestamp 1676037725
transform 1 0 48300 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_517
timestamp 1676037725
transform 1 0 48668 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_525
timestamp 1676037725
transform 1 0 49404 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1676037725
transform 1 0 1380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_21
timestamp 1676037725
transform 1 0 3036 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1676037725
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1676037725
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1676037725
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1676037725
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1676037725
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1676037725
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1676037725
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1676037725
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_97
timestamp 1676037725
transform 1 0 10028 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_123
timestamp 1676037725
transform 1 0 12420 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_127
timestamp 1676037725
transform 1 0 12788 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_131
timestamp 1676037725
transform 1 0 13156 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1676037725
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_141
timestamp 1676037725
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_163
timestamp 1676037725
transform 1 0 16100 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_167
timestamp 1676037725
transform 1 0 16468 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_171
timestamp 1676037725
transform 1 0 16836 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_179
timestamp 1676037725
transform 1 0 17572 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1676037725
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1676037725
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_202
timestamp 1676037725
transform 1 0 19688 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_228
timestamp 1676037725
transform 1 0 22080 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_235
timestamp 1676037725
transform 1 0 22724 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_250
timestamp 1676037725
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_253
timestamp 1676037725
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_258
timestamp 1676037725
transform 1 0 24840 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_271
timestamp 1676037725
transform 1 0 26036 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_279
timestamp 1676037725
transform 1 0 26772 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_28_302
timestamp 1676037725
transform 1 0 28888 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_28_309
timestamp 1676037725
transform 1 0 29532 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_315
timestamp 1676037725
transform 1 0 30084 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_327
timestamp 1676037725
transform 1 0 31188 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_340
timestamp 1676037725
transform 1 0 32384 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_353
timestamp 1676037725
transform 1 0 33580 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_361
timestamp 1676037725
transform 1 0 34316 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_365
timestamp 1676037725
transform 1 0 34684 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_370
timestamp 1676037725
transform 1 0 35144 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_376
timestamp 1676037725
transform 1 0 35696 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_397
timestamp 1676037725
transform 1 0 37628 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_410
timestamp 1676037725
transform 1 0 38824 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_418
timestamp 1676037725
transform 1 0 39560 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_421
timestamp 1676037725
transform 1 0 39836 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_427
timestamp 1676037725
transform 1 0 40388 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_437
timestamp 1676037725
transform 1 0 41308 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_449
timestamp 1676037725
transform 1 0 42412 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_461
timestamp 1676037725
transform 1 0 43516 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_473
timestamp 1676037725
transform 1 0 44620 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_477
timestamp 1676037725
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_489
timestamp 1676037725
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_501
timestamp 1676037725
transform 1 0 47196 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_513
timestamp 1676037725
transform 1 0 48300 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_525
timestamp 1676037725
transform 1 0 49404 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1676037725
transform 1 0 1380 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_21
timestamp 1676037725
transform 1 0 3036 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_43
timestamp 1676037725
transform 1 0 5060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1676037725
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1676037725
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_69
timestamp 1676037725
transform 1 0 7452 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_75
timestamp 1676037725
transform 1 0 8004 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_87
timestamp 1676037725
transform 1 0 9108 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_93
timestamp 1676037725
transform 1 0 9660 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_97
timestamp 1676037725
transform 1 0 10028 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_110
timestamp 1676037725
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_113
timestamp 1676037725
transform 1 0 11500 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_135
timestamp 1676037725
transform 1 0 13524 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_148
timestamp 1676037725
transform 1 0 14720 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_159
timestamp 1676037725
transform 1 0 15732 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1676037725
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1676037725
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_180
timestamp 1676037725
transform 1 0 17664 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_195
timestamp 1676037725
transform 1 0 19044 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_222
timestamp 1676037725
transform 1 0 21528 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_225
timestamp 1676037725
transform 1 0 21804 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_236
timestamp 1676037725
transform 1 0 22816 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_240
timestamp 1676037725
transform 1 0 23184 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_252
timestamp 1676037725
transform 1 0 24288 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_265
timestamp 1676037725
transform 1 0 25484 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_278
timestamp 1676037725
transform 1 0 26680 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_281
timestamp 1676037725
transform 1 0 26956 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_292
timestamp 1676037725
transform 1 0 27968 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_307
timestamp 1676037725
transform 1 0 29348 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_324
timestamp 1676037725
transform 1 0 30912 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_331
timestamp 1676037725
transform 1 0 31556 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1676037725
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_337
timestamp 1676037725
transform 1 0 32108 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_348
timestamp 1676037725
transform 1 0 33120 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_352
timestamp 1676037725
transform 1 0 33488 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_373
timestamp 1676037725
transform 1 0 35420 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_386
timestamp 1676037725
transform 1 0 36616 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_29_393
timestamp 1676037725
transform 1 0 37260 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_401
timestamp 1676037725
transform 1 0 37996 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_422
timestamp 1676037725
transform 1 0 39928 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_426
timestamp 1676037725
transform 1 0 40296 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_436
timestamp 1676037725
transform 1 0 41216 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_449
timestamp 1676037725
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_461
timestamp 1676037725
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_473
timestamp 1676037725
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_485
timestamp 1676037725
transform 1 0 45724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_497
timestamp 1676037725
transform 1 0 46828 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1676037725
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_505
timestamp 1676037725
transform 1 0 47564 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_517
timestamp 1676037725
transform 1 0 48668 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_525
timestamp 1676037725
transform 1 0 49404 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1676037725
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_21
timestamp 1676037725
transform 1 0 3036 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1676037725
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_29
timestamp 1676037725
transform 1 0 3772 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_47
timestamp 1676037725
transform 1 0 5428 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_59
timestamp 1676037725
transform 1 0 6532 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_71
timestamp 1676037725
transform 1 0 7636 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_75
timestamp 1676037725
transform 1 0 8004 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_80
timestamp 1676037725
transform 1 0 8464 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_85
timestamp 1676037725
transform 1 0 8924 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_108
timestamp 1676037725
transform 1 0 11040 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_116
timestamp 1676037725
transform 1 0 11776 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_120
timestamp 1676037725
transform 1 0 12144 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1676037725
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1676037725
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_141
timestamp 1676037725
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_163
timestamp 1676037725
transform 1 0 16100 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_169
timestamp 1676037725
transform 1 0 16652 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_179
timestamp 1676037725
transform 1 0 17572 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_192
timestamp 1676037725
transform 1 0 18768 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_197
timestamp 1676037725
transform 1 0 19228 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_212
timestamp 1676037725
transform 1 0 20608 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_216
timestamp 1676037725
transform 1 0 20976 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_226
timestamp 1676037725
transform 1 0 21896 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_250
timestamp 1676037725
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1676037725
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_264
timestamp 1676037725
transform 1 0 25392 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_288
timestamp 1676037725
transform 1 0 27600 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_300
timestamp 1676037725
transform 1 0 28704 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_306
timestamp 1676037725
transform 1 0 29256 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_309
timestamp 1676037725
transform 1 0 29532 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_320
timestamp 1676037725
transform 1 0 30544 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_328
timestamp 1676037725
transform 1 0 31280 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_339
timestamp 1676037725
transform 1 0 32292 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_352
timestamp 1676037725
transform 1 0 33488 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_365
timestamp 1676037725
transform 1 0 34684 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_391
timestamp 1676037725
transform 1 0 37076 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_397
timestamp 1676037725
transform 1 0 37628 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_410
timestamp 1676037725
transform 1 0 38824 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_418
timestamp 1676037725
transform 1 0 39560 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_421
timestamp 1676037725
transform 1 0 39836 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_443
timestamp 1676037725
transform 1 0 41860 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_455
timestamp 1676037725
transform 1 0 42964 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_467
timestamp 1676037725
transform 1 0 44068 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1676037725
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_477
timestamp 1676037725
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_489
timestamp 1676037725
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_501
timestamp 1676037725
transform 1 0 47196 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_513
timestamp 1676037725
transform 1 0 48300 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_517
timestamp 1676037725
transform 1 0 48668 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_525
timestamp 1676037725
transform 1 0 49404 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1676037725
transform 1 0 1380 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_21
timestamp 1676037725
transform 1 0 3036 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_41
timestamp 1676037725
transform 1 0 4876 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_49
timestamp 1676037725
transform 1 0 5612 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1676037725
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1676037725
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1676037725
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1676037725
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_96
timestamp 1676037725
transform 1 0 9936 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_103
timestamp 1676037725
transform 1 0 10580 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_110
timestamp 1676037725
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_113
timestamp 1676037725
transform 1 0 11500 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_117
timestamp 1676037725
transform 1 0 11868 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_122
timestamp 1676037725
transform 1 0 12328 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_146
timestamp 1676037725
transform 1 0 14536 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_154
timestamp 1676037725
transform 1 0 15272 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_158
timestamp 1676037725
transform 1 0 15640 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_166
timestamp 1676037725
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_169
timestamp 1676037725
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_180
timestamp 1676037725
transform 1 0 17664 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_207
timestamp 1676037725
transform 1 0 20148 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp 1676037725
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_225
timestamp 1676037725
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_238
timestamp 1676037725
transform 1 0 23000 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_262
timestamp 1676037725
transform 1 0 25208 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_31_277
timestamp 1676037725
transform 1 0 26588 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_281
timestamp 1676037725
transform 1 0 26956 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_289
timestamp 1676037725
transform 1 0 27692 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_293
timestamp 1676037725
transform 1 0 28060 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_306
timestamp 1676037725
transform 1 0 29256 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_319
timestamp 1676037725
transform 1 0 30452 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_334
timestamp 1676037725
transform 1 0 31832 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_337
timestamp 1676037725
transform 1 0 32108 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_348
timestamp 1676037725
transform 1 0 33120 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_361
timestamp 1676037725
transform 1 0 34316 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_374
timestamp 1676037725
transform 1 0 35512 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_387
timestamp 1676037725
transform 1 0 36708 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1676037725
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_393
timestamp 1676037725
transform 1 0 37260 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_399
timestamp 1676037725
transform 1 0 37812 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_420
timestamp 1676037725
transform 1 0 39744 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_433
timestamp 1676037725
transform 1 0 40940 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_445
timestamp 1676037725
transform 1 0 42044 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_449
timestamp 1676037725
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_461
timestamp 1676037725
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_473
timestamp 1676037725
transform 1 0 44620 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_485
timestamp 1676037725
transform 1 0 45724 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_497
timestamp 1676037725
transform 1 0 46828 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1676037725
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_505
timestamp 1676037725
transform 1 0 47564 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_517
timestamp 1676037725
transform 1 0 48668 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_525
timestamp 1676037725
transform 1 0 49404 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1676037725
transform 1 0 1380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_21
timestamp 1676037725
transform 1 0 3036 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1676037725
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_29
timestamp 1676037725
transform 1 0 3772 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_47
timestamp 1676037725
transform 1 0 5428 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_67
timestamp 1676037725
transform 1 0 7268 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_71
timestamp 1676037725
transform 1 0 7636 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_75
timestamp 1676037725
transform 1 0 8004 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1676037725
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_85
timestamp 1676037725
transform 1 0 8924 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_93
timestamp 1676037725
transform 1 0 9660 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_98
timestamp 1676037725
transform 1 0 10120 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_109
timestamp 1676037725
transform 1 0 11132 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_114
timestamp 1676037725
transform 1 0 11592 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_138
timestamp 1676037725
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_141
timestamp 1676037725
transform 1 0 14076 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_147
timestamp 1676037725
transform 1 0 14628 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_151
timestamp 1676037725
transform 1 0 14996 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_158
timestamp 1676037725
transform 1 0 15640 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_181
timestamp 1676037725
transform 1 0 17756 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1676037725
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_197
timestamp 1676037725
transform 1 0 19228 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_205
timestamp 1676037725
transform 1 0 19964 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_231
timestamp 1676037725
transform 1 0 22356 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_244
timestamp 1676037725
transform 1 0 23552 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_253
timestamp 1676037725
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_258
timestamp 1676037725
transform 1 0 24840 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_32_302
timestamp 1676037725
transform 1 0 28888 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_32_309
timestamp 1676037725
transform 1 0 29532 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_314
timestamp 1676037725
transform 1 0 29992 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_327
timestamp 1676037725
transform 1 0 31188 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_340
timestamp 1676037725
transform 1 0 32384 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_348
timestamp 1676037725
transform 1 0 33120 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_360
timestamp 1676037725
transform 1 0 34224 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_365
timestamp 1676037725
transform 1 0 34684 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_376
timestamp 1676037725
transform 1 0 35696 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_389
timestamp 1676037725
transform 1 0 36892 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_397
timestamp 1676037725
transform 1 0 37628 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_408
timestamp 1676037725
transform 1 0 38640 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_415
timestamp 1676037725
transform 1 0 39284 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 1676037725
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_421
timestamp 1676037725
transform 1 0 39836 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_432
timestamp 1676037725
transform 1 0 40848 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_445
timestamp 1676037725
transform 1 0 42044 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_457
timestamp 1676037725
transform 1 0 43148 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_469
timestamp 1676037725
transform 1 0 44252 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_475
timestamp 1676037725
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_477
timestamp 1676037725
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_489
timestamp 1676037725
transform 1 0 46092 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_501
timestamp 1676037725
transform 1 0 47196 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_513
timestamp 1676037725
transform 1 0 48300 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_525
timestamp 1676037725
transform 1 0 49404 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1676037725
transform 1 0 1380 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_21
timestamp 1676037725
transform 1 0 3036 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_41
timestamp 1676037725
transform 1 0 4876 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_48
timestamp 1676037725
transform 1 0 5520 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_57
timestamp 1676037725
transform 1 0 6348 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_75
timestamp 1676037725
transform 1 0 8004 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_82
timestamp 1676037725
transform 1 0 8648 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_86
timestamp 1676037725
transform 1 0 9016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_90
timestamp 1676037725
transform 1 0 9384 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_99
timestamp 1676037725
transform 1 0 10212 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_106
timestamp 1676037725
transform 1 0 10856 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_113
timestamp 1676037725
transform 1 0 11500 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_119
timestamp 1676037725
transform 1 0 12052 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_127
timestamp 1676037725
transform 1 0 12788 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_135
timestamp 1676037725
transform 1 0 13524 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_146
timestamp 1676037725
transform 1 0 14536 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_158
timestamp 1676037725
transform 1 0 15640 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_166
timestamp 1676037725
transform 1 0 16376 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_169
timestamp 1676037725
transform 1 0 16652 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_193
timestamp 1676037725
transform 1 0 18860 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_201
timestamp 1676037725
transform 1 0 19596 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_222
timestamp 1676037725
transform 1 0 21528 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_225
timestamp 1676037725
transform 1 0 21804 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_237
timestamp 1676037725
transform 1 0 22908 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_245
timestamp 1676037725
transform 1 0 23644 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_267
timestamp 1676037725
transform 1 0 25668 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_274
timestamp 1676037725
transform 1 0 26312 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_33_281
timestamp 1676037725
transform 1 0 26956 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_304
timestamp 1676037725
transform 1 0 29072 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_317
timestamp 1676037725
transform 1 0 30268 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_330
timestamp 1676037725
transform 1 0 31464 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_337
timestamp 1676037725
transform 1 0 32108 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_359
timestamp 1676037725
transform 1 0 34132 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_372
timestamp 1676037725
transform 1 0 35328 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_389
timestamp 1676037725
transform 1 0 36892 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_393
timestamp 1676037725
transform 1 0 37260 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_397
timestamp 1676037725
transform 1 0 37628 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_418
timestamp 1676037725
transform 1 0 39560 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_431
timestamp 1676037725
transform 1 0 40756 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_443
timestamp 1676037725
transform 1 0 41860 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1676037725
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_449
timestamp 1676037725
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_461
timestamp 1676037725
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_473
timestamp 1676037725
transform 1 0 44620 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_485
timestamp 1676037725
transform 1 0 45724 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_497
timestamp 1676037725
transform 1 0 46828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1676037725
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_505
timestamp 1676037725
transform 1 0 47564 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_513
timestamp 1676037725
transform 1 0 48300 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_517
timestamp 1676037725
transform 1 0 48668 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_525
timestamp 1676037725
transform 1 0 49404 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_3
timestamp 1676037725
transform 1 0 1380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_21
timestamp 1676037725
transform 1 0 3036 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1676037725
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_29
timestamp 1676037725
transform 1 0 3772 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_47
timestamp 1676037725
transform 1 0 5428 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_67
timestamp 1676037725
transform 1 0 7268 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_34_76
timestamp 1676037725
transform 1 0 8096 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_34_85
timestamp 1676037725
transform 1 0 8924 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_96
timestamp 1676037725
transform 1 0 9936 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_103
timestamp 1676037725
transform 1 0 10580 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_110
timestamp 1676037725
transform 1 0 11224 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_34_120
timestamp 1676037725
transform 1 0 12144 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_130
timestamp 1676037725
transform 1 0 13064 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_138
timestamp 1676037725
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_141
timestamp 1676037725
transform 1 0 14076 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_163
timestamp 1676037725
transform 1 0 16100 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_170
timestamp 1676037725
transform 1 0 16744 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_194
timestamp 1676037725
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_197
timestamp 1676037725
transform 1 0 19228 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_212
timestamp 1676037725
transform 1 0 20608 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_216
timestamp 1676037725
transform 1 0 20976 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_237
timestamp 1676037725
transform 1 0 22908 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_250
timestamp 1676037725
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_253
timestamp 1676037725
transform 1 0 24380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_264
timestamp 1676037725
transform 1 0 25392 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_268
timestamp 1676037725
transform 1 0 25760 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_278
timestamp 1676037725
transform 1 0 26680 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_285
timestamp 1676037725
transform 1 0 27324 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_292
timestamp 1676037725
transform 1 0 27968 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_34_305
timestamp 1676037725
transform 1 0 29164 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_309
timestamp 1676037725
transform 1 0 29532 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_314
timestamp 1676037725
transform 1 0 29992 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_322
timestamp 1676037725
transform 1 0 30728 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_332
timestamp 1676037725
transform 1 0 31648 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_339
timestamp 1676037725
transform 1 0 32292 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_347
timestamp 1676037725
transform 1 0 33028 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_358
timestamp 1676037725
transform 1 0 34040 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_34_365
timestamp 1676037725
transform 1 0 34684 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_387
timestamp 1676037725
transform 1 0 36708 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_394
timestamp 1676037725
transform 1 0 37352 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_418
timestamp 1676037725
transform 1 0 39560 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_421
timestamp 1676037725
transform 1 0 39836 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_432
timestamp 1676037725
transform 1 0 40848 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_445
timestamp 1676037725
transform 1 0 42044 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_457
timestamp 1676037725
transform 1 0 43148 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_469
timestamp 1676037725
transform 1 0 44252 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 1676037725
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_477
timestamp 1676037725
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_489
timestamp 1676037725
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_501
timestamp 1676037725
transform 1 0 47196 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_513
timestamp 1676037725
transform 1 0 48300 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_525
timestamp 1676037725
transform 1 0 49404 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1676037725
transform 1 0 1380 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_21
timestamp 1676037725
transform 1 0 3036 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_41
timestamp 1676037725
transform 1 0 4876 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_49
timestamp 1676037725
transform 1 0 5612 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_53
timestamp 1676037725
transform 1 0 5980 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_57
timestamp 1676037725
transform 1 0 6348 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_75
timestamp 1676037725
transform 1 0 8004 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_95
timestamp 1676037725
transform 1 0 9844 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_99
timestamp 1676037725
transform 1 0 10212 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_103
timestamp 1676037725
transform 1 0 10580 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_110
timestamp 1676037725
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_113
timestamp 1676037725
transform 1 0 11500 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_119
timestamp 1676037725
transform 1 0 12052 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_124
timestamp 1676037725
transform 1 0 12512 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_128
timestamp 1676037725
transform 1 0 12880 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_138
timestamp 1676037725
transform 1 0 13800 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_166
timestamp 1676037725
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_169
timestamp 1676037725
transform 1 0 16652 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_186
timestamp 1676037725
transform 1 0 18216 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_210
timestamp 1676037725
transform 1 0 20424 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_218
timestamp 1676037725
transform 1 0 21160 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_35_225
timestamp 1676037725
transform 1 0 21804 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_231
timestamp 1676037725
transform 1 0 22356 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_253
timestamp 1676037725
transform 1 0 24380 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_266
timestamp 1676037725
transform 1 0 25576 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_274
timestamp 1676037725
transform 1 0 26312 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_278
timestamp 1676037725
transform 1 0 26680 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_281
timestamp 1676037725
transform 1 0 26956 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_292
timestamp 1676037725
transform 1 0 27968 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_305
timestamp 1676037725
transform 1 0 29164 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_318
timestamp 1676037725
transform 1 0 30360 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_331
timestamp 1676037725
transform 1 0 31556 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1676037725
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_337
timestamp 1676037725
transform 1 0 32108 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_344
timestamp 1676037725
transform 1 0 32752 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_369
timestamp 1676037725
transform 1 0 35052 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_375
timestamp 1676037725
transform 1 0 35604 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1676037725
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1676037725
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_393
timestamp 1676037725
transform 1 0 37260 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_415
timestamp 1676037725
transform 1 0 39284 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_421
timestamp 1676037725
transform 1 0 39836 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_434
timestamp 1676037725
transform 1 0 41032 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_446
timestamp 1676037725
transform 1 0 42136 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_449
timestamp 1676037725
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_461
timestamp 1676037725
transform 1 0 43516 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_473
timestamp 1676037725
transform 1 0 44620 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_485
timestamp 1676037725
transform 1 0 45724 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_497
timestamp 1676037725
transform 1 0 46828 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 1676037725
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_505
timestamp 1676037725
transform 1 0 47564 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_517
timestamp 1676037725
transform 1 0 48668 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_525
timestamp 1676037725
transform 1 0 49404 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_3
timestamp 1676037725
transform 1 0 1380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_21
timestamp 1676037725
transform 1 0 3036 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1676037725
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_29
timestamp 1676037725
transform 1 0 3772 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_47
timestamp 1676037725
transform 1 0 5428 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_67
timestamp 1676037725
transform 1 0 7268 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_75
timestamp 1676037725
transform 1 0 8004 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_82
timestamp 1676037725
transform 1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_85
timestamp 1676037725
transform 1 0 8924 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_103
timestamp 1676037725
transform 1 0 10580 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_109
timestamp 1676037725
transform 1 0 11132 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_126
timestamp 1676037725
transform 1 0 12696 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_134
timestamp 1676037725
transform 1 0 13432 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_141
timestamp 1676037725
transform 1 0 14076 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_149
timestamp 1676037725
transform 1 0 14812 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_173
timestamp 1676037725
transform 1 0 17020 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_193
timestamp 1676037725
transform 1 0 18860 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_197
timestamp 1676037725
transform 1 0 19228 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_215
timestamp 1676037725
transform 1 0 20884 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_230
timestamp 1676037725
transform 1 0 22264 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_243
timestamp 1676037725
transform 1 0 23460 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1676037725
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_253
timestamp 1676037725
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_264
timestamp 1676037725
transform 1 0 25392 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_279
timestamp 1676037725
transform 1 0 26772 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_291
timestamp 1676037725
transform 1 0 27876 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_304
timestamp 1676037725
transform 1 0 29072 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_309
timestamp 1676037725
transform 1 0 29532 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_314
timestamp 1676037725
transform 1 0 29992 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_322
timestamp 1676037725
transform 1 0 30728 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_343
timestamp 1676037725
transform 1 0 32660 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_356
timestamp 1676037725
transform 1 0 33856 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_36_365
timestamp 1676037725
transform 1 0 34684 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_371
timestamp 1676037725
transform 1 0 35236 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_381
timestamp 1676037725
transform 1 0 36156 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_388
timestamp 1676037725
transform 1 0 36800 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_392
timestamp 1676037725
transform 1 0 37168 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_414
timestamp 1676037725
transform 1 0 39192 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_36_421
timestamp 1676037725
transform 1 0 39836 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_432
timestamp 1676037725
transform 1 0 40848 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_445
timestamp 1676037725
transform 1 0 42044 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_457
timestamp 1676037725
transform 1 0 43148 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_461
timestamp 1676037725
transform 1 0 43516 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_473
timestamp 1676037725
transform 1 0 44620 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_477
timestamp 1676037725
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_489
timestamp 1676037725
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_501
timestamp 1676037725
transform 1 0 47196 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_510
timestamp 1676037725
transform 1 0 48024 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_517
timestamp 1676037725
transform 1 0 48668 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_525
timestamp 1676037725
transform 1 0 49404 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1676037725
transform 1 0 1380 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_21
timestamp 1676037725
transform 1 0 3036 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_29
timestamp 1676037725
transform 1 0 3772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_34
timestamp 1676037725
transform 1 0 4232 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_54
timestamp 1676037725
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_57
timestamp 1676037725
transform 1 0 6348 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_37_63
timestamp 1676037725
transform 1 0 6900 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_37_85
timestamp 1676037725
transform 1 0 8924 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_93
timestamp 1676037725
transform 1 0 9660 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_110
timestamp 1676037725
transform 1 0 11224 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_113
timestamp 1676037725
transform 1 0 11500 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_117
timestamp 1676037725
transform 1 0 11868 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_121
timestamp 1676037725
transform 1 0 12236 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_141
timestamp 1676037725
transform 1 0 14076 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_149
timestamp 1676037725
transform 1 0 14812 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_166
timestamp 1676037725
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_169
timestamp 1676037725
transform 1 0 16652 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_191
timestamp 1676037725
transform 1 0 18676 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_220
timestamp 1676037725
transform 1 0 21344 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_225
timestamp 1676037725
transform 1 0 21804 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_248
timestamp 1676037725
transform 1 0 23920 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_256
timestamp 1676037725
transform 1 0 24656 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_278
timestamp 1676037725
transform 1 0 26680 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_281
timestamp 1676037725
transform 1 0 26956 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_286
timestamp 1676037725
transform 1 0 27416 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_292
timestamp 1676037725
transform 1 0 27968 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_313
timestamp 1676037725
transform 1 0 29900 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_326
timestamp 1676037725
transform 1 0 31096 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_37_333
timestamp 1676037725
transform 1 0 31740 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_337
timestamp 1676037725
transform 1 0 32108 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_368
timestamp 1676037725
transform 1 0 34960 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_374
timestamp 1676037725
transform 1 0 35512 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_387
timestamp 1676037725
transform 1 0 36708 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1676037725
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_393
timestamp 1676037725
transform 1 0 37260 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_415
timestamp 1676037725
transform 1 0 39284 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_443
timestamp 1676037725
transform 1 0 41860 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 1676037725
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_449
timestamp 1676037725
transform 1 0 42412 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_454
timestamp 1676037725
transform 1 0 42872 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_468
timestamp 1676037725
transform 1 0 44160 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_477
timestamp 1676037725
transform 1 0 44988 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_489
timestamp 1676037725
transform 1 0 46092 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_497
timestamp 1676037725
transform 1 0 46828 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_502
timestamp 1676037725
transform 1 0 47288 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_505
timestamp 1676037725
transform 1 0 47564 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_517
timestamp 1676037725
transform 1 0 48668 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_525
timestamp 1676037725
transform 1 0 49404 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_3
timestamp 1676037725
transform 1 0 1380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_21
timestamp 1676037725
transform 1 0 3036 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1676037725
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_38_29
timestamp 1676037725
transform 1 0 3772 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_35
timestamp 1676037725
transform 1 0 4324 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_42
timestamp 1676037725
transform 1 0 4968 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_62
timestamp 1676037725
transform 1 0 6808 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_82
timestamp 1676037725
transform 1 0 8648 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_85
timestamp 1676037725
transform 1 0 8924 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_91
timestamp 1676037725
transform 1 0 9476 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_98
timestamp 1676037725
transform 1 0 10120 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_118
timestamp 1676037725
transform 1 0 11960 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_138
timestamp 1676037725
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_141
timestamp 1676037725
transform 1 0 14076 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_150
timestamp 1676037725
transform 1 0 14904 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_170
timestamp 1676037725
transform 1 0 16744 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_194
timestamp 1676037725
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_197
timestamp 1676037725
transform 1 0 19228 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_205
timestamp 1676037725
transform 1 0 19964 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_229
timestamp 1676037725
transform 1 0 22172 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_233
timestamp 1676037725
transform 1 0 22540 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_237
timestamp 1676037725
transform 1 0 22908 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_250
timestamp 1676037725
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_253
timestamp 1676037725
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_259
timestamp 1676037725
transform 1 0 24932 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_287
timestamp 1676037725
transform 1 0 27508 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_300
timestamp 1676037725
transform 1 0 28704 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_309
timestamp 1676037725
transform 1 0 29532 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_320
timestamp 1676037725
transform 1 0 30544 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_328
timestamp 1676037725
transform 1 0 31280 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_350
timestamp 1676037725
transform 1 0 33304 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1676037725
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1676037725
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_365
timestamp 1676037725
transform 1 0 34684 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_389
timestamp 1676037725
transform 1 0 36892 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_413
timestamp 1676037725
transform 1 0 39100 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1676037725
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_421
timestamp 1676037725
transform 1 0 39836 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_432
timestamp 1676037725
transform 1 0 40848 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_473
timestamp 1676037725
transform 1 0 44620 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_484
timestamp 1676037725
transform 1 0 45632 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_488
timestamp 1676037725
transform 1 0 46000 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_492
timestamp 1676037725
transform 1 0 46368 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_498
timestamp 1676037725
transform 1 0 46920 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_502
timestamp 1676037725
transform 1 0 47288 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_509
timestamp 1676037725
transform 1 0 47932 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_517
timestamp 1676037725
transform 1 0 48668 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_525
timestamp 1676037725
transform 1 0 49404 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1676037725
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_15
timestamp 1676037725
transform 1 0 2484 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_34
timestamp 1676037725
transform 1 0 4232 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_54
timestamp 1676037725
transform 1 0 6072 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_57
timestamp 1676037725
transform 1 0 6348 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_62
timestamp 1676037725
transform 1 0 6808 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_66
timestamp 1676037725
transform 1 0 7176 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_70
timestamp 1676037725
transform 1 0 7544 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_90
timestamp 1676037725
transform 1 0 9384 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_110
timestamp 1676037725
transform 1 0 11224 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_113
timestamp 1676037725
transform 1 0 11500 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_126
timestamp 1676037725
transform 1 0 12696 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_148
timestamp 1676037725
transform 1 0 14720 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_166
timestamp 1676037725
transform 1 0 16376 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_169
timestamp 1676037725
transform 1 0 16652 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_188
timestamp 1676037725
transform 1 0 18400 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_212
timestamp 1676037725
transform 1 0 20608 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_218
timestamp 1676037725
transform 1 0 21160 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_222
timestamp 1676037725
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_225
timestamp 1676037725
transform 1 0 21804 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_242
timestamp 1676037725
transform 1 0 23368 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_250
timestamp 1676037725
transform 1 0 24104 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_278
timestamp 1676037725
transform 1 0 26680 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_281
timestamp 1676037725
transform 1 0 26956 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_287
timestamp 1676037725
transform 1 0 27508 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_294
timestamp 1676037725
transform 1 0 28152 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_301
timestamp 1676037725
transform 1 0 28796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_308
timestamp 1676037725
transform 1 0 29440 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_39_334
timestamp 1676037725
transform 1 0 31832 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_337
timestamp 1676037725
transform 1 0 32108 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_348
timestamp 1676037725
transform 1 0 33120 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_352
timestamp 1676037725
transform 1 0 33488 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_373
timestamp 1676037725
transform 1 0 35420 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_379
timestamp 1676037725
transform 1 0 35972 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_39_389
timestamp 1676037725
transform 1 0 36892 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_393
timestamp 1676037725
transform 1 0 37260 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_404
timestamp 1676037725
transform 1 0 38272 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_426
timestamp 1676037725
transform 1 0 40296 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_444
timestamp 1676037725
transform 1 0 41952 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_449
timestamp 1676037725
transform 1 0 42412 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_457
timestamp 1676037725
transform 1 0 43148 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_463
timestamp 1676037725
transform 1 0 43700 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_477
timestamp 1676037725
transform 1 0 44988 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_489
timestamp 1676037725
transform 1 0 46092 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_495
timestamp 1676037725
transform 1 0 46644 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_500
timestamp 1676037725
transform 1 0 47104 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_505
timestamp 1676037725
transform 1 0 47564 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_509
timestamp 1676037725
transform 1 0 47932 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_514
timestamp 1676037725
transform 1 0 48392 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_522
timestamp 1676037725
transform 1 0 49128 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_526
timestamp 1676037725
transform 1 0 49496 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_3
timestamp 1676037725
transform 1 0 1380 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_9
timestamp 1676037725
transform 1 0 1932 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_26
timestamp 1676037725
transform 1 0 3496 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_29
timestamp 1676037725
transform 1 0 3772 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_34
timestamp 1676037725
transform 1 0 4232 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_54
timestamp 1676037725
transform 1 0 6072 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_57
timestamp 1676037725
transform 1 0 6348 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_62
timestamp 1676037725
transform 1 0 6808 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_82
timestamp 1676037725
transform 1 0 8648 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_85
timestamp 1676037725
transform 1 0 8924 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_90
timestamp 1676037725
transform 1 0 9384 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_110
timestamp 1676037725
transform 1 0 11224 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_113
timestamp 1676037725
transform 1 0 11500 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_118
timestamp 1676037725
transform 1 0 11960 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_138
timestamp 1676037725
transform 1 0 13800 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_141
timestamp 1676037725
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_146
timestamp 1676037725
transform 1 0 14536 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_166
timestamp 1676037725
transform 1 0 16376 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_169
timestamp 1676037725
transform 1 0 16652 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_174
timestamp 1676037725
transform 1 0 17112 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_194
timestamp 1676037725
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_197
timestamp 1676037725
transform 1 0 19228 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_202
timestamp 1676037725
transform 1 0 19688 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_222
timestamp 1676037725
transform 1 0 21528 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_225
timestamp 1676037725
transform 1 0 21804 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_243
timestamp 1676037725
transform 1 0 23460 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_250
timestamp 1676037725
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_253
timestamp 1676037725
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_264
timestamp 1676037725
transform 1 0 25392 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_270
timestamp 1676037725
transform 1 0 25944 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_275
timestamp 1676037725
transform 1 0 26404 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_279
timestamp 1676037725
transform 1 0 26772 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_281
timestamp 1676037725
transform 1 0 26956 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_287
timestamp 1676037725
transform 1 0 27508 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_294
timestamp 1676037725
transform 1 0 28152 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1676037725
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1676037725
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_309
timestamp 1676037725
transform 1 0 29532 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_314
timestamp 1676037725
transform 1 0 29992 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_321
timestamp 1676037725
transform 1 0 30636 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_328
timestamp 1676037725
transform 1 0 31280 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_337
timestamp 1676037725
transform 1 0 32108 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_342
timestamp 1676037725
transform 1 0 32568 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_349
timestamp 1676037725
transform 1 0 33212 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_362
timestamp 1676037725
transform 1 0 34408 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_365
timestamp 1676037725
transform 1 0 34684 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_370
timestamp 1676037725
transform 1 0 35144 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_387
timestamp 1676037725
transform 1 0 36708 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_391
timestamp 1676037725
transform 1 0 37076 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_393
timestamp 1676037725
transform 1 0 37260 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_404
timestamp 1676037725
transform 1 0 38272 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_412
timestamp 1676037725
transform 1 0 39008 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_416
timestamp 1676037725
transform 1 0 39376 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_421
timestamp 1676037725
transform 1 0 39836 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_426
timestamp 1676037725
transform 1 0 40296 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_433
timestamp 1676037725
transform 1 0 40940 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_442
timestamp 1676037725
transform 1 0 41768 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_40_449
timestamp 1676037725
transform 1 0 42412 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_471
timestamp 1676037725
transform 1 0 44436 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 1676037725
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_477
timestamp 1676037725
transform 1 0 44988 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_483
timestamp 1676037725
transform 1 0 45540 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_491
timestamp 1676037725
transform 1 0 46276 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_499
timestamp 1676037725
transform 1 0 47012 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_503
timestamp 1676037725
transform 1 0 47380 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_505
timestamp 1676037725
transform 1 0 47564 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_525
timestamp 1676037725
transform 1 0 49404 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1676037725
transform 1 0 9660 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1676037725
transform 1 0 47012 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1676037725
transform 1 0 3036 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input4 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1564 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input5
timestamp 1676037725
transform 1 0 1564 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1676037725
transform 1 0 2300 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1676037725
transform 1 0 1564 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input8
timestamp 1676037725
transform 1 0 1564 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input9
timestamp 1676037725
transform 1 0 1564 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input10
timestamp 1676037725
transform 1 0 1564 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input11
timestamp 1676037725
transform 1 0 2300 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input12
timestamp 1676037725
transform 1 0 1564 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input13
timestamp 1676037725
transform 1 0 1564 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp 1676037725
transform 1 0 2300 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input15
timestamp 1676037725
transform 1 0 1564 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input16
timestamp 1676037725
transform 1 0 2300 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input17
timestamp 1676037725
transform 1 0 1564 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input18
timestamp 1676037725
transform 1 0 1564 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1676037725
transform 1 0 2300 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input20
timestamp 1676037725
transform 1 0 1564 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input21
timestamp 1676037725
transform 1 0 1564 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1676037725
transform 1 0 2852 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input23
timestamp 1676037725
transform 1 0 1564 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input24
timestamp 1676037725
transform 1 0 3404 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input25
timestamp 1676037725
transform 1 0 1564 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input26
timestamp 1676037725
transform 1 0 1564 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input27
timestamp 1676037725
transform 1 0 1564 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input28
timestamp 1676037725
transform 1 0 2300 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input29
timestamp 1676037725
transform 1 0 1564 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input30
timestamp 1676037725
transform 1 0 1564 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input31
timestamp 1676037725
transform 1 0 1564 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input32
timestamp 1676037725
transform 1 0 2300 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1676037725
transform 1 0 48392 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input34
timestamp 1676037725
transform 1 0 49036 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input35
timestamp 1676037725
transform 1 0 49036 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1676037725
transform 1 0 48392 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input37
timestamp 1676037725
transform 1 0 49036 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1676037725
transform 1 0 49036 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input39
timestamp 1676037725
transform 1 0 49036 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1676037725
transform 1 0 48392 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input41
timestamp 1676037725
transform 1 0 49036 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input42
timestamp 1676037725
transform 1 0 49036 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input43
timestamp 1676037725
transform 1 0 49036 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input44
timestamp 1676037725
transform 1 0 49036 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1676037725
transform 1 0 48392 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input46
timestamp 1676037725
transform 1 0 49036 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input47
timestamp 1676037725
transform 1 0 49036 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input48
timestamp 1676037725
transform 1 0 48300 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1676037725
transform 1 0 47656 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1676037725
transform 1 0 46092 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input51
timestamp 1676037725
transform 1 0 48300 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1676037725
transform 1 0 47748 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1676037725
transform 1 0 47012 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input54
timestamp 1676037725
transform 1 0 48484 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input55
timestamp 1676037725
transform 1 0 49036 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input56
timestamp 1676037725
transform 1 0 49036 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1676037725
transform 1 0 49128 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input58
timestamp 1676037725
transform 1 0 49036 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input59
timestamp 1676037725
transform 1 0 49036 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input60
timestamp 1676037725
transform 1 0 49036 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1676037725
transform 1 0 48392 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input62
timestamp 1676037725
transform 1 0 49036 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1676037725
transform 1 0 27048 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1676037725
transform 1 0 29716 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1676037725
transform 1 0 32292 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1676037725
transform 1 0 34868 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input67
timestamp 1676037725
transform 1 0 36524 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input68
timestamp 1676037725
transform 1 0 33672 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input69
timestamp 1676037725
transform 1 0 32016 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input70
timestamp 1676037725
transform 1 0 40020 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input71
timestamp 1676037725
transform 1 0 40664 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input72
timestamp 1676037725
transform 1 0 41492 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input73
timestamp 1676037725
transform 1 0 43700 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input74
timestamp 1676037725
transform 1 0 11776 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input75
timestamp 1676037725
transform 1 0 43240 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input76
timestamp 1676037725
transform 1 0 41032 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input77
timestamp 1676037725
transform 1 0 44068 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input78
timestamp 1676037725
transform 1 0 45172 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input79
timestamp 1676037725
transform 1 0 42596 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input80
timestamp 1676037725
transform 1 0 41308 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input81
timestamp 1676037725
transform 1 0 45356 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input82
timestamp 1676037725
transform 1 0 41584 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input83
timestamp 1676037725
transform 1 0 44712 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input84
timestamp 1676037725
transform 1 0 43240 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input85
timestamp 1676037725
transform 1 0 26036 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input86
timestamp 1676037725
transform 1 0 11776 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input87
timestamp 1676037725
transform 1 0 32936 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input88
timestamp 1676037725
transform 1 0 31004 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input89
timestamp 1676037725
transform 1 0 23828 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input90
timestamp 1676037725
transform 1 0 28520 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input91
timestamp 1676037725
transform 1 0 27876 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input92
timestamp 1676037725
transform 1 0 28520 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input93
timestamp 1676037725
transform 1 0 28980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input94
timestamp 1676037725
transform 1 0 30820 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input95
timestamp 1676037725
transform 1 0 32936 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input96
timestamp 1676037725
transform 1 0 35052 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input97
timestamp 1676037725
transform 1 0 37444 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_16  input98
timestamp 1676037725
transform 1 0 42596 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input99
timestamp 1676037725
transform 1 0 43516 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input100
timestamp 1676037725
transform 1 0 45356 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input101
timestamp 1676037725
transform 1 0 47196 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input102
timestamp 1676037725
transform 1 0 46460 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input103
timestamp 1676037725
transform 1 0 45908 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input104
timestamp 1676037725
transform 1 0 46644 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input105
timestamp 1676037725
transform 1 0 46736 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input106
timestamp 1676037725
transform 1 0 48116 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input107
timestamp 1676037725
transform 1 0 48024 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input108
timestamp 1676037725
transform 1 0 48760 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input109
timestamp 1676037725
transform 1 0 44988 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input110
timestamp 1676037725
transform 1 0 45172 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_12  output111 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 40664 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output112
timestamp 1676037725
transform 1 0 3404 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output113
timestamp 1676037725
transform 1 0 1564 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output114
timestamp 1676037725
transform 1 0 1564 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output115
timestamp 1676037725
transform 1 0 1564 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output116
timestamp 1676037725
transform 1 0 1564 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output117
timestamp 1676037725
transform 1 0 1564 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output118
timestamp 1676037725
transform 1 0 1564 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output119
timestamp 1676037725
transform 1 0 1564 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output120
timestamp 1676037725
transform 1 0 3404 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output121
timestamp 1676037725
transform 1 0 1564 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output122
timestamp 1676037725
transform 1 0 1564 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output123
timestamp 1676037725
transform 1 0 1564 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output124
timestamp 1676037725
transform 1 0 1564 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output125
timestamp 1676037725
transform 1 0 3956 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output126
timestamp 1676037725
transform 1 0 3956 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output127
timestamp 1676037725
transform 1 0 5796 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output128
timestamp 1676037725
transform 1 0 5796 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output129
timestamp 1676037725
transform 1 0 6532 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output130
timestamp 1676037725
transform 1 0 3956 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output131
timestamp 1676037725
transform 1 0 5796 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output132
timestamp 1676037725
transform 1 0 6532 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output133
timestamp 1676037725
transform 1 0 8372 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output134
timestamp 1676037725
transform 1 0 9108 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output135
timestamp 1676037725
transform 1 0 1564 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output136
timestamp 1676037725
transform 1 0 1564 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output137
timestamp 1676037725
transform 1 0 1564 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output138
timestamp 1676037725
transform 1 0 1564 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output139
timestamp 1676037725
transform 1 0 1564 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output140
timestamp 1676037725
transform 1 0 1564 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output141
timestamp 1676037725
transform 1 0 1564 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output142
timestamp 1676037725
transform 1 0 1564 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output143
timestamp 1676037725
transform 1 0 45816 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output144
timestamp 1676037725
transform 1 0 47932 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output145
timestamp 1676037725
transform 1 0 47932 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output146
timestamp 1676037725
transform 1 0 46092 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output147
timestamp 1676037725
transform 1 0 47932 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output148
timestamp 1676037725
transform 1 0 47932 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output149
timestamp 1676037725
transform 1 0 47932 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output150
timestamp 1676037725
transform 1 0 45816 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output151
timestamp 1676037725
transform 1 0 47932 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output152
timestamp 1676037725
transform 1 0 47932 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output153
timestamp 1676037725
transform 1 0 47932 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output154
timestamp 1676037725
transform 1 0 43976 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output155
timestamp 1676037725
transform 1 0 46092 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output156
timestamp 1676037725
transform 1 0 47932 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output157
timestamp 1676037725
transform 1 0 47932 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output158
timestamp 1676037725
transform 1 0 47932 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output159
timestamp 1676037725
transform 1 0 47932 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output160
timestamp 1676037725
transform 1 0 47932 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output161
timestamp 1676037725
transform 1 0 47932 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output162
timestamp 1676037725
transform 1 0 47932 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output163
timestamp 1676037725
transform 1 0 47932 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output164
timestamp 1676037725
transform 1 0 47932 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output165
timestamp 1676037725
transform 1 0 45816 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output166
timestamp 1676037725
transform 1 0 45816 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output167
timestamp 1676037725
transform 1 0 46092 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output168
timestamp 1676037725
transform 1 0 47932 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output169
timestamp 1676037725
transform 1 0 47932 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output170
timestamp 1676037725
transform 1 0 47932 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output171
timestamp 1676037725
transform 1 0 45816 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output172
timestamp 1676037725
transform 1 0 47932 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output173
timestamp 1676037725
transform 1 0 3956 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output174
timestamp 1676037725
transform 1 0 7176 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output175
timestamp 1676037725
transform 1 0 7912 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output176
timestamp 1676037725
transform 1 0 9752 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output177
timestamp 1676037725
transform 1 0 9752 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output178
timestamp 1676037725
transform 1 0 10488 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output179
timestamp 1676037725
transform 1 0 9752 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output180
timestamp 1676037725
transform 1 0 12604 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output181
timestamp 1676037725
transform 1 0 12328 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output182
timestamp 1676037725
transform 1 0 12328 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output183
timestamp 1676037725
transform 1 0 13248 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output184
timestamp 1676037725
transform 1 0 3404 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output185
timestamp 1676037725
transform 1 0 14904 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output186
timestamp 1676037725
transform 1 0 15272 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output187
timestamp 1676037725
transform 1 0 14904 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output188
timestamp 1676037725
transform 1 0 17388 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output189
timestamp 1676037725
transform 1 0 14904 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output190
timestamp 1676037725
transform 1 0 16928 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output191
timestamp 1676037725
transform 1 0 19412 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output192
timestamp 1676037725
transform 1 0 17480 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output193
timestamp 1676037725
transform 1 0 21988 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output194
timestamp 1676037725
transform 1 0 20056 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output195
timestamp 1676037725
transform 1 0 2024 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output196
timestamp 1676037725
transform 1 0 2760 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output197
timestamp 1676037725
transform 1 0 4600 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output198
timestamp 1676037725
transform 1 0 4600 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output199
timestamp 1676037725
transform 1 0 5336 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output200
timestamp 1676037725
transform 1 0 4600 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output201
timestamp 1676037725
transform 1 0 7452 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output202
timestamp 1676037725
transform 1 0 7176 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output203
timestamp 1676037725
transform 1 0 11776 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output204
timestamp 1676037725
transform 1 0 14260 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output205
timestamp 1676037725
transform 1 0 16836 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output206
timestamp 1676037725
transform 1 0 18124 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output207
timestamp 1676037725
transform 1 0 20056 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output208
timestamp 1676037725
transform 1 0 22356 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output209
timestamp 1676037725
transform 1 0 24564 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output210
timestamp 1676037725
transform 1 0 27140 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 49864 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 49864 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 49864 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 49864 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 49864 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 49864 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 49864 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 49864 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 49864 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 49864 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 49864 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1676037725
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1676037725
transform -1 0 49864 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1676037725
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1676037725
transform -1 0 49864 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1676037725
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1676037725
transform -1 0 49864 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1676037725
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1676037725
transform -1 0 49864 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1676037725
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1676037725
transform -1 0 49864 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1676037725
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1676037725
transform -1 0 49864 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1676037725
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1676037725
transform -1 0 49864 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1676037725
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1676037725
transform -1 0 49864 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1676037725
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1676037725
transform -1 0 49864 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1676037725
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1676037725
transform -1 0 49864 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1676037725
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1676037725
transform -1 0 49864 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1676037725
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1676037725
transform -1 0 49864 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1676037725
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1676037725
transform -1 0 49864 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1676037725
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1676037725
transform -1 0 49864 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1676037725
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1676037725
transform -1 0 49864 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1676037725
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1676037725
transform -1 0 49864 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1676037725
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1676037725
transform -1 0 49864 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1676037725
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1676037725
transform -1 0 49864 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1676037725
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1676037725
transform -1 0 49864 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1676037725
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1676037725
transform -1 0 49864 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1676037725
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1676037725
transform -1 0 49864 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1676037725
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1676037725
transform -1 0 49864 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1676037725
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1676037725
transform -1 0 49864 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1676037725
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1676037725
transform -1 0 49864 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1676037725
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1676037725
transform -1 0 49864 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1676037725
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1676037725
transform -1 0 49864 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1676037725
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1676037725
transform -1 0 49864 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1676037725
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1676037725
transform -1 0 49864 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1676037725
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1676037725
transform -1 0 49864 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1676037725
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1676037725
transform -1 0 49864 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  sb_1__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 26772 0 1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 24104 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 22724 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22264 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 20516 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 17020 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 18584 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 20240 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 17112 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19136 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 21988 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 19688 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21068 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 20976 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 19228 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19596 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19688 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 17112 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19412 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 20332 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 18768 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21988 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 23828 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 23368 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 25760 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 27048 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 25576 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 27232 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 28060 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 24840 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 25668 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 24840 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 21068 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22448 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 28520 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 30452 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 32292 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 32292 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 34868 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 35052 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 34868 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 36340 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_1__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 37444 0 1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 34868 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 35144 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_1__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 35788 0 1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 33856 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 34868 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 33764 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 32292 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 32108 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 31004 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 27968 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 29716 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 28428 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 26956 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 28796 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 30360 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 31096 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 32292 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 30728 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 29716 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 27508 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 26864 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_1__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 41584 0 1 22848
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 30820 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 29992 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 31372 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 33120 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 33580 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 35052 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 34868 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 32292 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 33120 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 37444 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 37260 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 37260 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 37444 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 37720 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 37720 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 35788 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 33580 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 35236 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 37904 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 38088 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 40020 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 38916 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 37720 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 38180 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 40020 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 37720 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 37444 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 37076 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 32292 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 29348 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 25024 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_22.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 24840 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_22.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 24012 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_24.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 24564 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_24.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 23920 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_26.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 24564 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_26.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 24564 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 23644 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22264 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21988 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19688 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19412 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19412 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19320 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 20240 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21988 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 20424 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_40.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 16836 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_40.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 12972 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 12880 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 14260 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 14260 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 12696 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11684 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 10580 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11960 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 14260 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 14536 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 15180 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_58.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 16836 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_58.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 17112 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_1.mux_l1_in_0_
timestamp 1676037725
transform 1 0 30728 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_1.mux_l1_in_1_
timestamp 1676037725
transform 1 0 27232 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_1.mux_l1_in_2_
timestamp 1676037725
transform 1 0 22632 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_1.mux_l1_in_3__258
timestamp 1676037725
transform 1 0 26036 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_1.mux_l1_in_3_
timestamp 1676037725
transform 1 0 22080 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_1.mux_l2_in_0_
timestamp 1676037725
transform 1 0 25852 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_1.mux_l2_in_1_
timestamp 1676037725
transform 1 0 22908 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_1.mux_l3_in_0_
timestamp 1676037725
transform 1 0 22080 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 17204 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_3.mux_l1_in_0_
timestamp 1676037725
transform 1 0 27048 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_3.mux_l1_in_1_
timestamp 1676037725
transform 1 0 24564 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_3.mux_l2_in_0_
timestamp 1676037725
transform 1 0 21436 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_3.mux_l2_in_1_
timestamp 1676037725
transform 1 0 17940 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_3.mux_l2_in_1__211
timestamp 1676037725
transform 1 0 16560 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_3.mux_l3_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 10580 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_5.mux_l1_in_0_
timestamp 1676037725
transform 1 0 25852 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_5.mux_l1_in_1_
timestamp 1676037725
transform 1 0 25208 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_5.mux_l2_in_0_
timestamp 1676037725
transform 1 0 21068 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_5.mux_l2_in_1__214
timestamp 1676037725
transform 1 0 19412 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_5.mux_l2_in_1_
timestamp 1676037725
transform 1 0 18308 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_5.mux_l3_in_0_
timestamp 1676037725
transform 1 0 17388 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 10948 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_7.mux_l1_in_0_
timestamp 1676037725
transform 1 0 27140 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_7.mux_l1_in_1_
timestamp 1676037725
transform 1 0 24656 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_7.mux_l1_in_2_
timestamp 1676037725
transform 1 0 19504 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_7.mux_l2_in_0_
timestamp 1676037725
transform 1 0 23092 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_7.mux_l2_in_1_
timestamp 1676037725
transform 1 0 19688 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_7.mux_l2_in_1__216
timestamp 1676037725
transform 1 0 18676 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_7.mux_l3_in_0_
timestamp 1676037725
transform 1 0 19872 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 16836 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_11.mux_l1_in_0_
timestamp 1676037725
transform 1 0 28060 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_11.mux_l1_in_1_
timestamp 1676037725
transform 1 0 25760 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_11.mux_l1_in_2_
timestamp 1676037725
transform 1 0 20884 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_11.mux_l1_in_3__259
timestamp 1676037725
transform 1 0 21988 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_11.mux_l1_in_3_
timestamp 1676037725
transform 1 0 20792 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_11.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24656 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_11.mux_l2_in_1_
timestamp 1676037725
transform 1 0 19504 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_11.mux_l3_in_0_
timestamp 1676037725
transform 1 0 18216 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 12328 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_13.mux_l1_in_0_
timestamp 1676037725
transform 1 0 27140 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_13.mux_l1_in_1_
timestamp 1676037725
transform 1 0 24748 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_13.mux_l1_in_2_
timestamp 1676037725
transform 1 0 21160 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_13.mux_l2_in_0_
timestamp 1676037725
transform 1 0 23276 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_13.mux_l2_in_1__260
timestamp 1676037725
transform 1 0 15364 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_13.mux_l2_in_1_
timestamp 1676037725
transform 1 0 19780 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_13.mux_l3_in_0_
timestamp 1676037725
transform 1 0 18124 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 11868 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_21.mux_l1_in_0_
timestamp 1676037725
transform 1 0 27876 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_21.mux_l1_in_1_
timestamp 1676037725
transform 1 0 24564 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_21.mux_l1_in_2_
timestamp 1676037725
transform 1 0 21988 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_21.mux_l2_in_0_
timestamp 1676037725
transform 1 0 22540 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_21.mux_l2_in_1__261
timestamp 1676037725
transform 1 0 16836 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_21.mux_l2_in_1_
timestamp 1676037725
transform 1 0 19780 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_21.mux_l3_in_0_
timestamp 1676037725
transform 1 0 17388 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 9844 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_29.mux_l1_in_0_
timestamp 1676037725
transform 1 0 29532 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_29.mux_l1_in_1_
timestamp 1676037725
transform 1 0 26404 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_29.mux_l1_in_2_
timestamp 1676037725
transform 1 0 24104 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_29.mux_l2_in_0_
timestamp 1676037725
transform 1 0 25576 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_29.mux_l2_in_1_
timestamp 1676037725
transform 1 0 23276 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_29.mux_l2_in_1__262
timestamp 1676037725
transform 1 0 24564 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_29.mux_l3_in_0_
timestamp 1676037725
transform 1 0 22724 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 15180 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_37.mux_l1_in_0_
timestamp 1676037725
transform 1 0 31556 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_37.mux_l1_in_1_
timestamp 1676037725
transform 1 0 29624 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_37.mux_l2_in_0_
timestamp 1676037725
transform 1 0 28520 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_37.mux_l2_in_1_
timestamp 1676037725
transform 1 0 25116 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_37.mux_l2_in_1__212
timestamp 1676037725
transform 1 0 23828 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_37.mux_l3_in_0_
timestamp 1676037725
transform 1 0 23276 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18400 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_45.mux_l1_in_0_
timestamp 1676037725
transform 1 0 32292 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_45.mux_l2_in_0_
timestamp 1676037725
transform 1 0 28244 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_45.mux_l2_in_1_
timestamp 1676037725
transform 1 0 28336 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_45.mux_l2_in_1__213
timestamp 1676037725
transform 1 0 27692 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_45.mux_l3_in_0_
timestamp 1676037725
transform 1 0 23276 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_45.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 10948 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_53.mux_l1_in_0_
timestamp 1676037725
transform 1 0 30268 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_53.mux_l2_in_0_
timestamp 1676037725
transform 1 0 25944 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_53.mux_l2_in_1_
timestamp 1676037725
transform 1 0 22632 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_53.mux_l2_in_1__215
timestamp 1676037725
transform 1 0 24564 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_53.mux_l3_in_0_
timestamp 1676037725
transform 1 0 20700 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_53.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 16468 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_0.mux_l1_in_0_
timestamp 1676037725
transform 1 0 29440 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_0.mux_l1_in_1_
timestamp 1676037725
transform 1 0 33304 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_0.mux_l1_in_2_
timestamp 1676037725
transform 1 0 27784 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_0.mux_l2_in_0_
timestamp 1676037725
transform 1 0 31004 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_0.mux_l2_in_1__217
timestamp 1676037725
transform 1 0 29808 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_0.mux_l2_in_1_
timestamp 1676037725
transform 1 0 29716 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_0.mux_l3_in_0_
timestamp 1676037725
transform 1 0 33488 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 39284 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_2.mux_l1_in_0_
timestamp 1676037725
transform 1 0 33212 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_2.mux_l1_in_1_
timestamp 1676037725
transform 1 0 32292 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_2.mux_l1_in_2_
timestamp 1676037725
transform 1 0 28336 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_2.mux_l2_in_0_
timestamp 1676037725
transform 1 0 35788 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_2.mux_l2_in_1__220
timestamp 1676037725
transform 1 0 33856 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_2.mux_l2_in_1_
timestamp 1676037725
transform 1 0 33488 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_2.mux_l3_in_0_
timestamp 1676037725
transform 1 0 37996 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 40848 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_4.mux_l1_in_0_
timestamp 1676037725
transform 1 0 35696 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_4.mux_l1_in_1_
timestamp 1676037725
transform 1 0 32752 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_4.mux_l1_in_2_
timestamp 1676037725
transform 1 0 30728 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_4.mux_l2_in_0_
timestamp 1676037725
transform 1 0 36248 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_4.mux_l2_in_1_
timestamp 1676037725
transform 1 0 35696 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_4.mux_l2_in_1__224
timestamp 1676037725
transform 1 0 31556 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_4.mux_l3_in_0_
timestamp 1676037725
transform 1 0 37444 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 41308 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_6.mux_l1_in_0_
timestamp 1676037725
transform 1 0 34868 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_6.mux_l1_in_1_
timestamp 1676037725
transform 1 0 33396 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_6.mux_l1_in_2_
timestamp 1676037725
transform 1 0 36064 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_6.mux_l1_in_3__227
timestamp 1676037725
transform 1 0 33764 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_6.mux_l1_in_3_
timestamp 1676037725
transform 1 0 32292 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_6.mux_l2_in_0_
timestamp 1676037725
transform 1 0 35880 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_6.mux_l2_in_1_
timestamp 1676037725
transform 1 0 38088 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_6.mux_l3_in_0_
timestamp 1676037725
transform 1 0 37260 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 41216 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_10.mux_l1_in_0_
timestamp 1676037725
transform 1 0 33396 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_10.mux_l1_in_1_
timestamp 1676037725
transform 1 0 32660 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_10.mux_l1_in_2_
timestamp 1676037725
transform 1 0 33304 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_10.mux_l1_in_3_
timestamp 1676037725
transform 1 0 31004 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_10.mux_l1_in_3__218
timestamp 1676037725
transform 1 0 30912 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_10.mux_l2_in_0_
timestamp 1676037725
transform 1 0 34500 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_10.mux_l2_in_1_
timestamp 1676037725
transform 1 0 37444 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_10.mux_l3_in_0_
timestamp 1676037725
transform 1 0 37444 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 40756 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_12.mux_l1_in_0_
timestamp 1676037725
transform 1 0 32292 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_12.mux_l1_in_1_
timestamp 1676037725
transform 1 0 32292 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_12.mux_l1_in_2_
timestamp 1676037725
transform 1 0 27140 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_12.mux_l2_in_0_
timestamp 1676037725
transform 1 0 32292 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_12.mux_l2_in_1_
timestamp 1676037725
transform 1 0 32292 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_12.mux_l2_in_1__219
timestamp 1676037725
transform 1 0 31372 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_12.mux_l3_in_0_
timestamp 1676037725
transform 1 0 35880 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 40204 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_20.mux_l1_in_0_
timestamp 1676037725
transform 1 0 30636 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_20.mux_l1_in_1_
timestamp 1676037725
transform 1 0 29808 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_20.mux_l1_in_2_
timestamp 1676037725
transform 1 0 27140 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_20.mux_l2_in_0_
timestamp 1676037725
transform 1 0 30636 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_20.mux_l2_in_1_
timestamp 1676037725
transform 1 0 30176 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_20.mux_l2_in_1__221
timestamp 1676037725
transform 1 0 27324 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_20.mux_l3_in_0_
timestamp 1676037725
transform 1 0 32200 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 38272 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_28.mux_l1_in_0_
timestamp 1676037725
transform 1 0 29716 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_28.mux_l1_in_1_
timestamp 1676037725
transform 1 0 29716 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_28.mux_l1_in_2_
timestamp 1676037725
transform 1 0 25668 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_28.mux_l2_in_0_
timestamp 1676037725
transform 1 0 29716 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_28.mux_l2_in_1_
timestamp 1676037725
transform 1 0 30176 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_28.mux_l2_in_1__222
timestamp 1676037725
transform 1 0 29716 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_28.mux_l3_in_0_
timestamp 1676037725
transform 1 0 32568 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 37628 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_36.mux_l1_in_0_
timestamp 1676037725
transform 1 0 31556 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_36.mux_l1_in_1_
timestamp 1676037725
transform 1 0 31004 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_36.mux_l2_in_0_
timestamp 1676037725
transform 1 0 33304 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_36.mux_l2_in_1__223
timestamp 1676037725
transform 1 0 29716 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_36.mux_l2_in_1_
timestamp 1676037725
transform 1 0 30544 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_36.mux_l3_in_0_
timestamp 1676037725
transform 1 0 34868 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 38916 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_44.mux_l1_in_0_
timestamp 1676037725
transform 1 0 29716 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_44.mux_l1_in_1__225
timestamp 1676037725
transform 1 0 29716 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_44.mux_l1_in_1_
timestamp 1676037725
transform 1 0 28152 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_44.mux_l2_in_0_
timestamp 1676037725
transform 1 0 32568 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_44.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 37444 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_52.mux_l1_in_0_
timestamp 1676037725
transform 1 0 28704 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_52.mux_l1_in_1_
timestamp 1676037725
transform 1 0 26956 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_52.mux_l1_in_1__226
timestamp 1676037725
transform 1 0 26404 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_52.mux_l2_in_0_
timestamp 1676037725
transform 1 0 29716 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_52.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 36616 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_0.mux_l1_in_0_
timestamp 1676037725
transform 1 0 35880 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_0.mux_l1_in_1_
timestamp 1676037725
transform 1 0 40480 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_0.mux_l1_in_2_
timestamp 1676037725
transform 1 0 24564 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_0.mux_l1_in_3__228
timestamp 1676037725
transform 1 0 29716 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_0.mux_l1_in_3_
timestamp 1676037725
transform 1 0 28428 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_0.mux_l2_in_0_
timestamp 1676037725
transform 1 0 35880 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_0.mux_l2_in_1_
timestamp 1676037725
transform 1 0 28336 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_0.mux_l3_in_0_
timestamp 1676037725
transform 1 0 29716 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 27876 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_2.mux_l1_in_0_
timestamp 1676037725
transform 1 0 37444 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_2.mux_l1_in_1_
timestamp 1676037725
transform 1 0 40020 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_2.mux_l1_in_2_
timestamp 1676037725
transform 1 0 30360 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_2.mux_l2_in_0_
timestamp 1676037725
transform 1 0 38640 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_2.mux_l2_in_1_
timestamp 1676037725
transform 1 0 33028 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_2.mux_l2_in_1__234
timestamp 1676037725
transform 1 0 32476 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_2.mux_l3_in_0_
timestamp 1676037725
transform 1 0 32292 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 29164 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_4.mux_l1_in_0_
timestamp 1676037725
transform 1 0 34500 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_4.mux_l1_in_1_
timestamp 1676037725
transform 1 0 40020 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_4.mux_l2_in_0_
timestamp 1676037725
transform 1 0 35328 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_4.mux_l2_in_1__244
timestamp 1676037725
transform 1 0 31280 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_4.mux_l2_in_1_
timestamp 1676037725
transform 1 0 30084 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_4.mux_l3_in_0_
timestamp 1676037725
transform 1 0 30820 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 27140 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_6.mux_l1_in_0_
timestamp 1676037725
transform 1 0 40204 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_6.mux_l1_in_1_
timestamp 1676037725
transform 1 0 41216 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_6.mux_l1_in_2_
timestamp 1676037725
transform 1 0 32660 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_6.mux_l2_in_0_
timestamp 1676037725
transform 1 0 39652 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_6.mux_l2_in_1_
timestamp 1676037725
transform 1 0 36064 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_6.mux_l2_in_1__252
timestamp 1676037725
transform 1 0 37076 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_6.mux_l3_in_0_
timestamp 1676037725
transform 1 0 33580 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 30360 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_8.mux_l1_in_0_
timestamp 1676037725
transform 1 0 39468 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_8.mux_l1_in_1_
timestamp 1676037725
transform 1 0 41216 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_8.mux_l1_in_2_
timestamp 1676037725
transform 1 0 33488 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_8.mux_l2_in_0_
timestamp 1676037725
transform 1 0 40020 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_8.mux_l2_in_1__253
timestamp 1676037725
transform 1 0 39008 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_8.mux_l2_in_1_
timestamp 1676037725
transform 1 0 40020 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_8.mux_l3_in_0_
timestamp 1676037725
transform 1 0 37444 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 31464 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_10.mux_l1_in_0_
timestamp 1676037725
transform 1 0 34684 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_10.mux_l1_in_1_
timestamp 1676037725
transform 1 0 41216 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_10.mux_l2_in_0_
timestamp 1676037725
transform 1 0 36064 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_10.mux_l2_in_1_
timestamp 1676037725
transform 1 0 30912 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_10.mux_l2_in_1__229
timestamp 1676037725
transform 1 0 28980 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_10.mux_l3_in_0_
timestamp 1676037725
transform 1 0 31464 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 26404 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_12.mux_l1_in_0_
timestamp 1676037725
transform 1 0 39928 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_12.mux_l2_in_0_
timestamp 1676037725
transform 1 0 40388 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_12.mux_l2_in_1__230
timestamp 1676037725
transform 1 0 34868 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_12.mux_l2_in_1_
timestamp 1676037725
transform 1 0 35972 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_12.mux_l3_in_0_
timestamp 1676037725
transform 1 0 36064 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 29716 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_14.mux_l1_in_0_
timestamp 1676037725
transform 1 0 40112 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_14.mux_l2_in_0_
timestamp 1676037725
transform 1 0 40480 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_14.mux_l2_in_1__231
timestamp 1676037725
transform 1 0 37076 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_14.mux_l2_in_1_
timestamp 1676037725
transform 1 0 34684 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_14.mux_l3_in_0_
timestamp 1676037725
transform 1 0 35880 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 29716 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_16.mux_l1_in_0_
timestamp 1676037725
transform 1 0 37812 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_16.mux_l2_in_0_
timestamp 1676037725
transform 1 0 40480 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_16.mux_l2_in_1__232
timestamp 1676037725
transform 1 0 38640 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_16.mux_l2_in_1_
timestamp 1676037725
transform 1 0 34868 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_16.mux_l3_in_0_
timestamp 1676037725
transform 1 0 37444 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 28980 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_18.mux_l1_in_0_
timestamp 1676037725
transform 1 0 37996 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_18.mux_l2_in_0_
timestamp 1676037725
transform 1 0 39652 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_18.mux_l2_in_1__233
timestamp 1676037725
transform 1 0 31372 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_18.mux_l2_in_1_
timestamp 1676037725
transform 1 0 32292 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_18.mux_l3_in_0_
timestamp 1676037725
transform 1 0 31004 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 24564 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_20.mux_l1_in_0_
timestamp 1676037725
transform 1 0 27324 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_20.mux_l1_in_1__235
timestamp 1676037725
transform 1 0 24748 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_20.mux_l1_in_1_
timestamp 1676037725
transform 1 0 24840 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_20.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24932 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 22448 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_22.mux_l1_in_0_
timestamp 1676037725
transform 1 0 25852 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_22.mux_l1_in_1__236
timestamp 1676037725
transform 1 0 24196 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_22.mux_l1_in_1_
timestamp 1676037725
transform 1 0 23276 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_22.mux_l2_in_0_
timestamp 1676037725
transform 1 0 23000 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 20056 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_24.mux_l1_in_0_
timestamp 1676037725
transform 1 0 27140 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_24.mux_l1_in_1_
timestamp 1676037725
transform 1 0 22724 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_24.mux_l1_in_1__237
timestamp 1676037725
transform 1 0 23828 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_24.mux_l2_in_0_
timestamp 1676037725
transform 1 0 23276 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 16100 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_26.mux_l1_in_0_
timestamp 1676037725
transform 1 0 27416 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_26.mux_l1_in_1__238
timestamp 1676037725
transform 1 0 25392 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_26.mux_l1_in_1_
timestamp 1676037725
transform 1 0 24196 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_26.mux_l2_in_0_
timestamp 1676037725
transform 1 0 22080 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19412 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_28.mux_l1_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_28.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20700 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_28.mux_l2_in_0__239
timestamp 1676037725
transform 1 0 19780 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 15456 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_30.mux_l1_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_30.mux_l2_in_0__240
timestamp 1676037725
transform 1 0 17204 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_30.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19412 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 13524 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_32.mux_l1_in_0_
timestamp 1676037725
transform 1 0 18952 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_32.mux_l2_in_0_
timestamp 1676037725
transform 1 0 16744 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_32.mux_l2_in_0__241
timestamp 1676037725
transform 1 0 17112 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 12880 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_34.mux_l1_in_0_
timestamp 1676037725
transform 1 0 22264 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_34.mux_l2_in_0_
timestamp 1676037725
transform 1 0 18860 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_34.mux_l2_in_0__242
timestamp 1676037725
transform 1 0 19504 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 14720 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_36.mux_l1_in_0_
timestamp 1676037725
transform 1 0 27140 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_36.mux_l1_in_1__243
timestamp 1676037725
transform 1 0 21620 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_36.mux_l1_in_1_
timestamp 1676037725
transform 1 0 21988 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_36.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20700 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 15364 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_40.mux_l1_in_0_
timestamp 1676037725
transform 1 0 12788 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_40.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11776 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_40.mux_l2_in_0__245
timestamp 1676037725
transform 1 0 13064 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_40.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 9752 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_42.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16744 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_42.mux_l2_in_0__246
timestamp 1676037725
transform 1 0 10856 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_42.mux_l2_in_0_
timestamp 1676037725
transform 1 0 13892 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_42.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 10304 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_44.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15548 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_44.mux_l2_in_0__247
timestamp 1676037725
transform 1 0 10304 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_44.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12512 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_44.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 9844 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_46.mux_l1_in_0_
timestamp 1676037725
transform 1 0 11868 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_46.mux_l2_in_0__248
timestamp 1676037725
transform 1 0 9660 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_46.mux_l2_in_0_
timestamp 1676037725
transform 1 0 10396 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_46.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 9108 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_48.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_48.mux_l2_in_0_
timestamp 1676037725
transform 1 0 13708 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_48.mux_l2_in_0__249
timestamp 1676037725
transform 1 0 10304 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_48.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 8372 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_50.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16928 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_50.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12972 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_50.mux_l2_in_0__250
timestamp 1676037725
transform 1 0 9660 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_50.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 9936 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_58.mux_l1_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_58.mux_l2_in_0__251
timestamp 1676037725
transform 1 0 11684 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_58.mux_l2_in_0_
timestamp 1676037725
transform 1 0 16744 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_58.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 9108 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1676037725
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1676037725
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1676037725
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1676037725
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1676037725
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1676037725
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1676037725
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1676037725
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1676037725
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1676037725
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1676037725
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1676037725
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1676037725
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1676037725
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1676037725
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1676037725
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1676037725
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1676037725
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1676037725
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1676037725
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1676037725
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1676037725
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1676037725
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1676037725
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1676037725
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1676037725
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1676037725
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1676037725
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1676037725
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1676037725
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1676037725
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1676037725
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1676037725
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1676037725
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1676037725
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1676037725
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1676037725
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1676037725
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1676037725
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1676037725
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1676037725
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1676037725
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1676037725
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1676037725
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1676037725
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1676037725
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1676037725
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1676037725
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1676037725
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1676037725
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1676037725
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1676037725
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1676037725
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1676037725
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1676037725
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1676037725
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1676037725
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1676037725
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1676037725
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1676037725
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1676037725
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1676037725
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1676037725
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1676037725
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1676037725
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1676037725
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1676037725
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1676037725
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1676037725
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1676037725
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1676037725
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1676037725
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1676037725
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1676037725
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1676037725
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1676037725
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1676037725
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1676037725
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1676037725
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1676037725
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1676037725
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1676037725
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1676037725
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1676037725
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1676037725
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1676037725
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1676037725
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1676037725
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1676037725
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1676037725
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1676037725
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1676037725
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1676037725
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1676037725
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1676037725
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1676037725
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1676037725
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1676037725
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1676037725
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1676037725
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1676037725
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1676037725
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1676037725
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1676037725
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1676037725
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1676037725
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1676037725
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1676037725
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1676037725
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1676037725
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1676037725
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1676037725
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1676037725
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1676037725
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1676037725
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1676037725
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1676037725
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1676037725
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1676037725
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1676037725
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1676037725
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1676037725
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1676037725
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1676037725
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1676037725
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1676037725
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1676037725
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1676037725
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1676037725
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1676037725
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1676037725
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1676037725
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1676037725
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1676037725
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1676037725
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1676037725
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1676037725
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1676037725
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1676037725
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1676037725
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1676037725
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1676037725
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1676037725
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1676037725
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1676037725
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1676037725
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1676037725
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1676037725
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1676037725
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1676037725
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1676037725
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1676037725
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1676037725
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1676037725
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1676037725
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1676037725
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1676037725
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1676037725
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1676037725
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1676037725
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1676037725
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1676037725
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1676037725
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1676037725
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1676037725
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1676037725
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1676037725
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1676037725
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1676037725
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1676037725
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1676037725
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1676037725
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1676037725
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1676037725
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1676037725
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1676037725
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1676037725
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1676037725
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1676037725
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1676037725
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1676037725
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1676037725
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1676037725
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1676037725
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1676037725
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1676037725
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1676037725
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1676037725
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1676037725
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1676037725
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1676037725
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1676037725
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1676037725
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1676037725
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1676037725
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1676037725
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1676037725
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1676037725
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1676037725
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1676037725
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1676037725
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1676037725
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1676037725
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1676037725
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1676037725
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1676037725
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1676037725
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1676037725
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1676037725
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1676037725
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1676037725
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1676037725
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1676037725
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1676037725
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1676037725
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1676037725
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1676037725
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1676037725
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1676037725
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1676037725
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1676037725
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1676037725
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1676037725
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1676037725
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1676037725
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1676037725
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1676037725
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1676037725
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1676037725
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1676037725
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1676037725
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1676037725
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1676037725
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1676037725
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1676037725
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1676037725
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1676037725
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1676037725
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1676037725
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1676037725
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1676037725
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1676037725
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1676037725
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1676037725
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1676037725
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1676037725
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1676037725
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1676037725
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1676037725
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1676037725
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1676037725
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1676037725
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1676037725
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1676037725
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1676037725
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1676037725
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1676037725
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1676037725
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1676037725
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1676037725
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1676037725
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1676037725
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1676037725
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1676037725
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1676037725
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1676037725
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1676037725
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1676037725
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1676037725
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1676037725
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1676037725
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1676037725
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1676037725
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1676037725
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1676037725
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1676037725
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1676037725
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1676037725
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1676037725
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1676037725
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1676037725
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1676037725
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1676037725
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1676037725
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1676037725
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1676037725
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1676037725
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1676037725
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1676037725
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1676037725
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1676037725
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1676037725
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1676037725
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1676037725
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1676037725
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1676037725
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1676037725
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1676037725
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1676037725
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1676037725
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1676037725
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1676037725
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1676037725
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1676037725
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1676037725
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1676037725
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1676037725
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1676037725
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1676037725
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1676037725
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1676037725
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1676037725
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1676037725
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1676037725
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1676037725
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1676037725
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1676037725
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1676037725
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1676037725
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1676037725
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1676037725
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1676037725
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1676037725
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1676037725
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1676037725
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1676037725
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1676037725
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1676037725
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1676037725
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1676037725
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1676037725
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1676037725
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1676037725
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1676037725
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1676037725
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1676037725
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1676037725
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1676037725
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1676037725
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1676037725
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1676037725
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1676037725
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1676037725
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1676037725
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1676037725
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1676037725
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1676037725
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1676037725
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1676037725
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1676037725
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1676037725
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1676037725
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1676037725
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1676037725
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1676037725
transform 1 0 6256 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1676037725
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1676037725
transform 1 0 11408 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1676037725
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1676037725
transform 1 0 16560 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1676037725
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1676037725
transform 1 0 21712 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1676037725
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1676037725
transform 1 0 26864 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1676037725
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1676037725
transform 1 0 32016 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1676037725
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1676037725
transform 1 0 37168 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1676037725
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1676037725
transform 1 0 42320 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1676037725
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1676037725
transform 1 0 47472 0 1 23936
box -38 -48 130 592
<< labels >>
flabel metal4 s 7944 2128 8264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 17944 2128 18264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 27944 2128 28264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 37944 2128 38264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 47944 2128 48264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2944 2128 3264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 12944 2128 13264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 22944 2128 23264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 32944 2128 33264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 42944 2128 43264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 9586 0 9642 800 0 FreeSans 224 90 0 0 ccff_head
port 2 nsew signal input
flabel metal2 s 49238 26200 49294 27000 0 FreeSans 224 90 0 0 ccff_head_1
port 3 nsew signal input
flabel metal2 s 41326 0 41382 800 0 FreeSans 224 90 0 0 ccff_tail
port 4 nsew signal tristate
flabel metal2 s 1582 26200 1638 27000 0 FreeSans 224 90 0 0 ccff_tail_0
port 5 nsew signal tristate
flabel metal3 s 0 1504 800 1624 0 FreeSans 480 0 0 0 chanx_left_in[0]
port 6 nsew signal input
flabel metal3 s 0 5584 800 5704 0 FreeSans 480 0 0 0 chanx_left_in[10]
port 7 nsew signal input
flabel metal3 s 0 5992 800 6112 0 FreeSans 480 0 0 0 chanx_left_in[11]
port 8 nsew signal input
flabel metal3 s 0 6400 800 6520 0 FreeSans 480 0 0 0 chanx_left_in[12]
port 9 nsew signal input
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 chanx_left_in[13]
port 10 nsew signal input
flabel metal3 s 0 7216 800 7336 0 FreeSans 480 0 0 0 chanx_left_in[14]
port 11 nsew signal input
flabel metal3 s 0 7624 800 7744 0 FreeSans 480 0 0 0 chanx_left_in[15]
port 12 nsew signal input
flabel metal3 s 0 8032 800 8152 0 FreeSans 480 0 0 0 chanx_left_in[16]
port 13 nsew signal input
flabel metal3 s 0 8440 800 8560 0 FreeSans 480 0 0 0 chanx_left_in[17]
port 14 nsew signal input
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 chanx_left_in[18]
port 15 nsew signal input
flabel metal3 s 0 9256 800 9376 0 FreeSans 480 0 0 0 chanx_left_in[19]
port 16 nsew signal input
flabel metal3 s 0 1912 800 2032 0 FreeSans 480 0 0 0 chanx_left_in[1]
port 17 nsew signal input
flabel metal3 s 0 9664 800 9784 0 FreeSans 480 0 0 0 chanx_left_in[20]
port 18 nsew signal input
flabel metal3 s 0 10072 800 10192 0 FreeSans 480 0 0 0 chanx_left_in[21]
port 19 nsew signal input
flabel metal3 s 0 10480 800 10600 0 FreeSans 480 0 0 0 chanx_left_in[22]
port 20 nsew signal input
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 chanx_left_in[23]
port 21 nsew signal input
flabel metal3 s 0 11296 800 11416 0 FreeSans 480 0 0 0 chanx_left_in[24]
port 22 nsew signal input
flabel metal3 s 0 11704 800 11824 0 FreeSans 480 0 0 0 chanx_left_in[25]
port 23 nsew signal input
flabel metal3 s 0 12112 800 12232 0 FreeSans 480 0 0 0 chanx_left_in[26]
port 24 nsew signal input
flabel metal3 s 0 12520 800 12640 0 FreeSans 480 0 0 0 chanx_left_in[27]
port 25 nsew signal input
flabel metal3 s 0 12928 800 13048 0 FreeSans 480 0 0 0 chanx_left_in[28]
port 26 nsew signal input
flabel metal3 s 0 13336 800 13456 0 FreeSans 480 0 0 0 chanx_left_in[29]
port 27 nsew signal input
flabel metal3 s 0 2320 800 2440 0 FreeSans 480 0 0 0 chanx_left_in[2]
port 28 nsew signal input
flabel metal3 s 0 2728 800 2848 0 FreeSans 480 0 0 0 chanx_left_in[3]
port 29 nsew signal input
flabel metal3 s 0 3136 800 3256 0 FreeSans 480 0 0 0 chanx_left_in[4]
port 30 nsew signal input
flabel metal3 s 0 3544 800 3664 0 FreeSans 480 0 0 0 chanx_left_in[5]
port 31 nsew signal input
flabel metal3 s 0 3952 800 4072 0 FreeSans 480 0 0 0 chanx_left_in[6]
port 32 nsew signal input
flabel metal3 s 0 4360 800 4480 0 FreeSans 480 0 0 0 chanx_left_in[7]
port 33 nsew signal input
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 chanx_left_in[8]
port 34 nsew signal input
flabel metal3 s 0 5176 800 5296 0 FreeSans 480 0 0 0 chanx_left_in[9]
port 35 nsew signal input
flabel metal3 s 0 13744 800 13864 0 FreeSans 480 0 0 0 chanx_left_out[0]
port 36 nsew signal tristate
flabel metal3 s 0 17824 800 17944 0 FreeSans 480 0 0 0 chanx_left_out[10]
port 37 nsew signal tristate
flabel metal3 s 0 18232 800 18352 0 FreeSans 480 0 0 0 chanx_left_out[11]
port 38 nsew signal tristate
flabel metal3 s 0 18640 800 18760 0 FreeSans 480 0 0 0 chanx_left_out[12]
port 39 nsew signal tristate
flabel metal3 s 0 19048 800 19168 0 FreeSans 480 0 0 0 chanx_left_out[13]
port 40 nsew signal tristate
flabel metal3 s 0 19456 800 19576 0 FreeSans 480 0 0 0 chanx_left_out[14]
port 41 nsew signal tristate
flabel metal3 s 0 19864 800 19984 0 FreeSans 480 0 0 0 chanx_left_out[15]
port 42 nsew signal tristate
flabel metal3 s 0 20272 800 20392 0 FreeSans 480 0 0 0 chanx_left_out[16]
port 43 nsew signal tristate
flabel metal3 s 0 20680 800 20800 0 FreeSans 480 0 0 0 chanx_left_out[17]
port 44 nsew signal tristate
flabel metal3 s 0 21088 800 21208 0 FreeSans 480 0 0 0 chanx_left_out[18]
port 45 nsew signal tristate
flabel metal3 s 0 21496 800 21616 0 FreeSans 480 0 0 0 chanx_left_out[19]
port 46 nsew signal tristate
flabel metal3 s 0 14152 800 14272 0 FreeSans 480 0 0 0 chanx_left_out[1]
port 47 nsew signal tristate
flabel metal3 s 0 21904 800 22024 0 FreeSans 480 0 0 0 chanx_left_out[20]
port 48 nsew signal tristate
flabel metal3 s 0 22312 800 22432 0 FreeSans 480 0 0 0 chanx_left_out[21]
port 49 nsew signal tristate
flabel metal3 s 0 22720 800 22840 0 FreeSans 480 0 0 0 chanx_left_out[22]
port 50 nsew signal tristate
flabel metal3 s 0 23128 800 23248 0 FreeSans 480 0 0 0 chanx_left_out[23]
port 51 nsew signal tristate
flabel metal3 s 0 23536 800 23656 0 FreeSans 480 0 0 0 chanx_left_out[24]
port 52 nsew signal tristate
flabel metal3 s 0 23944 800 24064 0 FreeSans 480 0 0 0 chanx_left_out[25]
port 53 nsew signal tristate
flabel metal3 s 0 24352 800 24472 0 FreeSans 480 0 0 0 chanx_left_out[26]
port 54 nsew signal tristate
flabel metal3 s 0 24760 800 24880 0 FreeSans 480 0 0 0 chanx_left_out[27]
port 55 nsew signal tristate
flabel metal3 s 0 25168 800 25288 0 FreeSans 480 0 0 0 chanx_left_out[28]
port 56 nsew signal tristate
flabel metal3 s 0 25576 800 25696 0 FreeSans 480 0 0 0 chanx_left_out[29]
port 57 nsew signal tristate
flabel metal3 s 0 14560 800 14680 0 FreeSans 480 0 0 0 chanx_left_out[2]
port 58 nsew signal tristate
flabel metal3 s 0 14968 800 15088 0 FreeSans 480 0 0 0 chanx_left_out[3]
port 59 nsew signal tristate
flabel metal3 s 0 15376 800 15496 0 FreeSans 480 0 0 0 chanx_left_out[4]
port 60 nsew signal tristate
flabel metal3 s 0 15784 800 15904 0 FreeSans 480 0 0 0 chanx_left_out[5]
port 61 nsew signal tristate
flabel metal3 s 0 16192 800 16312 0 FreeSans 480 0 0 0 chanx_left_out[6]
port 62 nsew signal tristate
flabel metal3 s 0 16600 800 16720 0 FreeSans 480 0 0 0 chanx_left_out[7]
port 63 nsew signal tristate
flabel metal3 s 0 17008 800 17128 0 FreeSans 480 0 0 0 chanx_left_out[8]
port 64 nsew signal tristate
flabel metal3 s 0 17416 800 17536 0 FreeSans 480 0 0 0 chanx_left_out[9]
port 65 nsew signal tristate
flabel metal3 s 50200 13608 51000 13728 0 FreeSans 480 0 0 0 chanx_right_in_0[0]
port 66 nsew signal input
flabel metal3 s 50200 17688 51000 17808 0 FreeSans 480 0 0 0 chanx_right_in_0[10]
port 67 nsew signal input
flabel metal3 s 50200 18096 51000 18216 0 FreeSans 480 0 0 0 chanx_right_in_0[11]
port 68 nsew signal input
flabel metal3 s 50200 18504 51000 18624 0 FreeSans 480 0 0 0 chanx_right_in_0[12]
port 69 nsew signal input
flabel metal3 s 50200 18912 51000 19032 0 FreeSans 480 0 0 0 chanx_right_in_0[13]
port 70 nsew signal input
flabel metal3 s 50200 19320 51000 19440 0 FreeSans 480 0 0 0 chanx_right_in_0[14]
port 71 nsew signal input
flabel metal3 s 50200 19728 51000 19848 0 FreeSans 480 0 0 0 chanx_right_in_0[15]
port 72 nsew signal input
flabel metal3 s 50200 20136 51000 20256 0 FreeSans 480 0 0 0 chanx_right_in_0[16]
port 73 nsew signal input
flabel metal3 s 50200 20544 51000 20664 0 FreeSans 480 0 0 0 chanx_right_in_0[17]
port 74 nsew signal input
flabel metal3 s 50200 20952 51000 21072 0 FreeSans 480 0 0 0 chanx_right_in_0[18]
port 75 nsew signal input
flabel metal3 s 50200 21360 51000 21480 0 FreeSans 480 0 0 0 chanx_right_in_0[19]
port 76 nsew signal input
flabel metal3 s 50200 14016 51000 14136 0 FreeSans 480 0 0 0 chanx_right_in_0[1]
port 77 nsew signal input
flabel metal3 s 50200 21768 51000 21888 0 FreeSans 480 0 0 0 chanx_right_in_0[20]
port 78 nsew signal input
flabel metal3 s 50200 22176 51000 22296 0 FreeSans 480 0 0 0 chanx_right_in_0[21]
port 79 nsew signal input
flabel metal3 s 50200 22584 51000 22704 0 FreeSans 480 0 0 0 chanx_right_in_0[22]
port 80 nsew signal input
flabel metal3 s 50200 22992 51000 23112 0 FreeSans 480 0 0 0 chanx_right_in_0[23]
port 81 nsew signal input
flabel metal3 s 50200 23400 51000 23520 0 FreeSans 480 0 0 0 chanx_right_in_0[24]
port 82 nsew signal input
flabel metal3 s 50200 23808 51000 23928 0 FreeSans 480 0 0 0 chanx_right_in_0[25]
port 83 nsew signal input
flabel metal3 s 50200 24216 51000 24336 0 FreeSans 480 0 0 0 chanx_right_in_0[26]
port 84 nsew signal input
flabel metal3 s 50200 24624 51000 24744 0 FreeSans 480 0 0 0 chanx_right_in_0[27]
port 85 nsew signal input
flabel metal3 s 50200 25032 51000 25152 0 FreeSans 480 0 0 0 chanx_right_in_0[28]
port 86 nsew signal input
flabel metal3 s 50200 25440 51000 25560 0 FreeSans 480 0 0 0 chanx_right_in_0[29]
port 87 nsew signal input
flabel metal3 s 50200 14424 51000 14544 0 FreeSans 480 0 0 0 chanx_right_in_0[2]
port 88 nsew signal input
flabel metal3 s 50200 14832 51000 14952 0 FreeSans 480 0 0 0 chanx_right_in_0[3]
port 89 nsew signal input
flabel metal3 s 50200 15240 51000 15360 0 FreeSans 480 0 0 0 chanx_right_in_0[4]
port 90 nsew signal input
flabel metal3 s 50200 15648 51000 15768 0 FreeSans 480 0 0 0 chanx_right_in_0[5]
port 91 nsew signal input
flabel metal3 s 50200 16056 51000 16176 0 FreeSans 480 0 0 0 chanx_right_in_0[6]
port 92 nsew signal input
flabel metal3 s 50200 16464 51000 16584 0 FreeSans 480 0 0 0 chanx_right_in_0[7]
port 93 nsew signal input
flabel metal3 s 50200 16872 51000 16992 0 FreeSans 480 0 0 0 chanx_right_in_0[8]
port 94 nsew signal input
flabel metal3 s 50200 17280 51000 17400 0 FreeSans 480 0 0 0 chanx_right_in_0[9]
port 95 nsew signal input
flabel metal3 s 50200 1368 51000 1488 0 FreeSans 480 0 0 0 chanx_right_out_0[0]
port 96 nsew signal tristate
flabel metal3 s 50200 5448 51000 5568 0 FreeSans 480 0 0 0 chanx_right_out_0[10]
port 97 nsew signal tristate
flabel metal3 s 50200 5856 51000 5976 0 FreeSans 480 0 0 0 chanx_right_out_0[11]
port 98 nsew signal tristate
flabel metal3 s 50200 6264 51000 6384 0 FreeSans 480 0 0 0 chanx_right_out_0[12]
port 99 nsew signal tristate
flabel metal3 s 50200 6672 51000 6792 0 FreeSans 480 0 0 0 chanx_right_out_0[13]
port 100 nsew signal tristate
flabel metal3 s 50200 7080 51000 7200 0 FreeSans 480 0 0 0 chanx_right_out_0[14]
port 101 nsew signal tristate
flabel metal3 s 50200 7488 51000 7608 0 FreeSans 480 0 0 0 chanx_right_out_0[15]
port 102 nsew signal tristate
flabel metal3 s 50200 7896 51000 8016 0 FreeSans 480 0 0 0 chanx_right_out_0[16]
port 103 nsew signal tristate
flabel metal3 s 50200 8304 51000 8424 0 FreeSans 480 0 0 0 chanx_right_out_0[17]
port 104 nsew signal tristate
flabel metal3 s 50200 8712 51000 8832 0 FreeSans 480 0 0 0 chanx_right_out_0[18]
port 105 nsew signal tristate
flabel metal3 s 50200 9120 51000 9240 0 FreeSans 480 0 0 0 chanx_right_out_0[19]
port 106 nsew signal tristate
flabel metal3 s 50200 1776 51000 1896 0 FreeSans 480 0 0 0 chanx_right_out_0[1]
port 107 nsew signal tristate
flabel metal3 s 50200 9528 51000 9648 0 FreeSans 480 0 0 0 chanx_right_out_0[20]
port 108 nsew signal tristate
flabel metal3 s 50200 9936 51000 10056 0 FreeSans 480 0 0 0 chanx_right_out_0[21]
port 109 nsew signal tristate
flabel metal3 s 50200 10344 51000 10464 0 FreeSans 480 0 0 0 chanx_right_out_0[22]
port 110 nsew signal tristate
flabel metal3 s 50200 10752 51000 10872 0 FreeSans 480 0 0 0 chanx_right_out_0[23]
port 111 nsew signal tristate
flabel metal3 s 50200 11160 51000 11280 0 FreeSans 480 0 0 0 chanx_right_out_0[24]
port 112 nsew signal tristate
flabel metal3 s 50200 11568 51000 11688 0 FreeSans 480 0 0 0 chanx_right_out_0[25]
port 113 nsew signal tristate
flabel metal3 s 50200 11976 51000 12096 0 FreeSans 480 0 0 0 chanx_right_out_0[26]
port 114 nsew signal tristate
flabel metal3 s 50200 12384 51000 12504 0 FreeSans 480 0 0 0 chanx_right_out_0[27]
port 115 nsew signal tristate
flabel metal3 s 50200 12792 51000 12912 0 FreeSans 480 0 0 0 chanx_right_out_0[28]
port 116 nsew signal tristate
flabel metal3 s 50200 13200 51000 13320 0 FreeSans 480 0 0 0 chanx_right_out_0[29]
port 117 nsew signal tristate
flabel metal3 s 50200 2184 51000 2304 0 FreeSans 480 0 0 0 chanx_right_out_0[2]
port 118 nsew signal tristate
flabel metal3 s 50200 2592 51000 2712 0 FreeSans 480 0 0 0 chanx_right_out_0[3]
port 119 nsew signal tristate
flabel metal3 s 50200 3000 51000 3120 0 FreeSans 480 0 0 0 chanx_right_out_0[4]
port 120 nsew signal tristate
flabel metal3 s 50200 3408 51000 3528 0 FreeSans 480 0 0 0 chanx_right_out_0[5]
port 121 nsew signal tristate
flabel metal3 s 50200 3816 51000 3936 0 FreeSans 480 0 0 0 chanx_right_out_0[6]
port 122 nsew signal tristate
flabel metal3 s 50200 4224 51000 4344 0 FreeSans 480 0 0 0 chanx_right_out_0[7]
port 123 nsew signal tristate
flabel metal3 s 50200 4632 51000 4752 0 FreeSans 480 0 0 0 chanx_right_out_0[8]
port 124 nsew signal tristate
flabel metal3 s 50200 5040 51000 5160 0 FreeSans 480 0 0 0 chanx_right_out_0[9]
port 125 nsew signal tristate
flabel metal2 s 21546 26200 21602 27000 0 FreeSans 224 90 0 0 chany_top_in[0]
port 126 nsew signal input
flabel metal2 s 27986 26200 28042 27000 0 FreeSans 224 90 0 0 chany_top_in[10]
port 127 nsew signal input
flabel metal2 s 28630 26200 28686 27000 0 FreeSans 224 90 0 0 chany_top_in[11]
port 128 nsew signal input
flabel metal2 s 29274 26200 29330 27000 0 FreeSans 224 90 0 0 chany_top_in[12]
port 129 nsew signal input
flabel metal2 s 29918 26200 29974 27000 0 FreeSans 224 90 0 0 chany_top_in[13]
port 130 nsew signal input
flabel metal2 s 30562 26200 30618 27000 0 FreeSans 224 90 0 0 chany_top_in[14]
port 131 nsew signal input
flabel metal2 s 31206 26200 31262 27000 0 FreeSans 224 90 0 0 chany_top_in[15]
port 132 nsew signal input
flabel metal2 s 31850 26200 31906 27000 0 FreeSans 224 90 0 0 chany_top_in[16]
port 133 nsew signal input
flabel metal2 s 32494 26200 32550 27000 0 FreeSans 224 90 0 0 chany_top_in[17]
port 134 nsew signal input
flabel metal2 s 33138 26200 33194 27000 0 FreeSans 224 90 0 0 chany_top_in[18]
port 135 nsew signal input
flabel metal2 s 33782 26200 33838 27000 0 FreeSans 224 90 0 0 chany_top_in[19]
port 136 nsew signal input
flabel metal2 s 22190 26200 22246 27000 0 FreeSans 224 90 0 0 chany_top_in[1]
port 137 nsew signal input
flabel metal2 s 34426 26200 34482 27000 0 FreeSans 224 90 0 0 chany_top_in[20]
port 138 nsew signal input
flabel metal2 s 35070 26200 35126 27000 0 FreeSans 224 90 0 0 chany_top_in[21]
port 139 nsew signal input
flabel metal2 s 35714 26200 35770 27000 0 FreeSans 224 90 0 0 chany_top_in[22]
port 140 nsew signal input
flabel metal2 s 36358 26200 36414 27000 0 FreeSans 224 90 0 0 chany_top_in[23]
port 141 nsew signal input
flabel metal2 s 37002 26200 37058 27000 0 FreeSans 224 90 0 0 chany_top_in[24]
port 142 nsew signal input
flabel metal2 s 37646 26200 37702 27000 0 FreeSans 224 90 0 0 chany_top_in[25]
port 143 nsew signal input
flabel metal2 s 38290 26200 38346 27000 0 FreeSans 224 90 0 0 chany_top_in[26]
port 144 nsew signal input
flabel metal2 s 38934 26200 38990 27000 0 FreeSans 224 90 0 0 chany_top_in[27]
port 145 nsew signal input
flabel metal2 s 39578 26200 39634 27000 0 FreeSans 224 90 0 0 chany_top_in[28]
port 146 nsew signal input
flabel metal2 s 40222 26200 40278 27000 0 FreeSans 224 90 0 0 chany_top_in[29]
port 147 nsew signal input
flabel metal2 s 22834 26200 22890 27000 0 FreeSans 224 90 0 0 chany_top_in[2]
port 148 nsew signal input
flabel metal2 s 23478 26200 23534 27000 0 FreeSans 224 90 0 0 chany_top_in[3]
port 149 nsew signal input
flabel metal2 s 24122 26200 24178 27000 0 FreeSans 224 90 0 0 chany_top_in[4]
port 150 nsew signal input
flabel metal2 s 24766 26200 24822 27000 0 FreeSans 224 90 0 0 chany_top_in[5]
port 151 nsew signal input
flabel metal2 s 25410 26200 25466 27000 0 FreeSans 224 90 0 0 chany_top_in[6]
port 152 nsew signal input
flabel metal2 s 26054 26200 26110 27000 0 FreeSans 224 90 0 0 chany_top_in[7]
port 153 nsew signal input
flabel metal2 s 26698 26200 26754 27000 0 FreeSans 224 90 0 0 chany_top_in[8]
port 154 nsew signal input
flabel metal2 s 27342 26200 27398 27000 0 FreeSans 224 90 0 0 chany_top_in[9]
port 155 nsew signal input
flabel metal2 s 2226 26200 2282 27000 0 FreeSans 224 90 0 0 chany_top_out[0]
port 156 nsew signal tristate
flabel metal2 s 8666 26200 8722 27000 0 FreeSans 224 90 0 0 chany_top_out[10]
port 157 nsew signal tristate
flabel metal2 s 9310 26200 9366 27000 0 FreeSans 224 90 0 0 chany_top_out[11]
port 158 nsew signal tristate
flabel metal2 s 9954 26200 10010 27000 0 FreeSans 224 90 0 0 chany_top_out[12]
port 159 nsew signal tristate
flabel metal2 s 10598 26200 10654 27000 0 FreeSans 224 90 0 0 chany_top_out[13]
port 160 nsew signal tristate
flabel metal2 s 11242 26200 11298 27000 0 FreeSans 224 90 0 0 chany_top_out[14]
port 161 nsew signal tristate
flabel metal2 s 11886 26200 11942 27000 0 FreeSans 224 90 0 0 chany_top_out[15]
port 162 nsew signal tristate
flabel metal2 s 12530 26200 12586 27000 0 FreeSans 224 90 0 0 chany_top_out[16]
port 163 nsew signal tristate
flabel metal2 s 13174 26200 13230 27000 0 FreeSans 224 90 0 0 chany_top_out[17]
port 164 nsew signal tristate
flabel metal2 s 13818 26200 13874 27000 0 FreeSans 224 90 0 0 chany_top_out[18]
port 165 nsew signal tristate
flabel metal2 s 14462 26200 14518 27000 0 FreeSans 224 90 0 0 chany_top_out[19]
port 166 nsew signal tristate
flabel metal2 s 2870 26200 2926 27000 0 FreeSans 224 90 0 0 chany_top_out[1]
port 167 nsew signal tristate
flabel metal2 s 15106 26200 15162 27000 0 FreeSans 224 90 0 0 chany_top_out[20]
port 168 nsew signal tristate
flabel metal2 s 15750 26200 15806 27000 0 FreeSans 224 90 0 0 chany_top_out[21]
port 169 nsew signal tristate
flabel metal2 s 16394 26200 16450 27000 0 FreeSans 224 90 0 0 chany_top_out[22]
port 170 nsew signal tristate
flabel metal2 s 17038 26200 17094 27000 0 FreeSans 224 90 0 0 chany_top_out[23]
port 171 nsew signal tristate
flabel metal2 s 17682 26200 17738 27000 0 FreeSans 224 90 0 0 chany_top_out[24]
port 172 nsew signal tristate
flabel metal2 s 18326 26200 18382 27000 0 FreeSans 224 90 0 0 chany_top_out[25]
port 173 nsew signal tristate
flabel metal2 s 18970 26200 19026 27000 0 FreeSans 224 90 0 0 chany_top_out[26]
port 174 nsew signal tristate
flabel metal2 s 19614 26200 19670 27000 0 FreeSans 224 90 0 0 chany_top_out[27]
port 175 nsew signal tristate
flabel metal2 s 20258 26200 20314 27000 0 FreeSans 224 90 0 0 chany_top_out[28]
port 176 nsew signal tristate
flabel metal2 s 20902 26200 20958 27000 0 FreeSans 224 90 0 0 chany_top_out[29]
port 177 nsew signal tristate
flabel metal2 s 3514 26200 3570 27000 0 FreeSans 224 90 0 0 chany_top_out[2]
port 178 nsew signal tristate
flabel metal2 s 4158 26200 4214 27000 0 FreeSans 224 90 0 0 chany_top_out[3]
port 179 nsew signal tristate
flabel metal2 s 4802 26200 4858 27000 0 FreeSans 224 90 0 0 chany_top_out[4]
port 180 nsew signal tristate
flabel metal2 s 5446 26200 5502 27000 0 FreeSans 224 90 0 0 chany_top_out[5]
port 181 nsew signal tristate
flabel metal2 s 6090 26200 6146 27000 0 FreeSans 224 90 0 0 chany_top_out[6]
port 182 nsew signal tristate
flabel metal2 s 6734 26200 6790 27000 0 FreeSans 224 90 0 0 chany_top_out[7]
port 183 nsew signal tristate
flabel metal2 s 7378 26200 7434 27000 0 FreeSans 224 90 0 0 chany_top_out[8]
port 184 nsew signal tristate
flabel metal2 s 8022 26200 8078 27000 0 FreeSans 224 90 0 0 chany_top_out[9]
port 185 nsew signal tristate
flabel metal2 s 11702 0 11758 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[0]
port 186 nsew signal tristate
flabel metal2 s 13818 0 13874 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[1]
port 187 nsew signal tristate
flabel metal2 s 15934 0 15990 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[2]
port 188 nsew signal tristate
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[3]
port 189 nsew signal tristate
flabel metal2 s 28630 0 28686 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[0]
port 190 nsew signal input
flabel metal2 s 30746 0 30802 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[1]
port 191 nsew signal input
flabel metal2 s 32862 0 32918 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[2]
port 192 nsew signal input
flabel metal2 s 34978 0 35034 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[3]
port 193 nsew signal input
flabel metal2 s 20166 0 20222 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[0]
port 194 nsew signal tristate
flabel metal2 s 22282 0 22338 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[1]
port 195 nsew signal tristate
flabel metal2 s 24398 0 24454 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[2]
port 196 nsew signal tristate
flabel metal2 s 26514 0 26570 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[3]
port 197 nsew signal tristate
flabel metal2 s 37094 0 37150 800 0 FreeSans 224 90 0 0 isol_n
port 198 nsew signal input
flabel metal2 s 39210 0 39266 800 0 FreeSans 224 90 0 0 prog_clk
port 199 nsew signal input
flabel metal2 s 42154 26200 42210 27000 0 FreeSans 224 90 0 0 prog_reset_top_in
port 200 nsew signal input
flabel metal2 s 42798 26200 42854 27000 0 FreeSans 224 90 0 0 reset_top_in
port 201 nsew signal input
flabel metal2 s 43442 0 43498 800 0 FreeSans 224 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
port 202 nsew signal input
flabel metal2 s 45558 0 45614 800 0 FreeSans 224 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
port 203 nsew signal input
flabel metal2 s 47674 0 47730 800 0 FreeSans 224 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
port 204 nsew signal input
flabel metal2 s 49790 0 49846 800 0 FreeSans 224 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
port 205 nsew signal input
flabel metal2 s 43442 26200 43498 27000 0 FreeSans 224 90 0 0 test_enable_top_in
port 206 nsew signal input
flabel metal2 s 45374 26200 45430 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_
port 207 nsew signal input
flabel metal2 s 46018 26200 46074 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_
port 208 nsew signal input
flabel metal2 s 46662 26200 46718 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_
port 209 nsew signal input
flabel metal2 s 47306 26200 47362 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_
port 210 nsew signal input
flabel metal2 s 47950 26200 48006 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_
port 211 nsew signal input
flabel metal2 s 48594 26200 48650 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_
port 212 nsew signal input
flabel metal2 s 44086 26200 44142 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_
port 213 nsew signal input
flabel metal2 s 44730 26200 44786 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_
port 214 nsew signal input
flabel metal2 s 1122 0 1178 800 0 FreeSans 224 90 0 0 top_width_0_height_0_subtile_0__pin_inpad_0_
port 215 nsew signal tristate
flabel metal2 s 3238 0 3294 800 0 FreeSans 224 90 0 0 top_width_0_height_0_subtile_1__pin_inpad_0_
port 216 nsew signal tristate
flabel metal2 s 5354 0 5410 800 0 FreeSans 224 90 0 0 top_width_0_height_0_subtile_2__pin_inpad_0_
port 217 nsew signal tristate
flabel metal2 s 7470 0 7526 800 0 FreeSans 224 90 0 0 top_width_0_height_0_subtile_3__pin_inpad_0_
port 218 nsew signal tristate
rlabel metal1 25484 23936 25484 23936 0 VGND
rlabel metal1 25484 24480 25484 24480 0 VPWR
rlabel metal2 21942 5644 21942 5644 0 cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_
rlabel metal2 20470 5916 20470 5916 0 cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_
rlabel metal2 18998 6494 18998 6494 0 cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_
rlabel metal1 17250 6290 17250 6290 0 cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_
rlabel metal1 21298 19244 21298 19244 0 cbx_1__0_.cbx_8__0_.ccff_head
rlabel metal2 18630 9044 18630 9044 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_0.ccff_tail
rlabel metal1 21298 14892 21298 14892 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[0\]
rlabel metal1 17020 13498 17020 13498 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[1\]
rlabel metal1 18354 10166 18354 10166 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[2\]
rlabel metal2 15318 9588 15318 9588 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_1.ccff_tail
rlabel metal2 17434 15045 17434 15045 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[0\]
rlabel metal1 16146 13804 16146 13804 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[1\]
rlabel metal2 13754 10625 13754 10625 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[2\]
rlabel metal2 12742 10370 12742 10370 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_2.ccff_tail
rlabel metal1 15180 9622 15180 9622 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[0\]
rlabel metal1 13754 13158 13754 13158 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[1\]
rlabel metal1 11270 11016 11270 11016 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[2\]
rlabel metal1 13655 14790 13655 14790 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[0\]
rlabel metal1 13754 15572 13754 15572 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[1\]
rlabel metal1 13064 15334 13064 15334 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[2\]
rlabel metal1 15548 13362 15548 13362 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18216 7854 18216 7854 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 19596 6766 19596 6766 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal2 15594 14450 15594 14450 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 17618 14994 17618 14994 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 17526 14450 17526 14450 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 15870 12614 15870 12614 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 15640 11186 15640 11186 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 16974 14042 16974 14042 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 18262 10132 18262 10132 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 18630 10030 18630 10030 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 17342 7922 17342 7922 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 12926 16150 12926 16150 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 14582 10778 14582 10778 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 16744 7378 16744 7378 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 13202 16218 13202 16218 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 17802 13974 17802 13974 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 15962 14416 15962 14416 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 18216 11254 18216 11254 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 12696 15878 12696 15878 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 15456 14042 15456 14042 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal2 14398 9894 14398 9894 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 17802 10744 17802 10744 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal2 16054 11594 16054 11594 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 9752 15062 9752 15062 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 12466 9894 12466 9894 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal2 12834 8636 12834 8636 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 9522 15130 9522 15130 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14766 14484 14766 14484 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 14904 14314 14904 14314 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 15548 10642 15548 10642 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 11546 12954 11546 12954 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 12190 12886 12190 12886 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal2 12098 10302 12098 10302 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 11868 14042 11868 14042 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 12604 9622 12604 9622 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 13524 15538 13524 15538 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 12834 14518 12834 14518 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal2 13478 14013 13478 14013 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 13984 15470 13984 15470 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 15870 15130 15870 15130 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 18216 14790 18216 14790 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 14858 11356 14858 11356 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 12282 15844 12282 15844 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 14674 15130 14674 15130 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 13616 14246 13616 14246 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 14306 14382 14306 14382 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 11684 16218 11684 16218 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 19550 3434 19550 3434 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.ccff_tail
rlabel metal1 20194 3060 20194 3060 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
rlabel metal1 26358 3026 26358 3026 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_out
rlabel metal1 27140 4182 27140 4182 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel via1 23322 3094 23322 3094 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.ccff_tail
rlabel metal1 19228 2414 19228 2414 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
rlabel metal2 21482 3740 21482 3740 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_out
rlabel metal1 24449 4522 24449 4522 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 27554 2958 27554 2958 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.ccff_tail
rlabel metal2 19182 4114 19182 4114 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
rlabel metal2 20838 4012 20838 4012 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_out
rlabel metal2 24334 4522 24334 4522 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 18308 6222 18308 6222 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
rlabel metal1 19182 6086 19182 6086 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_out
rlabel metal2 24794 3740 24794 3740 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal2 9614 1588 9614 1588 0 ccff_head
rlabel metal1 47242 23120 47242 23120 0 ccff_head_1
rlabel metal2 41354 1622 41354 1622 0 ccff_tail
rlabel metal1 2990 23222 2990 23222 0 ccff_tail_0
rlabel metal3 1004 1564 1004 1564 0 chanx_left_in[0]
rlabel metal3 820 5644 820 5644 0 chanx_left_in[10]
rlabel metal3 820 6052 820 6052 0 chanx_left_in[11]
rlabel metal3 1004 6460 1004 6460 0 chanx_left_in[12]
rlabel metal3 820 6868 820 6868 0 chanx_left_in[13]
rlabel metal3 820 7276 820 7276 0 chanx_left_in[14]
rlabel metal3 820 7684 820 7684 0 chanx_left_in[15]
rlabel metal3 1142 8092 1142 8092 0 chanx_left_in[16]
rlabel metal3 958 8500 958 8500 0 chanx_left_in[17]
rlabel metal3 820 8908 820 8908 0 chanx_left_in[18]
rlabel metal3 820 9316 820 9316 0 chanx_left_in[19]
rlabel metal3 958 1972 958 1972 0 chanx_left_in[1]
rlabel metal3 820 9724 820 9724 0 chanx_left_in[20]
rlabel metal3 958 10132 958 10132 0 chanx_left_in[21]
rlabel metal3 820 10540 820 10540 0 chanx_left_in[22]
rlabel metal3 1142 10948 1142 10948 0 chanx_left_in[23]
rlabel metal3 820 11356 820 11356 0 chanx_left_in[24]
rlabel metal3 820 11764 820 11764 0 chanx_left_in[25]
rlabel metal3 866 12172 866 12172 0 chanx_left_in[26]
rlabel metal3 1004 12580 1004 12580 0 chanx_left_in[27]
rlabel metal3 820 12988 820 12988 0 chanx_left_in[28]
rlabel metal2 3542 13651 3542 13651 0 chanx_left_in[29]
rlabel metal3 820 2380 820 2380 0 chanx_left_in[2]
rlabel metal3 820 2788 820 2788 0 chanx_left_in[3]
rlabel metal3 820 3196 820 3196 0 chanx_left_in[4]
rlabel metal3 820 3604 820 3604 0 chanx_left_in[5]
rlabel metal3 1188 4012 1188 4012 0 chanx_left_in[6]
rlabel metal3 820 4420 820 4420 0 chanx_left_in[7]
rlabel metal3 820 4828 820 4828 0 chanx_left_in[8]
rlabel metal3 1510 5236 1510 5236 0 chanx_left_in[9]
rlabel metal2 2806 13549 2806 13549 0 chanx_left_out[0]
rlabel metal3 1694 17884 1694 17884 0 chanx_left_out[10]
rlabel metal2 2898 18819 2898 18819 0 chanx_left_out[11]
rlabel metal3 1004 18700 1004 18700 0 chanx_left_out[12]
rlabel metal3 1004 19108 1004 19108 0 chanx_left_out[13]
rlabel metal3 1694 19516 1694 19516 0 chanx_left_out[14]
rlabel metal2 3358 20689 3358 20689 0 chanx_left_out[15]
rlabel via2 3910 20349 3910 20349 0 chanx_left_out[16]
rlabel metal3 1004 20740 1004 20740 0 chanx_left_out[17]
rlabel metal1 2852 22678 2852 22678 0 chanx_left_out[18]
rlabel metal3 1694 21556 1694 21556 0 chanx_left_out[19]
rlabel metal3 1004 14212 1004 14212 0 chanx_left_out[1]
rlabel metal2 3818 22015 3818 22015 0 chanx_left_out[20]
rlabel metal3 1579 22372 1579 22372 0 chanx_left_out[21]
rlabel metal3 2062 22780 2062 22780 0 chanx_left_out[22]
rlabel metal3 2016 23188 2016 23188 0 chanx_left_out[23]
rlabel metal3 2062 23596 2062 23596 0 chanx_left_out[24]
rlabel metal3 2200 24004 2200 24004 0 chanx_left_out[25]
rlabel metal3 1740 24412 1740 24412 0 chanx_left_out[26]
rlabel metal3 1924 24820 1924 24820 0 chanx_left_out[27]
rlabel metal3 2016 25228 2016 25228 0 chanx_left_out[28]
rlabel metal3 2062 25636 2062 25636 0 chanx_left_out[29]
rlabel metal3 1004 14620 1004 14620 0 chanx_left_out[2]
rlabel metal3 1004 15028 1004 15028 0 chanx_left_out[3]
rlabel metal3 1004 15436 1004 15436 0 chanx_left_out[4]
rlabel metal3 1004 15844 1004 15844 0 chanx_left_out[5]
rlabel metal3 1004 16252 1004 16252 0 chanx_left_out[6]
rlabel metal3 1004 16660 1004 16660 0 chanx_left_out[7]
rlabel metal3 958 17068 958 17068 0 chanx_left_out[8]
rlabel metal2 2806 17833 2806 17833 0 chanx_left_out[9]
rlabel metal1 48438 13906 48438 13906 0 chanx_right_in_0[0]
rlabel metal2 49082 18003 49082 18003 0 chanx_right_in_0[10]
rlabel metal1 49128 18734 49128 18734 0 chanx_right_in_0[11]
rlabel metal2 48622 18649 48622 18649 0 chanx_right_in_0[12]
rlabel metal2 49174 19159 49174 19159 0 chanx_right_in_0[13]
rlabel metal1 49266 19754 49266 19754 0 chanx_right_in_0[14]
rlabel metal2 49082 20111 49082 20111 0 chanx_right_in_0[15]
rlabel metal2 48622 20315 48622 20315 0 chanx_right_in_0[16]
rlabel metal2 49082 20757 49082 20757 0 chanx_right_in_0[17]
rlabel metal2 49082 21267 49082 21267 0 chanx_right_in_0[18]
rlabel metal2 49174 21675 49174 21675 0 chanx_right_in_0[19]
rlabel metal2 49174 14025 49174 14025 0 chanx_right_in_0[1]
rlabel metal2 48622 21913 48622 21913 0 chanx_right_in_0[20]
rlabel metal2 49082 22423 49082 22423 0 chanx_right_in_0[21]
rlabel metal1 49128 23086 49128 23086 0 chanx_right_in_0[22]
rlabel via2 48346 23069 48346 23069 0 chanx_right_in_0[23]
rlabel metal2 47886 23273 47886 23273 0 chanx_right_in_0[24]
rlabel metal2 46322 23409 46322 23409 0 chanx_right_in_0[25]
rlabel metal1 48392 22610 48392 22610 0 chanx_right_in_0[26]
rlabel metal1 47380 21998 47380 21998 0 chanx_right_in_0[27]
rlabel metal1 47012 22610 47012 22610 0 chanx_right_in_0[28]
rlabel metal1 48392 24242 48392 24242 0 chanx_right_in_0[29]
rlabel metal2 49082 14433 49082 14433 0 chanx_right_in_0[2]
rlabel metal2 49082 14943 49082 14943 0 chanx_right_in_0[3]
rlabel metal2 49358 15385 49358 15385 0 chanx_right_in_0[4]
rlabel metal2 49082 15895 49082 15895 0 chanx_right_in_0[5]
rlabel metal1 49128 16558 49128 16558 0 chanx_right_in_0[6]
rlabel metal1 48714 17238 48714 17238 0 chanx_right_in_0[7]
rlabel metal2 48622 17051 48622 17051 0 chanx_right_in_0[8]
rlabel metal2 49082 17493 49082 17493 0 chanx_right_in_0[9]
rlabel metal2 46690 2737 46690 2737 0 chanx_right_out_0[0]
rlabel metal1 49312 4658 49312 4658 0 chanx_right_out_0[10]
rlabel metal2 49174 5593 49174 5593 0 chanx_right_out_0[11]
rlabel metal3 49596 6324 49596 6324 0 chanx_right_out_0[12]
rlabel metal1 49312 5746 49312 5746 0 chanx_right_out_0[13]
rlabel metal1 49220 6358 49220 6358 0 chanx_right_out_0[14]
rlabel metal3 49734 7548 49734 7548 0 chanx_right_out_0[15]
rlabel metal2 46874 8177 46874 8177 0 chanx_right_out_0[16]
rlabel metal1 49266 7446 49266 7446 0 chanx_right_out_0[17]
rlabel metal1 49220 7922 49220 7922 0 chanx_right_out_0[18]
rlabel metal2 49174 8857 49174 8857 0 chanx_right_out_0[19]
rlabel metal2 46782 2397 46782 2397 0 chanx_right_out_0[1]
rlabel metal3 48814 9588 48814 9588 0 chanx_right_out_0[20]
rlabel metal1 49220 9010 49220 9010 0 chanx_right_out_0[21]
rlabel metal1 49266 9622 49266 9622 0 chanx_right_out_0[22]
rlabel metal2 49174 10455 49174 10455 0 chanx_right_out_0[23]
rlabel metal1 49220 10710 49220 10710 0 chanx_right_out_0[24]
rlabel metal2 49174 11407 49174 11407 0 chanx_right_out_0[25]
rlabel metal2 49174 11917 49174 11917 0 chanx_right_out_0[26]
rlabel metal2 49174 12359 49174 12359 0 chanx_right_out_0[27]
rlabel via2 49174 12835 49174 12835 0 chanx_right_out_0[28]
rlabel metal3 49734 13260 49734 13260 0 chanx_right_out_0[29]
rlabel metal3 49412 2244 49412 2244 0 chanx_right_out_0[2]
rlabel metal2 46874 2805 46874 2805 0 chanx_right_out_0[3]
rlabel metal3 49504 3060 49504 3060 0 chanx_right_out_0[4]
rlabel metal2 49174 2975 49174 2975 0 chanx_right_out_0[5]
rlabel metal1 49220 3094 49220 3094 0 chanx_right_out_0[6]
rlabel metal2 49174 3927 49174 3927 0 chanx_right_out_0[7]
rlabel metal1 47610 5134 47610 5134 0 chanx_right_out_0[8]
rlabel metal1 49266 4114 49266 4114 0 chanx_right_out_0[9]
rlabel metal2 21942 24701 21942 24701 0 chany_top_in[0]
rlabel metal1 29946 24208 29946 24208 0 chany_top_in[10]
rlabel metal1 31326 24242 31326 24242 0 chany_top_in[11]
rlabel metal2 35098 24412 35098 24412 0 chany_top_in[12]
rlabel via2 34178 21981 34178 21981 0 chany_top_in[13]
rlabel metal1 32890 23188 32890 23188 0 chany_top_in[14]
rlabel metal2 32246 21556 32246 21556 0 chany_top_in[15]
rlabel metal2 39238 24650 39238 24650 0 chany_top_in[16]
rlabel metal1 40894 24140 40894 24140 0 chany_top_in[17]
rlabel metal2 38686 24463 38686 24463 0 chany_top_in[18]
rlabel metal3 38318 21420 38318 21420 0 chany_top_in[19]
rlabel metal1 14858 23222 14858 23222 0 chany_top_in[1]
rlabel metal2 34507 26316 34507 26316 0 chany_top_in[20]
rlabel metal1 41078 23664 41078 23664 0 chany_top_in[21]
rlabel metal2 35742 25476 35742 25476 0 chany_top_in[22]
rlabel metal1 41354 23732 41354 23732 0 chany_top_in[23]
rlabel metal2 37030 24354 37030 24354 0 chany_top_in[24]
rlabel metal1 38916 22066 38916 22066 0 chany_top_in[25]
rlabel metal3 41170 21964 41170 21964 0 chany_top_in[26]
rlabel metal2 41814 23698 41814 23698 0 chany_top_in[27]
rlabel metal2 40342 22848 40342 22848 0 chany_top_in[28]
rlabel metal1 43194 21998 43194 21998 0 chany_top_in[29]
rlabel metal1 25898 20434 25898 20434 0 chany_top_in[2]
rlabel metal1 16054 23562 16054 23562 0 chany_top_in[3]
rlabel metal1 33166 24208 33166 24208 0 chany_top_in[4]
rlabel metal2 31234 24378 31234 24378 0 chany_top_in[5]
rlabel metal1 24748 24174 24748 24174 0 chany_top_in[6]
rlabel metal2 28750 24242 28750 24242 0 chany_top_in[7]
rlabel metal1 27416 24174 27416 24174 0 chany_top_in[8]
rlabel metal1 28750 23732 28750 23732 0 chany_top_in[9]
rlabel metal1 3588 22202 3588 22202 0 chany_top_out[0]
rlabel metal1 8464 24242 8464 24242 0 chany_top_out[10]
rlabel metal1 9246 23766 9246 23766 0 chany_top_out[11]
rlabel metal1 10166 22542 10166 22542 0 chany_top_out[12]
rlabel metal1 10672 23766 10672 23766 0 chany_top_out[13]
rlabel metal2 11270 24728 11270 24728 0 chany_top_out[14]
rlabel metal1 10994 24276 10994 24276 0 chany_top_out[15]
rlabel metal1 12834 22542 12834 22542 0 chany_top_out[16]
rlabel metal2 13386 24735 13386 24735 0 chany_top_out[17]
rlabel metal1 13708 24242 13708 24242 0 chany_top_out[18]
rlabel metal2 14398 24361 14398 24361 0 chany_top_out[19]
rlabel metal1 3542 23018 3542 23018 0 chany_top_out[1]
rlabel metal1 15226 22542 15226 22542 0 chany_top_out[20]
rlabel metal2 15778 24728 15778 24728 0 chany_top_out[21]
rlabel metal2 16146 25041 16146 25041 0 chany_top_out[22]
rlabel metal1 17618 22134 17618 22134 0 chany_top_out[23]
rlabel metal1 16928 24242 16928 24242 0 chany_top_out[24]
rlabel metal1 18262 23766 18262 23766 0 chany_top_out[25]
rlabel metal1 19458 22134 19458 22134 0 chany_top_out[26]
rlabel metal1 19136 24242 19136 24242 0 chany_top_out[27]
rlabel metal2 20562 25313 20562 25313 0 chany_top_out[28]
rlabel metal2 20930 25272 20930 25272 0 chany_top_out[29]
rlabel metal1 3404 24242 3404 24242 0 chany_top_out[2]
rlabel metal1 4094 23766 4094 23766 0 chany_top_out[3]
rlabel metal2 5106 24429 5106 24429 0 chany_top_out[4]
rlabel metal2 5474 24966 5474 24966 0 chany_top_out[5]
rlabel metal2 6118 24728 6118 24728 0 chany_top_out[6]
rlabel metal1 6302 24242 6302 24242 0 chany_top_out[7]
rlabel metal1 7682 22542 7682 22542 0 chany_top_out[8]
rlabel metal2 7866 23919 7866 23919 0 chany_top_out[9]
rlabel metal1 17848 12818 17848 12818 0 clknet_0_prog_clk
rlabel metal1 13570 8500 13570 8500 0 clknet_4_0_0_prog_clk
rlabel metal1 33672 10574 33672 10574 0 clknet_4_10_0_prog_clk
rlabel metal1 36110 13294 36110 13294 0 clknet_4_11_0_prog_clk
rlabel metal1 32338 17238 32338 17238 0 clknet_4_12_0_prog_clk
rlabel metal2 35282 19108 35282 19108 0 clknet_4_13_0_prog_clk
rlabel metal1 38962 17068 38962 17068 0 clknet_4_14_0_prog_clk
rlabel metal1 35788 17714 35788 17714 0 clknet_4_15_0_prog_clk
rlabel metal1 12098 11764 12098 11764 0 clknet_4_1_0_prog_clk
rlabel metal2 20930 3230 20930 3230 0 clknet_4_2_0_prog_clk
rlabel metal2 21482 11424 21482 11424 0 clknet_4_3_0_prog_clk
rlabel metal1 19964 16014 19964 16014 0 clknet_4_4_0_prog_clk
rlabel metal1 19642 18292 19642 18292 0 clknet_4_5_0_prog_clk
rlabel metal1 25760 18802 25760 18802 0 clknet_4_6_0_prog_clk
rlabel metal1 19688 20366 19688 20366 0 clknet_4_7_0_prog_clk
rlabel metal2 28842 5712 28842 5712 0 clknet_4_8_0_prog_clk
rlabel metal2 24886 14110 24886 14110 0 clknet_4_9_0_prog_clk
rlabel metal2 11730 1622 11730 1622 0 gfpga_pad_io_soc_dir[0]
rlabel metal2 13846 1622 13846 1622 0 gfpga_pad_io_soc_dir[1]
rlabel metal2 15962 1622 15962 1622 0 gfpga_pad_io_soc_dir[2]
rlabel metal2 18078 823 18078 823 0 gfpga_pad_io_soc_dir[3]
rlabel metal2 28658 1588 28658 1588 0 gfpga_pad_io_soc_in[0]
rlabel metal2 30774 1588 30774 1588 0 gfpga_pad_io_soc_in[1]
rlabel metal2 32890 1588 32890 1588 0 gfpga_pad_io_soc_in[2]
rlabel metal2 35006 1588 35006 1588 0 gfpga_pad_io_soc_in[3]
rlabel metal2 20194 1622 20194 1622 0 gfpga_pad_io_soc_out[0]
rlabel metal2 22310 1622 22310 1622 0 gfpga_pad_io_soc_out[1]
rlabel metal2 24426 1622 24426 1622 0 gfpga_pad_io_soc_out[2]
rlabel metal2 26542 1622 26542 1622 0 gfpga_pad_io_soc_out[3]
rlabel metal2 37122 1588 37122 1588 0 isol_n
rlabel metal1 10396 2550 10396 2550 0 net1
rlabel metal2 1886 10166 1886 10166 0 net10
rlabel metal2 45586 4896 45586 4896 0 net100
rlabel metal2 31786 15164 31786 15164 0 net101
rlabel metal1 33672 13294 33672 13294 0 net102
rlabel metal2 35190 18275 35190 18275 0 net103
rlabel metal1 18262 15674 18262 15674 0 net104
rlabel metal1 16330 17170 16330 17170 0 net105
rlabel via2 13202 15011 13202 15011 0 net106
rlabel metal1 18354 18122 18354 18122 0 net107
rlabel metal2 17434 19533 17434 19533 0 net108
rlabel metal1 40572 21454 40572 21454 0 net109
rlabel metal1 21114 14926 21114 14926 0 net11
rlabel metal1 40848 19482 40848 19482 0 net110
rlabel metal1 39422 2414 39422 2414 0 net111
rlabel metal2 10902 19176 10902 19176 0 net112
rlabel metal1 1794 13328 1794 13328 0 net113
rlabel metal1 1794 18768 1794 18768 0 net114
rlabel metal1 1794 19414 1794 19414 0 net115
rlabel metal1 14582 19992 14582 19992 0 net116
rlabel metal2 1794 19567 1794 19567 0 net117
rlabel metal1 4002 20876 4002 20876 0 net118
rlabel metal1 1794 21556 1794 21556 0 net119
rlabel metal2 12190 9248 12190 9248 0 net12
rlabel metal2 3634 20196 3634 20196 0 net120
rlabel metal1 1794 21930 1794 21930 0 net121
rlabel metal1 2300 22610 2300 22610 0 net122
rlabel metal1 1794 23120 1794 23120 0 net123
rlabel metal1 2277 13906 2277 13906 0 net124
rlabel metal2 4094 21828 4094 21828 0 net125
rlabel metal2 4094 21114 4094 21114 0 net126
rlabel metal2 6026 21556 6026 21556 0 net127
rlabel metal1 6026 20978 6026 20978 0 net128
rlabel metal1 5934 20570 5934 20570 0 net129
rlabel via2 1794 9435 1794 9435 0 net13
rlabel metal1 5934 18734 5934 18734 0 net130
rlabel metal1 6026 19754 6026 19754 0 net131
rlabel metal1 5290 22406 5290 22406 0 net132
rlabel metal1 7084 21386 7084 21386 0 net133
rlabel metal1 7912 22406 7912 22406 0 net134
rlabel metal1 5796 14382 5796 14382 0 net135
rlabel metal2 6670 15164 6670 15164 0 net136
rlabel metal2 10442 15028 10442 15028 0 net137
rlabel metal2 1794 15878 1794 15878 0 net138
rlabel metal2 6854 16796 6854 16796 0 net139
rlabel metal1 12512 2618 12512 2618 0 net14
rlabel metal2 8326 17884 8326 17884 0 net140
rlabel metal2 10534 17204 10534 17204 0 net141
rlabel metal1 2277 18258 2277 18258 0 net142
rlabel metal2 36570 3910 36570 3910 0 net143
rlabel metal1 47794 4590 47794 4590 0 net144
rlabel metal1 47886 5202 47886 5202 0 net145
rlabel metal2 40066 7276 40066 7276 0 net146
rlabel metal1 47840 5678 47840 5678 0 net147
rlabel metal1 47288 6290 47288 6290 0 net148
rlabel metal1 47932 6766 47932 6766 0 net149
rlabel metal2 11914 10268 11914 10268 0 net15
rlabel metal2 42734 9214 42734 9214 0 net150
rlabel metal2 42826 8636 42826 8636 0 net151
rlabel metal2 43746 9180 43746 9180 0 net152
rlabel metal2 46782 9214 46782 9214 0 net153
rlabel metal2 39882 3774 39882 3774 0 net154
rlabel metal2 45770 10540 45770 10540 0 net155
rlabel metal2 44206 10268 44206 10268 0 net156
rlabel metal2 47058 10846 47058 10846 0 net157
rlabel metal2 46690 10812 46690 10812 0 net158
rlabel metal1 47472 10642 47472 10642 0 net159
rlabel metal1 4715 10506 4715 10506 0 net16
rlabel metal2 42734 11934 42734 11934 0 net160
rlabel metal1 46966 11730 46966 11730 0 net161
rlabel metal2 47978 12410 47978 12410 0 net162
rlabel metal1 47518 12818 47518 12818 0 net163
rlabel metal2 46322 13566 46322 13566 0 net164
rlabel metal2 44666 3434 44666 3434 0 net165
rlabel metal2 45862 4318 45862 4318 0 net166
rlabel metal1 46138 3536 46138 3536 0 net167
rlabel metal2 47150 3604 47150 3604 0 net168
rlabel metal2 47242 4454 47242 4454 0 net169
rlabel metal1 4347 10778 4347 10778 0 net17
rlabel metal2 47058 4828 47058 4828 0 net170
rlabel metal1 45816 5202 45816 5202 0 net171
rlabel metal1 47472 4114 47472 4114 0 net172
rlabel metal1 5014 19822 5014 19822 0 net173
rlabel metal1 7452 24174 7452 24174 0 net174
rlabel metal1 8142 23766 8142 23766 0 net175
rlabel metal1 9982 22542 9982 22542 0 net176
rlabel metal1 10764 23698 10764 23698 0 net177
rlabel metal1 10856 21658 10856 21658 0 net178
rlabel metal1 10856 24174 10856 24174 0 net179
rlabel metal1 4347 11254 4347 11254 0 net18
rlabel metal2 12834 22780 12834 22780 0 net180
rlabel metal1 15318 20570 15318 20570 0 net181
rlabel metal1 13662 21862 13662 21862 0 net182
rlabel metal2 13478 23868 13478 23868 0 net183
rlabel metal1 3864 22950 3864 22950 0 net184
rlabel metal1 15134 22678 15134 22678 0 net185
rlabel metal1 17480 19958 17480 19958 0 net186
rlabel metal1 15134 23664 15134 23664 0 net187
rlabel metal1 17618 21964 17618 21964 0 net188
rlabel metal1 15870 24174 15870 24174 0 net189
rlabel metal1 3266 11526 3266 11526 0 net19
rlabel metal1 17940 23698 17940 23698 0 net190
rlabel metal1 20470 21998 20470 21998 0 net191
rlabel metal2 17618 24412 17618 24412 0 net192
rlabel metal1 22448 23290 22448 23290 0 net193
rlabel metal1 20102 24106 20102 24106 0 net194
rlabel metal1 2300 24174 2300 24174 0 net195
rlabel metal1 3266 23698 3266 23698 0 net196
rlabel metal2 4830 23052 4830 23052 0 net197
rlabel metal2 4646 23868 4646 23868 0 net198
rlabel metal1 5382 23018 5382 23018 0 net199
rlabel metal1 47058 23188 47058 23188 0 net2
rlabel metal1 3634 12274 3634 12274 0 net20
rlabel metal2 6578 24004 6578 24004 0 net200
rlabel metal2 7498 23324 7498 23324 0 net201
rlabel metal1 7866 23086 7866 23086 0 net202
rlabel metal1 12282 2414 12282 2414 0 net203
rlabel metal1 15456 2414 15456 2414 0 net204
rlabel metal1 17894 2414 17894 2414 0 net205
rlabel metal1 18354 2958 18354 2958 0 net206
rlabel metal1 20102 2482 20102 2482 0 net207
rlabel metal1 21528 2890 21528 2890 0 net208
rlabel metal2 23138 3026 23138 3026 0 net209
rlabel metal1 4347 11594 4347 11594 0 net21
rlabel metal1 26772 2822 26772 2822 0 net210
rlabel metal1 17572 17850 17572 17850 0 net211
rlabel metal1 24794 14586 24794 14586 0 net212
rlabel metal2 27922 21318 27922 21318 0 net213
rlabel metal1 19182 14042 19182 14042 0 net214
rlabel metal1 23828 19958 23828 19958 0 net215
rlabel metal2 20102 13124 20102 13124 0 net216
rlabel metal1 30084 14382 30084 14382 0 net217
rlabel metal1 31280 7378 31280 7378 0 net218
rlabel metal1 32154 10642 32154 10642 0 net219
rlabel metal1 4370 23086 4370 23086 0 net22
rlabel metal1 33994 15130 33994 15130 0 net220
rlabel metal1 28428 12614 28428 12614 0 net221
rlabel metal2 29946 9350 29946 9350 0 net222
rlabel metal1 30774 7854 30774 7854 0 net223
rlabel metal1 31786 13974 31786 13974 0 net224
rlabel metal1 29256 8942 29256 8942 0 net225
rlabel metal1 27002 11730 27002 11730 0 net226
rlabel metal2 32706 8313 32706 8313 0 net227
rlabel metal2 28842 19652 28842 19652 0 net228
rlabel metal1 30268 15674 30268 15674 0 net229
rlabel metal2 13754 23120 13754 23120 0 net23
rlabel metal1 35742 17306 35742 17306 0 net230
rlabel metal1 35144 15130 35144 15130 0 net231
rlabel metal1 35512 13294 35512 13294 0 net232
rlabel metal1 32430 11798 32430 11798 0 net233
rlabel metal1 32706 21556 32706 21556 0 net234
rlabel metal1 25116 13294 25116 13294 0 net235
rlabel metal1 24058 13838 24058 13838 0 net236
rlabel metal1 23690 10234 23690 10234 0 net237
rlabel metal1 25116 10642 25116 10642 0 net238
rlabel metal1 20102 11322 20102 11322 0 net239
rlabel metal1 14904 16626 14904 16626 0 net24
rlabel metal1 17848 12614 17848 12614 0 net240
rlabel metal1 17158 10642 17158 10642 0 net241
rlabel metal1 19504 10234 19504 10234 0 net242
rlabel metal1 22310 7854 22310 7854 0 net243
rlabel metal1 31004 18258 31004 18258 0 net244
rlabel metal1 12972 13498 12972 13498 0 net245
rlabel metal1 13478 18394 13478 18394 0 net246
rlabel metal1 12098 18632 12098 18632 0 net247
rlabel metal1 10626 18394 10626 18394 0 net248
rlabel metal1 13892 20570 13892 20570 0 net249
rlabel metal1 4370 2414 4370 2414 0 net25
rlabel metal2 12650 21318 12650 21318 0 net250
rlabel metal1 11914 24208 11914 24208 0 net251
rlabel metal1 37352 21114 37352 21114 0 net252
rlabel metal1 40388 19754 40388 19754 0 net253
rlabel metal1 18952 9146 18952 9146 0 net254
rlabel metal1 19228 8466 19228 8466 0 net255
rlabel metal1 11638 13906 11638 13906 0 net256
rlabel metal1 16468 14382 16468 14382 0 net257
rlabel metal1 25944 13294 25944 13294 0 net258
rlabel metal1 21712 12206 21712 12206 0 net259
rlabel metal1 14628 10642 14628 10642 0 net26
rlabel metal1 19320 18734 19320 18734 0 net260
rlabel metal1 19872 20910 19872 20910 0 net261
rlabel metal1 24242 16762 24242 16762 0 net262
rlabel metal1 17112 15334 17112 15334 0 net27
rlabel metal2 16974 6902 16974 6902 0 net28
rlabel metal2 1886 5100 1886 5100 0 net29
rlabel metal1 4991 2550 4991 2550 0 net3
rlabel metal1 4393 4658 4393 4658 0 net30
rlabel metal1 15870 17170 15870 17170 0 net31
rlabel metal1 17204 12070 17204 12070 0 net32
rlabel metal2 48438 14484 48438 14484 0 net33
rlabel metal1 47426 18054 47426 18054 0 net34
rlabel metal2 41446 17799 41446 17799 0 net35
rlabel metal2 48438 18462 48438 18462 0 net36
rlabel metal2 47426 18870 47426 18870 0 net37
rlabel metal2 16514 18819 16514 18819 0 net38
rlabel metal1 45540 20332 45540 20332 0 net39
rlabel metal1 1794 5576 1794 5576 0 net4
rlabel metal2 48438 19992 48438 19992 0 net40
rlabel metal2 43654 21250 43654 21250 0 net41
rlabel metal1 41676 19890 41676 19890 0 net42
rlabel metal2 48714 20621 48714 20621 0 net43
rlabel metal2 48530 14535 48530 14535 0 net44
rlabel metal2 48438 21352 48438 21352 0 net45
rlabel via2 16054 16541 16054 16541 0 net46
rlabel metal1 18630 14246 18630 14246 0 net47
rlabel metal2 19366 19244 19366 19244 0 net48
rlabel metal1 44666 21930 44666 21930 0 net49
rlabel metal1 15962 12818 15962 12818 0 net5
rlabel metal1 44252 22066 44252 22066 0 net50
rlabel metal2 12466 21369 12466 21369 0 net51
rlabel metal1 44988 22202 44988 22202 0 net52
rlabel metal1 43976 22746 43976 22746 0 net53
rlabel metal2 24978 24225 24978 24225 0 net54
rlabel metal2 49266 14297 49266 14297 0 net55
rlabel via2 48346 14875 48346 14875 0 net56
rlabel metal1 49082 15674 49082 15674 0 net57
rlabel metal2 46874 13345 46874 13345 0 net58
rlabel metal2 49266 15929 49266 15929 0 net59
rlabel metal2 2346 10744 2346 10744 0 net6
rlabel metal2 49266 16864 49266 16864 0 net60
rlabel metal2 48438 17442 48438 17442 0 net61
rlabel metal2 47426 17272 47426 17272 0 net62
rlabel metal1 26266 19244 26266 19244 0 net63
rlabel metal1 27600 18394 27600 18394 0 net64
rlabel metal2 31970 18462 31970 18462 0 net65
rlabel metal2 34822 23120 34822 23120 0 net66
rlabel metal2 36570 21624 36570 21624 0 net67
rlabel metal2 32706 20434 32706 20434 0 net68
rlabel metal1 32016 19822 32016 19822 0 net69
rlabel metal2 38778 8381 38778 8381 0 net7
rlabel metal1 35190 19754 35190 19754 0 net70
rlabel metal1 36202 21590 36202 21590 0 net71
rlabel metal1 34178 20910 34178 20910 0 net72
rlabel metal2 29946 20825 29946 20825 0 net73
rlabel via2 12098 21981 12098 21981 0 net74
rlabel metal3 37651 20876 37651 20876 0 net75
rlabel metal1 41308 23630 41308 23630 0 net76
rlabel metal2 32246 18819 32246 18819 0 net77
rlabel metal3 29601 19244 29601 19244 0 net78
rlabel metal3 41561 20332 41561 20332 0 net79
rlabel metal1 4347 7514 4347 7514 0 net8
rlabel metal2 32522 21709 32522 21709 0 net80
rlabel metal1 33994 19822 33994 19822 0 net81
rlabel metal1 35328 19890 35328 19890 0 net82
rlabel metal3 36156 22168 36156 22168 0 net83
rlabel metal2 43286 21624 43286 21624 0 net84
rlabel metal2 26128 19278 26128 19278 0 net85
rlabel metal2 12098 23137 12098 23137 0 net86
rlabel metal1 32108 16218 32108 16218 0 net87
rlabel metal2 32246 14110 32246 14110 0 net88
rlabel metal2 33304 17714 33304 17714 0 net89
rlabel metal1 4347 7718 4347 7718 0 net9
rlabel metal1 32798 18156 32798 18156 0 net90
rlabel metal1 27830 24038 27830 24038 0 net91
rlabel metal1 28796 21318 28796 21318 0 net92
rlabel metal1 28980 2618 28980 2618 0 net93
rlabel metal1 27508 2550 27508 2550 0 net94
rlabel metal1 30866 2278 30866 2278 0 net95
rlabel metal1 34776 2618 34776 2618 0 net96
rlabel metal1 37306 2482 37306 2482 0 net97
rlabel metal2 12282 11628 12282 11628 0 net98
rlabel metal1 43838 2516 43838 2516 0 net99
rlabel metal2 39238 2064 39238 2064 0 prog_clk
rlabel metal1 42412 24174 42412 24174 0 prog_reset_top_in
rlabel metal2 43470 1588 43470 1588 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal2 45586 2132 45586 2132 0 right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal2 47702 2642 47702 2642 0 right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal2 49818 2608 49818 2608 0 right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal1 27876 13362 27876 13362 0 sb_1__0_.mem_left_track_1.ccff_head
rlabel metal1 22678 20332 22678 20332 0 sb_1__0_.mem_left_track_1.ccff_tail
rlabel metal1 28796 13362 28796 13362 0 sb_1__0_.mem_left_track_1.mem_out\[0\]
rlabel metal1 25944 16218 25944 16218 0 sb_1__0_.mem_left_track_1.mem_out\[1\]
rlabel metal2 21390 14994 21390 14994 0 sb_1__0_.mem_left_track_11.ccff_head
rlabel metal1 20424 18190 20424 18190 0 sb_1__0_.mem_left_track_11.ccff_tail
rlabel metal2 21482 12818 21482 12818 0 sb_1__0_.mem_left_track_11.mem_out\[0\]
rlabel metal2 20102 16014 20102 16014 0 sb_1__0_.mem_left_track_11.mem_out\[1\]
rlabel metal1 18860 19890 18860 19890 0 sb_1__0_.mem_left_track_13.ccff_tail
rlabel metal1 21436 18054 21436 18054 0 sb_1__0_.mem_left_track_13.mem_out\[0\]
rlabel metal1 21252 20570 21252 20570 0 sb_1__0_.mem_left_track_13.mem_out\[1\]
rlabel metal1 18078 21556 18078 21556 0 sb_1__0_.mem_left_track_21.ccff_tail
rlabel metal1 25714 22066 25714 22066 0 sb_1__0_.mem_left_track_21.mem_out\[0\]
rlabel metal2 19090 24242 19090 24242 0 sb_1__0_.mem_left_track_21.mem_out\[1\]
rlabel metal2 25162 19686 25162 19686 0 sb_1__0_.mem_left_track_29.ccff_tail
rlabel metal2 24150 17646 24150 17646 0 sb_1__0_.mem_left_track_29.mem_out\[0\]
rlabel metal2 23690 18496 23690 18496 0 sb_1__0_.mem_left_track_29.mem_out\[1\]
rlabel metal2 18814 19686 18814 19686 0 sb_1__0_.mem_left_track_3.ccff_tail
rlabel metal1 21459 19890 21459 19890 0 sb_1__0_.mem_left_track_3.mem_out\[0\]
rlabel metal2 21850 20009 21850 20009 0 sb_1__0_.mem_left_track_3.mem_out\[1\]
rlabel metal2 27370 18632 27370 18632 0 sb_1__0_.mem_left_track_37.ccff_tail
rlabel metal2 32154 19584 32154 19584 0 sb_1__0_.mem_left_track_37.mem_out\[0\]
rlabel metal2 25898 15776 25898 15776 0 sb_1__0_.mem_left_track_37.mem_out\[1\]
rlabel metal1 26312 23154 26312 23154 0 sb_1__0_.mem_left_track_45.ccff_tail
rlabel metal1 32430 22508 32430 22508 0 sb_1__0_.mem_left_track_45.mem_out\[0\]
rlabel metal1 28428 22066 28428 22066 0 sb_1__0_.mem_left_track_45.mem_out\[1\]
rlabel metal2 18906 16286 18906 16286 0 sb_1__0_.mem_left_track_5.ccff_tail
rlabel metal1 20332 21318 20332 21318 0 sb_1__0_.mem_left_track_5.mem_out\[0\]
rlabel metal1 17979 16762 17979 16762 0 sb_1__0_.mem_left_track_5.mem_out\[1\]
rlabel metal1 27462 22984 27462 22984 0 sb_1__0_.mem_left_track_53.mem_out\[0\]
rlabel metal1 21889 21114 21889 21114 0 sb_1__0_.mem_left_track_53.mem_out\[1\]
rlabel metal1 25668 15538 25668 15538 0 sb_1__0_.mem_left_track_7.mem_out\[0\]
rlabel metal2 23782 13923 23782 13923 0 sb_1__0_.mem_left_track_7.mem_out\[1\]
rlabel metal1 18676 18666 18676 18666 0 sb_1__0_.mem_right_track_0.ccff_head
rlabel metal1 32430 17102 32430 17102 0 sb_1__0_.mem_right_track_0.ccff_tail
rlabel via2 33902 13379 33902 13379 0 sb_1__0_.mem_right_track_0.mem_out\[0\]
rlabel metal1 30406 16218 30406 16218 0 sb_1__0_.mem_right_track_0.mem_out\[1\]
rlabel metal1 36524 11526 36524 11526 0 sb_1__0_.mem_right_track_10.ccff_head
rlabel metal1 35788 10234 35788 10234 0 sb_1__0_.mem_right_track_10.ccff_tail
rlabel metal1 33718 19890 33718 19890 0 sb_1__0_.mem_right_track_10.mem_out\[0\]
rlabel metal1 35098 13770 35098 13770 0 sb_1__0_.mem_right_track_10.mem_out\[1\]
rlabel metal2 33902 12818 33902 12818 0 sb_1__0_.mem_right_track_12.ccff_tail
rlabel metal2 32890 17646 32890 17646 0 sb_1__0_.mem_right_track_12.mem_out\[0\]
rlabel metal1 32476 12138 32476 12138 0 sb_1__0_.mem_right_track_12.mem_out\[1\]
rlabel metal1 37030 15674 37030 15674 0 sb_1__0_.mem_right_track_2.ccff_tail
rlabel metal1 33764 20978 33764 20978 0 sb_1__0_.mem_right_track_2.mem_out\[0\]
rlabel metal1 35781 15674 35781 15674 0 sb_1__0_.mem_right_track_2.mem_out\[1\]
rlabel metal2 31786 12104 31786 12104 0 sb_1__0_.mem_right_track_20.ccff_tail
rlabel metal2 31878 13124 31878 13124 0 sb_1__0_.mem_right_track_20.mem_out\[0\]
rlabel metal1 31050 12750 31050 12750 0 sb_1__0_.mem_right_track_20.mem_out\[1\]
rlabel metal1 32430 9486 32430 9486 0 sb_1__0_.mem_right_track_28.ccff_tail
rlabel metal1 30360 14926 30360 14926 0 sb_1__0_.mem_right_track_28.mem_out\[0\]
rlabel metal1 30774 10608 30774 10608 0 sb_1__0_.mem_right_track_28.mem_out\[1\]
rlabel metal2 34086 8772 34086 8772 0 sb_1__0_.mem_right_track_36.ccff_tail
rlabel metal1 31464 14450 31464 14450 0 sb_1__0_.mem_right_track_36.mem_out\[0\]
rlabel metal2 32614 8228 32614 8228 0 sb_1__0_.mem_right_track_36.mem_out\[1\]
rlabel metal1 37996 13362 37996 13362 0 sb_1__0_.mem_right_track_4.ccff_tail
rlabel metal1 36892 15946 36892 15946 0 sb_1__0_.mem_right_track_4.mem_out\[0\]
rlabel metal1 36754 14586 36754 14586 0 sb_1__0_.mem_right_track_4.mem_out\[1\]
rlabel metal2 32430 9724 32430 9724 0 sb_1__0_.mem_right_track_44.ccff_tail
rlabel metal2 29992 15572 29992 15572 0 sb_1__0_.mem_right_track_44.mem_out\[0\]
rlabel metal1 29210 17034 29210 17034 0 sb_1__0_.mem_right_track_52.mem_out\[0\]
rlabel metal1 34408 14450 34408 14450 0 sb_1__0_.mem_right_track_6.mem_out\[0\]
rlabel metal1 36708 12070 36708 12070 0 sb_1__0_.mem_right_track_6.mem_out\[1\]
rlabel metal1 31050 23154 31050 23154 0 sb_1__0_.mem_top_track_0.ccff_tail
rlabel metal2 36478 22593 36478 22593 0 sb_1__0_.mem_top_track_0.mem_out\[0\]
rlabel metal1 32522 22066 32522 22066 0 sb_1__0_.mem_top_track_0.mem_out\[1\]
rlabel metal1 38180 20502 38180 20502 0 sb_1__0_.mem_top_track_10.ccff_head
rlabel metal1 33856 18666 33856 18666 0 sb_1__0_.mem_top_track_10.ccff_tail
rlabel metal1 41814 19958 41814 19958 0 sb_1__0_.mem_top_track_10.mem_out\[0\]
rlabel metal1 37030 19890 37030 19890 0 sb_1__0_.mem_top_track_10.mem_out\[1\]
rlabel metal1 39008 18666 39008 18666 0 sb_1__0_.mem_top_track_12.ccff_tail
rlabel metal1 38725 19142 38725 19142 0 sb_1__0_.mem_top_track_12.mem_out\[0\]
rlabel metal1 37996 18190 37996 18190 0 sb_1__0_.mem_top_track_12.mem_out\[1\]
rlabel metal1 38180 16150 38180 16150 0 sb_1__0_.mem_top_track_14.ccff_tail
rlabel metal2 41814 19074 41814 19074 0 sb_1__0_.mem_top_track_14.mem_out\[0\]
rlabel metal1 37628 16626 37628 16626 0 sb_1__0_.mem_top_track_14.mem_out\[1\]
rlabel metal1 37720 15062 37720 15062 0 sb_1__0_.mem_top_track_16.ccff_tail
rlabel metal1 39330 15878 39330 15878 0 sb_1__0_.mem_top_track_16.mem_out\[0\]
rlabel metal2 41814 15844 41814 15844 0 sb_1__0_.mem_top_track_16.mem_out\[1\]
rlabel metal2 34086 14280 34086 14280 0 sb_1__0_.mem_top_track_18.ccff_tail
rlabel metal2 38318 16864 38318 16864 0 sb_1__0_.mem_top_track_18.mem_out\[0\]
rlabel metal1 39100 14518 39100 14518 0 sb_1__0_.mem_top_track_18.mem_out\[1\]
rlabel metal1 34178 23494 34178 23494 0 sb_1__0_.mem_top_track_2.ccff_tail
rlabel metal1 38272 24242 38272 24242 0 sb_1__0_.mem_top_track_2.mem_out\[0\]
rlabel metal1 35098 22542 35098 22542 0 sb_1__0_.mem_top_track_2.mem_out\[1\]
rlabel metal1 25208 13974 25208 13974 0 sb_1__0_.mem_top_track_20.ccff_tail
rlabel metal2 25530 13600 25530 13600 0 sb_1__0_.mem_top_track_20.mem_out\[0\]
rlabel metal1 25438 12954 25438 12954 0 sb_1__0_.mem_top_track_22.ccff_tail
rlabel metal1 26542 14042 26542 14042 0 sb_1__0_.mem_top_track_22.mem_out\[0\]
rlabel metal1 24426 13362 24426 13362 0 sb_1__0_.mem_top_track_24.ccff_tail
rlabel metal1 27278 15946 27278 15946 0 sb_1__0_.mem_top_track_24.mem_out\[0\]
rlabel metal1 23184 13362 23184 13362 0 sb_1__0_.mem_top_track_26.ccff_tail
rlabel metal1 27278 15538 27278 15538 0 sb_1__0_.mem_top_track_26.mem_out\[0\]
rlabel metal1 21390 11628 21390 11628 0 sb_1__0_.mem_top_track_28.ccff_tail
rlabel metal1 23874 9010 23874 9010 0 sb_1__0_.mem_top_track_28.mem_out\[0\]
rlabel metal1 19872 7786 19872 7786 0 sb_1__0_.mem_top_track_30.ccff_tail
rlabel metal1 21045 8398 21045 8398 0 sb_1__0_.mem_top_track_30.mem_out\[0\]
rlabel metal2 19642 10472 19642 10472 0 sb_1__0_.mem_top_track_32.ccff_tail
rlabel metal2 19734 8466 19734 8466 0 sb_1__0_.mem_top_track_32.mem_out\[0\]
rlabel metal1 21896 10234 21896 10234 0 sb_1__0_.mem_top_track_34.ccff_tail
rlabel metal1 20976 9486 20976 9486 0 sb_1__0_.mem_top_track_34.mem_out\[0\]
rlabel metal1 20286 11288 20286 11288 0 sb_1__0_.mem_top_track_36.ccff_tail
rlabel metal1 22034 11016 22034 11016 0 sb_1__0_.mem_top_track_36.mem_out\[0\]
rlabel metal2 33442 21012 33442 21012 0 sb_1__0_.mem_top_track_4.ccff_tail
rlabel metal1 40618 22100 40618 22100 0 sb_1__0_.mem_top_track_4.mem_out\[0\]
rlabel metal1 32568 20502 32568 20502 0 sb_1__0_.mem_top_track_4.mem_out\[1\]
rlabel metal1 13432 13838 13432 13838 0 sb_1__0_.mem_top_track_40.ccff_tail
rlabel metal1 13340 12750 13340 12750 0 sb_1__0_.mem_top_track_40.mem_out\[0\]
rlabel metal1 15318 18190 15318 18190 0 sb_1__0_.mem_top_track_42.ccff_tail
rlabel metal1 14628 14042 14628 14042 0 sb_1__0_.mem_top_track_42.mem_out\[0\]
rlabel metal1 13294 18802 13294 18802 0 sb_1__0_.mem_top_track_44.ccff_tail
rlabel metal1 16008 18938 16008 18938 0 sb_1__0_.mem_top_track_44.mem_out\[0\]
rlabel metal1 12328 17850 12328 17850 0 sb_1__0_.mem_top_track_46.ccff_tail
rlabel metal2 12742 17782 12742 17782 0 sb_1__0_.mem_top_track_46.mem_out\[0\]
rlabel metal2 14858 20978 14858 20978 0 sb_1__0_.mem_top_track_48.ccff_tail
rlabel metal1 13800 19686 13800 19686 0 sb_1__0_.mem_top_track_48.mem_out\[0\]
rlabel metal1 13662 21488 13662 21488 0 sb_1__0_.mem_top_track_50.ccff_tail
rlabel metal2 16330 20604 16330 20604 0 sb_1__0_.mem_top_track_50.mem_out\[0\]
rlabel metal1 17480 23018 17480 23018 0 sb_1__0_.mem_top_track_58.mem_out\[0\]
rlabel metal1 38870 23290 38870 23290 0 sb_1__0_.mem_top_track_6.ccff_tail
rlabel metal1 36340 21658 36340 21658 0 sb_1__0_.mem_top_track_6.mem_out\[0\]
rlabel metal1 37168 23018 37168 23018 0 sb_1__0_.mem_top_track_6.mem_out\[1\]
rlabel metal1 41814 21012 41814 21012 0 sb_1__0_.mem_top_track_8.mem_out\[0\]
rlabel metal2 39238 21148 39238 21148 0 sb_1__0_.mem_top_track_8.mem_out\[1\]
rlabel metal1 6854 22644 6854 22644 0 sb_1__0_.mux_left_track_1.out
rlabel metal1 26358 18292 26358 18292 0 sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 26772 18394 26772 18394 0 sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 22678 13770 22678 13770 0 sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 22724 14994 22724 14994 0 sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 24840 18122 24840 18122 0 sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 22770 15130 22770 15130 0 sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 21942 19040 21942 19040 0 sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 7360 16218 7360 16218 0 sb_1__0_.mux_left_track_11.out
rlabel metal1 25714 18258 25714 18258 0 sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 25438 18394 25438 18394 0 sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 20930 14246 20930 14246 0 sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 20378 15062 20378 15062 0 sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 21712 18394 21712 18394 0 sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 19550 16694 19550 16694 0 sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 13984 16558 13984 16558 0 sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 15686 16218 15686 16218 0 sb_1__0_.mux_left_track_13.out
rlabel metal2 23782 21114 23782 21114 0 sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 24242 20910 24242 20910 0 sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20838 15674 20838 15674 0 sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 18630 19958 18630 19958 0 sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 19182 18938 19182 18938 0 sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 15870 18802 15870 18802 0 sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 8832 23222 8832 23222 0 sb_1__0_.mux_left_track_21.out
rlabel via2 27922 23307 27922 23307 0 sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 24058 21862 24058 21862 0 sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 22034 19414 22034 19414 0 sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 17848 21658 17848 21658 0 sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 19320 21046 19320 21046 0 sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 10074 23188 10074 23188 0 sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 15502 15674 15502 15674 0 sb_1__0_.mux_left_track_29.out
rlabel metal1 27416 19822 27416 19822 0 sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 26220 19754 26220 19754 0 sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 23966 15130 23966 15130 0 sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 24426 19686 24426 19686 0 sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 23092 17850 23092 17850 0 sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 15686 18003 15686 18003 0 sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 10534 20570 10534 20570 0 sb_1__0_.mux_left_track_3.out
rlabel metal1 22126 21930 22126 21930 0 sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 24610 20502 24610 20502 0 sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20378 21862 20378 21862 0 sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 17618 18938 17618 18938 0 sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 16882 19890 16882 19890 0 sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 17848 15334 17848 15334 0 sb_1__0_.mux_left_track_37.out
rlabel metal2 29026 19142 29026 19142 0 sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 29302 18394 29302 18394 0 sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 23782 16660 23782 16660 0 sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 25162 15810 25162 15810 0 sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 22862 15946 22862 15946 0 sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 8050 18734 8050 18734 0 sb_1__0_.mux_left_track_45.out
rlabel metal1 29578 21930 29578 21930 0 sb_1__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 28060 22202 28060 22202 0 sb_1__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 28106 21658 28106 21658 0 sb_1__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 11178 20961 11178 20961 0 sb_1__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 5750 22610 5750 22610 0 sb_1__0_.mux_left_track_5.out
rlabel metal1 21574 18870 21574 18870 0 sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 24564 17850 24564 17850 0 sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 17940 16014 17940 16014 0 sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 18124 14042 18124 14042 0 sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 16100 15878 16100 15878 0 sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_4_X
rlabel via2 16514 20757 16514 20757 0 sb_1__0_.mux_left_track_53.out
rlabel metal3 28382 22236 28382 22236 0 sb_1__0_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22586 19482 22586 19482 0 sb_1__0_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21344 19346 21344 19346 0 sb_1__0_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 20792 19482 20792 19482 0 sb_1__0_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 9522 17884 9522 17884 0 sb_1__0_.mux_left_track_7.out
rlabel metal1 24150 15470 24150 15470 0 sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 23506 15368 23506 15368 0 sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 20194 12585 20194 12585 0 sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 21229 15402 21229 15402 0 sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 19872 12954 19872 12954 0 sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 19550 15674 19550 15674 0 sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 45034 14110 45034 14110 0 sb_1__0_.mux_right_track_0.out
rlabel metal1 31050 17102 31050 17102 0 sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 33626 13498 33626 13498 0 sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 29026 14314 29026 14314 0 sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 33994 16490 33994 16490 0 sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 33350 15334 33350 15334 0 sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 39514 14484 39514 14484 0 sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 45540 11152 45540 11152 0 sb_1__0_.mux_right_track_10.out
rlabel metal1 34868 13838 34868 13838 0 sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 34868 14042 34868 14042 0 sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 35328 9146 35328 9146 0 sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 32706 10302 32706 10302 0 sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 37582 13124 37582 13124 0 sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 37858 10234 37858 10234 0 sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 39238 10234 39238 10234 0 sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal2 40250 11934 40250 11934 0 sb_1__0_.mux_right_track_12.out
rlabel metal1 32706 15062 32706 15062 0 sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 32522 15130 32522 15130 0 sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 32292 10574 32292 10574 0 sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 36064 12954 36064 12954 0 sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 33120 10506 33120 10506 0 sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 39330 12444 39330 12444 0 sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 45862 14348 45862 14348 0 sb_1__0_.mux_right_track_2.out
rlabel metal2 36294 19754 36294 19754 0 sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 34270 18394 34270 18394 0 sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 29486 14807 29486 14807 0 sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 38502 17884 38502 17884 0 sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 33626 15130 33626 15130 0 sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 40986 14994 40986 14994 0 sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 43516 10030 43516 10030 0 sb_1__0_.mux_right_track_20.out
rlabel metal2 31142 18224 31142 18224 0 sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 31004 16218 31004 16218 0 sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 29164 12954 29164 12954 0 sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 32522 14450 32522 14450 0 sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 30314 12682 30314 12682 0 sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 32384 14246 32384 14246 0 sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 44298 8670 44298 8670 0 sb_1__0_.mux_right_track_28.out
rlabel metal1 30038 13362 30038 13362 0 sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 29946 13294 29946 13294 0 sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 25714 9656 25714 9656 0 sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 32798 9554 32798 9554 0 sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 32614 9622 32614 9622 0 sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 37858 8976 37858 8976 0 sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 40158 7888 40158 7888 0 sb_1__0_.mux_right_track_36.out
rlabel metal2 33810 10999 33810 10999 0 sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 33672 11050 33672 11050 0 sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 34914 9010 34914 9010 0 sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 35282 8432 35282 8432 0 sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 39146 8500 39146 8500 0 sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 46138 12988 46138 12988 0 sb_1__0_.mux_right_track_4.out
rlabel metal1 36754 16660 36754 16660 0 sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 36340 16558 36340 16558 0 sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 36110 13838 36110 13838 0 sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 37122 13974 37122 13974 0 sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 36800 14042 36800 14042 0 sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 41538 13668 41538 13668 0 sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 40250 7480 40250 7480 0 sb_1__0_.mux_right_track_44.out
rlabel metal1 32338 16490 32338 16490 0 sb_1__0_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 32706 9520 32706 9520 0 sb_1__0_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 36018 8466 36018 8466 0 sb_1__0_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 43746 6289 43746 6289 0 sb_1__0_.mux_right_track_52.out
rlabel metal1 29486 11186 29486 11186 0 sb_1__0_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 29348 11050 29348 11050 0 sb_1__0_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 32798 11271 32798 11271 0 sb_1__0_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 45540 12274 45540 12274 0 sb_1__0_.mux_right_track_6.out
rlabel metal1 36570 15062 36570 15062 0 sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 33442 14790 33442 14790 0 sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 36570 10778 36570 10778 0 sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 35374 7990 35374 7990 0 sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 36616 14790 36616 14790 0 sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 37904 11866 37904 11866 0 sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 41446 12240 41446 12240 0 sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 19642 24276 19642 24276 0 sb_1__0_.mux_top_track_0.out
rlabel metal1 36156 22746 36156 22746 0 sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 39836 22474 39836 22474 0 sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 26726 20842 26726 20842 0 sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 28612 19482 28612 19482 0 sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 30268 23154 30268 23154 0 sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 29256 21114 29256 21114 0 sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 29762 23460 29762 23460 0 sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 26864 21658 26864 21658 0 sb_1__0_.mux_top_track_10.out
rlabel metal1 35650 19482 35650 19482 0 sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 39974 19584 39974 19584 0 sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 36064 19686 36064 19686 0 sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 31878 17544 31878 17544 0 sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 30636 18938 30636 18938 0 sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 26450 23528 26450 23528 0 sb_1__0_.mux_top_track_12.out
rlabel metal2 40894 19312 40894 19312 0 sb_1__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 40434 18360 40434 18360 0 sb_1__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 36064 17034 36064 17034 0 sb_1__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 33902 20264 33902 20264 0 sb_1__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 20838 22950 20838 22950 0 sb_1__0_.mux_top_track_14.out
rlabel metal1 40572 17714 40572 17714 0 sb_1__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 38870 17850 38870 17850 0 sb_1__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 35696 14858 35696 14858 0 sb_1__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 35926 19278 35926 19278 0 sb_1__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 21344 19686 21344 19686 0 sb_1__0_.mux_top_track_16.out
rlabel metal2 40986 17952 40986 17952 0 sb_1__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 39698 16218 39698 16218 0 sb_1__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 36662 13498 36662 13498 0 sb_1__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 36984 17306 36984 17306 0 sb_1__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 21666 19652 21666 19652 0 sb_1__0_.mux_top_track_18.out
rlabel metal1 40112 15130 40112 15130 0 sb_1__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 32522 15028 32522 15028 0 sb_1__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 32062 14756 32062 14756 0 sb_1__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 30590 14790 30590 14790 0 sb_1__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 23920 23086 23920 23086 0 sb_1__0_.mux_top_track_2.out
rlabel metal1 38318 23834 38318 23834 0 sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 40066 23528 40066 23528 0 sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 32614 21896 32614 21896 0 sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 37214 23562 37214 23562 0 sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 32890 21862 32890 21862 0 sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 29394 23766 29394 23766 0 sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 15594 17238 15594 17238 0 sb_1__0_.mux_top_track_20.out
rlabel metal1 26404 17306 26404 17306 0 sb_1__0_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 25116 13498 25116 13498 0 sb_1__0_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 23828 17306 23828 17306 0 sb_1__0_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 19964 16422 19964 16422 0 sb_1__0_.mux_top_track_22.out
rlabel metal1 24702 15674 24702 15674 0 sb_1__0_.mux_top_track_22.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 23368 12070 23368 12070 0 sb_1__0_.mux_top_track_22.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 20286 16388 20286 16388 0 sb_1__0_.mux_top_track_22.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 16146 19414 16146 19414 0 sb_1__0_.mux_top_track_24.out
rlabel metal1 23828 13362 23828 13362 0 sb_1__0_.mux_top_track_24.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 23598 13158 23598 13158 0 sb_1__0_.mux_top_track_24.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21022 13770 21022 13770 0 sb_1__0_.mux_top_track_24.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 17710 17782 17710 17782 0 sb_1__0_.mux_top_track_26.out
rlabel metal1 22586 13396 22586 13396 0 sb_1__0_.mux_top_track_26.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 23368 13226 23368 13226 0 sb_1__0_.mux_top_track_26.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21850 17544 21850 17544 0 sb_1__0_.mux_top_track_26.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 15502 19856 15502 19856 0 sb_1__0_.mux_top_track_28.out
rlabel metal1 24242 9078 24242 9078 0 sb_1__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20700 11526 20700 11526 0 sb_1__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 13064 17782 13064 17782 0 sb_1__0_.mux_top_track_30.out
rlabel metal1 21620 7514 21620 7514 0 sb_1__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal3 14582 12580 14582 12580 0 sb_1__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 12880 17850 12880 17850 0 sb_1__0_.mux_top_track_32.out
rlabel metal2 18998 10914 18998 10914 0 sb_1__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 14904 17510 14904 17510 0 sb_1__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 12190 22542 12190 22542 0 sb_1__0_.mux_top_track_34.out
rlabel metal1 20056 12818 20056 12818 0 sb_1__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17572 12954 17572 12954 0 sb_1__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 15364 19482 15364 19482 0 sb_1__0_.mux_top_track_36.out
rlabel metal1 21206 12716 21206 12716 0 sb_1__0_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21528 12818 21528 12818 0 sb_1__0_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19826 12682 19826 12682 0 sb_1__0_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 27186 23086 27186 23086 0 sb_1__0_.mux_top_track_4.out
rlabel metal1 35190 20570 35190 20570 0 sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 40066 21896 40066 21896 0 sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 35098 21862 35098 21862 0 sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 30682 18394 30682 18394 0 sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 30590 21114 30590 21114 0 sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 9798 19380 9798 19380 0 sb_1__0_.mux_top_track_40.out
rlabel metal1 12696 10234 12696 10234 0 sb_1__0_.mux_top_track_40.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 11546 14586 11546 14586 0 sb_1__0_.mux_top_track_40.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 6831 24174 6831 24174 0 sb_1__0_.mux_top_track_42.out
rlabel metal2 16790 16898 16790 16898 0 sb_1__0_.mux_top_track_42.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13938 18156 13938 18156 0 sb_1__0_.mux_top_track_42.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 7038 23698 7038 23698 0 sb_1__0_.mux_top_track_44.out
rlabel metal2 15594 17952 15594 17952 0 sb_1__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 12190 19312 12190 19312 0 sb_1__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_1_X
rlabel via1 5474 23035 5474 23035 0 sb_1__0_.mux_top_track_46.out
rlabel metal1 11684 15130 11684 15130 0 sb_1__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 10258 18122 10258 18122 0 sb_1__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 4462 24174 4462 24174 0 sb_1__0_.mux_top_track_48.out
rlabel metal1 16836 18394 16836 18394 0 sb_1__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 12650 20264 12650 20264 0 sb_1__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 8556 23630 8556 23630 0 sb_1__0_.mux_top_track_50.out
rlabel metal1 16698 20026 16698 20026 0 sb_1__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 11270 20944 11270 20944 0 sb_1__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 9200 23086 9200 23086 0 sb_1__0_.mux_top_track_58.out
rlabel metal1 17250 18836 17250 18836 0 sb_1__0_.mux_top_track_58.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 9706 23834 9706 23834 0 sb_1__0_.mux_top_track_58.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 21482 24140 21482 24140 0 sb_1__0_.mux_top_track_6.out
rlabel metal1 40204 21658 40204 21658 0 sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 40664 22202 40664 22202 0 sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 32752 18938 32752 18938 0 sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 39698 23528 39698 23528 0 sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 35052 23834 35052 23834 0 sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 33626 24072 33626 24072 0 sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_5_X
rlabel via2 31510 22389 31510 22389 0 sb_1__0_.mux_top_track_8.out
rlabel metal1 40020 23494 40020 23494 0 sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 40848 20774 40848 20774 0 sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 33534 19720 33534 19720 0 sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 39422 21114 39422 21114 0 sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 38962 20026 38962 20026 0 sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 35466 23137 35466 23137 0 sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 45770 24174 45770 24174 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_
rlabel metal1 46414 24174 46414 24174 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_
rlabel metal2 46874 25041 46874 25041 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_
rlabel metal1 47748 24174 47748 24174 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_
rlabel metal1 48024 23766 48024 23766 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_
rlabel metal2 48806 25007 48806 25007 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_
rlabel metal1 44620 23086 44620 23086 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_
rlabel metal1 45034 24174 45034 24174 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_
rlabel metal2 1150 2115 1150 2115 0 top_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal2 3266 1299 3266 1299 0 top_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal2 5382 2183 5382 2183 0 top_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal2 7498 1962 7498 1962 0 top_width_0_height_0_subtile_3__pin_inpad_0_
<< properties >>
string FIXED_BBOX 0 0 51000 27000
<< end >>
