magic
tech sky130A
magscale 1 2
timestamp 1656240930
<< viali >>
rect 4997 14569 5031 14603
rect 6469 14569 6503 14603
rect 10609 14569 10643 14603
rect 18337 14569 18371 14603
rect 2237 14433 2271 14467
rect 3157 14433 3191 14467
rect 4629 14433 4663 14467
rect 5181 14433 5215 14467
rect 8769 14433 8803 14467
rect 10333 14433 10367 14467
rect 13921 14433 13955 14467
rect 14197 14433 14231 14467
rect 1961 14365 1995 14399
rect 2881 14365 2915 14399
rect 3525 14365 3559 14399
rect 4353 14365 4387 14399
rect 4905 14365 4939 14399
rect 6653 14365 6687 14399
rect 10077 14365 10111 14399
rect 10425 14365 10459 14399
rect 10977 14365 11011 14399
rect 11253 14365 11287 14399
rect 12909 14365 12943 14399
rect 13645 14365 13679 14399
rect 14381 14365 14415 14399
rect 14657 14365 14691 14399
rect 16313 14365 16347 14399
rect 16681 14365 16715 14399
rect 16948 14365 16982 14399
rect 5549 14297 5583 14331
rect 12664 14297 12698 14331
rect 16046 14297 16080 14331
rect 18429 14297 18463 14331
rect 3341 14229 3375 14263
rect 4721 14229 4755 14263
rect 5365 14229 5399 14263
rect 8953 14229 8987 14263
rect 11161 14229 11195 14263
rect 11529 14229 11563 14263
rect 14933 14229 14967 14263
rect 16405 14229 16439 14263
rect 18061 14229 18095 14263
rect 4169 14025 4203 14059
rect 4445 14025 4479 14059
rect 4905 14025 4939 14059
rect 8217 14025 8251 14059
rect 9873 14025 9907 14059
rect 15117 14025 15151 14059
rect 5549 13957 5583 13991
rect 8576 13957 8610 13991
rect 14841 13957 14875 13991
rect 16230 13957 16264 13991
rect 1961 13889 1995 13923
rect 2237 13889 2271 13923
rect 2881 13889 2915 13923
rect 3525 13889 3559 13923
rect 3617 13889 3651 13923
rect 4353 13889 4387 13923
rect 4629 13889 4663 13923
rect 4721 13889 4755 13923
rect 5089 13889 5123 13923
rect 5273 13889 5307 13923
rect 6837 13889 6871 13923
rect 7104 13889 7138 13923
rect 11078 13889 11112 13923
rect 11345 13889 11379 13923
rect 12642 13889 12676 13923
rect 13349 13889 13383 13923
rect 16497 13889 16531 13923
rect 16681 13889 16715 13923
rect 16937 13889 16971 13923
rect 18429 13889 18463 13923
rect 3157 13821 3191 13855
rect 3341 13821 3375 13855
rect 5365 13821 5399 13855
rect 8309 13821 8343 13855
rect 12909 13821 12943 13855
rect 13093 13821 13127 13855
rect 14657 13821 14691 13855
rect 18245 13821 18279 13855
rect 9965 13753 9999 13787
rect 11529 13753 11563 13787
rect 14473 13753 14507 13787
rect 3985 13685 4019 13719
rect 9689 13685 9723 13719
rect 18061 13685 18095 13719
rect 3065 13481 3099 13515
rect 5549 13481 5583 13515
rect 11805 13481 11839 13515
rect 18337 13481 18371 13515
rect 3249 13413 3283 13447
rect 1961 13345 1995 13379
rect 2513 13345 2547 13379
rect 4537 13345 4571 13379
rect 12081 13345 12115 13379
rect 17141 13345 17175 13379
rect 17601 13345 17635 13379
rect 2237 13277 2271 13311
rect 3433 13277 3467 13311
rect 4077 13277 4111 13311
rect 4169 13277 4203 13311
rect 5181 13277 5215 13311
rect 8769 13277 8803 13311
rect 11621 13277 11655 13311
rect 13654 13277 13688 13311
rect 13921 13277 13955 13311
rect 15218 13277 15252 13311
rect 15485 13277 15519 13311
rect 17233 13277 17267 13311
rect 18521 13277 18555 13311
rect 2605 13209 2639 13243
rect 8502 13209 8536 13243
rect 11354 13209 11388 13243
rect 11989 13209 12023 13243
rect 12265 13209 12299 13243
rect 15577 13209 15611 13243
rect 16874 13209 16908 13243
rect 2697 13141 2731 13175
rect 3525 13141 3559 13175
rect 3893 13141 3927 13175
rect 4353 13141 4387 13175
rect 4997 13141 5031 13175
rect 5273 13141 5307 13175
rect 7389 13141 7423 13175
rect 10241 13141 10275 13175
rect 12541 13141 12575 13175
rect 14105 13141 14139 13175
rect 15761 13141 15795 13175
rect 2329 12937 2363 12971
rect 2789 12937 2823 12971
rect 3525 12937 3559 12971
rect 3985 12937 4019 12971
rect 4353 12937 4387 12971
rect 4813 12937 4847 12971
rect 10977 12937 11011 12971
rect 11345 12937 11379 12971
rect 2697 12869 2731 12903
rect 5825 12869 5859 12903
rect 9842 12869 9876 12903
rect 16497 12869 16531 12903
rect 18245 12869 18279 12903
rect 18429 12869 18463 12903
rect 3433 12801 3467 12835
rect 4997 12801 5031 12835
rect 5273 12801 5307 12835
rect 5549 12801 5583 12835
rect 5641 12801 5675 12835
rect 9249 12801 9283 12835
rect 9505 12801 9539 12835
rect 9597 12801 9631 12835
rect 12642 12801 12676 12835
rect 12909 12801 12943 12835
rect 13185 12801 13219 12835
rect 14585 12801 14619 12835
rect 14841 12801 14875 12835
rect 16046 12801 16080 12835
rect 16681 12801 16715 12835
rect 16948 12801 16982 12835
rect 1961 12733 1995 12767
rect 2237 12733 2271 12767
rect 2973 12733 3007 12767
rect 3249 12733 3283 12767
rect 4445 12733 4479 12767
rect 4629 12733 4663 12767
rect 16313 12733 16347 12767
rect 8125 12665 8159 12699
rect 13461 12665 13495 12699
rect 3893 12597 3927 12631
rect 5089 12597 5123 12631
rect 5365 12597 5399 12631
rect 11529 12597 11563 12631
rect 13093 12597 13127 12631
rect 14933 12597 14967 12631
rect 18061 12597 18095 12631
rect 3433 12393 3467 12427
rect 3617 12393 3651 12427
rect 4537 12393 4571 12427
rect 4629 12393 4663 12427
rect 13461 12393 13495 12427
rect 14105 12393 14139 12427
rect 15761 12393 15795 12427
rect 5549 12325 5583 12359
rect 10057 12325 10091 12359
rect 13829 12325 13863 12359
rect 2881 12257 2915 12291
rect 3985 12257 4019 12291
rect 5273 12257 5307 12291
rect 11437 12257 11471 12291
rect 11529 12257 11563 12291
rect 17141 12257 17175 12291
rect 17969 12257 18003 12291
rect 1961 12189 1995 12223
rect 2237 12189 2271 12223
rect 3157 12189 3191 12223
rect 3249 12189 3283 12223
rect 4169 12189 4203 12223
rect 4997 12189 5031 12223
rect 6009 12189 6043 12223
rect 11796 12189 11830 12223
rect 15218 12189 15252 12223
rect 15485 12189 15519 12223
rect 17693 12189 17727 12223
rect 5825 12121 5859 12155
rect 11192 12121 11226 12155
rect 13553 12121 13587 12155
rect 16874 12121 16908 12155
rect 17509 12121 17543 12155
rect 4077 12053 4111 12087
rect 5089 12053 5123 12087
rect 5641 12053 5675 12087
rect 12909 12053 12943 12087
rect 13093 12053 13127 12087
rect 13277 12053 13311 12087
rect 17417 12053 17451 12087
rect 3065 11849 3099 11883
rect 3341 11849 3375 11883
rect 5641 11849 5675 11883
rect 8585 11849 8619 11883
rect 10057 11849 10091 11883
rect 13553 11849 13587 11883
rect 4169 11781 4203 11815
rect 8922 11781 8956 11815
rect 18245 11781 18279 11815
rect 18429 11781 18463 11815
rect 2605 11713 2639 11747
rect 2697 11713 2731 11747
rect 3157 11713 3191 11747
rect 4261 11713 4295 11747
rect 5089 11713 5123 11747
rect 5825 11713 5859 11747
rect 7205 11713 7239 11747
rect 7461 11713 7495 11747
rect 8677 11713 8711 11747
rect 13194 11713 13228 11747
rect 13461 11713 13495 11747
rect 14666 11713 14700 11747
rect 14933 11713 14967 11747
rect 16138 11713 16172 11747
rect 16405 11713 16439 11747
rect 17805 11713 17839 11747
rect 18061 11713 18095 11747
rect 1961 11645 1995 11679
rect 2237 11645 2271 11679
rect 2513 11645 2547 11679
rect 3617 11645 3651 11679
rect 3985 11645 4019 11679
rect 5181 11645 5215 11679
rect 5365 11645 5399 11679
rect 5917 11577 5951 11611
rect 11897 11577 11931 11611
rect 3525 11509 3559 11543
rect 4629 11509 4663 11543
rect 4721 11509 4755 11543
rect 11621 11509 11655 11543
rect 12081 11509 12115 11543
rect 15025 11509 15059 11543
rect 16681 11509 16715 11543
rect 2881 11305 2915 11339
rect 6193 11305 6227 11339
rect 10885 11305 10919 11339
rect 14381 11305 14415 11339
rect 2605 11237 2639 11271
rect 2789 11237 2823 11271
rect 4813 11237 4847 11271
rect 8953 11237 8987 11271
rect 14473 11237 14507 11271
rect 15945 11237 15979 11271
rect 17601 11237 17635 11271
rect 1961 11169 1995 11203
rect 3525 11169 3559 11203
rect 4261 11169 4295 11203
rect 5549 11169 5583 11203
rect 2237 11101 2271 11135
rect 3249 11101 3283 11135
rect 4353 11101 4387 11135
rect 5733 11101 5767 11135
rect 10333 11101 10367 11135
rect 12265 11101 12299 11135
rect 12357 11101 12391 11135
rect 13921 11101 13955 11135
rect 15853 11101 15887 11135
rect 17325 11101 17359 11135
rect 17417 11101 17451 11135
rect 17693 11101 17727 11135
rect 17969 11101 18003 11135
rect 2421 11033 2455 11067
rect 5089 11033 5123 11067
rect 10066 11033 10100 11067
rect 11998 11033 12032 11067
rect 12624 11033 12658 11067
rect 14197 11033 14231 11067
rect 15586 11033 15620 11067
rect 17080 11033 17114 11067
rect 3341 10965 3375 10999
rect 3893 10965 3927 10999
rect 4445 10965 4479 10999
rect 4997 10965 5031 10999
rect 5641 10965 5675 10999
rect 6101 10965 6135 10999
rect 13737 10965 13771 10999
rect 3525 10761 3559 10795
rect 4813 10761 4847 10795
rect 6193 10761 6227 10795
rect 6837 10761 6871 10795
rect 9413 10761 9447 10795
rect 16681 10761 16715 10795
rect 2605 10693 2639 10727
rect 3065 10693 3099 10727
rect 15577 10693 15611 10727
rect 17509 10693 17543 10727
rect 2421 10625 2455 10659
rect 3157 10625 3191 10659
rect 3985 10625 4019 10659
rect 5733 10625 5767 10659
rect 5825 10625 5859 10659
rect 6745 10625 6779 10659
rect 8300 10625 8334 10659
rect 11078 10625 11112 10659
rect 11345 10625 11379 10659
rect 13654 10625 13688 10659
rect 13921 10625 13955 10659
rect 15126 10625 15160 10659
rect 15393 10625 15427 10659
rect 16037 10625 16071 10659
rect 16313 10625 16347 10659
rect 16865 10625 16899 10659
rect 17141 10625 17175 10659
rect 1961 10557 1995 10591
rect 2237 10557 2271 10591
rect 2881 10557 2915 10591
rect 3709 10557 3743 10591
rect 3893 10557 3927 10591
rect 4905 10557 4939 10591
rect 5089 10557 5123 10591
rect 5641 10557 5675 10591
rect 7021 10557 7055 10591
rect 8033 10557 8067 10591
rect 15761 10557 15795 10591
rect 17693 10557 17727 10591
rect 17969 10557 18003 10591
rect 4353 10489 4387 10523
rect 16497 10489 16531 10523
rect 16957 10489 16991 10523
rect 4445 10421 4479 10455
rect 5273 10421 5307 10455
rect 6377 10421 6411 10455
rect 9965 10421 9999 10455
rect 12541 10421 12575 10455
rect 14013 10421 14047 10455
rect 15945 10421 15979 10455
rect 16221 10421 16255 10455
rect 17417 10421 17451 10455
rect 4169 10217 4203 10251
rect 13369 10217 13403 10251
rect 14473 10217 14507 10251
rect 4997 10149 5031 10183
rect 5273 10149 5307 10183
rect 13461 10149 13495 10183
rect 14565 10149 14599 10183
rect 16037 10149 16071 10183
rect 17601 10149 17635 10183
rect 2513 10081 2547 10115
rect 2605 10081 2639 10115
rect 3893 10081 3927 10115
rect 4721 10081 4755 10115
rect 5549 10081 5583 10115
rect 6377 10081 6411 10115
rect 11989 10081 12023 10115
rect 17969 10081 18003 10115
rect 1409 10013 1443 10047
rect 1685 10013 1719 10047
rect 3157 10013 3191 10047
rect 4537 10013 4571 10047
rect 6561 10013 6595 10047
rect 7389 10013 7423 10047
rect 7656 10013 7690 10047
rect 10149 10013 10183 10047
rect 10405 10013 10439 10047
rect 14289 10013 14323 10047
rect 15945 10013 15979 10047
rect 17417 10013 17451 10047
rect 17693 10013 17727 10047
rect 5641 9945 5675 9979
rect 12234 9945 12268 9979
rect 13737 9945 13771 9979
rect 15678 9945 15712 9979
rect 17150 9945 17184 9979
rect 2697 9877 2731 9911
rect 3065 9877 3099 9911
rect 3341 9877 3375 9911
rect 3617 9877 3651 9911
rect 4629 9877 4663 9911
rect 5733 9877 5767 9911
rect 6101 9877 6135 9911
rect 6469 9877 6503 9911
rect 6929 9877 6963 9911
rect 8769 9877 8803 9911
rect 11529 9877 11563 9911
rect 13921 9877 13955 9911
rect 3249 9673 3283 9707
rect 4077 9673 4111 9707
rect 4445 9673 4479 9707
rect 4537 9673 4571 9707
rect 4997 9673 5031 9707
rect 6377 9673 6411 9707
rect 16773 9673 16807 9707
rect 17693 9673 17727 9707
rect 18061 9673 18095 9707
rect 5825 9605 5859 9639
rect 6745 9605 6779 9639
rect 11078 9605 11112 9639
rect 11713 9605 11747 9639
rect 13820 9605 13854 9639
rect 18429 9605 18463 9639
rect 2237 9537 2271 9571
rect 3433 9537 3467 9571
rect 3985 9537 4019 9571
rect 4905 9537 4939 9571
rect 5457 9537 5491 9571
rect 9054 9537 9088 9571
rect 9321 9537 9355 9571
rect 11345 9537 11379 9571
rect 12081 9537 12115 9571
rect 12337 9537 12371 9571
rect 16138 9537 16172 9571
rect 17141 9537 17175 9571
rect 17601 9537 17635 9571
rect 1961 9469 1995 9503
rect 2881 9469 2915 9503
rect 3157 9469 3191 9503
rect 3893 9469 3927 9503
rect 5181 9469 5215 9503
rect 6837 9469 6871 9503
rect 7021 9469 7055 9503
rect 9689 9469 9723 9503
rect 11897 9469 11931 9503
rect 13553 9469 13587 9503
rect 16405 9469 16439 9503
rect 17877 9469 17911 9503
rect 5549 9401 5583 9435
rect 7941 9401 7975 9435
rect 11529 9401 11563 9435
rect 17233 9401 17267 9435
rect 3617 9333 3651 9367
rect 9965 9333 9999 9367
rect 13461 9333 13495 9367
rect 14933 9333 14967 9367
rect 15025 9333 15059 9367
rect 16957 9333 16991 9367
rect 18337 9333 18371 9367
rect 3801 9129 3835 9163
rect 4721 9129 4755 9163
rect 7021 9129 7055 9163
rect 13369 9129 13403 9163
rect 16957 9129 16991 9163
rect 3065 9061 3099 9095
rect 10333 9061 10367 9095
rect 2513 8993 2547 9027
rect 2605 8993 2639 9027
rect 4445 8993 4479 9027
rect 5917 8993 5951 9027
rect 6469 8993 6503 9027
rect 11805 8993 11839 9027
rect 11989 8993 12023 9027
rect 13829 8993 13863 9027
rect 17049 8993 17083 9027
rect 1961 8925 1995 8959
rect 2237 8925 2271 8959
rect 3433 8925 3467 8959
rect 4169 8925 4203 8959
rect 5733 8925 5767 8959
rect 7389 8925 7423 8959
rect 7645 8925 7679 8959
rect 8953 8925 8987 8959
rect 14105 8925 14139 8959
rect 15577 8925 15611 8959
rect 3249 8857 3283 8891
rect 3525 8857 3559 8891
rect 4997 8857 5031 8891
rect 5641 8857 5675 8891
rect 9198 8857 9232 8891
rect 11538 8857 11572 8891
rect 12234 8857 12268 8891
rect 14350 8857 14384 8891
rect 15822 8857 15856 8891
rect 17294 8857 17328 8891
rect 2697 8789 2731 8823
rect 4261 8789 4295 8823
rect 4905 8789 4939 8823
rect 5273 8789 5307 8823
rect 6101 8789 6135 8823
rect 6561 8789 6595 8823
rect 6653 8789 6687 8823
rect 7113 8789 7147 8823
rect 8769 8789 8803 8823
rect 10425 8789 10459 8823
rect 13461 8789 13495 8823
rect 13645 8789 13679 8823
rect 15485 8789 15519 8823
rect 18429 8789 18463 8823
rect 2927 8585 2961 8619
rect 4445 8585 4479 8619
rect 5917 8585 5951 8619
rect 7481 8585 7515 8619
rect 7941 8585 7975 8619
rect 11345 8585 11379 8619
rect 12725 8585 12759 8619
rect 14381 8585 14415 8619
rect 16037 8585 16071 8619
rect 17969 8585 18003 8619
rect 18429 8585 18463 8619
rect 6377 8517 6411 8551
rect 1961 8449 1995 8483
rect 3341 8449 3375 8483
rect 4077 8449 4111 8483
rect 5089 8449 5123 8483
rect 5181 8449 5215 8483
rect 7113 8449 7147 8483
rect 9617 8449 9651 8483
rect 9873 8449 9907 8483
rect 9965 8449 9999 8483
rect 10232 8449 10266 8483
rect 11897 8449 11931 8483
rect 13838 8449 13872 8483
rect 14105 8449 14139 8483
rect 14197 8449 14231 8483
rect 14565 8449 14599 8483
rect 14832 8449 14866 8483
rect 16497 8449 16531 8483
rect 17049 8449 17083 8483
rect 17509 8449 17543 8483
rect 18153 8449 18187 8483
rect 18245 8449 18279 8483
rect 2237 8381 2271 8415
rect 3157 8381 3191 8415
rect 3801 8381 3835 8415
rect 3985 8381 4019 8415
rect 5365 8381 5399 8415
rect 6929 8381 6963 8415
rect 7021 8381 7055 8415
rect 8033 8381 8067 8415
rect 8125 8381 8159 8415
rect 11989 8381 12023 8415
rect 12081 8381 12115 8415
rect 12541 8381 12575 8415
rect 17233 8381 17267 8415
rect 17417 8381 17451 8415
rect 4721 8313 4755 8347
rect 6101 8313 6135 8347
rect 7573 8313 7607 8347
rect 8493 8313 8527 8347
rect 11529 8313 11563 8347
rect 15945 8313 15979 8347
rect 16313 8313 16347 8347
rect 16865 8313 16899 8347
rect 3433 8245 3467 8279
rect 4537 8245 4571 8279
rect 5549 8245 5583 8279
rect 5733 8245 5767 8279
rect 17877 8245 17911 8279
rect 3433 8041 3467 8075
rect 8953 8041 8987 8075
rect 10517 8041 10551 8075
rect 11713 8041 11747 8075
rect 12541 8041 12575 8075
rect 18429 8041 18463 8075
rect 3065 7973 3099 8007
rect 7113 7973 7147 8007
rect 15025 7973 15059 8007
rect 1961 7905 1995 7939
rect 2237 7905 2271 7939
rect 2513 7905 2547 7939
rect 4353 7905 4387 7939
rect 5181 7905 5215 7939
rect 5273 7905 5307 7939
rect 5733 7905 5767 7939
rect 6561 7905 6595 7939
rect 7849 7905 7883 7939
rect 8217 7905 8251 7939
rect 11345 7905 11379 7939
rect 12173 7905 12207 7939
rect 12357 7905 12391 7939
rect 13185 7905 13219 7939
rect 14289 7905 14323 7939
rect 16405 7905 16439 7939
rect 16681 7905 16715 7939
rect 17785 7905 17819 7939
rect 17877 7905 17911 7939
rect 2697 7837 2731 7871
rect 3617 7837 3651 7871
rect 6653 7837 6687 7871
rect 10333 7837 10367 7871
rect 12909 7837 12943 7871
rect 13737 7837 13771 7871
rect 14381 7837 14415 7871
rect 18245 7837 18279 7871
rect 3157 7769 3191 7803
rect 4261 7769 4295 7803
rect 6745 7769 6779 7803
rect 8401 7769 8435 7803
rect 10066 7769 10100 7803
rect 10609 7769 10643 7803
rect 13001 7769 13035 7803
rect 14473 7769 14507 7803
rect 16138 7769 16172 7803
rect 2605 7701 2639 7735
rect 3801 7701 3835 7735
rect 4169 7701 4203 7735
rect 4721 7701 4755 7735
rect 5089 7701 5123 7735
rect 5825 7701 5859 7735
rect 5917 7701 5951 7735
rect 6285 7701 6319 7735
rect 7205 7701 7239 7735
rect 7573 7701 7607 7735
rect 7665 7701 7699 7735
rect 8309 7701 8343 7735
rect 8769 7701 8803 7735
rect 10793 7701 10827 7735
rect 11161 7701 11195 7735
rect 11253 7701 11287 7735
rect 12081 7701 12115 7735
rect 13369 7701 13403 7735
rect 13921 7701 13955 7735
rect 14841 7701 14875 7735
rect 16773 7701 16807 7735
rect 16865 7701 16899 7735
rect 17233 7701 17267 7735
rect 17325 7701 17359 7735
rect 17693 7701 17727 7735
rect 1409 7497 1443 7531
rect 2329 7497 2363 7531
rect 2789 7497 2823 7531
rect 3433 7497 3467 7531
rect 4905 7497 4939 7531
rect 4997 7497 5031 7531
rect 5365 7497 5399 7531
rect 6193 7497 6227 7531
rect 7757 7497 7791 7531
rect 8125 7497 8159 7531
rect 8953 7497 8987 7531
rect 9781 7497 9815 7531
rect 10149 7497 10183 7531
rect 10977 7497 11011 7531
rect 11345 7497 11379 7531
rect 11897 7497 11931 7531
rect 13093 7497 13127 7531
rect 13461 7497 13495 7531
rect 13921 7497 13955 7531
rect 14749 7497 14783 7531
rect 16037 7497 16071 7531
rect 16405 7497 16439 7531
rect 16681 7497 16715 7531
rect 17141 7497 17175 7531
rect 17969 7497 18003 7531
rect 18337 7497 18371 7531
rect 7389 7429 7423 7463
rect 9321 7429 9355 7463
rect 12357 7429 12391 7463
rect 13001 7429 13035 7463
rect 1961 7361 1995 7395
rect 2881 7361 2915 7395
rect 3249 7361 3283 7395
rect 3709 7361 3743 7395
rect 4169 7361 4203 7395
rect 5825 7361 5859 7395
rect 8493 7361 8527 7395
rect 8585 7361 8619 7395
rect 14013 7361 14047 7395
rect 15577 7361 15611 7395
rect 16221 7361 16255 7395
rect 17049 7361 17083 7395
rect 17877 7361 17911 7395
rect 18521 7361 18555 7395
rect 1685 7293 1719 7327
rect 1869 7293 1903 7327
rect 2973 7293 3007 7327
rect 3893 7293 3927 7327
rect 4077 7293 4111 7327
rect 4813 7293 4847 7327
rect 5641 7293 5675 7327
rect 5733 7293 5767 7327
rect 6653 7293 6687 7327
rect 6929 7293 6963 7327
rect 7113 7293 7147 7327
rect 7297 7293 7331 7327
rect 8033 7293 8067 7327
rect 8769 7293 8803 7327
rect 9413 7293 9447 7327
rect 9597 7293 9631 7327
rect 10241 7293 10275 7327
rect 10333 7293 10367 7327
rect 10701 7293 10735 7327
rect 10885 7293 10919 7327
rect 11989 7293 12023 7327
rect 12081 7293 12115 7327
rect 12909 7293 12943 7327
rect 14105 7293 14139 7327
rect 14841 7293 14875 7327
rect 15025 7293 15059 7327
rect 15669 7293 15703 7327
rect 15761 7293 15795 7327
rect 17325 7293 17359 7327
rect 18153 7293 18187 7327
rect 3525 7225 3559 7259
rect 4537 7225 4571 7259
rect 17509 7225 17543 7259
rect 2421 7157 2455 7191
rect 11529 7157 11563 7191
rect 13553 7157 13587 7191
rect 14381 7157 14415 7191
rect 15209 7157 15243 7191
rect 2789 6953 2823 6987
rect 3617 6953 3651 6987
rect 4905 6953 4939 6987
rect 5733 6953 5767 6987
rect 6929 6953 6963 6987
rect 7941 6953 7975 6987
rect 9505 6953 9539 6987
rect 11437 6953 11471 6987
rect 16681 6953 16715 6987
rect 17509 6953 17543 6987
rect 2237 6817 2271 6851
rect 3065 6817 3099 6851
rect 4721 6817 4755 6851
rect 5549 6817 5583 6851
rect 6377 6817 6411 6851
rect 7757 6817 7791 6851
rect 8585 6817 8619 6851
rect 9965 6817 9999 6851
rect 10149 6817 10183 6851
rect 10885 6817 10919 6851
rect 11897 6817 11931 6851
rect 11989 6817 12023 6851
rect 12817 6817 12851 6851
rect 13645 6817 13679 6851
rect 14381 6817 14415 6851
rect 15117 6817 15151 6851
rect 16313 6817 16347 6851
rect 16497 6817 16531 6851
rect 17233 6817 17267 6851
rect 17969 6817 18003 6851
rect 18153 6817 18187 6851
rect 1685 6749 1719 6783
rect 1961 6749 1995 6783
rect 2421 6749 2455 6783
rect 3985 6749 4019 6783
rect 4445 6749 4479 6783
rect 4537 6749 4571 6783
rect 6745 6749 6779 6783
rect 7481 6749 7515 6783
rect 8309 6749 8343 6783
rect 8401 6749 8435 6783
rect 9321 6749 9355 6783
rect 9873 6749 9907 6783
rect 11161 6749 11195 6783
rect 13461 6749 13495 6783
rect 14473 6749 14507 6783
rect 16221 6749 16255 6783
rect 18521 6749 18555 6783
rect 3249 6681 3283 6715
rect 5365 6681 5399 6715
rect 10793 6681 10827 6715
rect 12633 6681 12667 6715
rect 12725 6681 12759 6715
rect 14565 6681 14599 6715
rect 15301 6681 15335 6715
rect 17049 6681 17083 6715
rect 1501 6613 1535 6647
rect 1777 6613 1811 6647
rect 2329 6613 2363 6647
rect 3157 6613 3191 6647
rect 3801 6613 3835 6647
rect 4077 6613 4111 6647
rect 5273 6613 5307 6647
rect 6101 6613 6135 6647
rect 6193 6613 6227 6647
rect 6561 6613 6595 6647
rect 7113 6613 7147 6647
rect 7573 6613 7607 6647
rect 8953 6613 8987 6647
rect 10333 6613 10367 6647
rect 10701 6613 10735 6647
rect 11345 6613 11379 6647
rect 11805 6613 11839 6647
rect 12265 6613 12299 6647
rect 13093 6613 13127 6647
rect 13553 6613 13587 6647
rect 14933 6613 14967 6647
rect 15393 6613 15427 6647
rect 15761 6613 15795 6647
rect 15853 6613 15887 6647
rect 17141 6613 17175 6647
rect 17877 6613 17911 6647
rect 18337 6613 18371 6647
rect 2237 6409 2271 6443
rect 2421 6409 2455 6443
rect 3249 6409 3283 6443
rect 3801 6409 3835 6443
rect 4169 6409 4203 6443
rect 4261 6409 4295 6443
rect 4629 6409 4663 6443
rect 5089 6409 5123 6443
rect 5825 6409 5859 6443
rect 6193 6409 6227 6443
rect 6837 6409 6871 6443
rect 8033 6409 8067 6443
rect 9229 6409 9263 6443
rect 9597 6409 9631 6443
rect 9689 6409 9723 6443
rect 10471 6409 10505 6443
rect 13553 6409 13587 6443
rect 14013 6409 14047 6443
rect 14473 6409 14507 6443
rect 15209 6409 15243 6443
rect 16037 6409 16071 6443
rect 17417 6409 17451 6443
rect 1777 6341 1811 6375
rect 3341 6341 3375 6375
rect 4997 6341 5031 6375
rect 7205 6341 7239 6375
rect 7297 6341 7331 6375
rect 17049 6341 17083 6375
rect 18337 6341 18371 6375
rect 1869 6273 1903 6307
rect 2605 6273 2639 6307
rect 2697 6273 2731 6307
rect 8861 6273 8895 6307
rect 10241 6273 10275 6307
rect 11345 6273 11379 6307
rect 11897 6273 11931 6307
rect 12633 6273 12667 6307
rect 12725 6273 12759 6307
rect 14381 6273 14415 6307
rect 15301 6273 15335 6307
rect 17877 6273 17911 6307
rect 1685 6205 1719 6239
rect 3157 6205 3191 6239
rect 4353 6205 4387 6239
rect 5181 6205 5215 6239
rect 5549 6205 5583 6239
rect 5733 6205 5767 6239
rect 6745 6205 6779 6239
rect 7389 6205 7423 6239
rect 7849 6205 7883 6239
rect 7941 6205 7975 6239
rect 8585 6205 8619 6239
rect 8769 6205 8803 6239
rect 9505 6205 9539 6239
rect 11989 6205 12023 6239
rect 12081 6205 12115 6239
rect 12541 6205 12575 6239
rect 13277 6205 13311 6239
rect 13461 6205 13495 6239
rect 14657 6205 14691 6239
rect 15485 6205 15519 6239
rect 16129 6205 16163 6239
rect 16221 6205 16255 6239
rect 16865 6205 16899 6239
rect 16957 6205 16991 6239
rect 17969 6205 18003 6239
rect 18061 6205 18095 6239
rect 6561 6137 6595 6171
rect 10057 6137 10091 6171
rect 14841 6137 14875 6171
rect 2881 6069 2915 6103
rect 3709 6069 3743 6103
rect 8401 6069 8435 6103
rect 11161 6069 11195 6103
rect 11529 6069 11563 6103
rect 13093 6069 13127 6103
rect 13921 6069 13955 6103
rect 15669 6069 15703 6103
rect 17509 6069 17543 6103
rect 1593 5865 1627 5899
rect 3985 5865 4019 5899
rect 5641 5865 5675 5899
rect 6469 5865 6503 5899
rect 6745 5865 6779 5899
rect 12633 5865 12667 5899
rect 13645 5865 13679 5899
rect 13737 5865 13771 5899
rect 15761 5865 15795 5899
rect 18337 5865 18371 5899
rect 4077 5797 4111 5831
rect 7941 5797 7975 5831
rect 15853 5797 15887 5831
rect 17509 5797 17543 5831
rect 1501 5729 1535 5763
rect 2237 5729 2271 5763
rect 2881 5729 2915 5763
rect 3065 5729 3099 5763
rect 5089 5729 5123 5763
rect 5917 5729 5951 5763
rect 7205 5729 7239 5763
rect 8677 5729 8711 5763
rect 9229 5729 9263 5763
rect 9965 5729 9999 5763
rect 10241 5729 10275 5763
rect 12449 5729 12483 5763
rect 13093 5729 13127 5763
rect 13185 5729 13219 5763
rect 14381 5729 14415 5763
rect 15209 5729 15243 5763
rect 15301 5729 15335 5763
rect 16497 5729 16531 5763
rect 17325 5729 17359 5763
rect 18061 5729 18095 5763
rect 3249 5661 3283 5695
rect 3617 5661 3651 5695
rect 3801 5661 3835 5695
rect 4269 5661 4303 5695
rect 4537 5661 4571 5695
rect 4813 5661 4847 5695
rect 6561 5661 6595 5695
rect 7297 5661 7331 5695
rect 7389 5661 7423 5695
rect 8493 5661 8527 5695
rect 8953 5661 8987 5695
rect 9505 5661 9539 5695
rect 10885 5661 10919 5695
rect 11161 5661 11195 5695
rect 12265 5661 12299 5695
rect 13461 5661 13495 5695
rect 13921 5661 13955 5695
rect 14105 5661 14139 5695
rect 16221 5661 16255 5695
rect 18521 5661 18555 5695
rect 1961 5593 1995 5627
rect 2789 5593 2823 5627
rect 6837 5593 6871 5627
rect 8401 5593 8435 5627
rect 13001 5593 13035 5627
rect 15393 5593 15427 5627
rect 17141 5593 17175 5627
rect 17969 5593 18003 5627
rect 2053 5525 2087 5559
rect 2421 5525 2455 5559
rect 3433 5525 3467 5559
rect 4353 5525 4387 5559
rect 5181 5525 5215 5559
rect 5273 5525 5307 5559
rect 6009 5525 6043 5559
rect 6101 5525 6135 5559
rect 7757 5525 7791 5559
rect 8033 5525 8067 5559
rect 9413 5525 9447 5559
rect 9873 5525 9907 5559
rect 11805 5525 11839 5559
rect 12173 5525 12207 5559
rect 16313 5525 16347 5559
rect 16681 5525 16715 5559
rect 17049 5525 17083 5559
rect 17877 5525 17911 5559
rect 1501 5321 1535 5355
rect 1869 5321 1903 5355
rect 2329 5321 2363 5355
rect 2789 5321 2823 5355
rect 3065 5321 3099 5355
rect 3985 5321 4019 5355
rect 4445 5321 4479 5355
rect 4813 5321 4847 5355
rect 5457 5321 5491 5355
rect 5917 5321 5951 5355
rect 6561 5321 6595 5355
rect 7389 5321 7423 5355
rect 7849 5321 7883 5355
rect 8309 5321 8343 5355
rect 8769 5321 8803 5355
rect 10057 5321 10091 5355
rect 10793 5321 10827 5355
rect 10885 5321 10919 5355
rect 11529 5321 11563 5355
rect 12633 5321 12667 5355
rect 13185 5321 13219 5355
rect 13553 5321 13587 5355
rect 13645 5321 13679 5355
rect 15853 5321 15887 5355
rect 16313 5321 16347 5355
rect 18061 5321 18095 5355
rect 2237 5253 2271 5287
rect 4905 5253 4939 5287
rect 6745 5253 6779 5287
rect 8217 5253 8251 5287
rect 9965 5253 9999 5287
rect 11897 5253 11931 5287
rect 14381 5253 14415 5287
rect 15761 5253 15795 5287
rect 18521 5253 18555 5287
rect 1685 5185 1719 5219
rect 2973 5185 3007 5219
rect 3249 5185 3283 5219
rect 3525 5185 3559 5219
rect 4169 5185 4203 5219
rect 5825 5185 5859 5219
rect 6377 5185 6411 5219
rect 9137 5185 9171 5219
rect 12725 5185 12759 5219
rect 15025 5185 15059 5219
rect 15117 5185 15151 5219
rect 16681 5185 16715 5219
rect 17969 5185 18003 5219
rect 2513 5117 2547 5151
rect 5365 5117 5399 5151
rect 6009 5117 6043 5151
rect 7113 5117 7147 5151
rect 7297 5117 7331 5151
rect 8401 5117 8435 5151
rect 9229 5117 9263 5151
rect 9413 5117 9447 5151
rect 10149 5117 10183 5151
rect 10701 5117 10735 5151
rect 11989 5117 12023 5151
rect 12173 5117 12207 5151
rect 12449 5117 12483 5151
rect 13737 5117 13771 5151
rect 14473 5117 14507 5151
rect 14565 5117 14599 5151
rect 15669 5117 15703 5151
rect 16957 5117 16991 5151
rect 18153 5117 18187 5151
rect 3341 5049 3375 5083
rect 3617 5049 3651 5083
rect 5181 5049 5215 5083
rect 14841 5049 14875 5083
rect 3801 4981 3835 5015
rect 4353 4981 4387 5015
rect 6837 4981 6871 5015
rect 7757 4981 7791 5015
rect 9597 4981 9631 5015
rect 11253 4981 11287 5015
rect 13093 4981 13127 5015
rect 14013 4981 14047 5015
rect 15301 4981 15335 5015
rect 16221 4981 16255 5015
rect 17601 4981 17635 5015
rect 1501 4777 1535 4811
rect 1869 4777 1903 4811
rect 2237 4777 2271 4811
rect 4169 4777 4203 4811
rect 4353 4777 4387 4811
rect 4537 4777 4571 4811
rect 4813 4777 4847 4811
rect 5641 4777 5675 4811
rect 9873 4777 9907 4811
rect 11805 4777 11839 4811
rect 17693 4777 17727 4811
rect 18061 4777 18095 4811
rect 18429 4777 18463 4811
rect 3985 4709 4019 4743
rect 6469 4709 6503 4743
rect 11713 4709 11747 4743
rect 16589 4709 16623 4743
rect 6101 4641 6135 4675
rect 6193 4641 6227 4675
rect 7297 4641 7331 4675
rect 8033 4641 8067 4675
rect 9597 4641 9631 4675
rect 10517 4641 10551 4675
rect 10793 4641 10827 4675
rect 10977 4641 11011 4675
rect 12817 4641 12851 4675
rect 13461 4641 13495 4675
rect 13645 4641 13679 4675
rect 14657 4641 14691 4675
rect 15025 4641 15059 4675
rect 15209 4641 15243 4675
rect 16313 4641 16347 4675
rect 17233 4641 17267 4675
rect 1685 4573 1719 4607
rect 2053 4573 2087 4607
rect 2421 4573 2455 4607
rect 2789 4573 2823 4607
rect 3065 4573 3099 4607
rect 3341 4573 3375 4607
rect 3617 4573 3651 4607
rect 3801 4573 3835 4607
rect 4997 4573 5031 4607
rect 6009 4573 6043 4607
rect 9413 4573 9447 4607
rect 9505 4573 9539 4607
rect 10333 4573 10367 4607
rect 11069 4573 11103 4607
rect 11989 4573 12023 4607
rect 12541 4573 12575 4607
rect 14473 4573 14507 4607
rect 16129 4573 16163 4607
rect 16957 4573 16991 4607
rect 17509 4573 17543 4607
rect 17877 4573 17911 4607
rect 18245 4573 18279 4607
rect 7849 4505 7883 4539
rect 8309 4505 8343 4539
rect 13369 4505 13403 4539
rect 14565 4505 14599 4539
rect 16221 4505 16255 4539
rect 2605 4437 2639 4471
rect 2881 4437 2915 4471
rect 3157 4437 3191 4471
rect 3433 4437 3467 4471
rect 5181 4437 5215 4471
rect 6653 4437 6687 4471
rect 7021 4437 7055 4471
rect 7113 4437 7147 4471
rect 7481 4437 7515 4471
rect 7941 4437 7975 4471
rect 8585 4437 8619 4471
rect 9045 4437 9079 4471
rect 10241 4437 10275 4471
rect 11437 4437 11471 4471
rect 12173 4437 12207 4471
rect 12633 4437 12667 4471
rect 13001 4437 13035 4471
rect 13829 4437 13863 4471
rect 14105 4437 14139 4471
rect 15301 4437 15335 4471
rect 15669 4437 15703 4471
rect 15761 4437 15795 4471
rect 17049 4437 17083 4471
rect 1501 4233 1535 4267
rect 1869 4233 1903 4267
rect 3709 4233 3743 4267
rect 3893 4233 3927 4267
rect 6377 4233 6411 4267
rect 6561 4233 6595 4267
rect 7021 4233 7055 4267
rect 7389 4233 7423 4267
rect 7481 4233 7515 4267
rect 8769 4233 8803 4267
rect 9321 4233 9355 4267
rect 9413 4233 9447 4267
rect 10793 4233 10827 4267
rect 13277 4233 13311 4267
rect 13737 4233 13771 4267
rect 14105 4233 14139 4267
rect 15117 4233 15151 4267
rect 15577 4233 15611 4267
rect 15945 4233 15979 4267
rect 17693 4233 17727 4267
rect 6929 4165 6963 4199
rect 7849 4165 7883 4199
rect 10425 4165 10459 4199
rect 15209 4165 15243 4199
rect 1685 4097 1719 4131
rect 2053 4097 2087 4131
rect 2421 4097 2455 4131
rect 2697 4097 2731 4131
rect 2973 4097 3007 4131
rect 3249 4097 3283 4131
rect 3433 4097 3467 4131
rect 3617 4097 3651 4131
rect 4169 4097 4203 4131
rect 4353 4097 4387 4131
rect 10609 4097 10643 4131
rect 11529 4097 11563 4131
rect 12265 4097 12299 4131
rect 12909 4097 12943 4131
rect 14197 4097 14231 4131
rect 14473 4097 14507 4131
rect 16037 4097 16071 4131
rect 16773 4097 16807 4131
rect 17141 4097 17175 4131
rect 17509 4097 17543 4131
rect 17877 4097 17911 4131
rect 18245 4097 18279 4131
rect 7665 4029 7699 4063
rect 8401 4029 8435 4063
rect 9505 4029 9539 4063
rect 11989 4029 12023 4063
rect 12633 4029 12667 4063
rect 12817 4029 12851 4063
rect 13553 4029 13587 4063
rect 13645 4029 13679 4063
rect 15301 4029 15335 4063
rect 16129 4029 16163 4063
rect 2513 3961 2547 3995
rect 4537 3961 4571 3995
rect 8953 3961 8987 3995
rect 12173 3961 12207 3995
rect 14657 3961 14691 3995
rect 16957 3961 16991 3995
rect 17325 3961 17359 3995
rect 18061 3961 18095 3995
rect 18429 3961 18463 3995
rect 2237 3893 2271 3927
rect 2789 3893 2823 3927
rect 3065 3893 3099 3927
rect 8125 3893 8159 3927
rect 10333 3893 10367 3927
rect 11713 3893 11747 3927
rect 12449 3893 12483 3927
rect 14381 3893 14415 3927
rect 14749 3893 14783 3927
rect 16405 3893 16439 3927
rect 1501 3689 1535 3723
rect 2145 3689 2179 3723
rect 2697 3689 2731 3723
rect 3249 3689 3283 3723
rect 3525 3689 3559 3723
rect 4169 3689 4203 3723
rect 10793 3689 10827 3723
rect 12541 3689 12575 3723
rect 15485 3689 15519 3723
rect 16497 3689 16531 3723
rect 17693 3689 17727 3723
rect 18061 3689 18095 3723
rect 18429 3689 18463 3723
rect 6837 3621 6871 3655
rect 12725 3621 12759 3655
rect 13553 3621 13587 3655
rect 13737 3621 13771 3655
rect 13921 3621 13955 3655
rect 14197 3621 14231 3655
rect 14657 3621 14691 3655
rect 15761 3621 15795 3655
rect 17325 3621 17359 3655
rect 13001 3553 13035 3587
rect 1685 3485 1719 3519
rect 1777 3485 1811 3519
rect 2329 3485 2363 3519
rect 2605 3485 2639 3519
rect 2881 3485 2915 3519
rect 3157 3501 3191 3535
rect 3985 3485 4019 3519
rect 4353 3485 4387 3519
rect 6653 3485 6687 3519
rect 7573 3485 7607 3519
rect 7849 3485 7883 3519
rect 10977 3485 11011 3519
rect 14749 3485 14783 3519
rect 15025 3485 15059 3519
rect 15301 3485 15335 3519
rect 15577 3485 15611 3519
rect 16221 3485 16255 3519
rect 16681 3485 16715 3519
rect 16773 3485 16807 3519
rect 17141 3485 17175 3519
rect 17509 3485 17543 3519
rect 17877 3485 17911 3519
rect 18245 3485 18279 3519
rect 12909 3417 12943 3451
rect 14473 3417 14507 3451
rect 1961 3349 1995 3383
rect 2421 3349 2455 3383
rect 2973 3349 3007 3383
rect 3801 3349 3835 3383
rect 7757 3349 7791 3383
rect 8033 3349 8067 3383
rect 11161 3349 11195 3383
rect 13369 3349 13403 3383
rect 14933 3349 14967 3383
rect 15209 3349 15243 3383
rect 16129 3349 16163 3383
rect 16405 3349 16439 3383
rect 16957 3349 16991 3383
rect 1501 3145 1535 3179
rect 3893 3145 3927 3179
rect 12541 3145 12575 3179
rect 12909 3145 12943 3179
rect 13185 3145 13219 3179
rect 16221 3145 16255 3179
rect 16497 3145 16531 3179
rect 17049 3145 17083 3179
rect 18061 3145 18095 3179
rect 18429 3145 18463 3179
rect 12725 3077 12759 3111
rect 1685 3009 1719 3043
rect 2053 3009 2087 3043
rect 2421 3009 2455 3043
rect 2789 3009 2823 3043
rect 3065 3009 3099 3043
rect 3341 3009 3375 3043
rect 5549 3009 5583 3043
rect 7021 3009 7055 3043
rect 7481 3009 7515 3043
rect 11345 3009 11379 3043
rect 11713 3009 11747 3043
rect 11805 3009 11839 3043
rect 13553 3009 13587 3043
rect 13829 3009 13863 3043
rect 14013 3009 14047 3043
rect 14105 3009 14139 3043
rect 14473 3009 14507 3043
rect 15025 3009 15059 3043
rect 15209 3009 15243 3043
rect 15485 3009 15519 3043
rect 15761 3009 15795 3043
rect 16037 3009 16071 3043
rect 16313 3009 16347 3043
rect 16865 3009 16899 3043
rect 17141 3009 17175 3043
rect 17509 3009 17543 3043
rect 17877 3009 17911 3043
rect 18245 3009 18279 3043
rect 3617 2941 3651 2975
rect 1869 2873 1903 2907
rect 2881 2873 2915 2907
rect 7297 2873 7331 2907
rect 13093 2873 13127 2907
rect 13461 2873 13495 2907
rect 14657 2873 14691 2907
rect 15393 2873 15427 2907
rect 15945 2873 15979 2907
rect 16681 2873 16715 2907
rect 2237 2805 2271 2839
rect 2605 2805 2639 2839
rect 3157 2805 3191 2839
rect 3525 2805 3559 2839
rect 5365 2805 5399 2839
rect 7205 2805 7239 2839
rect 11161 2805 11195 2839
rect 11529 2805 11563 2839
rect 11989 2805 12023 2839
rect 14289 2805 14323 2839
rect 14841 2805 14875 2839
rect 15669 2805 15703 2839
rect 17325 2805 17359 2839
rect 17693 2805 17727 2839
rect 1501 2601 1535 2635
rect 15025 2601 15059 2635
rect 15301 2601 15335 2635
rect 18429 2601 18463 2635
rect 14197 2533 14231 2567
rect 15945 2533 15979 2567
rect 16497 2533 16531 2567
rect 1685 2397 1719 2431
rect 2053 2397 2087 2431
rect 2421 2397 2455 2431
rect 2789 2397 2823 2431
rect 3249 2397 3283 2431
rect 3341 2397 3375 2431
rect 3801 2397 3835 2431
rect 4905 2397 4939 2431
rect 5457 2397 5491 2431
rect 6653 2397 6687 2431
rect 7389 2397 7423 2431
rect 7941 2397 7975 2431
rect 8953 2397 8987 2431
rect 9597 2397 9631 2431
rect 10701 2397 10735 2431
rect 11529 2397 11563 2431
rect 12081 2397 12115 2431
rect 12909 2397 12943 2431
rect 13369 2397 13403 2431
rect 13737 2397 13771 2431
rect 14381 2397 14415 2431
rect 14841 2397 14875 2431
rect 15393 2397 15427 2431
rect 15761 2397 15795 2431
rect 16221 2397 16255 2431
rect 16313 2397 16347 2431
rect 16773 2397 16807 2431
rect 17049 2397 17083 2431
rect 17509 2397 17543 2431
rect 17877 2397 17911 2431
rect 18245 2397 18279 2431
rect 4169 2329 4203 2363
rect 12633 2329 12667 2363
rect 1869 2261 1903 2295
rect 2237 2261 2271 2295
rect 2605 2261 2639 2295
rect 3065 2261 3099 2295
rect 3525 2261 3559 2295
rect 3985 2261 4019 2295
rect 4721 2261 4755 2295
rect 5641 2261 5675 2295
rect 6469 2261 6503 2295
rect 7205 2261 7239 2295
rect 8125 2261 8159 2295
rect 9137 2261 9171 2295
rect 9781 2261 9815 2295
rect 10517 2261 10551 2295
rect 11713 2261 11747 2295
rect 12265 2261 12299 2295
rect 12725 2261 12759 2295
rect 13093 2261 13127 2295
rect 13553 2261 13587 2295
rect 13921 2261 13955 2295
rect 14657 2261 14691 2295
rect 15577 2261 15611 2295
rect 16037 2261 16071 2295
rect 16957 2261 16991 2295
rect 17233 2261 17267 2295
rect 17693 2261 17727 2295
rect 18061 2261 18095 2295
<< metal1 >>
rect 2130 15172 2136 15224
rect 2188 15212 2194 15224
rect 4522 15212 4528 15224
rect 2188 15184 4528 15212
rect 2188 15172 2194 15184
rect 4522 15172 4528 15184
rect 4580 15172 4586 15224
rect 11790 14900 11796 14952
rect 11848 14940 11854 14952
rect 18322 14940 18328 14952
rect 11848 14912 18328 14940
rect 11848 14900 11854 14912
rect 18322 14900 18328 14912
rect 18380 14900 18386 14952
rect 6270 14832 6276 14884
rect 6328 14872 6334 14884
rect 11514 14872 11520 14884
rect 6328 14844 11520 14872
rect 6328 14832 6334 14844
rect 11514 14832 11520 14844
rect 11572 14872 11578 14884
rect 12618 14872 12624 14884
rect 11572 14844 12624 14872
rect 11572 14832 11578 14844
rect 12618 14832 12624 14844
rect 12676 14832 12682 14884
rect 1854 14764 1860 14816
rect 1912 14804 1918 14816
rect 5810 14804 5816 14816
rect 1912 14776 5816 14804
rect 1912 14764 1918 14776
rect 5810 14764 5816 14776
rect 5868 14764 5874 14816
rect 8570 14764 8576 14816
rect 8628 14804 8634 14816
rect 13262 14804 13268 14816
rect 8628 14776 13268 14804
rect 8628 14764 8634 14776
rect 13262 14764 13268 14776
rect 13320 14764 13326 14816
rect 1104 14714 18860 14736
rect 1104 14662 3174 14714
rect 3226 14662 3238 14714
rect 3290 14662 3302 14714
rect 3354 14662 3366 14714
rect 3418 14662 3430 14714
rect 3482 14662 7622 14714
rect 7674 14662 7686 14714
rect 7738 14662 7750 14714
rect 7802 14662 7814 14714
rect 7866 14662 7878 14714
rect 7930 14662 12070 14714
rect 12122 14662 12134 14714
rect 12186 14662 12198 14714
rect 12250 14662 12262 14714
rect 12314 14662 12326 14714
rect 12378 14662 16518 14714
rect 16570 14662 16582 14714
rect 16634 14662 16646 14714
rect 16698 14662 16710 14714
rect 16762 14662 16774 14714
rect 16826 14662 18860 14714
rect 1104 14640 18860 14662
rect 2038 14560 2044 14612
rect 2096 14600 2102 14612
rect 4985 14603 5043 14609
rect 4985 14600 4997 14603
rect 2096 14572 4997 14600
rect 2096 14560 2102 14572
rect 4985 14569 4997 14572
rect 5031 14569 5043 14603
rect 4985 14563 5043 14569
rect 2240 14504 2774 14532
rect 2240 14476 2268 14504
rect 2222 14464 2228 14476
rect 2135 14436 2228 14464
rect 2222 14424 2228 14436
rect 2280 14424 2286 14476
rect 1946 14396 1952 14408
rect 1907 14368 1952 14396
rect 1946 14356 1952 14368
rect 2004 14356 2010 14408
rect 2746 14328 2774 14504
rect 3050 14492 3056 14544
rect 3108 14532 3114 14544
rect 4798 14532 4804 14544
rect 3108 14504 4804 14532
rect 3108 14492 3114 14504
rect 3160 14473 3188 14504
rect 4798 14492 4804 14504
rect 4856 14492 4862 14544
rect 5000 14532 5028 14563
rect 5994 14560 6000 14612
rect 6052 14600 6058 14612
rect 6457 14603 6515 14609
rect 6457 14600 6469 14603
rect 6052 14572 6469 14600
rect 6052 14560 6058 14572
rect 6457 14569 6469 14572
rect 6503 14569 6515 14603
rect 6457 14563 6515 14569
rect 9950 14560 9956 14612
rect 10008 14600 10014 14612
rect 10597 14603 10655 14609
rect 10597 14600 10609 14603
rect 10008 14572 10609 14600
rect 10008 14560 10014 14572
rect 10597 14569 10609 14572
rect 10643 14569 10655 14603
rect 15930 14600 15936 14612
rect 10597 14563 10655 14569
rect 11532 14572 15936 14600
rect 5000 14504 5304 14532
rect 3145 14467 3203 14473
rect 3145 14433 3157 14467
rect 3191 14433 3203 14467
rect 3145 14427 3203 14433
rect 4062 14424 4068 14476
rect 4120 14464 4126 14476
rect 4617 14467 4675 14473
rect 4617 14464 4629 14467
rect 4120 14436 4629 14464
rect 4120 14424 4126 14436
rect 4617 14433 4629 14436
rect 4663 14464 4675 14467
rect 5169 14467 5227 14473
rect 5169 14464 5181 14467
rect 4663 14436 5181 14464
rect 4663 14433 4675 14436
rect 4617 14427 4675 14433
rect 5169 14433 5181 14436
rect 5215 14433 5227 14467
rect 5169 14427 5227 14433
rect 2869 14399 2927 14405
rect 2869 14365 2881 14399
rect 2915 14396 2927 14399
rect 3050 14396 3056 14408
rect 2915 14368 3056 14396
rect 2915 14365 2927 14368
rect 2869 14359 2927 14365
rect 3050 14356 3056 14368
rect 3108 14356 3114 14408
rect 3513 14399 3571 14405
rect 3513 14365 3525 14399
rect 3559 14396 3571 14399
rect 4154 14396 4160 14408
rect 3559 14368 4160 14396
rect 3559 14365 3571 14368
rect 3513 14359 3571 14365
rect 4154 14356 4160 14368
rect 4212 14356 4218 14408
rect 4338 14396 4344 14408
rect 4299 14368 4344 14396
rect 4338 14356 4344 14368
rect 4396 14356 4402 14408
rect 4893 14399 4951 14405
rect 4893 14365 4905 14399
rect 4939 14396 4951 14399
rect 5276 14396 5304 14504
rect 8478 14464 8484 14476
rect 6656 14436 8484 14464
rect 6656 14405 6684 14436
rect 8478 14424 8484 14436
rect 8536 14424 8542 14476
rect 8754 14464 8760 14476
rect 8715 14436 8760 14464
rect 8754 14424 8760 14436
rect 8812 14424 8818 14476
rect 10321 14467 10379 14473
rect 10321 14433 10333 14467
rect 10367 14464 10379 14467
rect 11330 14464 11336 14476
rect 10367 14436 11336 14464
rect 10367 14433 10379 14436
rect 10321 14427 10379 14433
rect 11330 14424 11336 14436
rect 11388 14424 11394 14476
rect 4939 14368 5304 14396
rect 6641 14399 6699 14405
rect 4939 14365 4951 14368
rect 4893 14359 4951 14365
rect 6641 14365 6653 14399
rect 6687 14365 6699 14399
rect 6641 14359 6699 14365
rect 10065 14399 10123 14405
rect 10065 14365 10077 14399
rect 10111 14396 10123 14399
rect 10226 14396 10232 14408
rect 10111 14368 10232 14396
rect 10111 14365 10123 14368
rect 10065 14359 10123 14365
rect 10226 14356 10232 14368
rect 10284 14356 10290 14408
rect 10413 14399 10471 14405
rect 10413 14365 10425 14399
rect 10459 14365 10471 14399
rect 10413 14359 10471 14365
rect 10965 14399 11023 14405
rect 10965 14365 10977 14399
rect 11011 14396 11023 14399
rect 11241 14399 11299 14405
rect 11241 14396 11253 14399
rect 11011 14368 11253 14396
rect 11011 14365 11023 14368
rect 10965 14359 11023 14365
rect 11241 14365 11253 14368
rect 11287 14396 11299 14399
rect 11532 14396 11560 14572
rect 15930 14560 15936 14572
rect 15988 14560 15994 14612
rect 18322 14600 18328 14612
rect 18283 14572 18328 14600
rect 18322 14560 18328 14572
rect 18380 14560 18386 14612
rect 13909 14467 13967 14473
rect 13909 14433 13921 14467
rect 13955 14464 13967 14467
rect 14185 14467 14243 14473
rect 14185 14464 14197 14467
rect 13955 14436 14197 14464
rect 13955 14433 13967 14436
rect 13909 14427 13967 14433
rect 14185 14433 14197 14436
rect 14231 14464 14243 14467
rect 15286 14464 15292 14476
rect 14231 14436 15292 14464
rect 14231 14433 14243 14436
rect 14185 14427 14243 14433
rect 15286 14424 15292 14436
rect 15344 14424 15350 14476
rect 11287 14368 11560 14396
rect 12897 14399 12955 14405
rect 11287 14365 11299 14368
rect 11241 14359 11299 14365
rect 12897 14365 12909 14399
rect 12943 14396 12955 14399
rect 12986 14396 12992 14408
rect 12943 14368 12992 14396
rect 12943 14365 12955 14368
rect 12897 14359 12955 14365
rect 5537 14331 5595 14337
rect 5537 14328 5549 14331
rect 2746 14300 5549 14328
rect 5537 14297 5549 14300
rect 5583 14297 5595 14331
rect 5537 14291 5595 14297
rect 5718 14288 5724 14340
rect 5776 14328 5782 14340
rect 10428 14328 10456 14359
rect 12986 14356 12992 14368
rect 13044 14356 13050 14408
rect 13354 14356 13360 14408
rect 13412 14396 13418 14408
rect 13633 14399 13691 14405
rect 13633 14396 13645 14399
rect 13412 14368 13645 14396
rect 13412 14356 13418 14368
rect 13633 14365 13645 14368
rect 13679 14365 13691 14399
rect 13633 14359 13691 14365
rect 13998 14356 14004 14408
rect 14056 14396 14062 14408
rect 14369 14399 14427 14405
rect 14369 14396 14381 14399
rect 14056 14368 14381 14396
rect 14056 14356 14062 14368
rect 14369 14365 14381 14368
rect 14415 14365 14427 14399
rect 14369 14359 14427 14365
rect 14645 14399 14703 14405
rect 14645 14365 14657 14399
rect 14691 14396 14703 14399
rect 14691 14368 16252 14396
rect 14691 14365 14703 14368
rect 14645 14359 14703 14365
rect 5776 14300 10456 14328
rect 12652 14331 12710 14337
rect 5776 14288 5782 14300
rect 12652 14297 12664 14331
rect 12698 14328 12710 14331
rect 13906 14328 13912 14340
rect 12698 14300 13912 14328
rect 12698 14297 12710 14300
rect 12652 14291 12710 14297
rect 13906 14288 13912 14300
rect 13964 14288 13970 14340
rect 14384 14328 14412 14359
rect 14384 14300 15056 14328
rect 2866 14220 2872 14272
rect 2924 14260 2930 14272
rect 3329 14263 3387 14269
rect 3329 14260 3341 14263
rect 2924 14232 3341 14260
rect 2924 14220 2930 14232
rect 3329 14229 3341 14232
rect 3375 14229 3387 14263
rect 3329 14223 3387 14229
rect 3786 14220 3792 14272
rect 3844 14260 3850 14272
rect 4709 14263 4767 14269
rect 4709 14260 4721 14263
rect 3844 14232 4721 14260
rect 3844 14220 3850 14232
rect 4709 14229 4721 14232
rect 4755 14229 4767 14263
rect 4709 14223 4767 14229
rect 4798 14220 4804 14272
rect 4856 14260 4862 14272
rect 5353 14263 5411 14269
rect 5353 14260 5365 14263
rect 4856 14232 5365 14260
rect 4856 14220 4862 14232
rect 5353 14229 5365 14232
rect 5399 14229 5411 14263
rect 5353 14223 5411 14229
rect 8754 14220 8760 14272
rect 8812 14260 8818 14272
rect 8941 14263 8999 14269
rect 8941 14260 8953 14263
rect 8812 14232 8953 14260
rect 8812 14220 8818 14232
rect 8941 14229 8953 14232
rect 8987 14229 8999 14263
rect 8941 14223 8999 14229
rect 9122 14220 9128 14272
rect 9180 14260 9186 14272
rect 11149 14263 11207 14269
rect 11149 14260 11161 14263
rect 9180 14232 11161 14260
rect 9180 14220 9186 14232
rect 11149 14229 11161 14232
rect 11195 14229 11207 14263
rect 11514 14260 11520 14272
rect 11475 14232 11520 14260
rect 11149 14223 11207 14229
rect 11514 14220 11520 14232
rect 11572 14220 11578 14272
rect 12434 14220 12440 14272
rect 12492 14260 12498 14272
rect 14734 14260 14740 14272
rect 12492 14232 14740 14260
rect 12492 14220 12498 14232
rect 14734 14220 14740 14232
rect 14792 14220 14798 14272
rect 14918 14260 14924 14272
rect 14879 14232 14924 14260
rect 14918 14220 14924 14232
rect 14976 14220 14982 14272
rect 15028 14260 15056 14300
rect 15654 14288 15660 14340
rect 15712 14328 15718 14340
rect 16034 14331 16092 14337
rect 16034 14328 16046 14331
rect 15712 14300 16046 14328
rect 15712 14288 15718 14300
rect 16034 14297 16046 14300
rect 16080 14297 16092 14331
rect 16224 14328 16252 14368
rect 16298 14356 16304 14408
rect 16356 14396 16362 14408
rect 16669 14399 16727 14405
rect 16669 14396 16681 14399
rect 16356 14368 16681 14396
rect 16356 14356 16362 14368
rect 16669 14365 16681 14368
rect 16715 14365 16727 14399
rect 16669 14359 16727 14365
rect 16936 14399 16994 14405
rect 16936 14365 16948 14399
rect 16982 14396 16994 14399
rect 18690 14396 18696 14408
rect 16982 14368 18696 14396
rect 16982 14365 16994 14368
rect 16936 14359 16994 14365
rect 18690 14356 18696 14368
rect 18748 14356 18754 14408
rect 16224 14300 16896 14328
rect 16034 14291 16092 14297
rect 16390 14260 16396 14272
rect 15028 14232 16396 14260
rect 16390 14220 16396 14232
rect 16448 14220 16454 14272
rect 16868 14260 16896 14300
rect 17586 14288 17592 14340
rect 17644 14328 17650 14340
rect 17644 14300 18092 14328
rect 17644 14288 17650 14300
rect 17770 14260 17776 14272
rect 16868 14232 17776 14260
rect 17770 14220 17776 14232
rect 17828 14220 17834 14272
rect 18064 14269 18092 14300
rect 18138 14288 18144 14340
rect 18196 14328 18202 14340
rect 18417 14331 18475 14337
rect 18417 14328 18429 14331
rect 18196 14300 18429 14328
rect 18196 14288 18202 14300
rect 18417 14297 18429 14300
rect 18463 14328 18475 14331
rect 18598 14328 18604 14340
rect 18463 14300 18604 14328
rect 18463 14297 18475 14300
rect 18417 14291 18475 14297
rect 18598 14288 18604 14300
rect 18656 14288 18662 14340
rect 18049 14263 18107 14269
rect 18049 14229 18061 14263
rect 18095 14229 18107 14263
rect 18049 14223 18107 14229
rect 1104 14170 18860 14192
rect 1104 14118 5398 14170
rect 5450 14118 5462 14170
rect 5514 14118 5526 14170
rect 5578 14118 5590 14170
rect 5642 14118 5654 14170
rect 5706 14118 9846 14170
rect 9898 14118 9910 14170
rect 9962 14118 9974 14170
rect 10026 14118 10038 14170
rect 10090 14118 10102 14170
rect 10154 14118 14294 14170
rect 14346 14118 14358 14170
rect 14410 14118 14422 14170
rect 14474 14118 14486 14170
rect 14538 14118 14550 14170
rect 14602 14118 18860 14170
rect 1104 14096 18860 14118
rect 3418 14016 3424 14068
rect 3476 14056 3482 14068
rect 4157 14059 4215 14065
rect 4157 14056 4169 14059
rect 3476 14028 4169 14056
rect 3476 14016 3482 14028
rect 4157 14025 4169 14028
rect 4203 14025 4215 14059
rect 4157 14019 4215 14025
rect 4433 14059 4491 14065
rect 4433 14025 4445 14059
rect 4479 14025 4491 14059
rect 4433 14019 4491 14025
rect 4893 14059 4951 14065
rect 4893 14025 4905 14059
rect 4939 14056 4951 14059
rect 5718 14056 5724 14068
rect 4939 14028 5724 14056
rect 4939 14025 4951 14028
rect 4893 14019 4951 14025
rect 3970 13988 3976 14000
rect 2884 13960 3976 13988
rect 1946 13920 1952 13932
rect 1907 13892 1952 13920
rect 1946 13880 1952 13892
rect 2004 13880 2010 13932
rect 2130 13880 2136 13932
rect 2188 13920 2194 13932
rect 2884 13929 2912 13960
rect 3970 13948 3976 13960
rect 4028 13948 4034 14000
rect 2225 13923 2283 13929
rect 2225 13920 2237 13923
rect 2188 13892 2237 13920
rect 2188 13880 2194 13892
rect 2225 13889 2237 13892
rect 2271 13889 2283 13923
rect 2225 13883 2283 13889
rect 2869 13923 2927 13929
rect 2869 13889 2881 13923
rect 2915 13889 2927 13923
rect 3510 13920 3516 13932
rect 3471 13892 3516 13920
rect 2869 13883 2927 13889
rect 3510 13880 3516 13892
rect 3568 13880 3574 13932
rect 3605 13923 3663 13929
rect 3605 13889 3617 13923
rect 3651 13920 3663 13923
rect 4246 13920 4252 13932
rect 3651 13892 4252 13920
rect 3651 13889 3663 13892
rect 3605 13883 3663 13889
rect 4246 13880 4252 13892
rect 4304 13880 4310 13932
rect 4341 13923 4399 13929
rect 4341 13889 4353 13923
rect 4387 13920 4399 13923
rect 4448 13920 4476 14019
rect 5718 14016 5724 14028
rect 5776 14016 5782 14068
rect 8110 14056 8116 14068
rect 6840 14028 8116 14056
rect 4522 13948 4528 14000
rect 4580 13988 4586 14000
rect 5537 13991 5595 13997
rect 5537 13988 5549 13991
rect 4580 13960 5549 13988
rect 4580 13948 4586 13960
rect 5537 13957 5549 13960
rect 5583 13957 5595 13991
rect 5537 13951 5595 13957
rect 4614 13920 4620 13932
rect 4387 13892 4476 13920
rect 4575 13892 4620 13920
rect 4387 13889 4399 13892
rect 4341 13883 4399 13889
rect 4614 13880 4620 13892
rect 4672 13880 4678 13932
rect 4709 13923 4767 13929
rect 4709 13889 4721 13923
rect 4755 13920 4767 13923
rect 5074 13920 5080 13932
rect 4755 13892 5080 13920
rect 4755 13889 4767 13892
rect 4709 13883 4767 13889
rect 5074 13880 5080 13892
rect 5132 13880 5138 13932
rect 5258 13920 5264 13932
rect 5219 13892 5264 13920
rect 5258 13880 5264 13892
rect 5316 13880 5322 13932
rect 6840 13929 6868 14028
rect 8110 14016 8116 14028
rect 8168 14016 8174 14068
rect 8205 14059 8263 14065
rect 8205 14025 8217 14059
rect 8251 14056 8263 14059
rect 9766 14056 9772 14068
rect 8251 14028 9772 14056
rect 8251 14025 8263 14028
rect 8205 14019 8263 14025
rect 9766 14016 9772 14028
rect 9824 14016 9830 14068
rect 9861 14059 9919 14065
rect 9861 14025 9873 14059
rect 9907 14056 9919 14059
rect 12434 14056 12440 14068
rect 9907 14028 12440 14056
rect 9907 14025 9919 14028
rect 9861 14019 9919 14025
rect 12434 14016 12440 14028
rect 12492 14016 12498 14068
rect 12802 14016 12808 14068
rect 12860 14056 12866 14068
rect 15105 14059 15163 14065
rect 15105 14056 15117 14059
rect 12860 14028 15117 14056
rect 12860 14016 12866 14028
rect 15105 14025 15117 14028
rect 15151 14025 15163 14059
rect 15105 14019 15163 14025
rect 16298 14016 16304 14068
rect 16356 14056 16362 14068
rect 16356 14028 16712 14056
rect 16356 14016 16362 14028
rect 7282 13948 7288 14000
rect 7340 13988 7346 14000
rect 8570 13997 8576 14000
rect 8564 13988 8576 13997
rect 7340 13960 8340 13988
rect 8531 13960 8576 13988
rect 7340 13948 7346 13960
rect 6825 13923 6883 13929
rect 6825 13889 6837 13923
rect 6871 13889 6883 13923
rect 6825 13883 6883 13889
rect 7092 13923 7150 13929
rect 7092 13889 7104 13923
rect 7138 13920 7150 13923
rect 8202 13920 8208 13932
rect 7138 13892 8208 13920
rect 7138 13889 7150 13892
rect 7092 13883 7150 13889
rect 8202 13880 8208 13892
rect 8260 13880 8266 13932
rect 8312 13920 8340 13960
rect 8564 13951 8576 13960
rect 8570 13948 8576 13951
rect 8628 13948 8634 14000
rect 9306 13948 9312 14000
rect 9364 13988 9370 14000
rect 9364 13960 11284 13988
rect 9364 13948 9370 13960
rect 11054 13920 11060 13932
rect 11112 13929 11118 13932
rect 8312 13892 9996 13920
rect 11024 13892 11060 13920
rect 2958 13812 2964 13864
rect 3016 13852 3022 13864
rect 3145 13855 3203 13861
rect 3145 13852 3157 13855
rect 3016 13824 3157 13852
rect 3016 13812 3022 13824
rect 3145 13821 3157 13824
rect 3191 13852 3203 13855
rect 3191 13824 3280 13852
rect 3191 13821 3203 13824
rect 3145 13815 3203 13821
rect 3252 13784 3280 13824
rect 3326 13812 3332 13864
rect 3384 13852 3390 13864
rect 5353 13855 5411 13861
rect 5353 13852 5365 13855
rect 3384 13824 3429 13852
rect 3620 13824 5365 13852
rect 3384 13812 3390 13824
rect 3620 13784 3648 13824
rect 5353 13821 5365 13824
rect 5399 13821 5411 13855
rect 5353 13815 5411 13821
rect 8110 13812 8116 13864
rect 8168 13852 8174 13864
rect 8297 13855 8355 13861
rect 8297 13852 8309 13855
rect 8168 13824 8309 13852
rect 8168 13812 8174 13824
rect 8297 13821 8309 13824
rect 8343 13821 8355 13855
rect 8297 13815 8355 13821
rect 9490 13812 9496 13864
rect 9548 13852 9554 13864
rect 9548 13824 9904 13852
rect 9548 13812 9554 13824
rect 3252 13756 3648 13784
rect 3973 13719 4031 13725
rect 3973 13685 3985 13719
rect 4019 13716 4031 13719
rect 4338 13716 4344 13728
rect 4019 13688 4344 13716
rect 4019 13685 4031 13688
rect 3973 13679 4031 13685
rect 4338 13676 4344 13688
rect 4396 13676 4402 13728
rect 9582 13676 9588 13728
rect 9640 13716 9646 13728
rect 9677 13719 9735 13725
rect 9677 13716 9689 13719
rect 9640 13688 9689 13716
rect 9640 13676 9646 13688
rect 9677 13685 9689 13688
rect 9723 13685 9735 13719
rect 9876 13716 9904 13824
rect 9968 13793 9996 13892
rect 11054 13880 11060 13892
rect 11112 13883 11124 13929
rect 11112 13880 11118 13883
rect 11256 13852 11284 13960
rect 13722 13948 13728 14000
rect 13780 13988 13786 14000
rect 14829 13991 14887 13997
rect 13780 13960 14780 13988
rect 13780 13948 13786 13960
rect 11330 13880 11336 13932
rect 11388 13920 11394 13932
rect 12630 13923 12688 13929
rect 12630 13920 12642 13923
rect 11388 13892 11433 13920
rect 11624 13892 12642 13920
rect 11388 13880 11394 13892
rect 11256 13824 11560 13852
rect 11532 13793 11560 13824
rect 9953 13787 10011 13793
rect 9953 13753 9965 13787
rect 9999 13753 10011 13787
rect 9953 13747 10011 13753
rect 11517 13787 11575 13793
rect 11517 13753 11529 13787
rect 11563 13753 11575 13787
rect 11517 13747 11575 13753
rect 11624 13716 11652 13892
rect 12630 13889 12642 13892
rect 12676 13920 12688 13923
rect 12802 13920 12808 13932
rect 12676 13892 12808 13920
rect 12676 13889 12688 13892
rect 12630 13883 12688 13889
rect 12802 13880 12808 13892
rect 12860 13880 12866 13932
rect 13170 13880 13176 13932
rect 13228 13920 13234 13932
rect 13337 13923 13395 13929
rect 13337 13920 13349 13923
rect 13228 13892 13349 13920
rect 13228 13880 13234 13892
rect 13337 13889 13349 13892
rect 13383 13889 13395 13923
rect 14752 13920 14780 13960
rect 14829 13957 14841 13991
rect 14875 13988 14887 13991
rect 15194 13988 15200 14000
rect 14875 13960 15200 13988
rect 14875 13957 14887 13960
rect 14829 13951 14887 13957
rect 15194 13948 15200 13960
rect 15252 13948 15258 14000
rect 16206 13948 16212 14000
rect 16264 13997 16270 14000
rect 16264 13988 16276 13997
rect 16264 13960 16309 13988
rect 16264 13951 16276 13960
rect 16264 13948 16270 13951
rect 16684 13929 16712 14028
rect 16485 13923 16543 13929
rect 14752 13892 16436 13920
rect 13337 13883 13395 13889
rect 12897 13855 12955 13861
rect 12897 13821 12909 13855
rect 12943 13852 12955 13855
rect 12986 13852 12992 13864
rect 12943 13824 12992 13852
rect 12943 13821 12955 13824
rect 12897 13815 12955 13821
rect 12986 13812 12992 13824
rect 13044 13852 13050 13864
rect 13081 13855 13139 13861
rect 13081 13852 13093 13855
rect 13044 13824 13093 13852
rect 13044 13812 13050 13824
rect 13081 13821 13093 13824
rect 13127 13821 13139 13855
rect 13081 13815 13139 13821
rect 14182 13812 14188 13864
rect 14240 13852 14246 13864
rect 14642 13852 14648 13864
rect 14240 13824 14504 13852
rect 14603 13824 14648 13852
rect 14240 13812 14246 13824
rect 14476 13793 14504 13824
rect 14642 13812 14648 13824
rect 14700 13812 14706 13864
rect 16408 13852 16436 13892
rect 16485 13889 16497 13923
rect 16531 13920 16543 13923
rect 16669 13923 16727 13929
rect 16669 13920 16681 13923
rect 16531 13892 16681 13920
rect 16531 13889 16543 13892
rect 16485 13883 16543 13889
rect 16669 13889 16681 13892
rect 16715 13889 16727 13923
rect 16925 13923 16983 13929
rect 16925 13920 16937 13923
rect 16669 13883 16727 13889
rect 16776 13892 16937 13920
rect 16776 13852 16804 13892
rect 16925 13889 16937 13892
rect 16971 13889 16983 13923
rect 18414 13920 18420 13932
rect 16925 13883 16983 13889
rect 17972 13892 18420 13920
rect 17972 13852 18000 13892
rect 18414 13880 18420 13892
rect 18472 13880 18478 13932
rect 16408 13824 16804 13852
rect 17696 13824 18000 13852
rect 18233 13855 18291 13861
rect 14461 13787 14519 13793
rect 14461 13753 14473 13787
rect 14507 13753 14519 13787
rect 14461 13747 14519 13753
rect 14734 13744 14740 13796
rect 14792 13784 14798 13796
rect 14792 13756 15608 13784
rect 14792 13744 14798 13756
rect 9876 13688 11652 13716
rect 9677 13679 9735 13685
rect 11698 13676 11704 13728
rect 11756 13716 11762 13728
rect 12710 13716 12716 13728
rect 11756 13688 12716 13716
rect 11756 13676 11762 13688
rect 12710 13676 12716 13688
rect 12768 13676 12774 13728
rect 12894 13676 12900 13728
rect 12952 13716 12958 13728
rect 14918 13716 14924 13728
rect 12952 13688 14924 13716
rect 12952 13676 12958 13688
rect 14918 13676 14924 13688
rect 14976 13676 14982 13728
rect 15580 13716 15608 13756
rect 17696 13716 17724 13824
rect 18233 13821 18245 13855
rect 18279 13852 18291 13855
rect 18322 13852 18328 13864
rect 18279 13824 18328 13852
rect 18279 13821 18291 13824
rect 18233 13815 18291 13821
rect 18322 13812 18328 13824
rect 18380 13812 18386 13864
rect 18046 13716 18052 13728
rect 15580 13688 17724 13716
rect 18007 13688 18052 13716
rect 18046 13676 18052 13688
rect 18104 13676 18110 13728
rect 1104 13626 18860 13648
rect 1104 13574 3174 13626
rect 3226 13574 3238 13626
rect 3290 13574 3302 13626
rect 3354 13574 3366 13626
rect 3418 13574 3430 13626
rect 3482 13574 7622 13626
rect 7674 13574 7686 13626
rect 7738 13574 7750 13626
rect 7802 13574 7814 13626
rect 7866 13574 7878 13626
rect 7930 13574 12070 13626
rect 12122 13574 12134 13626
rect 12186 13574 12198 13626
rect 12250 13574 12262 13626
rect 12314 13574 12326 13626
rect 12378 13574 16518 13626
rect 16570 13574 16582 13626
rect 16634 13574 16646 13626
rect 16698 13574 16710 13626
rect 16762 13574 16774 13626
rect 16826 13574 18860 13626
rect 1104 13552 18860 13574
rect 3053 13515 3111 13521
rect 3053 13481 3065 13515
rect 3099 13512 3111 13515
rect 4982 13512 4988 13524
rect 3099 13484 4988 13512
rect 3099 13481 3111 13484
rect 3053 13475 3111 13481
rect 4982 13472 4988 13484
rect 5040 13472 5046 13524
rect 5537 13515 5595 13521
rect 5537 13481 5549 13515
rect 5583 13512 5595 13515
rect 5810 13512 5816 13524
rect 5583 13484 5816 13512
rect 5583 13481 5595 13484
rect 5537 13475 5595 13481
rect 5810 13472 5816 13484
rect 5868 13472 5874 13524
rect 9398 13472 9404 13524
rect 9456 13512 9462 13524
rect 11793 13515 11851 13521
rect 9456 13484 11652 13512
rect 9456 13472 9462 13484
rect 2774 13404 2780 13456
rect 2832 13444 2838 13456
rect 3237 13447 3295 13453
rect 3237 13444 3249 13447
rect 2832 13416 3249 13444
rect 2832 13404 2838 13416
rect 3237 13413 3249 13416
rect 3283 13413 3295 13447
rect 3510 13444 3516 13456
rect 3237 13407 3295 13413
rect 3344 13416 3516 13444
rect 1946 13376 1952 13388
rect 1907 13348 1952 13376
rect 1946 13336 1952 13348
rect 2004 13336 2010 13388
rect 2501 13379 2559 13385
rect 2501 13345 2513 13379
rect 2547 13376 2559 13379
rect 3344 13376 3372 13416
rect 3510 13404 3516 13416
rect 3568 13444 3574 13456
rect 4062 13444 4068 13456
rect 3568 13416 4068 13444
rect 3568 13404 3574 13416
rect 4062 13404 4068 13416
rect 4120 13404 4126 13456
rect 11624 13444 11652 13484
rect 11793 13481 11805 13515
rect 11839 13512 11851 13515
rect 13998 13512 14004 13524
rect 11839 13484 14004 13512
rect 11839 13481 11851 13484
rect 11793 13475 11851 13481
rect 13998 13472 14004 13484
rect 14056 13472 14062 13524
rect 16390 13472 16396 13524
rect 16448 13512 16454 13524
rect 16448 13484 17264 13512
rect 16448 13472 16454 13484
rect 11624 13416 12434 13444
rect 2547 13348 3372 13376
rect 2547 13345 2559 13348
rect 2501 13339 2559 13345
rect 3602 13336 3608 13388
rect 3660 13376 3666 13388
rect 3660 13348 4200 13376
rect 3660 13336 3666 13348
rect 1854 13268 1860 13320
rect 1912 13308 1918 13320
rect 2225 13311 2283 13317
rect 2225 13308 2237 13311
rect 1912 13280 2237 13308
rect 1912 13268 1918 13280
rect 2225 13277 2237 13280
rect 2271 13277 2283 13311
rect 2225 13271 2283 13277
rect 3421 13311 3479 13317
rect 3421 13277 3433 13311
rect 3467 13308 3479 13311
rect 3510 13308 3516 13320
rect 3467 13280 3516 13308
rect 3467 13277 3479 13280
rect 3421 13271 3479 13277
rect 3510 13268 3516 13280
rect 3568 13268 3574 13320
rect 4172 13317 4200 13348
rect 4246 13336 4252 13388
rect 4304 13376 4310 13388
rect 4525 13379 4583 13385
rect 4525 13376 4537 13379
rect 4304 13348 4537 13376
rect 4304 13336 4310 13348
rect 4525 13345 4537 13348
rect 4571 13345 4583 13379
rect 4525 13339 4583 13345
rect 11974 13336 11980 13388
rect 12032 13376 12038 13388
rect 12069 13379 12127 13385
rect 12069 13376 12081 13379
rect 12032 13348 12081 13376
rect 12032 13336 12038 13348
rect 12069 13345 12081 13348
rect 12115 13345 12127 13379
rect 12406 13376 12434 13416
rect 12894 13376 12900 13388
rect 12406 13348 12900 13376
rect 12069 13339 12127 13345
rect 12894 13336 12900 13348
rect 12952 13336 12958 13388
rect 17126 13376 17132 13388
rect 17087 13348 17132 13376
rect 17126 13336 17132 13348
rect 17184 13336 17190 13388
rect 4065 13311 4123 13317
rect 4065 13277 4077 13311
rect 4111 13277 4123 13311
rect 4065 13271 4123 13277
rect 4157 13311 4215 13317
rect 4157 13277 4169 13311
rect 4203 13277 4215 13311
rect 4157 13271 4215 13277
rect 2593 13243 2651 13249
rect 2593 13209 2605 13243
rect 2639 13240 2651 13243
rect 2958 13240 2964 13252
rect 2639 13212 2964 13240
rect 2639 13209 2651 13212
rect 2593 13203 2651 13209
rect 2958 13200 2964 13212
rect 3016 13200 3022 13252
rect 4080 13240 4108 13271
rect 4614 13268 4620 13320
rect 4672 13308 4678 13320
rect 4672 13280 4936 13308
rect 4672 13268 4678 13280
rect 4798 13240 4804 13252
rect 4080 13212 4804 13240
rect 4798 13200 4804 13212
rect 4856 13200 4862 13252
rect 4908 13240 4936 13280
rect 5166 13268 5172 13320
rect 5224 13308 5230 13320
rect 5224 13280 5269 13308
rect 5224 13268 5230 13280
rect 8110 13268 8116 13320
rect 8168 13308 8174 13320
rect 8757 13311 8815 13317
rect 8757 13308 8769 13311
rect 8168 13280 8769 13308
rect 8168 13268 8174 13280
rect 8757 13277 8769 13280
rect 8803 13277 8815 13311
rect 8757 13271 8815 13277
rect 9214 13268 9220 13320
rect 9272 13308 9278 13320
rect 9272 13280 11468 13308
rect 9272 13268 9278 13280
rect 8478 13240 8484 13252
rect 8536 13249 8542 13252
rect 4908 13212 8484 13240
rect 8478 13200 8484 13212
rect 8536 13203 8548 13249
rect 11342 13243 11400 13249
rect 11342 13240 11354 13243
rect 8588 13212 11354 13240
rect 8536 13200 8542 13203
rect 2682 13172 2688 13184
rect 2643 13144 2688 13172
rect 2682 13132 2688 13144
rect 2740 13132 2746 13184
rect 3326 13132 3332 13184
rect 3384 13172 3390 13184
rect 3513 13175 3571 13181
rect 3513 13172 3525 13175
rect 3384 13144 3525 13172
rect 3384 13132 3390 13144
rect 3513 13141 3525 13144
rect 3559 13141 3571 13175
rect 3878 13172 3884 13184
rect 3839 13144 3884 13172
rect 3513 13135 3571 13141
rect 3878 13132 3884 13144
rect 3936 13132 3942 13184
rect 3970 13132 3976 13184
rect 4028 13172 4034 13184
rect 4341 13175 4399 13181
rect 4341 13172 4353 13175
rect 4028 13144 4353 13172
rect 4028 13132 4034 13144
rect 4341 13141 4353 13144
rect 4387 13141 4399 13175
rect 4341 13135 4399 13141
rect 4985 13175 5043 13181
rect 4985 13141 4997 13175
rect 5031 13172 5043 13175
rect 5074 13172 5080 13184
rect 5031 13144 5080 13172
rect 5031 13141 5043 13144
rect 4985 13135 5043 13141
rect 5074 13132 5080 13144
rect 5132 13132 5138 13184
rect 5258 13172 5264 13184
rect 5219 13144 5264 13172
rect 5258 13132 5264 13144
rect 5316 13132 5322 13184
rect 7374 13172 7380 13184
rect 7335 13144 7380 13172
rect 7374 13132 7380 13144
rect 7432 13132 7438 13184
rect 7466 13132 7472 13184
rect 7524 13172 7530 13184
rect 8588 13172 8616 13212
rect 11342 13209 11354 13212
rect 11388 13209 11400 13243
rect 11440 13240 11468 13280
rect 11514 13268 11520 13320
rect 11572 13308 11578 13320
rect 11609 13311 11667 13317
rect 11609 13308 11621 13311
rect 11572 13280 11621 13308
rect 11572 13268 11578 13280
rect 11609 13277 11621 13280
rect 11655 13277 11667 13311
rect 11609 13271 11667 13277
rect 13078 13268 13084 13320
rect 13136 13308 13142 13320
rect 13136 13280 13584 13308
rect 13136 13268 13142 13280
rect 11790 13240 11796 13252
rect 11440 13212 11796 13240
rect 11342 13203 11400 13209
rect 11790 13200 11796 13212
rect 11848 13200 11854 13252
rect 11977 13243 12035 13249
rect 11977 13209 11989 13243
rect 12023 13240 12035 13243
rect 12253 13243 12311 13249
rect 12253 13240 12265 13243
rect 12023 13212 12265 13240
rect 12023 13209 12035 13212
rect 11977 13203 12035 13209
rect 12253 13209 12265 13212
rect 12299 13240 12311 13243
rect 13446 13240 13452 13252
rect 12299 13212 13452 13240
rect 12299 13209 12311 13212
rect 12253 13203 12311 13209
rect 13446 13200 13452 13212
rect 13504 13200 13510 13252
rect 13556 13240 13584 13280
rect 13630 13268 13636 13320
rect 13688 13317 13694 13320
rect 13688 13308 13700 13317
rect 13909 13311 13967 13317
rect 13688 13280 13733 13308
rect 13688 13271 13700 13280
rect 13909 13277 13921 13311
rect 13955 13277 13967 13311
rect 13909 13271 13967 13277
rect 13688 13268 13694 13271
rect 13924 13240 13952 13271
rect 14182 13268 14188 13320
rect 14240 13308 14246 13320
rect 15206 13311 15264 13317
rect 15206 13308 15218 13311
rect 14240 13280 15218 13308
rect 14240 13268 14246 13280
rect 15206 13277 15218 13280
rect 15252 13277 15264 13311
rect 15470 13308 15476 13320
rect 15431 13280 15476 13308
rect 15206 13271 15264 13277
rect 15470 13268 15476 13280
rect 15528 13268 15534 13320
rect 17236 13317 17264 13484
rect 17862 13472 17868 13524
rect 17920 13512 17926 13524
rect 18325 13515 18383 13521
rect 18325 13512 18337 13515
rect 17920 13484 18337 13512
rect 17920 13472 17926 13484
rect 18325 13481 18337 13484
rect 18371 13481 18383 13515
rect 18325 13475 18383 13481
rect 17402 13336 17408 13388
rect 17460 13376 17466 13388
rect 17589 13379 17647 13385
rect 17589 13376 17601 13379
rect 17460 13348 17601 13376
rect 17460 13336 17466 13348
rect 17589 13345 17601 13348
rect 17635 13345 17647 13379
rect 17589 13339 17647 13345
rect 17221 13311 17279 13317
rect 17221 13277 17233 13311
rect 17267 13277 17279 13311
rect 17221 13271 17279 13277
rect 17770 13268 17776 13320
rect 17828 13308 17834 13320
rect 18509 13311 18567 13317
rect 18509 13308 18521 13311
rect 17828 13280 18521 13308
rect 17828 13268 17834 13280
rect 18509 13277 18521 13280
rect 18555 13277 18567 13311
rect 18509 13271 18567 13277
rect 15565 13243 15623 13249
rect 15565 13240 15577 13243
rect 13556 13212 13952 13240
rect 14016 13212 15577 13240
rect 7524 13144 8616 13172
rect 10229 13175 10287 13181
rect 7524 13132 7530 13144
rect 10229 13141 10241 13175
rect 10275 13172 10287 13175
rect 10778 13172 10784 13184
rect 10275 13144 10784 13172
rect 10275 13141 10287 13144
rect 10229 13135 10287 13141
rect 10778 13132 10784 13144
rect 10836 13132 10842 13184
rect 12066 13132 12072 13184
rect 12124 13172 12130 13184
rect 12529 13175 12587 13181
rect 12529 13172 12541 13175
rect 12124 13144 12541 13172
rect 12124 13132 12130 13144
rect 12529 13141 12541 13144
rect 12575 13141 12587 13175
rect 12529 13135 12587 13141
rect 12710 13132 12716 13184
rect 12768 13172 12774 13184
rect 14016 13172 14044 13212
rect 15565 13209 15577 13212
rect 15611 13240 15623 13243
rect 16206 13240 16212 13252
rect 15611 13212 16212 13240
rect 15611 13209 15623 13212
rect 15565 13203 15623 13209
rect 16206 13200 16212 13212
rect 16264 13200 16270 13252
rect 16850 13240 16856 13252
rect 16908 13249 16914 13252
rect 16820 13212 16856 13240
rect 16850 13200 16856 13212
rect 16908 13203 16920 13249
rect 16908 13200 16914 13203
rect 12768 13144 14044 13172
rect 12768 13132 12774 13144
rect 14090 13132 14096 13184
rect 14148 13172 14154 13184
rect 15749 13175 15807 13181
rect 14148 13144 14193 13172
rect 14148 13132 14154 13144
rect 15749 13141 15761 13175
rect 15795 13172 15807 13175
rect 17770 13172 17776 13184
rect 15795 13144 17776 13172
rect 15795 13141 15807 13144
rect 15749 13135 15807 13141
rect 17770 13132 17776 13144
rect 17828 13132 17834 13184
rect 1104 13082 18860 13104
rect 1104 13030 5398 13082
rect 5450 13030 5462 13082
rect 5514 13030 5526 13082
rect 5578 13030 5590 13082
rect 5642 13030 5654 13082
rect 5706 13030 9846 13082
rect 9898 13030 9910 13082
rect 9962 13030 9974 13082
rect 10026 13030 10038 13082
rect 10090 13030 10102 13082
rect 10154 13030 14294 13082
rect 14346 13030 14358 13082
rect 14410 13030 14422 13082
rect 14474 13030 14486 13082
rect 14538 13030 14550 13082
rect 14602 13030 18860 13082
rect 1104 13008 18860 13030
rect 2314 12968 2320 12980
rect 2275 12940 2320 12968
rect 2314 12928 2320 12940
rect 2372 12928 2378 12980
rect 2777 12971 2835 12977
rect 2777 12937 2789 12971
rect 2823 12968 2835 12971
rect 3513 12971 3571 12977
rect 2823 12940 3464 12968
rect 2823 12937 2835 12940
rect 2777 12931 2835 12937
rect 2685 12903 2743 12909
rect 2685 12869 2697 12903
rect 2731 12900 2743 12903
rect 2866 12900 2872 12912
rect 2731 12872 2872 12900
rect 2731 12869 2743 12872
rect 2685 12863 2743 12869
rect 2866 12860 2872 12872
rect 2924 12860 2930 12912
rect 3436 12900 3464 12940
rect 3513 12937 3525 12971
rect 3559 12968 3571 12971
rect 3973 12971 4031 12977
rect 3973 12968 3985 12971
rect 3559 12940 3985 12968
rect 3559 12937 3571 12940
rect 3513 12931 3571 12937
rect 3973 12937 3985 12940
rect 4019 12937 4031 12971
rect 4338 12968 4344 12980
rect 4299 12940 4344 12968
rect 3973 12931 4031 12937
rect 4338 12928 4344 12940
rect 4396 12928 4402 12980
rect 4798 12968 4804 12980
rect 4759 12940 4804 12968
rect 4798 12928 4804 12940
rect 4856 12928 4862 12980
rect 5074 12928 5080 12980
rect 5132 12968 5138 12980
rect 5258 12968 5264 12980
rect 5132 12940 5264 12968
rect 5132 12928 5138 12940
rect 5258 12928 5264 12940
rect 5316 12968 5322 12980
rect 5316 12940 5948 12968
rect 5316 12928 5322 12940
rect 3694 12900 3700 12912
rect 3436 12872 3700 12900
rect 3694 12860 3700 12872
rect 3752 12860 3758 12912
rect 3878 12860 3884 12912
rect 3936 12900 3942 12912
rect 5813 12903 5871 12909
rect 5813 12900 5825 12903
rect 3936 12872 5825 12900
rect 3936 12860 3942 12872
rect 5813 12869 5825 12872
rect 5859 12869 5871 12903
rect 5813 12863 5871 12869
rect 1762 12792 1768 12844
rect 1820 12832 1826 12844
rect 3326 12832 3332 12844
rect 1820 12804 3332 12832
rect 1820 12792 1826 12804
rect 1949 12767 2007 12773
rect 1949 12733 1961 12767
rect 1995 12764 2007 12767
rect 2130 12764 2136 12776
rect 1995 12736 2136 12764
rect 1995 12733 2007 12736
rect 1949 12727 2007 12733
rect 2130 12724 2136 12736
rect 2188 12724 2194 12776
rect 2976 12773 3004 12804
rect 3326 12792 3332 12804
rect 3384 12792 3390 12844
rect 3421 12835 3479 12841
rect 3421 12801 3433 12835
rect 3467 12832 3479 12835
rect 4706 12832 4712 12844
rect 3467 12804 4712 12832
rect 3467 12801 3479 12804
rect 3421 12795 3479 12801
rect 4706 12792 4712 12804
rect 4764 12792 4770 12844
rect 4985 12835 5043 12841
rect 4985 12801 4997 12835
rect 5031 12801 5043 12835
rect 5258 12832 5264 12844
rect 5219 12804 5264 12832
rect 4985 12795 5043 12801
rect 2225 12767 2283 12773
rect 2225 12733 2237 12767
rect 2271 12733 2283 12767
rect 2225 12727 2283 12733
rect 2961 12767 3019 12773
rect 2961 12733 2973 12767
rect 3007 12733 3019 12767
rect 3234 12764 3240 12776
rect 3195 12736 3240 12764
rect 2961 12727 3019 12733
rect 2240 12696 2268 12727
rect 3234 12724 3240 12736
rect 3292 12724 3298 12776
rect 3878 12724 3884 12776
rect 3936 12724 3942 12776
rect 4430 12764 4436 12776
rect 4391 12736 4436 12764
rect 4430 12724 4436 12736
rect 4488 12724 4494 12776
rect 4614 12764 4620 12776
rect 4575 12736 4620 12764
rect 4614 12724 4620 12736
rect 4672 12724 4678 12776
rect 5000 12764 5028 12795
rect 5258 12792 5264 12804
rect 5316 12792 5322 12844
rect 5534 12832 5540 12844
rect 5495 12804 5540 12832
rect 5534 12792 5540 12804
rect 5592 12832 5598 12844
rect 5629 12835 5687 12841
rect 5629 12832 5641 12835
rect 5592 12804 5641 12832
rect 5592 12792 5598 12804
rect 5629 12801 5641 12804
rect 5675 12801 5687 12835
rect 5920 12832 5948 12940
rect 6178 12928 6184 12980
rect 6236 12968 6242 12980
rect 10965 12971 11023 12977
rect 10965 12968 10977 12971
rect 6236 12940 10977 12968
rect 6236 12928 6242 12940
rect 10965 12937 10977 12940
rect 11011 12937 11023 12971
rect 10965 12931 11023 12937
rect 11333 12971 11391 12977
rect 11333 12937 11345 12971
rect 11379 12968 11391 12971
rect 11379 12940 18460 12968
rect 11379 12937 11391 12940
rect 11333 12931 11391 12937
rect 8110 12860 8116 12912
rect 8168 12900 8174 12912
rect 8168 12872 9536 12900
rect 8168 12860 8174 12872
rect 8846 12832 8852 12844
rect 5920 12804 8852 12832
rect 5629 12795 5687 12801
rect 8846 12792 8852 12804
rect 8904 12792 8910 12844
rect 9237 12835 9295 12841
rect 9237 12801 9249 12835
rect 9283 12832 9295 12835
rect 9398 12832 9404 12844
rect 9283 12804 9404 12832
rect 9283 12801 9295 12804
rect 9237 12795 9295 12801
rect 9398 12792 9404 12804
rect 9456 12792 9462 12844
rect 9508 12841 9536 12872
rect 9674 12860 9680 12912
rect 9732 12900 9738 12912
rect 9830 12903 9888 12909
rect 9830 12900 9842 12903
rect 9732 12872 9842 12900
rect 9732 12860 9738 12872
rect 9830 12869 9842 12872
rect 9876 12869 9888 12903
rect 10980 12900 11008 12931
rect 11698 12900 11704 12912
rect 10980 12872 11704 12900
rect 9830 12863 9888 12869
rect 11698 12860 11704 12872
rect 11756 12860 11762 12912
rect 12986 12900 12992 12912
rect 12544 12872 12992 12900
rect 9493 12835 9551 12841
rect 9493 12801 9505 12835
rect 9539 12832 9551 12835
rect 9585 12835 9643 12841
rect 9585 12832 9597 12835
rect 9539 12804 9597 12832
rect 9539 12801 9551 12804
rect 9493 12795 9551 12801
rect 9585 12801 9597 12804
rect 9631 12832 9643 12835
rect 11422 12832 11428 12844
rect 9631 12804 11428 12832
rect 9631 12801 9643 12804
rect 9585 12795 9643 12801
rect 11422 12792 11428 12804
rect 11480 12832 11486 12844
rect 12544 12832 12572 12872
rect 11480 12804 12572 12832
rect 11480 12792 11486 12804
rect 12618 12792 12624 12844
rect 12676 12841 12682 12844
rect 12912 12841 12940 12872
rect 12986 12860 12992 12872
rect 13044 12900 13050 12912
rect 13044 12872 14872 12900
rect 13044 12860 13050 12872
rect 12676 12832 12688 12841
rect 12897 12835 12955 12841
rect 12676 12804 12721 12832
rect 12676 12795 12688 12804
rect 12897 12801 12909 12835
rect 12943 12801 12955 12835
rect 12897 12795 12955 12801
rect 13173 12835 13231 12841
rect 13173 12801 13185 12835
rect 13219 12832 13231 12835
rect 13446 12832 13452 12844
rect 13219 12804 13452 12832
rect 13219 12801 13231 12804
rect 13173 12795 13231 12801
rect 12676 12792 12682 12795
rect 13446 12792 13452 12804
rect 13504 12792 13510 12844
rect 14844 12841 14872 12872
rect 15470 12860 15476 12912
rect 15528 12900 15534 12912
rect 16298 12900 16304 12912
rect 15528 12872 16304 12900
rect 15528 12860 15534 12872
rect 14573 12835 14631 12841
rect 14573 12801 14585 12835
rect 14619 12832 14631 12835
rect 14829 12835 14887 12841
rect 14619 12804 14780 12832
rect 14619 12801 14631 12804
rect 14573 12795 14631 12801
rect 5166 12764 5172 12776
rect 5000 12736 5172 12764
rect 5166 12724 5172 12736
rect 5224 12724 5230 12776
rect 7466 12724 7472 12776
rect 7524 12764 7530 12776
rect 14752 12764 14780 12804
rect 14829 12801 14841 12835
rect 14875 12801 14887 12835
rect 14829 12795 14887 12801
rect 16022 12792 16028 12844
rect 16080 12841 16086 12844
rect 16080 12832 16092 12841
rect 16233 12832 16261 12872
rect 16298 12860 16304 12872
rect 16356 12860 16362 12912
rect 16482 12900 16488 12912
rect 16443 12872 16488 12900
rect 16482 12860 16488 12872
rect 16540 12860 16546 12912
rect 17126 12900 17132 12912
rect 16684 12872 17132 12900
rect 16684 12841 16712 12872
rect 17126 12860 17132 12872
rect 17184 12900 17190 12912
rect 17402 12900 17408 12912
rect 17184 12872 17408 12900
rect 17184 12860 17190 12872
rect 17402 12860 17408 12872
rect 17460 12860 17466 12912
rect 18230 12900 18236 12912
rect 18191 12872 18236 12900
rect 18230 12860 18236 12872
rect 18288 12860 18294 12912
rect 18432 12909 18460 12940
rect 18417 12903 18475 12909
rect 18417 12869 18429 12903
rect 18463 12900 18475 12903
rect 18506 12900 18512 12912
rect 18463 12872 18512 12900
rect 18463 12869 18475 12872
rect 18417 12863 18475 12869
rect 18506 12860 18512 12872
rect 18564 12860 18570 12912
rect 16669 12835 16727 12841
rect 16669 12832 16681 12835
rect 16080 12804 16125 12832
rect 16233 12804 16681 12832
rect 16080 12795 16092 12804
rect 16080 12792 16086 12795
rect 15010 12764 15016 12776
rect 7524 12736 8156 12764
rect 14752 12736 15016 12764
rect 7524 12724 7530 12736
rect 3050 12696 3056 12708
rect 2240 12668 3056 12696
rect 3050 12656 3056 12668
rect 3108 12696 3114 12708
rect 3896 12696 3924 12724
rect 3108 12668 3924 12696
rect 3108 12656 3114 12668
rect 4154 12656 4160 12708
rect 4212 12656 4218 12708
rect 8128 12705 8156 12736
rect 15010 12724 15016 12736
rect 15068 12724 15074 12776
rect 16316 12773 16344 12804
rect 16669 12801 16681 12804
rect 16715 12801 16727 12835
rect 16669 12795 16727 12801
rect 16936 12835 16994 12841
rect 16936 12801 16948 12835
rect 16982 12832 16994 12835
rect 17310 12832 17316 12844
rect 16982 12804 17316 12832
rect 16982 12801 16994 12804
rect 16936 12795 16994 12801
rect 17310 12792 17316 12804
rect 17368 12792 17374 12844
rect 16301 12767 16359 12773
rect 16301 12733 16313 12767
rect 16347 12764 16359 12767
rect 16347 12736 16381 12764
rect 16347 12733 16359 12736
rect 16301 12727 16359 12733
rect 8113 12699 8171 12705
rect 8113 12665 8125 12699
rect 8159 12665 8171 12699
rect 8113 12659 8171 12665
rect 10594 12656 10600 12708
rect 10652 12696 10658 12708
rect 10652 12668 11192 12696
rect 10652 12656 10658 12668
rect 1302 12588 1308 12640
rect 1360 12628 1366 12640
rect 3881 12631 3939 12637
rect 3881 12628 3893 12631
rect 1360 12600 3893 12628
rect 1360 12588 1366 12600
rect 3881 12597 3893 12600
rect 3927 12597 3939 12631
rect 4172 12628 4200 12656
rect 5077 12631 5135 12637
rect 5077 12628 5089 12631
rect 4172 12600 5089 12628
rect 3881 12591 3939 12597
rect 5077 12597 5089 12600
rect 5123 12597 5135 12631
rect 5350 12628 5356 12640
rect 5311 12600 5356 12628
rect 5077 12591 5135 12597
rect 5350 12588 5356 12600
rect 5408 12588 5414 12640
rect 6914 12588 6920 12640
rect 6972 12628 6978 12640
rect 7374 12628 7380 12640
rect 6972 12600 7380 12628
rect 6972 12588 6978 12600
rect 7374 12588 7380 12600
rect 7432 12628 7438 12640
rect 11054 12628 11060 12640
rect 7432 12600 11060 12628
rect 7432 12588 7438 12600
rect 11054 12588 11060 12600
rect 11112 12588 11118 12640
rect 11164 12628 11192 12668
rect 11238 12656 11244 12708
rect 11296 12696 11302 12708
rect 11296 12668 11652 12696
rect 11296 12656 11302 12668
rect 11517 12631 11575 12637
rect 11517 12628 11529 12631
rect 11164 12600 11529 12628
rect 11517 12597 11529 12600
rect 11563 12597 11575 12631
rect 11624 12628 11652 12668
rect 11698 12656 11704 12708
rect 11756 12696 11762 12708
rect 11882 12696 11888 12708
rect 11756 12668 11888 12696
rect 11756 12656 11762 12668
rect 11882 12656 11888 12668
rect 11940 12656 11946 12708
rect 13262 12656 13268 12708
rect 13320 12696 13326 12708
rect 13449 12699 13507 12705
rect 13449 12696 13461 12699
rect 13320 12668 13461 12696
rect 13320 12656 13326 12668
rect 13449 12665 13461 12668
rect 13495 12665 13507 12699
rect 15286 12696 15292 12708
rect 13449 12659 13507 12665
rect 14844 12668 15292 12696
rect 13081 12631 13139 12637
rect 13081 12628 13093 12631
rect 11624 12600 13093 12628
rect 11517 12591 11575 12597
rect 13081 12597 13093 12600
rect 13127 12597 13139 12631
rect 13081 12591 13139 12597
rect 13538 12588 13544 12640
rect 13596 12628 13602 12640
rect 14844 12628 14872 12668
rect 15286 12656 15292 12668
rect 15344 12656 15350 12708
rect 13596 12600 14872 12628
rect 14921 12631 14979 12637
rect 13596 12588 13602 12600
rect 14921 12597 14933 12631
rect 14967 12628 14979 12631
rect 15102 12628 15108 12640
rect 14967 12600 15108 12628
rect 14967 12597 14979 12600
rect 14921 12591 14979 12597
rect 15102 12588 15108 12600
rect 15160 12588 15166 12640
rect 16022 12588 16028 12640
rect 16080 12628 16086 12640
rect 17034 12628 17040 12640
rect 16080 12600 17040 12628
rect 16080 12588 16086 12600
rect 17034 12588 17040 12600
rect 17092 12628 17098 12640
rect 18049 12631 18107 12637
rect 18049 12628 18061 12631
rect 17092 12600 18061 12628
rect 17092 12588 17098 12600
rect 18049 12597 18061 12600
rect 18095 12597 18107 12631
rect 18049 12591 18107 12597
rect 1104 12538 18860 12560
rect 1104 12486 3174 12538
rect 3226 12486 3238 12538
rect 3290 12486 3302 12538
rect 3354 12486 3366 12538
rect 3418 12486 3430 12538
rect 3482 12486 7622 12538
rect 7674 12486 7686 12538
rect 7738 12486 7750 12538
rect 7802 12486 7814 12538
rect 7866 12486 7878 12538
rect 7930 12486 12070 12538
rect 12122 12486 12134 12538
rect 12186 12486 12198 12538
rect 12250 12486 12262 12538
rect 12314 12486 12326 12538
rect 12378 12486 16518 12538
rect 16570 12486 16582 12538
rect 16634 12486 16646 12538
rect 16698 12486 16710 12538
rect 16762 12486 16774 12538
rect 16826 12486 18860 12538
rect 1104 12464 18860 12486
rect 3326 12424 3332 12436
rect 2884 12396 3332 12424
rect 2884 12297 2912 12396
rect 3326 12384 3332 12396
rect 3384 12384 3390 12436
rect 3421 12427 3479 12433
rect 3421 12393 3433 12427
rect 3467 12424 3479 12427
rect 3510 12424 3516 12436
rect 3467 12396 3516 12424
rect 3467 12393 3479 12396
rect 3421 12387 3479 12393
rect 3510 12384 3516 12396
rect 3568 12384 3574 12436
rect 3605 12427 3663 12433
rect 3605 12393 3617 12427
rect 3651 12424 3663 12427
rect 4062 12424 4068 12436
rect 3651 12396 4068 12424
rect 3651 12393 3663 12396
rect 3605 12387 3663 12393
rect 4062 12384 4068 12396
rect 4120 12384 4126 12436
rect 4430 12384 4436 12436
rect 4488 12424 4494 12436
rect 4525 12427 4583 12433
rect 4525 12424 4537 12427
rect 4488 12396 4537 12424
rect 4488 12384 4494 12396
rect 4525 12393 4537 12396
rect 4571 12393 4583 12427
rect 4525 12387 4583 12393
rect 4617 12427 4675 12433
rect 4617 12393 4629 12427
rect 4663 12424 4675 12427
rect 4706 12424 4712 12436
rect 4663 12396 4712 12424
rect 4663 12393 4675 12396
rect 4617 12387 4675 12393
rect 4706 12384 4712 12396
rect 4764 12384 4770 12436
rect 4798 12384 4804 12436
rect 4856 12424 4862 12436
rect 4856 12396 5488 12424
rect 4856 12384 4862 12396
rect 5350 12356 5356 12368
rect 3896 12328 5356 12356
rect 2869 12291 2927 12297
rect 2869 12257 2881 12291
rect 2915 12257 2927 12291
rect 3896 12288 3924 12328
rect 5350 12316 5356 12328
rect 5408 12316 5414 12368
rect 2869 12251 2927 12257
rect 3252 12260 3924 12288
rect 1949 12223 2007 12229
rect 1949 12189 1961 12223
rect 1995 12189 2007 12223
rect 1949 12183 2007 12189
rect 2225 12223 2283 12229
rect 2225 12189 2237 12223
rect 2271 12220 2283 12223
rect 2774 12220 2780 12232
rect 2271 12192 2780 12220
rect 2271 12189 2283 12192
rect 2225 12183 2283 12189
rect 1964 12152 1992 12183
rect 2774 12180 2780 12192
rect 2832 12180 2838 12232
rect 3142 12220 3148 12232
rect 3068 12192 3148 12220
rect 2406 12152 2412 12164
rect 1964 12124 2412 12152
rect 2406 12112 2412 12124
rect 2464 12112 2470 12164
rect 3068 12152 3096 12192
rect 3142 12180 3148 12192
rect 3200 12180 3206 12232
rect 3252 12229 3280 12260
rect 3970 12248 3976 12300
rect 4028 12288 4034 12300
rect 4028 12260 4073 12288
rect 4028 12248 4034 12260
rect 4246 12248 4252 12300
rect 4304 12288 4310 12300
rect 5261 12291 5319 12297
rect 4304 12260 5120 12288
rect 4304 12248 4310 12260
rect 3237 12223 3295 12229
rect 3237 12189 3249 12223
rect 3283 12189 3295 12223
rect 3237 12183 3295 12189
rect 3326 12180 3332 12232
rect 3384 12220 3390 12232
rect 4157 12223 4215 12229
rect 4157 12220 4169 12223
rect 3384 12192 4169 12220
rect 3384 12180 3390 12192
rect 4157 12189 4169 12192
rect 4203 12220 4215 12223
rect 4798 12220 4804 12232
rect 4203 12192 4804 12220
rect 4203 12189 4215 12192
rect 4157 12183 4215 12189
rect 4798 12180 4804 12192
rect 4856 12180 4862 12232
rect 4982 12220 4988 12232
rect 4943 12192 4988 12220
rect 4982 12180 4988 12192
rect 5040 12180 5046 12232
rect 5092 12220 5120 12260
rect 5261 12257 5273 12291
rect 5307 12288 5319 12291
rect 5460 12288 5488 12396
rect 8570 12384 8576 12436
rect 8628 12424 8634 12436
rect 13446 12424 13452 12436
rect 8628 12396 13308 12424
rect 13407 12396 13452 12424
rect 8628 12384 8634 12396
rect 5537 12359 5595 12365
rect 5537 12325 5549 12359
rect 5583 12356 5595 12359
rect 5994 12356 6000 12368
rect 5583 12328 6000 12356
rect 5583 12325 5595 12328
rect 5537 12319 5595 12325
rect 5994 12316 6000 12328
rect 6052 12316 6058 12368
rect 8386 12316 8392 12368
rect 8444 12356 8450 12368
rect 10045 12359 10103 12365
rect 10045 12356 10057 12359
rect 8444 12328 10057 12356
rect 8444 12316 8450 12328
rect 10045 12325 10057 12328
rect 10091 12325 10103 12359
rect 13280 12356 13308 12396
rect 13446 12384 13452 12396
rect 13504 12384 13510 12436
rect 14090 12424 14096 12436
rect 14051 12396 14096 12424
rect 14090 12384 14096 12396
rect 14148 12384 14154 12436
rect 14734 12384 14740 12436
rect 14792 12424 14798 12436
rect 15749 12427 15807 12433
rect 15749 12424 15761 12427
rect 14792 12396 15761 12424
rect 14792 12384 14798 12396
rect 15749 12393 15761 12396
rect 15795 12393 15807 12427
rect 18046 12424 18052 12436
rect 15749 12387 15807 12393
rect 16132 12396 18052 12424
rect 13817 12359 13875 12365
rect 13817 12356 13829 12359
rect 13280 12328 13829 12356
rect 10045 12319 10103 12325
rect 13817 12325 13829 12328
rect 13863 12325 13875 12359
rect 13817 12319 13875 12325
rect 8202 12288 8208 12300
rect 5307 12260 8208 12288
rect 5307 12257 5319 12260
rect 5261 12251 5319 12257
rect 8202 12248 8208 12260
rect 8260 12248 8266 12300
rect 5997 12223 6055 12229
rect 5997 12220 6009 12223
rect 5092 12192 6009 12220
rect 5997 12189 6009 12192
rect 6043 12189 6055 12223
rect 5997 12183 6055 12189
rect 6086 12180 6092 12232
rect 6144 12220 6150 12232
rect 9214 12220 9220 12232
rect 6144 12192 9220 12220
rect 6144 12180 6150 12192
rect 9214 12180 9220 12192
rect 9272 12180 9278 12232
rect 10069 12220 10097 12319
rect 11422 12288 11428 12300
rect 11383 12260 11428 12288
rect 11422 12248 11428 12260
rect 11480 12288 11486 12300
rect 11517 12291 11575 12297
rect 11517 12288 11529 12291
rect 11480 12260 11529 12288
rect 11480 12248 11486 12260
rect 11517 12257 11529 12260
rect 11563 12257 11575 12291
rect 11517 12251 11575 12257
rect 10686 12220 10692 12232
rect 10069 12192 10692 12220
rect 10686 12180 10692 12192
rect 10744 12180 10750 12232
rect 11330 12220 11336 12232
rect 11072 12192 11336 12220
rect 5813 12155 5871 12161
rect 5813 12152 5825 12155
rect 3068 12124 5825 12152
rect 5813 12121 5825 12124
rect 5859 12121 5871 12155
rect 5813 12115 5871 12121
rect 5902 12112 5908 12164
rect 5960 12152 5966 12164
rect 11072 12152 11100 12192
rect 11330 12180 11336 12192
rect 11388 12180 11394 12232
rect 11790 12229 11796 12232
rect 11784 12183 11796 12229
rect 11848 12220 11854 12232
rect 11848 12192 11884 12220
rect 11790 12180 11796 12183
rect 11848 12180 11854 12192
rect 12066 12180 12072 12232
rect 12124 12220 12130 12232
rect 13832 12220 13860 12319
rect 16132 12288 16160 12396
rect 18046 12384 18052 12396
rect 18104 12384 18110 12436
rect 17310 12316 17316 12368
rect 17368 12356 17374 12368
rect 17586 12356 17592 12368
rect 17368 12328 17592 12356
rect 17368 12316 17374 12328
rect 17586 12316 17592 12328
rect 17644 12316 17650 12368
rect 17126 12288 17132 12300
rect 15396 12260 16160 12288
rect 17087 12260 17132 12288
rect 15206 12223 15264 12229
rect 15206 12220 15218 12223
rect 12124 12192 13676 12220
rect 13832 12192 15218 12220
rect 12124 12180 12130 12192
rect 5960 12124 11100 12152
rect 11180 12155 11238 12161
rect 5960 12112 5966 12124
rect 11180 12121 11192 12155
rect 11226 12152 11238 12155
rect 12802 12152 12808 12164
rect 11226 12124 12808 12152
rect 11226 12121 11238 12124
rect 11180 12115 11238 12121
rect 12802 12112 12808 12124
rect 12860 12112 12866 12164
rect 13541 12155 13599 12161
rect 13541 12152 13553 12155
rect 12912 12124 13553 12152
rect 12912 12096 12940 12124
rect 13541 12121 13553 12124
rect 13587 12121 13599 12155
rect 13541 12115 13599 12121
rect 1854 12044 1860 12096
rect 1912 12084 1918 12096
rect 3878 12084 3884 12096
rect 1912 12056 3884 12084
rect 1912 12044 1918 12056
rect 3878 12044 3884 12056
rect 3936 12044 3942 12096
rect 4065 12087 4123 12093
rect 4065 12053 4077 12087
rect 4111 12084 4123 12087
rect 4154 12084 4160 12096
rect 4111 12056 4160 12084
rect 4111 12053 4123 12056
rect 4065 12047 4123 12053
rect 4154 12044 4160 12056
rect 4212 12044 4218 12096
rect 4798 12044 4804 12096
rect 4856 12084 4862 12096
rect 5077 12087 5135 12093
rect 5077 12084 5089 12087
rect 4856 12056 5089 12084
rect 4856 12044 4862 12056
rect 5077 12053 5089 12056
rect 5123 12053 5135 12087
rect 5077 12047 5135 12053
rect 5166 12044 5172 12096
rect 5224 12084 5230 12096
rect 5626 12084 5632 12096
rect 5224 12056 5632 12084
rect 5224 12044 5230 12056
rect 5626 12044 5632 12056
rect 5684 12044 5690 12096
rect 5718 12044 5724 12096
rect 5776 12084 5782 12096
rect 12894 12084 12900 12096
rect 5776 12056 12900 12084
rect 5776 12044 5782 12056
rect 12894 12044 12900 12056
rect 12952 12044 12958 12096
rect 13078 12084 13084 12096
rect 13039 12056 13084 12084
rect 13078 12044 13084 12056
rect 13136 12044 13142 12096
rect 13265 12087 13323 12093
rect 13265 12053 13277 12087
rect 13311 12084 13323 12087
rect 13648 12084 13676 12192
rect 15206 12189 15218 12192
rect 15252 12189 15264 12223
rect 15396 12220 15424 12260
rect 17126 12248 17132 12260
rect 17184 12248 17190 12300
rect 17957 12291 18015 12297
rect 17236 12260 17816 12288
rect 15206 12183 15264 12189
rect 15304 12192 15424 12220
rect 14090 12112 14096 12164
rect 14148 12152 14154 12164
rect 14550 12152 14556 12164
rect 14148 12124 14556 12152
rect 14148 12112 14154 12124
rect 14550 12112 14556 12124
rect 14608 12112 14614 12164
rect 14642 12112 14648 12164
rect 14700 12152 14706 12164
rect 15304 12152 15332 12192
rect 15470 12180 15476 12232
rect 15528 12220 15534 12232
rect 17236 12220 17264 12260
rect 17678 12220 17684 12232
rect 15528 12192 15573 12220
rect 16684 12192 17264 12220
rect 17639 12192 17684 12220
rect 15528 12180 15534 12192
rect 16684 12152 16712 12192
rect 17678 12180 17684 12192
rect 17736 12180 17742 12232
rect 17788 12220 17816 12260
rect 17957 12257 17969 12291
rect 18003 12288 18015 12291
rect 18138 12288 18144 12300
rect 18003 12260 18144 12288
rect 18003 12257 18015 12260
rect 17957 12251 18015 12257
rect 18138 12248 18144 12260
rect 18196 12248 18202 12300
rect 18230 12220 18236 12232
rect 17788 12192 18236 12220
rect 18230 12180 18236 12192
rect 18288 12180 18294 12232
rect 14700 12124 15332 12152
rect 15396 12124 16712 12152
rect 14700 12112 14706 12124
rect 14182 12084 14188 12096
rect 13311 12056 14188 12084
rect 13311 12053 13323 12056
rect 13265 12047 13323 12053
rect 14182 12044 14188 12056
rect 14240 12044 14246 12096
rect 14734 12044 14740 12096
rect 14792 12084 14798 12096
rect 15396 12084 15424 12124
rect 16758 12112 16764 12164
rect 16816 12152 16822 12164
rect 16862 12155 16920 12161
rect 16862 12152 16874 12155
rect 16816 12124 16874 12152
rect 16816 12112 16822 12124
rect 16862 12121 16874 12124
rect 16908 12121 16920 12155
rect 17497 12155 17555 12161
rect 17497 12152 17509 12155
rect 16862 12115 16920 12121
rect 17052 12124 17509 12152
rect 14792 12056 15424 12084
rect 14792 12044 14798 12056
rect 15470 12044 15476 12096
rect 15528 12084 15534 12096
rect 17052 12084 17080 12124
rect 17497 12121 17509 12124
rect 17543 12152 17555 12155
rect 17586 12152 17592 12164
rect 17543 12124 17592 12152
rect 17543 12121 17555 12124
rect 17497 12115 17555 12121
rect 17586 12112 17592 12124
rect 17644 12112 17650 12164
rect 15528 12056 17080 12084
rect 15528 12044 15534 12056
rect 17126 12044 17132 12096
rect 17184 12084 17190 12096
rect 17405 12087 17463 12093
rect 17405 12084 17417 12087
rect 17184 12056 17417 12084
rect 17184 12044 17190 12056
rect 17405 12053 17417 12056
rect 17451 12053 17463 12087
rect 17405 12047 17463 12053
rect 1104 11994 18860 12016
rect 1104 11942 5398 11994
rect 5450 11942 5462 11994
rect 5514 11942 5526 11994
rect 5578 11942 5590 11994
rect 5642 11942 5654 11994
rect 5706 11942 9846 11994
rect 9898 11942 9910 11994
rect 9962 11942 9974 11994
rect 10026 11942 10038 11994
rect 10090 11942 10102 11994
rect 10154 11942 14294 11994
rect 14346 11942 14358 11994
rect 14410 11942 14422 11994
rect 14474 11942 14486 11994
rect 14538 11942 14550 11994
rect 14602 11942 18860 11994
rect 1104 11920 18860 11942
rect 2958 11840 2964 11892
rect 3016 11880 3022 11892
rect 3053 11883 3111 11889
rect 3053 11880 3065 11883
rect 3016 11852 3065 11880
rect 3016 11840 3022 11852
rect 3053 11849 3065 11852
rect 3099 11849 3111 11883
rect 3053 11843 3111 11849
rect 3329 11883 3387 11889
rect 3329 11849 3341 11883
rect 3375 11880 3387 11883
rect 3602 11880 3608 11892
rect 3375 11852 3608 11880
rect 3375 11849 3387 11852
rect 3329 11843 3387 11849
rect 3602 11840 3608 11852
rect 3660 11840 3666 11892
rect 3970 11840 3976 11892
rect 4028 11880 4034 11892
rect 5626 11880 5632 11892
rect 4028 11852 5396 11880
rect 5539 11852 5632 11880
rect 4028 11840 4034 11852
rect 4154 11812 4160 11824
rect 4115 11784 4160 11812
rect 4154 11772 4160 11784
rect 4212 11772 4218 11824
rect 2038 11704 2044 11756
rect 2096 11744 2102 11756
rect 2593 11747 2651 11753
rect 2593 11744 2605 11747
rect 2096 11716 2605 11744
rect 2096 11704 2102 11716
rect 2593 11713 2605 11716
rect 2639 11713 2651 11747
rect 2593 11707 2651 11713
rect 2685 11747 2743 11753
rect 2685 11713 2697 11747
rect 2731 11744 2743 11747
rect 2958 11744 2964 11756
rect 2731 11716 2964 11744
rect 2731 11713 2743 11716
rect 2685 11707 2743 11713
rect 2958 11704 2964 11716
rect 3016 11704 3022 11756
rect 3145 11747 3203 11753
rect 3145 11713 3157 11747
rect 3191 11744 3203 11747
rect 4062 11744 4068 11756
rect 3191 11716 4068 11744
rect 3191 11713 3203 11716
rect 3145 11707 3203 11713
rect 4062 11704 4068 11716
rect 4120 11704 4126 11756
rect 4249 11747 4307 11753
rect 4249 11740 4261 11747
rect 4295 11740 4307 11747
rect 5074 11744 5080 11756
rect 4246 11688 4252 11740
rect 4304 11688 4310 11740
rect 5035 11716 5080 11744
rect 5074 11704 5080 11716
rect 5132 11704 5138 11756
rect 1946 11676 1952 11688
rect 1907 11648 1952 11676
rect 1946 11636 1952 11648
rect 2004 11636 2010 11688
rect 2222 11676 2228 11688
rect 2183 11648 2228 11676
rect 2222 11636 2228 11648
rect 2280 11636 2286 11688
rect 2498 11676 2504 11688
rect 2459 11648 2504 11676
rect 2498 11636 2504 11648
rect 2556 11636 2562 11688
rect 3602 11676 3608 11688
rect 3563 11648 3608 11676
rect 3602 11636 3608 11648
rect 3660 11636 3666 11688
rect 3970 11676 3976 11688
rect 3931 11648 3976 11676
rect 3970 11636 3976 11648
rect 4028 11636 4034 11688
rect 5166 11676 5172 11688
rect 5127 11648 5172 11676
rect 5166 11636 5172 11648
rect 5224 11636 5230 11688
rect 5368 11685 5396 11852
rect 5626 11840 5632 11852
rect 5684 11880 5690 11892
rect 6086 11880 6092 11892
rect 5684 11852 6092 11880
rect 5684 11840 5690 11852
rect 6086 11840 6092 11852
rect 6144 11840 6150 11892
rect 8294 11880 8300 11892
rect 6932 11852 8300 11880
rect 5810 11744 5816 11756
rect 5771 11716 5816 11744
rect 5810 11704 5816 11716
rect 5868 11704 5874 11756
rect 5353 11679 5411 11685
rect 5353 11645 5365 11679
rect 5399 11676 5411 11679
rect 6932 11676 6960 11852
rect 8294 11840 8300 11852
rect 8352 11840 8358 11892
rect 8570 11880 8576 11892
rect 8531 11852 8576 11880
rect 8570 11840 8576 11852
rect 8628 11840 8634 11892
rect 9674 11840 9680 11892
rect 9732 11880 9738 11892
rect 10045 11883 10103 11889
rect 10045 11880 10057 11883
rect 9732 11852 10057 11880
rect 9732 11840 9738 11852
rect 10045 11849 10057 11852
rect 10091 11849 10103 11883
rect 10045 11843 10103 11849
rect 13541 11883 13599 11889
rect 13541 11849 13553 11883
rect 13587 11880 13599 11883
rect 13814 11880 13820 11892
rect 13587 11852 13820 11880
rect 13587 11849 13599 11852
rect 13541 11843 13599 11849
rect 13814 11840 13820 11852
rect 13872 11840 13878 11892
rect 15746 11840 15752 11892
rect 15804 11880 15810 11892
rect 15804 11852 18460 11880
rect 15804 11840 15810 11852
rect 18432 11824 18460 11852
rect 8110 11812 8116 11824
rect 7208 11784 8116 11812
rect 7208 11756 7236 11784
rect 8110 11772 8116 11784
rect 8168 11772 8174 11824
rect 8202 11772 8208 11824
rect 8260 11812 8266 11824
rect 8910 11815 8968 11821
rect 8910 11812 8922 11815
rect 8260 11784 8922 11812
rect 8260 11772 8266 11784
rect 8910 11781 8922 11784
rect 8956 11781 8968 11815
rect 8910 11775 8968 11781
rect 12986 11772 12992 11824
rect 13044 11812 13050 11824
rect 15378 11812 15384 11824
rect 13044 11784 15384 11812
rect 13044 11772 13050 11784
rect 7190 11744 7196 11756
rect 7151 11716 7196 11744
rect 7190 11704 7196 11716
rect 7248 11704 7254 11756
rect 7449 11747 7507 11753
rect 7449 11744 7461 11747
rect 7300 11716 7461 11744
rect 7300 11676 7328 11716
rect 7449 11713 7461 11716
rect 7495 11713 7507 11747
rect 8128 11744 8156 11772
rect 8665 11747 8723 11753
rect 8665 11744 8677 11747
rect 8128 11716 8677 11744
rect 7449 11707 7507 11713
rect 8665 11713 8677 11716
rect 8711 11713 8723 11747
rect 8665 11707 8723 11713
rect 9214 11704 9220 11756
rect 9272 11744 9278 11756
rect 12066 11744 12072 11756
rect 9272 11716 12072 11744
rect 9272 11704 9278 11716
rect 12066 11704 12072 11716
rect 12124 11704 12130 11756
rect 12894 11704 12900 11756
rect 12952 11744 12958 11756
rect 13464 11753 13492 11784
rect 13182 11747 13240 11753
rect 13182 11744 13194 11747
rect 12952 11716 13194 11744
rect 12952 11704 12958 11716
rect 13182 11713 13194 11716
rect 13228 11713 13240 11747
rect 13182 11707 13240 11713
rect 13449 11747 13507 11753
rect 13449 11713 13461 11747
rect 13495 11713 13507 11747
rect 14642 11744 14648 11756
rect 14700 11753 14706 11756
rect 14936 11753 14964 11784
rect 15378 11772 15384 11784
rect 15436 11812 15442 11824
rect 18230 11812 18236 11824
rect 15436 11784 18092 11812
rect 18191 11784 18236 11812
rect 15436 11772 15442 11784
rect 14612 11716 14648 11744
rect 13449 11707 13507 11713
rect 14642 11704 14648 11716
rect 14700 11707 14712 11753
rect 14921 11747 14979 11753
rect 14921 11713 14933 11747
rect 14967 11713 14979 11747
rect 16114 11744 16120 11756
rect 16172 11753 16178 11756
rect 16408 11753 16436 11784
rect 16084 11716 16120 11744
rect 14921 11707 14979 11713
rect 14700 11704 14706 11707
rect 16114 11704 16120 11716
rect 16172 11707 16184 11753
rect 16393 11747 16451 11753
rect 16393 11713 16405 11747
rect 16439 11713 16451 11747
rect 16393 11707 16451 11713
rect 16172 11704 16178 11707
rect 16942 11704 16948 11756
rect 17000 11744 17006 11756
rect 17310 11744 17316 11756
rect 17000 11716 17316 11744
rect 17000 11704 17006 11716
rect 17310 11704 17316 11716
rect 17368 11704 17374 11756
rect 17770 11704 17776 11756
rect 17828 11753 17834 11756
rect 18064 11753 18092 11784
rect 18230 11772 18236 11784
rect 18288 11772 18294 11824
rect 18414 11812 18420 11824
rect 18327 11784 18420 11812
rect 18414 11772 18420 11784
rect 18472 11772 18478 11824
rect 17828 11747 17851 11753
rect 17839 11713 17851 11747
rect 17828 11707 17851 11713
rect 18049 11747 18107 11753
rect 18049 11713 18061 11747
rect 18095 11713 18107 11747
rect 18049 11707 18107 11713
rect 17828 11704 17834 11707
rect 5399 11648 6960 11676
rect 7208 11648 7328 11676
rect 5399 11645 5411 11648
rect 5353 11639 5411 11645
rect 5902 11608 5908 11620
rect 5863 11580 5908 11608
rect 5902 11568 5908 11580
rect 5960 11568 5966 11620
rect 5994 11568 6000 11620
rect 6052 11608 6058 11620
rect 7208 11608 7236 11648
rect 13538 11636 13544 11688
rect 13596 11676 13602 11688
rect 13722 11676 13728 11688
rect 13596 11648 13728 11676
rect 13596 11636 13602 11648
rect 13722 11636 13728 11648
rect 13780 11636 13786 11688
rect 11885 11611 11943 11617
rect 6052 11580 7236 11608
rect 6052 11568 6058 11580
rect 2406 11500 2412 11552
rect 2464 11540 2470 11552
rect 3513 11543 3571 11549
rect 3513 11540 3525 11543
rect 2464 11512 3525 11540
rect 2464 11500 2470 11512
rect 3513 11509 3525 11512
rect 3559 11540 3571 11543
rect 4246 11540 4252 11552
rect 3559 11512 4252 11540
rect 3559 11509 3571 11512
rect 3513 11503 3571 11509
rect 4246 11500 4252 11512
rect 4304 11500 4310 11552
rect 4338 11500 4344 11552
rect 4396 11540 4402 11552
rect 4617 11543 4675 11549
rect 4617 11540 4629 11543
rect 4396 11512 4629 11540
rect 4396 11500 4402 11512
rect 4617 11509 4629 11512
rect 4663 11509 4675 11543
rect 4617 11503 4675 11509
rect 4709 11543 4767 11549
rect 4709 11509 4721 11543
rect 4755 11540 4767 11543
rect 4798 11540 4804 11552
rect 4755 11512 4804 11540
rect 4755 11509 4767 11512
rect 4709 11503 4767 11509
rect 4798 11500 4804 11512
rect 4856 11500 4862 11552
rect 7208 11540 7236 11580
rect 9600 11580 11744 11608
rect 9600 11540 9628 11580
rect 11606 11540 11612 11552
rect 7208 11512 9628 11540
rect 11567 11512 11612 11540
rect 11606 11500 11612 11512
rect 11664 11500 11670 11552
rect 11716 11540 11744 11580
rect 11885 11577 11897 11611
rect 11931 11608 11943 11611
rect 11931 11580 12434 11608
rect 11931 11577 11943 11580
rect 11885 11571 11943 11577
rect 12069 11543 12127 11549
rect 12069 11540 12081 11543
rect 11716 11512 12081 11540
rect 12069 11509 12081 11512
rect 12115 11509 12127 11543
rect 12406 11540 12434 11580
rect 14936 11580 15240 11608
rect 14936 11540 14964 11580
rect 12406 11512 14964 11540
rect 15013 11543 15071 11549
rect 12069 11503 12127 11509
rect 15013 11509 15025 11543
rect 15059 11540 15071 11543
rect 15102 11540 15108 11552
rect 15059 11512 15108 11540
rect 15059 11509 15071 11512
rect 15013 11503 15071 11509
rect 15102 11500 15108 11512
rect 15160 11500 15166 11552
rect 15212 11540 15240 11580
rect 16500 11580 16804 11608
rect 16500 11540 16528 11580
rect 15212 11512 16528 11540
rect 16574 11500 16580 11552
rect 16632 11540 16638 11552
rect 16669 11543 16727 11549
rect 16669 11540 16681 11543
rect 16632 11512 16681 11540
rect 16632 11500 16638 11512
rect 16669 11509 16681 11512
rect 16715 11509 16727 11543
rect 16776 11540 16804 11580
rect 17678 11540 17684 11552
rect 16776 11512 17684 11540
rect 16669 11503 16727 11509
rect 17678 11500 17684 11512
rect 17736 11500 17742 11552
rect 1104 11450 18860 11472
rect 1104 11398 3174 11450
rect 3226 11398 3238 11450
rect 3290 11398 3302 11450
rect 3354 11398 3366 11450
rect 3418 11398 3430 11450
rect 3482 11398 7622 11450
rect 7674 11398 7686 11450
rect 7738 11398 7750 11450
rect 7802 11398 7814 11450
rect 7866 11398 7878 11450
rect 7930 11398 12070 11450
rect 12122 11398 12134 11450
rect 12186 11398 12198 11450
rect 12250 11398 12262 11450
rect 12314 11398 12326 11450
rect 12378 11398 16518 11450
rect 16570 11398 16582 11450
rect 16634 11398 16646 11450
rect 16698 11398 16710 11450
rect 16762 11398 16774 11450
rect 16826 11398 18860 11450
rect 1104 11376 18860 11398
rect 2866 11336 2872 11348
rect 2827 11308 2872 11336
rect 2866 11296 2872 11308
rect 2924 11296 2930 11348
rect 6181 11339 6239 11345
rect 6181 11336 6193 11339
rect 3344 11308 6193 11336
rect 2222 11228 2228 11280
rect 2280 11268 2286 11280
rect 2590 11268 2596 11280
rect 2280 11240 2452 11268
rect 2551 11240 2596 11268
rect 2280 11228 2286 11240
rect 1949 11203 2007 11209
rect 1949 11169 1961 11203
rect 1995 11200 2007 11203
rect 2424 11200 2452 11240
rect 2590 11228 2596 11240
rect 2648 11228 2654 11280
rect 2774 11228 2780 11280
rect 2832 11268 2838 11280
rect 2958 11268 2964 11280
rect 2832 11240 2964 11268
rect 2832 11228 2838 11240
rect 2958 11228 2964 11240
rect 3016 11228 3022 11280
rect 3344 11200 3372 11308
rect 6181 11305 6193 11308
rect 6227 11305 6239 11339
rect 6181 11299 6239 11305
rect 7190 11296 7196 11348
rect 7248 11336 7254 11348
rect 7374 11336 7380 11348
rect 7248 11308 7380 11336
rect 7248 11296 7254 11308
rect 7374 11296 7380 11308
rect 7432 11296 7438 11348
rect 8110 11296 8116 11348
rect 8168 11336 8174 11348
rect 10873 11339 10931 11345
rect 8168 11308 10364 11336
rect 8168 11296 8174 11308
rect 4801 11271 4859 11277
rect 4801 11237 4813 11271
rect 4847 11268 4859 11271
rect 8938 11268 8944 11280
rect 4847 11240 5764 11268
rect 8899 11240 8944 11268
rect 4847 11237 4859 11240
rect 4801 11231 4859 11237
rect 1995 11172 2360 11200
rect 2424 11172 3372 11200
rect 3513 11203 3571 11209
rect 1995 11169 2007 11172
rect 1949 11163 2007 11169
rect 2222 11132 2228 11144
rect 2183 11104 2228 11132
rect 2222 11092 2228 11104
rect 2280 11092 2286 11144
rect 2332 11132 2360 11172
rect 3513 11169 3525 11203
rect 3559 11200 3571 11203
rect 3878 11200 3884 11212
rect 3559 11172 3884 11200
rect 3559 11169 3571 11172
rect 3513 11163 3571 11169
rect 3878 11160 3884 11172
rect 3936 11200 3942 11212
rect 4062 11200 4068 11212
rect 3936 11172 4068 11200
rect 3936 11160 3942 11172
rect 4062 11160 4068 11172
rect 4120 11160 4126 11212
rect 4154 11160 4160 11212
rect 4212 11200 4218 11212
rect 4249 11203 4307 11209
rect 4249 11200 4261 11203
rect 4212 11172 4261 11200
rect 4212 11160 4218 11172
rect 4249 11169 4261 11172
rect 4295 11169 4307 11203
rect 4249 11163 4307 11169
rect 5537 11203 5595 11209
rect 5537 11169 5549 11203
rect 5583 11169 5595 11203
rect 5537 11163 5595 11169
rect 3142 11132 3148 11144
rect 2332 11104 3148 11132
rect 3142 11092 3148 11104
rect 3200 11092 3206 11144
rect 3237 11135 3295 11141
rect 3237 11101 3249 11135
rect 3283 11132 3295 11135
rect 3602 11132 3608 11144
rect 3283 11104 3608 11132
rect 3283 11101 3295 11104
rect 3237 11095 3295 11101
rect 3602 11092 3608 11104
rect 3660 11092 3666 11144
rect 4338 11132 4344 11144
rect 4299 11104 4344 11132
rect 4338 11092 4344 11104
rect 4396 11092 4402 11144
rect 2409 11067 2467 11073
rect 2409 11033 2421 11067
rect 2455 11064 2467 11067
rect 2866 11064 2872 11076
rect 2455 11036 2872 11064
rect 2455 11033 2467 11036
rect 2409 11027 2467 11033
rect 2866 11024 2872 11036
rect 2924 11064 2930 11076
rect 5077 11067 5135 11073
rect 5077 11064 5089 11067
rect 2924 11036 5089 11064
rect 2924 11024 2930 11036
rect 5077 11033 5089 11036
rect 5123 11033 5135 11067
rect 5552 11064 5580 11163
rect 5736 11141 5764 11240
rect 8938 11228 8944 11240
rect 8996 11228 9002 11280
rect 10336 11268 10364 11308
rect 10873 11305 10885 11339
rect 10919 11336 10931 11339
rect 11146 11336 11152 11348
rect 10919 11308 11152 11336
rect 10919 11305 10931 11308
rect 10873 11299 10931 11305
rect 11146 11296 11152 11308
rect 11204 11296 11210 11348
rect 11974 11336 11980 11348
rect 11256 11308 11980 11336
rect 11256 11268 11284 11308
rect 11974 11296 11980 11308
rect 12032 11296 12038 11348
rect 12066 11296 12072 11348
rect 12124 11336 12130 11348
rect 13998 11336 14004 11348
rect 12124 11308 14004 11336
rect 12124 11296 12130 11308
rect 13998 11296 14004 11308
rect 14056 11296 14062 11348
rect 14369 11339 14427 11345
rect 14369 11305 14381 11339
rect 14415 11336 14427 11339
rect 14415 11308 17356 11336
rect 14415 11305 14427 11308
rect 14369 11299 14427 11305
rect 10336 11240 11284 11268
rect 13722 11228 13728 11280
rect 13780 11268 13786 11280
rect 13906 11268 13912 11280
rect 13780 11240 13912 11268
rect 13780 11228 13786 11240
rect 13906 11228 13912 11240
rect 13964 11268 13970 11280
rect 14461 11271 14519 11277
rect 14461 11268 14473 11271
rect 13964 11240 14473 11268
rect 13964 11228 13970 11240
rect 14461 11237 14473 11240
rect 14507 11237 14519 11271
rect 14461 11231 14519 11237
rect 15933 11271 15991 11277
rect 15933 11237 15945 11271
rect 15979 11268 15991 11271
rect 16114 11268 16120 11280
rect 15979 11240 16120 11268
rect 15979 11237 15991 11240
rect 15933 11231 15991 11237
rect 16114 11228 16120 11240
rect 16172 11228 16178 11280
rect 6638 11160 6644 11212
rect 6696 11200 6702 11212
rect 9214 11200 9220 11212
rect 6696 11172 9220 11200
rect 6696 11160 6702 11172
rect 9214 11160 9220 11172
rect 9272 11160 9278 11212
rect 14734 11200 14740 11212
rect 13372 11172 14740 11200
rect 5721 11135 5779 11141
rect 5721 11101 5733 11135
rect 5767 11101 5779 11135
rect 5721 11095 5779 11101
rect 9674 11092 9680 11144
rect 9732 11132 9738 11144
rect 10321 11135 10379 11141
rect 10321 11132 10333 11135
rect 9732 11104 10333 11132
rect 9732 11092 9738 11104
rect 10321 11101 10333 11104
rect 10367 11101 10379 11135
rect 12253 11135 12311 11141
rect 12253 11132 12265 11135
rect 10321 11095 10379 11101
rect 11808 11104 12265 11132
rect 11808 11076 11836 11104
rect 12253 11101 12265 11104
rect 12299 11132 12311 11135
rect 12345 11135 12403 11141
rect 12345 11132 12357 11135
rect 12299 11104 12357 11132
rect 12299 11101 12311 11104
rect 12253 11095 12311 11101
rect 12345 11101 12357 11104
rect 12391 11101 12403 11135
rect 12345 11095 12403 11101
rect 13078 11092 13084 11144
rect 13136 11132 13142 11144
rect 13372 11132 13400 11172
rect 14734 11160 14740 11172
rect 14792 11160 14798 11212
rect 17328 11200 17356 11308
rect 17589 11271 17647 11277
rect 17589 11237 17601 11271
rect 17635 11268 17647 11271
rect 18230 11268 18236 11280
rect 17635 11240 18236 11268
rect 17635 11237 17647 11240
rect 17589 11231 17647 11237
rect 18230 11228 18236 11240
rect 18288 11228 18294 11280
rect 17328 11172 17724 11200
rect 17696 11144 17724 11172
rect 13136 11104 13400 11132
rect 13909 11135 13967 11141
rect 13136 11092 13142 11104
rect 13909 11101 13921 11135
rect 13955 11132 13967 11135
rect 15746 11132 15752 11144
rect 13955 11104 15752 11132
rect 13955 11101 13967 11104
rect 13909 11095 13967 11101
rect 15746 11092 15752 11104
rect 15804 11092 15810 11144
rect 15841 11135 15899 11141
rect 15841 11101 15853 11135
rect 15887 11132 15899 11135
rect 16206 11132 16212 11144
rect 15887 11104 16212 11132
rect 15887 11101 15899 11104
rect 15841 11095 15899 11101
rect 16206 11092 16212 11104
rect 16264 11132 16270 11144
rect 17313 11135 17371 11141
rect 17313 11132 17325 11135
rect 16264 11104 17325 11132
rect 16264 11092 16270 11104
rect 17313 11101 17325 11104
rect 17359 11101 17371 11135
rect 17313 11095 17371 11101
rect 17405 11135 17463 11141
rect 17405 11101 17417 11135
rect 17451 11101 17463 11135
rect 17678 11132 17684 11144
rect 17639 11104 17684 11132
rect 17405 11095 17463 11101
rect 9398 11064 9404 11076
rect 5552 11036 9404 11064
rect 5077 11027 5135 11033
rect 9398 11024 9404 11036
rect 9456 11024 9462 11076
rect 9582 11024 9588 11076
rect 9640 11064 9646 11076
rect 10054 11067 10112 11073
rect 10054 11064 10066 11067
rect 9640 11036 10066 11064
rect 9640 11024 9646 11036
rect 10054 11033 10066 11036
rect 10100 11064 10112 11067
rect 11422 11064 11428 11076
rect 10100 11036 11428 11064
rect 10100 11033 10112 11036
rect 10054 11027 10112 11033
rect 11422 11024 11428 11036
rect 11480 11024 11486 11076
rect 11790 11024 11796 11076
rect 11848 11024 11854 11076
rect 11974 11024 11980 11076
rect 12032 11073 12038 11076
rect 12032 11064 12044 11073
rect 12612 11067 12670 11073
rect 12032 11036 12077 11064
rect 12032 11027 12044 11036
rect 12612 11033 12624 11067
rect 12658 11064 12670 11067
rect 12710 11064 12716 11076
rect 12658 11036 12716 11064
rect 12658 11033 12670 11036
rect 12612 11027 12670 11033
rect 12032 11024 12038 11027
rect 12710 11024 12716 11036
rect 12768 11024 12774 11076
rect 13538 11024 13544 11076
rect 13596 11064 13602 11076
rect 14185 11067 14243 11073
rect 13596 11036 13768 11064
rect 13596 11024 13602 11036
rect 3050 10956 3056 11008
rect 3108 10996 3114 11008
rect 3329 10999 3387 11005
rect 3329 10996 3341 10999
rect 3108 10968 3341 10996
rect 3108 10956 3114 10968
rect 3329 10965 3341 10968
rect 3375 10965 3387 10999
rect 3878 10996 3884 11008
rect 3839 10968 3884 10996
rect 3329 10959 3387 10965
rect 3878 10956 3884 10968
rect 3936 10956 3942 11008
rect 4430 10996 4436 11008
rect 4391 10968 4436 10996
rect 4430 10956 4436 10968
rect 4488 10956 4494 11008
rect 4982 10996 4988 11008
rect 4943 10968 4988 10996
rect 4982 10956 4988 10968
rect 5040 10956 5046 11008
rect 5629 10999 5687 11005
rect 5629 10965 5641 10999
rect 5675 10996 5687 10999
rect 5810 10996 5816 11008
rect 5675 10968 5816 10996
rect 5675 10965 5687 10968
rect 5629 10959 5687 10965
rect 5810 10956 5816 10968
rect 5868 10956 5874 11008
rect 6086 10996 6092 11008
rect 6047 10968 6092 10996
rect 6086 10956 6092 10968
rect 6144 10956 6150 11008
rect 10410 10956 10416 11008
rect 10468 10996 10474 11008
rect 11698 10996 11704 11008
rect 10468 10968 11704 10996
rect 10468 10956 10474 10968
rect 11698 10956 11704 10968
rect 11756 10956 11762 11008
rect 13740 11005 13768 11036
rect 14185 11033 14197 11067
rect 14231 11064 14243 11067
rect 15470 11064 15476 11076
rect 14231 11036 15476 11064
rect 14231 11033 14243 11036
rect 14185 11027 14243 11033
rect 15470 11024 15476 11036
rect 15528 11024 15534 11076
rect 15562 11024 15568 11076
rect 15620 11073 15626 11076
rect 15620 11064 15632 11073
rect 15620 11036 15665 11064
rect 15620 11027 15632 11036
rect 15620 11024 15626 11027
rect 15930 11024 15936 11076
rect 15988 11064 15994 11076
rect 16390 11064 16396 11076
rect 15988 11036 16396 11064
rect 15988 11024 15994 11036
rect 16390 11024 16396 11036
rect 16448 11024 16454 11076
rect 16942 11024 16948 11076
rect 17000 11064 17006 11076
rect 17126 11073 17132 11076
rect 17068 11067 17132 11073
rect 17068 11064 17080 11067
rect 17000 11036 17080 11064
rect 17000 11024 17006 11036
rect 17068 11033 17080 11036
rect 17114 11033 17132 11067
rect 17068 11027 17132 11033
rect 17126 11024 17132 11027
rect 17184 11024 17190 11076
rect 13725 10999 13783 11005
rect 13725 10965 13737 10999
rect 13771 10965 13783 10999
rect 13725 10959 13783 10965
rect 15654 10956 15660 11008
rect 15712 10996 15718 11008
rect 17420 10996 17448 11095
rect 17678 11092 17684 11104
rect 17736 11092 17742 11144
rect 17957 11135 18015 11141
rect 17957 11101 17969 11135
rect 18003 11132 18015 11135
rect 18598 11132 18604 11144
rect 18003 11104 18604 11132
rect 18003 11101 18015 11104
rect 17957 11095 18015 11101
rect 18598 11092 18604 11104
rect 18656 11092 18662 11144
rect 18046 11024 18052 11076
rect 18104 11064 18110 11076
rect 18506 11064 18512 11076
rect 18104 11036 18512 11064
rect 18104 11024 18110 11036
rect 18506 11024 18512 11036
rect 18564 11024 18570 11076
rect 18966 10996 18972 11008
rect 15712 10968 18972 10996
rect 15712 10956 15718 10968
rect 18966 10956 18972 10968
rect 19024 10956 19030 11008
rect 1104 10906 18860 10928
rect 1104 10854 5398 10906
rect 5450 10854 5462 10906
rect 5514 10854 5526 10906
rect 5578 10854 5590 10906
rect 5642 10854 5654 10906
rect 5706 10854 9846 10906
rect 9898 10854 9910 10906
rect 9962 10854 9974 10906
rect 10026 10854 10038 10906
rect 10090 10854 10102 10906
rect 10154 10854 14294 10906
rect 14346 10854 14358 10906
rect 14410 10854 14422 10906
rect 14474 10854 14486 10906
rect 14538 10854 14550 10906
rect 14602 10854 18860 10906
rect 1104 10832 18860 10854
rect 3513 10795 3571 10801
rect 3513 10761 3525 10795
rect 3559 10792 3571 10795
rect 4430 10792 4436 10804
rect 3559 10764 4436 10792
rect 3559 10761 3571 10764
rect 3513 10755 3571 10761
rect 4430 10752 4436 10764
rect 4488 10752 4494 10804
rect 4801 10795 4859 10801
rect 4801 10761 4813 10795
rect 4847 10792 4859 10795
rect 4982 10792 4988 10804
rect 4847 10764 4988 10792
rect 4847 10761 4859 10764
rect 4801 10755 4859 10761
rect 4982 10752 4988 10764
rect 5040 10792 5046 10804
rect 6181 10795 6239 10801
rect 5040 10764 6040 10792
rect 5040 10752 5046 10764
rect 2593 10727 2651 10733
rect 2593 10693 2605 10727
rect 2639 10724 2651 10727
rect 2682 10724 2688 10736
rect 2639 10696 2688 10724
rect 2639 10693 2651 10696
rect 2593 10687 2651 10693
rect 2682 10684 2688 10696
rect 2740 10684 2746 10736
rect 3053 10727 3111 10733
rect 3053 10693 3065 10727
rect 3099 10724 3111 10727
rect 3878 10724 3884 10736
rect 3099 10696 3884 10724
rect 3099 10693 3111 10696
rect 3053 10687 3111 10693
rect 3878 10684 3884 10696
rect 3936 10684 3942 10736
rect 4062 10684 4068 10736
rect 4120 10724 4126 10736
rect 5902 10724 5908 10736
rect 4120 10696 5908 10724
rect 4120 10684 4126 10696
rect 2406 10656 2412 10668
rect 2367 10628 2412 10656
rect 2406 10616 2412 10628
rect 2464 10656 2470 10668
rect 2958 10656 2964 10668
rect 2464 10628 2964 10656
rect 2464 10616 2470 10628
rect 2958 10616 2964 10628
rect 3016 10616 3022 10668
rect 3145 10659 3203 10665
rect 3145 10625 3157 10659
rect 3191 10656 3203 10659
rect 3786 10656 3792 10668
rect 3191 10628 3792 10656
rect 3191 10625 3203 10628
rect 3145 10619 3203 10625
rect 3786 10616 3792 10628
rect 3844 10616 3850 10668
rect 3973 10659 4031 10665
rect 3973 10625 3985 10659
rect 4019 10656 4031 10659
rect 4154 10656 4160 10668
rect 4019 10628 4160 10656
rect 4019 10625 4031 10628
rect 3973 10619 4031 10625
rect 4154 10616 4160 10628
rect 4212 10616 4218 10668
rect 1946 10588 1952 10600
rect 1907 10560 1952 10588
rect 1946 10548 1952 10560
rect 2004 10548 2010 10600
rect 2225 10591 2283 10597
rect 2225 10557 2237 10591
rect 2271 10588 2283 10591
rect 2774 10588 2780 10600
rect 2271 10560 2780 10588
rect 2271 10557 2283 10560
rect 2225 10551 2283 10557
rect 2774 10548 2780 10560
rect 2832 10548 2838 10600
rect 2869 10591 2927 10597
rect 2869 10557 2881 10591
rect 2915 10557 2927 10591
rect 2869 10551 2927 10557
rect 2884 10520 2912 10551
rect 3602 10548 3608 10600
rect 3660 10588 3666 10600
rect 3697 10591 3755 10597
rect 3697 10588 3709 10591
rect 3660 10560 3709 10588
rect 3660 10548 3666 10560
rect 3697 10557 3709 10560
rect 3743 10557 3755 10591
rect 3878 10588 3884 10600
rect 3839 10560 3884 10588
rect 3697 10551 3755 10557
rect 3878 10548 3884 10560
rect 3936 10548 3942 10600
rect 4706 10588 4712 10600
rect 3988 10560 4712 10588
rect 3988 10520 4016 10560
rect 4706 10548 4712 10560
rect 4764 10548 4770 10600
rect 4893 10591 4951 10597
rect 4893 10557 4905 10591
rect 4939 10588 4951 10591
rect 4982 10588 4988 10600
rect 4939 10560 4988 10588
rect 4939 10557 4951 10560
rect 4893 10551 4951 10557
rect 4982 10548 4988 10560
rect 5040 10548 5046 10600
rect 5077 10591 5135 10597
rect 5077 10557 5089 10591
rect 5123 10588 5135 10591
rect 5460 10588 5488 10696
rect 5902 10684 5908 10696
rect 5960 10684 5966 10736
rect 6012 10724 6040 10764
rect 6181 10761 6193 10795
rect 6227 10792 6239 10795
rect 6825 10795 6883 10801
rect 6825 10792 6837 10795
rect 6227 10764 6837 10792
rect 6227 10761 6239 10764
rect 6181 10755 6239 10761
rect 6825 10761 6837 10764
rect 6871 10761 6883 10795
rect 9398 10792 9404 10804
rect 9359 10764 9404 10792
rect 6825 10755 6883 10761
rect 9398 10752 9404 10764
rect 9456 10752 9462 10804
rect 9582 10752 9588 10804
rect 9640 10792 9646 10804
rect 11146 10792 11152 10804
rect 9640 10764 11152 10792
rect 9640 10752 9646 10764
rect 11146 10752 11152 10764
rect 11204 10752 11210 10804
rect 12802 10752 12808 10804
rect 12860 10792 12866 10804
rect 16022 10792 16028 10804
rect 12860 10764 16028 10792
rect 12860 10752 12866 10764
rect 16022 10752 16028 10764
rect 16080 10752 16086 10804
rect 16669 10795 16727 10801
rect 16669 10761 16681 10795
rect 16715 10792 16727 10795
rect 17770 10792 17776 10804
rect 16715 10764 17776 10792
rect 16715 10761 16727 10764
rect 16669 10755 16727 10761
rect 17770 10752 17776 10764
rect 17828 10752 17834 10804
rect 9306 10724 9312 10736
rect 6012 10696 9312 10724
rect 9306 10684 9312 10696
rect 9364 10684 9370 10736
rect 9674 10684 9680 10736
rect 9732 10724 9738 10736
rect 11790 10724 11796 10736
rect 9732 10696 11796 10724
rect 9732 10684 9738 10696
rect 5718 10656 5724 10668
rect 5679 10628 5724 10656
rect 5718 10616 5724 10628
rect 5776 10616 5782 10668
rect 5813 10659 5871 10665
rect 5813 10625 5825 10659
rect 5859 10656 5871 10659
rect 6178 10656 6184 10668
rect 5859 10628 6184 10656
rect 5859 10625 5871 10628
rect 5813 10619 5871 10625
rect 6178 10616 6184 10628
rect 6236 10616 6242 10668
rect 6733 10659 6791 10665
rect 6733 10625 6745 10659
rect 6779 10656 6791 10659
rect 7098 10656 7104 10668
rect 6779 10628 7104 10656
rect 6779 10625 6791 10628
rect 6733 10619 6791 10625
rect 7098 10616 7104 10628
rect 7156 10616 7162 10668
rect 8288 10659 8346 10665
rect 8288 10625 8300 10659
rect 8334 10656 8346 10659
rect 10594 10656 10600 10668
rect 8334 10628 10600 10656
rect 8334 10625 8346 10628
rect 8288 10619 8346 10625
rect 5626 10588 5632 10600
rect 5123 10560 5488 10588
rect 5587 10560 5632 10588
rect 5123 10557 5135 10560
rect 5077 10551 5135 10557
rect 5626 10548 5632 10560
rect 5684 10548 5690 10600
rect 6270 10548 6276 10600
rect 6328 10588 6334 10600
rect 7009 10591 7067 10597
rect 7009 10588 7021 10591
rect 6328 10560 7021 10588
rect 6328 10548 6334 10560
rect 7009 10557 7021 10560
rect 7055 10588 7067 10591
rect 7190 10588 7196 10600
rect 7055 10560 7196 10588
rect 7055 10557 7067 10560
rect 7009 10551 7067 10557
rect 7190 10548 7196 10560
rect 7248 10548 7254 10600
rect 7374 10548 7380 10600
rect 7432 10588 7438 10600
rect 8021 10591 8079 10597
rect 8021 10588 8033 10591
rect 7432 10560 8033 10588
rect 7432 10548 7438 10560
rect 8021 10557 8033 10560
rect 8067 10557 8079 10591
rect 8021 10551 8079 10557
rect 2884 10492 4016 10520
rect 4341 10523 4399 10529
rect 4341 10489 4353 10523
rect 4387 10520 4399 10523
rect 5810 10520 5816 10532
rect 4387 10492 5816 10520
rect 4387 10489 4399 10492
rect 4341 10483 4399 10489
rect 5810 10480 5816 10492
rect 5868 10480 5874 10532
rect 5920 10492 6684 10520
rect 3510 10412 3516 10464
rect 3568 10452 3574 10464
rect 4433 10455 4491 10461
rect 4433 10452 4445 10455
rect 3568 10424 4445 10452
rect 3568 10412 3574 10424
rect 4433 10421 4445 10424
rect 4479 10421 4491 10455
rect 4433 10415 4491 10421
rect 4982 10412 4988 10464
rect 5040 10452 5046 10464
rect 5261 10455 5319 10461
rect 5261 10452 5273 10455
rect 5040 10424 5273 10452
rect 5040 10412 5046 10424
rect 5261 10421 5273 10424
rect 5307 10421 5319 10455
rect 5261 10415 5319 10421
rect 5350 10412 5356 10464
rect 5408 10452 5414 10464
rect 5920 10452 5948 10492
rect 5408 10424 5948 10452
rect 6365 10455 6423 10461
rect 5408 10412 5414 10424
rect 6365 10421 6377 10455
rect 6411 10452 6423 10455
rect 6546 10452 6552 10464
rect 6411 10424 6552 10452
rect 6411 10421 6423 10424
rect 6365 10415 6423 10421
rect 6546 10412 6552 10424
rect 6604 10412 6610 10464
rect 6656 10452 6684 10492
rect 9048 10452 9076 10628
rect 10594 10616 10600 10628
rect 10652 10616 10658 10668
rect 11054 10616 11060 10668
rect 11112 10665 11118 10668
rect 11348 10665 11376 10696
rect 11790 10684 11796 10696
rect 11848 10684 11854 10736
rect 15565 10727 15623 10733
rect 13924 10696 15424 10724
rect 11112 10656 11124 10665
rect 11333 10659 11391 10665
rect 11112 10628 11157 10656
rect 11112 10619 11124 10628
rect 11333 10625 11345 10659
rect 11379 10625 11391 10659
rect 11333 10619 11391 10625
rect 11112 10616 11118 10619
rect 11698 10616 11704 10668
rect 11756 10656 11762 10668
rect 13924 10665 13952 10696
rect 15396 10668 15424 10696
rect 15565 10693 15577 10727
rect 15611 10724 15623 10727
rect 15654 10724 15660 10736
rect 15611 10696 15660 10724
rect 15611 10693 15623 10696
rect 15565 10687 15623 10693
rect 15654 10684 15660 10696
rect 15712 10684 15718 10736
rect 16206 10724 16212 10736
rect 15856 10696 16212 10724
rect 13642 10659 13700 10665
rect 13642 10656 13654 10659
rect 11756 10628 13654 10656
rect 11756 10616 11762 10628
rect 13642 10625 13654 10628
rect 13688 10625 13700 10659
rect 13642 10619 13700 10625
rect 13909 10659 13967 10665
rect 13909 10625 13921 10659
rect 13955 10625 13967 10659
rect 13909 10619 13967 10625
rect 14550 10616 14556 10668
rect 14608 10656 14614 10668
rect 15114 10659 15172 10665
rect 15114 10656 15126 10659
rect 14608 10628 15126 10656
rect 14608 10616 14614 10628
rect 15114 10625 15126 10628
rect 15160 10625 15172 10659
rect 15378 10656 15384 10668
rect 15291 10628 15384 10656
rect 15114 10619 15172 10625
rect 15378 10616 15384 10628
rect 15436 10656 15442 10668
rect 15856 10656 15884 10696
rect 16206 10684 16212 10696
rect 16264 10684 16270 10736
rect 17494 10724 17500 10736
rect 17455 10696 17500 10724
rect 17494 10684 17500 10696
rect 17552 10684 17558 10736
rect 15436 10628 15884 10656
rect 15436 10616 15442 10628
rect 15930 10616 15936 10668
rect 15988 10656 15994 10668
rect 16025 10659 16083 10665
rect 16025 10656 16037 10659
rect 15988 10628 16037 10656
rect 15988 10616 15994 10628
rect 16025 10625 16037 10628
rect 16071 10625 16083 10659
rect 16298 10656 16304 10668
rect 16259 10628 16304 10656
rect 16025 10619 16083 10625
rect 16298 10616 16304 10628
rect 16356 10616 16362 10668
rect 16853 10659 16911 10665
rect 16853 10625 16865 10659
rect 16899 10625 16911 10659
rect 16853 10619 16911 10625
rect 17129 10659 17187 10665
rect 17129 10625 17141 10659
rect 17175 10656 17187 10659
rect 17218 10656 17224 10668
rect 17175 10628 17224 10656
rect 17175 10625 17187 10628
rect 17129 10619 17187 10625
rect 15749 10591 15807 10597
rect 15749 10557 15761 10591
rect 15795 10588 15807 10591
rect 16316 10588 16344 10616
rect 15795 10560 16344 10588
rect 16868 10588 16896 10619
rect 17218 10616 17224 10628
rect 17276 10656 17282 10668
rect 18046 10656 18052 10668
rect 17276 10628 18052 10656
rect 17276 10616 17282 10628
rect 18046 10616 18052 10628
rect 18104 10616 18110 10668
rect 17586 10588 17592 10600
rect 16868 10560 17592 10588
rect 15795 10557 15807 10560
rect 15749 10551 15807 10557
rect 17586 10548 17592 10560
rect 17644 10548 17650 10600
rect 17678 10548 17684 10600
rect 17736 10588 17742 10600
rect 17957 10591 18015 10597
rect 17736 10560 17781 10588
rect 17736 10548 17742 10560
rect 17957 10557 17969 10591
rect 18003 10588 18015 10591
rect 18138 10588 18144 10600
rect 18003 10560 18144 10588
rect 18003 10557 18015 10560
rect 17957 10551 18015 10557
rect 18138 10548 18144 10560
rect 18196 10548 18202 10600
rect 9766 10480 9772 10532
rect 9824 10520 9830 10532
rect 16485 10523 16543 10529
rect 9824 10492 10456 10520
rect 9824 10480 9830 10492
rect 10428 10464 10456 10492
rect 16485 10489 16497 10523
rect 16531 10489 16543 10523
rect 16942 10520 16948 10532
rect 16903 10492 16948 10520
rect 16485 10483 16543 10489
rect 6656 10424 9076 10452
rect 9122 10412 9128 10464
rect 9180 10452 9186 10464
rect 9953 10455 10011 10461
rect 9953 10452 9965 10455
rect 9180 10424 9965 10452
rect 9180 10412 9186 10424
rect 9953 10421 9965 10424
rect 9999 10421 10011 10455
rect 9953 10415 10011 10421
rect 10410 10412 10416 10464
rect 10468 10412 10474 10464
rect 12434 10412 12440 10464
rect 12492 10452 12498 10464
rect 12529 10455 12587 10461
rect 12529 10452 12541 10455
rect 12492 10424 12541 10452
rect 12492 10412 12498 10424
rect 12529 10421 12541 10424
rect 12575 10421 12587 10455
rect 12529 10415 12587 10421
rect 14001 10455 14059 10461
rect 14001 10421 14013 10455
rect 14047 10452 14059 10455
rect 14182 10452 14188 10464
rect 14047 10424 14188 10452
rect 14047 10421 14059 10424
rect 14001 10415 14059 10421
rect 14182 10412 14188 10424
rect 14240 10412 14246 10464
rect 15930 10452 15936 10464
rect 15891 10424 15936 10452
rect 15930 10412 15936 10424
rect 15988 10412 15994 10464
rect 16206 10452 16212 10464
rect 16167 10424 16212 10452
rect 16206 10412 16212 10424
rect 16264 10412 16270 10464
rect 16500 10452 16528 10483
rect 16942 10480 16948 10492
rect 17000 10480 17006 10532
rect 17126 10452 17132 10464
rect 16500 10424 17132 10452
rect 17126 10412 17132 10424
rect 17184 10412 17190 10464
rect 17405 10455 17463 10461
rect 17405 10421 17417 10455
rect 17451 10452 17463 10455
rect 18690 10452 18696 10464
rect 17451 10424 18696 10452
rect 17451 10421 17463 10424
rect 17405 10415 17463 10421
rect 18690 10412 18696 10424
rect 18748 10412 18754 10464
rect 1104 10362 18860 10384
rect 1104 10310 3174 10362
rect 3226 10310 3238 10362
rect 3290 10310 3302 10362
rect 3354 10310 3366 10362
rect 3418 10310 3430 10362
rect 3482 10310 7622 10362
rect 7674 10310 7686 10362
rect 7738 10310 7750 10362
rect 7802 10310 7814 10362
rect 7866 10310 7878 10362
rect 7930 10310 12070 10362
rect 12122 10310 12134 10362
rect 12186 10310 12198 10362
rect 12250 10310 12262 10362
rect 12314 10310 12326 10362
rect 12378 10310 16518 10362
rect 16570 10310 16582 10362
rect 16634 10310 16646 10362
rect 16698 10310 16710 10362
rect 16762 10310 16774 10362
rect 16826 10310 18860 10362
rect 1104 10288 18860 10310
rect 2866 10208 2872 10260
rect 2924 10248 2930 10260
rect 3510 10248 3516 10260
rect 2924 10220 3516 10248
rect 2924 10208 2930 10220
rect 3510 10208 3516 10220
rect 3568 10208 3574 10260
rect 4154 10248 4160 10260
rect 4115 10220 4160 10248
rect 4154 10208 4160 10220
rect 4212 10208 4218 10260
rect 5626 10208 5632 10260
rect 5684 10248 5690 10260
rect 6822 10248 6828 10260
rect 5684 10220 6828 10248
rect 5684 10208 5690 10220
rect 6822 10208 6828 10220
rect 6880 10208 6886 10260
rect 7190 10208 7196 10260
rect 7248 10248 7254 10260
rect 13357 10251 13415 10257
rect 13357 10248 13369 10251
rect 7248 10220 13369 10248
rect 7248 10208 7254 10220
rect 13357 10217 13369 10220
rect 13403 10248 13415 10251
rect 13630 10248 13636 10260
rect 13403 10220 13636 10248
rect 13403 10217 13415 10220
rect 13357 10211 13415 10217
rect 13630 10208 13636 10220
rect 13688 10208 13694 10260
rect 14461 10251 14519 10257
rect 14461 10217 14473 10251
rect 14507 10248 14519 10251
rect 17678 10248 17684 10260
rect 14507 10220 17684 10248
rect 14507 10217 14519 10220
rect 14461 10211 14519 10217
rect 17678 10208 17684 10220
rect 17736 10208 17742 10260
rect 2774 10140 2780 10192
rect 2832 10180 2838 10192
rect 4985 10183 5043 10189
rect 4985 10180 4997 10183
rect 2832 10152 4997 10180
rect 2832 10140 2838 10152
rect 4985 10149 4997 10152
rect 5031 10149 5043 10183
rect 4985 10143 5043 10149
rect 5261 10183 5319 10189
rect 5261 10149 5273 10183
rect 5307 10180 5319 10183
rect 6178 10180 6184 10192
rect 5307 10152 6184 10180
rect 5307 10149 5319 10152
rect 5261 10143 5319 10149
rect 2498 10112 2504 10124
rect 2459 10084 2504 10112
rect 2498 10072 2504 10084
rect 2556 10072 2562 10124
rect 2593 10115 2651 10121
rect 2593 10081 2605 10115
rect 2639 10112 2651 10115
rect 3602 10112 3608 10124
rect 2639 10084 3608 10112
rect 2639 10081 2651 10084
rect 2593 10075 2651 10081
rect 3602 10072 3608 10084
rect 3660 10072 3666 10124
rect 3786 10072 3792 10124
rect 3844 10112 3850 10124
rect 3881 10115 3939 10121
rect 3881 10112 3893 10115
rect 3844 10084 3893 10112
rect 3844 10072 3850 10084
rect 3881 10081 3893 10084
rect 3927 10081 3939 10115
rect 4706 10112 4712 10124
rect 4667 10084 4712 10112
rect 3881 10075 3939 10081
rect 4706 10072 4712 10084
rect 4764 10072 4770 10124
rect 4798 10072 4804 10124
rect 4856 10112 4862 10124
rect 5276 10112 5304 10143
rect 6178 10140 6184 10152
rect 6236 10140 6242 10192
rect 13446 10180 13452 10192
rect 13407 10152 13452 10180
rect 13446 10140 13452 10152
rect 13504 10140 13510 10192
rect 13998 10140 14004 10192
rect 14056 10180 14062 10192
rect 14550 10180 14556 10192
rect 14056 10152 14556 10180
rect 14056 10140 14062 10152
rect 14550 10140 14556 10152
rect 14608 10140 14614 10192
rect 16022 10180 16028 10192
rect 15983 10152 16028 10180
rect 16022 10140 16028 10152
rect 16080 10140 16086 10192
rect 17586 10180 17592 10192
rect 17547 10152 17592 10180
rect 17586 10140 17592 10152
rect 17644 10140 17650 10192
rect 4856 10084 5304 10112
rect 5537 10115 5595 10121
rect 4856 10072 4862 10084
rect 5537 10081 5549 10115
rect 5583 10112 5595 10115
rect 6270 10112 6276 10124
rect 5583 10084 6276 10112
rect 5583 10081 5595 10084
rect 5537 10075 5595 10081
rect 6270 10072 6276 10084
rect 6328 10072 6334 10124
rect 6365 10115 6423 10121
rect 6365 10081 6377 10115
rect 6411 10112 6423 10115
rect 7282 10112 7288 10124
rect 6411 10084 7288 10112
rect 6411 10081 6423 10084
rect 6365 10075 6423 10081
rect 7282 10072 7288 10084
rect 7340 10072 7346 10124
rect 8938 10072 8944 10124
rect 8996 10112 9002 10124
rect 9950 10112 9956 10124
rect 8996 10084 9956 10112
rect 8996 10072 9002 10084
rect 9950 10072 9956 10084
rect 10008 10072 10014 10124
rect 11790 10072 11796 10124
rect 11848 10112 11854 10124
rect 11977 10115 12035 10121
rect 11977 10112 11989 10115
rect 11848 10084 11989 10112
rect 11848 10072 11854 10084
rect 11977 10081 11989 10084
rect 12023 10081 12035 10115
rect 17954 10112 17960 10124
rect 17915 10084 17960 10112
rect 11977 10075 12035 10081
rect 17954 10072 17960 10084
rect 18012 10072 18018 10124
rect 1394 10044 1400 10056
rect 1355 10016 1400 10044
rect 1394 10004 1400 10016
rect 1452 10004 1458 10056
rect 1673 10047 1731 10053
rect 1673 10013 1685 10047
rect 1719 10044 1731 10047
rect 2866 10044 2872 10056
rect 1719 10016 2872 10044
rect 1719 10013 1731 10016
rect 1673 10007 1731 10013
rect 2866 10004 2872 10016
rect 2924 10004 2930 10056
rect 3145 10047 3203 10053
rect 3145 10013 3157 10047
rect 3191 10044 3203 10047
rect 3694 10044 3700 10056
rect 3191 10016 3700 10044
rect 3191 10013 3203 10016
rect 3145 10007 3203 10013
rect 3694 10004 3700 10016
rect 3752 10004 3758 10056
rect 4062 10004 4068 10056
rect 4120 10044 4126 10056
rect 4525 10047 4583 10053
rect 4525 10044 4537 10047
rect 4120 10016 4537 10044
rect 4120 10004 4126 10016
rect 4525 10013 4537 10016
rect 4571 10044 4583 10047
rect 6178 10044 6184 10056
rect 4571 10016 6184 10044
rect 4571 10013 4583 10016
rect 4525 10007 4583 10013
rect 6178 10004 6184 10016
rect 6236 10004 6242 10056
rect 6546 10044 6552 10056
rect 6507 10016 6552 10044
rect 6546 10004 6552 10016
rect 6604 10004 6610 10056
rect 7374 10044 7380 10056
rect 7335 10016 7380 10044
rect 7374 10004 7380 10016
rect 7432 10004 7438 10056
rect 7650 10053 7656 10056
rect 7644 10044 7656 10053
rect 7563 10016 7656 10044
rect 7644 10007 7656 10016
rect 7708 10044 7714 10056
rect 9214 10044 9220 10056
rect 7708 10016 9220 10044
rect 7650 10004 7656 10007
rect 7708 10004 7714 10016
rect 9214 10004 9220 10016
rect 9272 10004 9278 10056
rect 9766 10004 9772 10056
rect 9824 10044 9830 10056
rect 10137 10047 10195 10053
rect 10137 10044 10149 10047
rect 9824 10016 10149 10044
rect 9824 10004 9830 10016
rect 10137 10013 10149 10016
rect 10183 10013 10195 10047
rect 10393 10047 10451 10053
rect 10393 10044 10405 10047
rect 10137 10007 10195 10013
rect 10244 10016 10405 10044
rect 5074 9976 5080 9988
rect 3068 9948 5080 9976
rect 2685 9911 2743 9917
rect 2685 9877 2697 9911
rect 2731 9908 2743 9911
rect 2774 9908 2780 9920
rect 2731 9880 2780 9908
rect 2731 9877 2743 9880
rect 2685 9871 2743 9877
rect 2774 9868 2780 9880
rect 2832 9868 2838 9920
rect 3068 9917 3096 9948
rect 5074 9936 5080 9948
rect 5132 9936 5138 9988
rect 5629 9979 5687 9985
rect 5629 9945 5641 9979
rect 5675 9976 5687 9979
rect 7466 9976 7472 9988
rect 5675 9948 7472 9976
rect 5675 9945 5687 9948
rect 5629 9939 5687 9945
rect 7466 9936 7472 9948
rect 7524 9936 7530 9988
rect 9858 9936 9864 9988
rect 9916 9976 9922 9988
rect 10244 9976 10272 10016
rect 10393 10013 10405 10016
rect 10439 10013 10451 10047
rect 10393 10007 10451 10013
rect 14277 10047 14335 10053
rect 14277 10013 14289 10047
rect 14323 10044 14335 10047
rect 15286 10044 15292 10056
rect 14323 10016 15292 10044
rect 14323 10013 14335 10016
rect 14277 10007 14335 10013
rect 15286 10004 15292 10016
rect 15344 10004 15350 10056
rect 15378 10004 15384 10056
rect 15436 10044 15442 10056
rect 15933 10047 15991 10053
rect 15933 10044 15945 10047
rect 15436 10016 15945 10044
rect 15436 10004 15442 10016
rect 15933 10013 15945 10016
rect 15979 10044 15991 10047
rect 17310 10044 17316 10056
rect 15979 10016 17316 10044
rect 15979 10013 15991 10016
rect 15933 10007 15991 10013
rect 17310 10004 17316 10016
rect 17368 10044 17374 10056
rect 17405 10047 17463 10053
rect 17405 10044 17417 10047
rect 17368 10016 17417 10044
rect 17368 10004 17374 10016
rect 17405 10013 17417 10016
rect 17451 10013 17463 10047
rect 17681 10047 17739 10053
rect 17681 10044 17693 10047
rect 17405 10007 17463 10013
rect 17512 10016 17693 10044
rect 9916 9948 10272 9976
rect 9916 9936 9922 9948
rect 10594 9936 10600 9988
rect 10652 9976 10658 9988
rect 12222 9979 12280 9985
rect 12222 9976 12234 9979
rect 10652 9948 12234 9976
rect 10652 9936 10658 9948
rect 12222 9945 12234 9948
rect 12268 9945 12280 9979
rect 12222 9939 12280 9945
rect 13725 9979 13783 9985
rect 13725 9945 13737 9979
rect 13771 9976 13783 9979
rect 15194 9976 15200 9988
rect 13771 9948 15200 9976
rect 13771 9945 13783 9948
rect 13725 9939 13783 9945
rect 15194 9936 15200 9948
rect 15252 9936 15258 9988
rect 15654 9976 15660 9988
rect 15712 9985 15718 9988
rect 15624 9948 15660 9976
rect 15654 9936 15660 9948
rect 15712 9939 15724 9985
rect 17138 9979 17196 9985
rect 17138 9976 17150 9979
rect 15856 9948 17150 9976
rect 15712 9936 15718 9939
rect 3053 9911 3111 9917
rect 3053 9877 3065 9911
rect 3099 9877 3111 9911
rect 3326 9908 3332 9920
rect 3287 9880 3332 9908
rect 3053 9871 3111 9877
rect 3326 9868 3332 9880
rect 3384 9868 3390 9920
rect 3510 9868 3516 9920
rect 3568 9908 3574 9920
rect 3605 9911 3663 9917
rect 3605 9908 3617 9911
rect 3568 9880 3617 9908
rect 3568 9868 3574 9880
rect 3605 9877 3617 9880
rect 3651 9908 3663 9911
rect 4062 9908 4068 9920
rect 3651 9880 4068 9908
rect 3651 9877 3663 9880
rect 3605 9871 3663 9877
rect 4062 9868 4068 9880
rect 4120 9868 4126 9920
rect 4614 9868 4620 9920
rect 4672 9908 4678 9920
rect 4672 9880 4717 9908
rect 4672 9868 4678 9880
rect 5718 9868 5724 9920
rect 5776 9908 5782 9920
rect 6089 9911 6147 9917
rect 5776 9880 5821 9908
rect 5776 9868 5782 9880
rect 6089 9877 6101 9911
rect 6135 9908 6147 9911
rect 6457 9911 6515 9917
rect 6457 9908 6469 9911
rect 6135 9880 6469 9908
rect 6135 9877 6147 9880
rect 6089 9871 6147 9877
rect 6457 9877 6469 9880
rect 6503 9877 6515 9911
rect 6914 9908 6920 9920
rect 6875 9880 6920 9908
rect 6457 9871 6515 9877
rect 6914 9868 6920 9880
rect 6972 9868 6978 9920
rect 8386 9868 8392 9920
rect 8444 9908 8450 9920
rect 8757 9911 8815 9917
rect 8757 9908 8769 9911
rect 8444 9880 8769 9908
rect 8444 9868 8450 9880
rect 8757 9877 8769 9880
rect 8803 9877 8815 9911
rect 8757 9871 8815 9877
rect 9398 9868 9404 9920
rect 9456 9908 9462 9920
rect 9950 9908 9956 9920
rect 9456 9880 9956 9908
rect 9456 9868 9462 9880
rect 9950 9868 9956 9880
rect 10008 9868 10014 9920
rect 11517 9911 11575 9917
rect 11517 9877 11529 9911
rect 11563 9908 11575 9911
rect 11698 9908 11704 9920
rect 11563 9880 11704 9908
rect 11563 9877 11575 9880
rect 11517 9871 11575 9877
rect 11698 9868 11704 9880
rect 11756 9868 11762 9920
rect 13906 9908 13912 9920
rect 13867 9880 13912 9908
rect 13906 9868 13912 9880
rect 13964 9868 13970 9920
rect 14642 9868 14648 9920
rect 14700 9908 14706 9920
rect 15102 9908 15108 9920
rect 14700 9880 15108 9908
rect 14700 9868 14706 9880
rect 15102 9868 15108 9880
rect 15160 9908 15166 9920
rect 15856 9908 15884 9948
rect 17138 9945 17150 9948
rect 17184 9945 17196 9979
rect 17138 9939 17196 9945
rect 15160 9880 15884 9908
rect 15160 9868 15166 9880
rect 16482 9868 16488 9920
rect 16540 9908 16546 9920
rect 17512 9908 17540 10016
rect 17681 10013 17693 10016
rect 17727 10044 17739 10047
rect 17862 10044 17868 10056
rect 17727 10016 17868 10044
rect 17727 10013 17739 10016
rect 17681 10007 17739 10013
rect 17862 10004 17868 10016
rect 17920 10004 17926 10056
rect 16540 9880 17540 9908
rect 16540 9868 16546 9880
rect 1104 9818 18860 9840
rect 1104 9766 5398 9818
rect 5450 9766 5462 9818
rect 5514 9766 5526 9818
rect 5578 9766 5590 9818
rect 5642 9766 5654 9818
rect 5706 9766 9846 9818
rect 9898 9766 9910 9818
rect 9962 9766 9974 9818
rect 10026 9766 10038 9818
rect 10090 9766 10102 9818
rect 10154 9766 14294 9818
rect 14346 9766 14358 9818
rect 14410 9766 14422 9818
rect 14474 9766 14486 9818
rect 14538 9766 14550 9818
rect 14602 9766 18860 9818
rect 1104 9744 18860 9766
rect 2958 9664 2964 9716
rect 3016 9704 3022 9716
rect 3237 9707 3295 9713
rect 3237 9704 3249 9707
rect 3016 9676 3249 9704
rect 3016 9664 3022 9676
rect 3237 9673 3249 9676
rect 3283 9673 3295 9707
rect 3237 9667 3295 9673
rect 3326 9664 3332 9716
rect 3384 9704 3390 9716
rect 4062 9704 4068 9716
rect 3384 9676 4068 9704
rect 3384 9664 3390 9676
rect 4062 9664 4068 9676
rect 4120 9664 4126 9716
rect 4154 9664 4160 9716
rect 4212 9704 4218 9716
rect 4433 9707 4491 9713
rect 4433 9704 4445 9707
rect 4212 9676 4445 9704
rect 4212 9664 4218 9676
rect 4433 9673 4445 9676
rect 4479 9673 4491 9707
rect 4433 9667 4491 9673
rect 4525 9707 4583 9713
rect 4525 9673 4537 9707
rect 4571 9704 4583 9707
rect 4614 9704 4620 9716
rect 4571 9676 4620 9704
rect 4571 9673 4583 9676
rect 4525 9667 4583 9673
rect 4614 9664 4620 9676
rect 4672 9664 4678 9716
rect 4890 9664 4896 9716
rect 4948 9704 4954 9716
rect 4985 9707 5043 9713
rect 4985 9704 4997 9707
rect 4948 9676 4997 9704
rect 4948 9664 4954 9676
rect 4985 9673 4997 9676
rect 5031 9673 5043 9707
rect 4985 9667 5043 9673
rect 5718 9664 5724 9716
rect 5776 9704 5782 9716
rect 6365 9707 6423 9713
rect 6365 9704 6377 9707
rect 5776 9676 6377 9704
rect 5776 9664 5782 9676
rect 6365 9673 6377 9676
rect 6411 9673 6423 9707
rect 6365 9667 6423 9673
rect 6454 9664 6460 9716
rect 6512 9704 6518 9716
rect 7650 9704 7656 9716
rect 6512 9676 7656 9704
rect 6512 9664 6518 9676
rect 7650 9664 7656 9676
rect 7708 9664 7714 9716
rect 8386 9664 8392 9716
rect 8444 9704 8450 9716
rect 11238 9704 11244 9716
rect 8444 9676 11244 9704
rect 8444 9664 8450 9676
rect 11238 9664 11244 9676
rect 11296 9664 11302 9716
rect 12618 9704 12624 9716
rect 11992 9676 12624 9704
rect 5813 9639 5871 9645
rect 5813 9636 5825 9639
rect 2240 9608 5825 9636
rect 2240 9580 2268 9608
rect 5813 9605 5825 9608
rect 5859 9605 5871 9639
rect 6730 9636 6736 9648
rect 6691 9608 6736 9636
rect 5813 9599 5871 9605
rect 6730 9596 6736 9608
rect 6788 9596 6794 9648
rect 9766 9636 9772 9648
rect 8036 9608 9772 9636
rect 8036 9580 8064 9608
rect 2222 9568 2228 9580
rect 2183 9540 2228 9568
rect 2222 9528 2228 9540
rect 2280 9528 2286 9580
rect 2774 9528 2780 9580
rect 2832 9568 2838 9580
rect 3326 9568 3332 9580
rect 2832 9540 3332 9568
rect 2832 9528 2838 9540
rect 3326 9528 3332 9540
rect 3384 9528 3390 9580
rect 3421 9571 3479 9577
rect 3421 9537 3433 9571
rect 3467 9537 3479 9571
rect 3421 9531 3479 9537
rect 1946 9500 1952 9512
rect 1907 9472 1952 9500
rect 1946 9460 1952 9472
rect 2004 9460 2010 9512
rect 2866 9500 2872 9512
rect 2827 9472 2872 9500
rect 2866 9460 2872 9472
rect 2924 9460 2930 9512
rect 3145 9503 3203 9509
rect 3145 9469 3157 9503
rect 3191 9469 3203 9503
rect 3436 9500 3464 9531
rect 3602 9528 3608 9580
rect 3660 9568 3666 9580
rect 3973 9571 4031 9577
rect 3973 9568 3985 9571
rect 3660 9540 3985 9568
rect 3660 9528 3666 9540
rect 3973 9537 3985 9540
rect 4019 9537 4031 9571
rect 3973 9531 4031 9537
rect 4893 9571 4951 9577
rect 4893 9537 4905 9571
rect 4939 9568 4951 9571
rect 5350 9568 5356 9580
rect 4939 9540 5356 9568
rect 4939 9537 4951 9540
rect 4893 9531 4951 9537
rect 5350 9528 5356 9540
rect 5408 9568 5414 9580
rect 5445 9571 5503 9577
rect 5445 9568 5457 9571
rect 5408 9540 5457 9568
rect 5408 9528 5414 9540
rect 5445 9537 5457 9540
rect 5491 9568 5503 9571
rect 6546 9568 6552 9580
rect 5491 9540 6552 9568
rect 5491 9537 5503 9540
rect 5445 9531 5503 9537
rect 6546 9528 6552 9540
rect 6604 9528 6610 9580
rect 7374 9528 7380 9580
rect 7432 9568 7438 9580
rect 8018 9568 8024 9580
rect 7432 9540 8024 9568
rect 7432 9528 7438 9540
rect 8018 9528 8024 9540
rect 8076 9528 8082 9580
rect 8294 9528 8300 9580
rect 8352 9568 8358 9580
rect 9324 9577 9352 9608
rect 9766 9596 9772 9608
rect 9824 9596 9830 9648
rect 9858 9596 9864 9648
rect 9916 9636 9922 9648
rect 10778 9636 10784 9648
rect 9916 9608 10784 9636
rect 9916 9596 9922 9608
rect 10778 9596 10784 9608
rect 10836 9596 10842 9648
rect 11054 9636 11060 9648
rect 11112 9645 11118 9648
rect 11024 9608 11060 9636
rect 11054 9596 11060 9608
rect 11112 9599 11124 9645
rect 11701 9639 11759 9645
rect 11701 9605 11713 9639
rect 11747 9636 11759 9639
rect 11992 9636 12020 9676
rect 12618 9664 12624 9676
rect 12676 9664 12682 9716
rect 14090 9664 14096 9716
rect 14148 9704 14154 9716
rect 14918 9704 14924 9716
rect 14148 9676 14924 9704
rect 14148 9664 14154 9676
rect 14918 9664 14924 9676
rect 14976 9664 14982 9716
rect 15286 9664 15292 9716
rect 15344 9704 15350 9716
rect 16482 9704 16488 9716
rect 15344 9676 16488 9704
rect 15344 9664 15350 9676
rect 16482 9664 16488 9676
rect 16540 9664 16546 9716
rect 16761 9707 16819 9713
rect 16761 9673 16773 9707
rect 16807 9704 16819 9707
rect 17494 9704 17500 9716
rect 16807 9676 17500 9704
rect 16807 9673 16819 9676
rect 16761 9667 16819 9673
rect 17494 9664 17500 9676
rect 17552 9664 17558 9716
rect 17681 9707 17739 9713
rect 17681 9673 17693 9707
rect 17727 9704 17739 9707
rect 17862 9704 17868 9716
rect 17727 9676 17868 9704
rect 17727 9673 17739 9676
rect 17681 9667 17739 9673
rect 17862 9664 17868 9676
rect 17920 9664 17926 9716
rect 18046 9704 18052 9716
rect 18007 9676 18052 9704
rect 18046 9664 18052 9676
rect 18104 9664 18110 9716
rect 13814 9645 13820 9648
rect 13808 9636 13820 9645
rect 11747 9608 12020 9636
rect 12084 9608 13584 9636
rect 13775 9608 13820 9636
rect 11747 9605 11759 9608
rect 11701 9599 11759 9605
rect 11112 9596 11118 9599
rect 9042 9571 9100 9577
rect 9042 9568 9054 9571
rect 8352 9540 9054 9568
rect 8352 9528 8358 9540
rect 9042 9537 9054 9540
rect 9088 9568 9100 9571
rect 9309 9571 9367 9577
rect 9088 9540 9260 9568
rect 9088 9537 9100 9540
rect 9042 9531 9100 9537
rect 3786 9500 3792 9512
rect 3436 9472 3792 9500
rect 3145 9463 3203 9469
rect 2958 9392 2964 9444
rect 3016 9432 3022 9444
rect 3160 9432 3188 9463
rect 3786 9460 3792 9472
rect 3844 9460 3850 9512
rect 3881 9503 3939 9509
rect 3881 9469 3893 9503
rect 3927 9500 3939 9503
rect 4338 9500 4344 9512
rect 3927 9472 4344 9500
rect 3927 9469 3939 9472
rect 3881 9463 3939 9469
rect 4338 9460 4344 9472
rect 4396 9500 4402 9512
rect 5169 9503 5227 9509
rect 5169 9500 5181 9503
rect 4396 9472 5181 9500
rect 4396 9460 4402 9472
rect 5169 9469 5181 9472
rect 5215 9500 5227 9503
rect 5258 9500 5264 9512
rect 5215 9472 5264 9500
rect 5215 9469 5227 9472
rect 5169 9463 5227 9469
rect 5258 9460 5264 9472
rect 5316 9460 5322 9512
rect 6822 9500 6828 9512
rect 6783 9472 6828 9500
rect 6822 9460 6828 9472
rect 6880 9460 6886 9512
rect 6914 9460 6920 9512
rect 6972 9500 6978 9512
rect 7009 9503 7067 9509
rect 7009 9500 7021 9503
rect 6972 9472 7021 9500
rect 6972 9460 6978 9472
rect 7009 9469 7021 9472
rect 7055 9500 7067 9503
rect 8110 9500 8116 9512
rect 7055 9472 8116 9500
rect 7055 9469 7067 9472
rect 7009 9463 7067 9469
rect 8110 9460 8116 9472
rect 8168 9460 8174 9512
rect 9232 9500 9260 9540
rect 9309 9537 9321 9571
rect 9355 9537 9367 9571
rect 9309 9531 9367 9537
rect 9398 9528 9404 9580
rect 9456 9568 9462 9580
rect 10042 9568 10048 9580
rect 9456 9540 10048 9568
rect 9456 9528 9462 9540
rect 10042 9528 10048 9540
rect 10100 9528 10106 9580
rect 11333 9571 11391 9577
rect 11333 9537 11345 9571
rect 11379 9568 11391 9571
rect 11790 9568 11796 9580
rect 11379 9540 11796 9568
rect 11379 9537 11391 9540
rect 11333 9531 11391 9537
rect 11790 9528 11796 9540
rect 11848 9568 11854 9580
rect 12084 9577 12112 9608
rect 12069 9571 12127 9577
rect 12069 9568 12081 9571
rect 11848 9540 12081 9568
rect 11848 9528 11854 9540
rect 12069 9537 12081 9540
rect 12115 9537 12127 9571
rect 12325 9571 12383 9577
rect 12325 9568 12337 9571
rect 12069 9531 12127 9537
rect 12176 9540 12337 9568
rect 9674 9500 9680 9512
rect 9232 9472 9352 9500
rect 9635 9472 9680 9500
rect 5537 9435 5595 9441
rect 5537 9432 5549 9435
rect 3016 9404 5549 9432
rect 3016 9392 3022 9404
rect 5537 9401 5549 9404
rect 5583 9401 5595 9435
rect 5537 9395 5595 9401
rect 6454 9392 6460 9444
rect 6512 9432 6518 9444
rect 7558 9432 7564 9444
rect 6512 9404 7564 9432
rect 6512 9392 6518 9404
rect 7558 9392 7564 9404
rect 7616 9392 7622 9444
rect 7929 9435 7987 9441
rect 7929 9401 7941 9435
rect 7975 9432 7987 9435
rect 8202 9432 8208 9444
rect 7975 9404 8208 9432
rect 7975 9401 7987 9404
rect 7929 9395 7987 9401
rect 8202 9392 8208 9404
rect 8260 9392 8266 9444
rect 9324 9432 9352 9472
rect 9674 9460 9680 9472
rect 9732 9460 9738 9512
rect 11885 9503 11943 9509
rect 11885 9500 11897 9503
rect 11348 9472 11897 9500
rect 11348 9444 11376 9472
rect 11885 9469 11897 9472
rect 11931 9469 11943 9503
rect 12176 9500 12204 9540
rect 12325 9537 12337 9540
rect 12371 9537 12383 9571
rect 12325 9531 12383 9537
rect 12618 9528 12624 9580
rect 12676 9568 12682 9580
rect 13354 9568 13360 9580
rect 12676 9540 13360 9568
rect 12676 9528 12682 9540
rect 13354 9528 13360 9540
rect 13412 9528 13418 9580
rect 13556 9512 13584 9608
rect 13808 9599 13820 9608
rect 13814 9596 13820 9599
rect 13872 9596 13878 9648
rect 13906 9596 13912 9648
rect 13964 9636 13970 9648
rect 18414 9636 18420 9648
rect 13964 9608 18420 9636
rect 13964 9596 13970 9608
rect 18414 9596 18420 9608
rect 18472 9596 18478 9648
rect 13832 9568 13860 9596
rect 14734 9568 14740 9580
rect 13832 9540 14740 9568
rect 14734 9528 14740 9540
rect 14792 9528 14798 9580
rect 14918 9528 14924 9580
rect 14976 9568 14982 9580
rect 16126 9571 16184 9577
rect 16126 9568 16138 9571
rect 14976 9540 16138 9568
rect 14976 9528 14982 9540
rect 16126 9537 16138 9540
rect 16172 9537 16184 9571
rect 16126 9531 16184 9537
rect 17129 9571 17187 9577
rect 17129 9537 17141 9571
rect 17175 9568 17187 9571
rect 17175 9540 17540 9568
rect 17175 9537 17187 9540
rect 17129 9531 17187 9537
rect 13538 9500 13544 9512
rect 11885 9463 11943 9469
rect 11992 9472 12204 9500
rect 13499 9472 13544 9500
rect 9324 9404 10456 9432
rect 3605 9367 3663 9373
rect 3605 9333 3617 9367
rect 3651 9364 3663 9367
rect 5258 9364 5264 9376
rect 3651 9336 5264 9364
rect 3651 9333 3663 9336
rect 3605 9327 3663 9333
rect 5258 9324 5264 9336
rect 5316 9324 5322 9376
rect 6730 9324 6736 9376
rect 6788 9364 6794 9376
rect 8570 9364 8576 9376
rect 6788 9336 8576 9364
rect 6788 9324 6794 9336
rect 8570 9324 8576 9336
rect 8628 9324 8634 9376
rect 9950 9364 9956 9376
rect 9911 9336 9956 9364
rect 9950 9324 9956 9336
rect 10008 9324 10014 9376
rect 10428 9364 10456 9404
rect 11330 9392 11336 9444
rect 11388 9392 11394 9444
rect 11514 9432 11520 9444
rect 11475 9404 11520 9432
rect 11514 9392 11520 9404
rect 11572 9392 11578 9444
rect 10594 9364 10600 9376
rect 10428 9336 10600 9364
rect 10594 9324 10600 9336
rect 10652 9324 10658 9376
rect 10962 9324 10968 9376
rect 11020 9364 11026 9376
rect 11992 9364 12020 9472
rect 13538 9460 13544 9472
rect 13596 9460 13602 9512
rect 16393 9503 16451 9509
rect 16393 9469 16405 9503
rect 16439 9500 16451 9503
rect 17310 9500 17316 9512
rect 16439 9472 17316 9500
rect 16439 9469 16451 9472
rect 16393 9463 16451 9469
rect 17310 9460 17316 9472
rect 17368 9460 17374 9512
rect 15378 9432 15384 9444
rect 14476 9404 15384 9432
rect 13446 9364 13452 9376
rect 11020 9336 12020 9364
rect 13359 9336 13452 9364
rect 11020 9324 11026 9336
rect 13446 9324 13452 9336
rect 13504 9364 13510 9376
rect 14476 9364 14504 9404
rect 15378 9392 15384 9404
rect 15436 9392 15442 9444
rect 17221 9435 17279 9441
rect 17221 9432 17233 9435
rect 16408 9404 17233 9432
rect 14918 9364 14924 9376
rect 13504 9336 14504 9364
rect 14879 9336 14924 9364
rect 13504 9324 13510 9336
rect 14918 9324 14924 9336
rect 14976 9324 14982 9376
rect 15010 9324 15016 9376
rect 15068 9364 15074 9376
rect 15068 9336 15113 9364
rect 15068 9324 15074 9336
rect 15286 9324 15292 9376
rect 15344 9364 15350 9376
rect 16408 9364 16436 9404
rect 17221 9401 17233 9404
rect 17267 9401 17279 9435
rect 17512 9432 17540 9540
rect 17586 9528 17592 9580
rect 17644 9568 17650 9580
rect 17644 9540 17689 9568
rect 17644 9528 17650 9540
rect 17862 9500 17868 9512
rect 17823 9472 17868 9500
rect 17862 9460 17868 9472
rect 17920 9460 17926 9512
rect 17954 9432 17960 9444
rect 17512 9404 17960 9432
rect 17221 9395 17279 9401
rect 17954 9392 17960 9404
rect 18012 9392 18018 9444
rect 16942 9364 16948 9376
rect 15344 9336 16436 9364
rect 16903 9336 16948 9364
rect 15344 9324 15350 9336
rect 16942 9324 16948 9336
rect 17000 9324 17006 9376
rect 17494 9324 17500 9376
rect 17552 9364 17558 9376
rect 18325 9367 18383 9373
rect 18325 9364 18337 9367
rect 17552 9336 18337 9364
rect 17552 9324 17558 9336
rect 18325 9333 18337 9336
rect 18371 9333 18383 9367
rect 18325 9327 18383 9333
rect 1104 9274 18860 9296
rect 1104 9222 3174 9274
rect 3226 9222 3238 9274
rect 3290 9222 3302 9274
rect 3354 9222 3366 9274
rect 3418 9222 3430 9274
rect 3482 9222 7622 9274
rect 7674 9222 7686 9274
rect 7738 9222 7750 9274
rect 7802 9222 7814 9274
rect 7866 9222 7878 9274
rect 7930 9222 12070 9274
rect 12122 9222 12134 9274
rect 12186 9222 12198 9274
rect 12250 9222 12262 9274
rect 12314 9222 12326 9274
rect 12378 9222 16518 9274
rect 16570 9222 16582 9274
rect 16634 9222 16646 9274
rect 16698 9222 16710 9274
rect 16762 9222 16774 9274
rect 16826 9222 18860 9274
rect 1104 9200 18860 9222
rect 3694 9160 3700 9172
rect 2700 9132 3700 9160
rect 2700 9092 2728 9132
rect 3694 9120 3700 9132
rect 3752 9120 3758 9172
rect 3789 9163 3847 9169
rect 3789 9129 3801 9163
rect 3835 9160 3847 9163
rect 3878 9160 3884 9172
rect 3835 9132 3884 9160
rect 3835 9129 3847 9132
rect 3789 9123 3847 9129
rect 3878 9120 3884 9132
rect 3936 9120 3942 9172
rect 4709 9163 4767 9169
rect 4709 9129 4721 9163
rect 4755 9160 4767 9163
rect 4890 9160 4896 9172
rect 4755 9132 4896 9160
rect 4755 9129 4767 9132
rect 4709 9123 4767 9129
rect 4890 9120 4896 9132
rect 4948 9120 4954 9172
rect 6270 9120 6276 9172
rect 6328 9160 6334 9172
rect 6638 9160 6644 9172
rect 6328 9132 6644 9160
rect 6328 9120 6334 9132
rect 6638 9120 6644 9132
rect 6696 9120 6702 9172
rect 6822 9120 6828 9172
rect 6880 9160 6886 9172
rect 7009 9163 7067 9169
rect 7009 9160 7021 9163
rect 6880 9132 7021 9160
rect 6880 9120 6886 9132
rect 7009 9129 7021 9132
rect 7055 9129 7067 9163
rect 7009 9123 7067 9129
rect 7116 9132 10548 9160
rect 2608 9064 2728 9092
rect 3053 9095 3111 9101
rect 2498 9024 2504 9036
rect 2459 8996 2504 9024
rect 2498 8984 2504 8996
rect 2556 8984 2562 9036
rect 2608 9033 2636 9064
rect 3053 9061 3065 9095
rect 3099 9092 3111 9095
rect 5166 9092 5172 9104
rect 3099 9064 5172 9092
rect 3099 9061 3111 9064
rect 3053 9055 3111 9061
rect 5166 9052 5172 9064
rect 5224 9052 5230 9104
rect 7116 9092 7144 9132
rect 5920 9064 7144 9092
rect 2593 9027 2651 9033
rect 2593 8993 2605 9027
rect 2639 8993 2651 9027
rect 2774 9024 2780 9036
rect 2593 8987 2651 8993
rect 2746 8984 2780 9024
rect 2832 9024 2838 9036
rect 4433 9027 4491 9033
rect 2832 8996 4292 9024
rect 2832 8984 2838 8996
rect 1946 8956 1952 8968
rect 1907 8928 1952 8956
rect 1946 8916 1952 8928
rect 2004 8916 2010 8968
rect 2225 8959 2283 8965
rect 2225 8925 2237 8959
rect 2271 8956 2283 8959
rect 2746 8956 2774 8984
rect 2271 8928 2774 8956
rect 3421 8959 3479 8965
rect 2271 8925 2283 8928
rect 2225 8919 2283 8925
rect 3421 8925 3433 8959
rect 3467 8956 3479 8959
rect 3786 8956 3792 8968
rect 3467 8928 3792 8956
rect 3467 8925 3479 8928
rect 3421 8919 3479 8925
rect 3786 8916 3792 8928
rect 3844 8916 3850 8968
rect 4154 8956 4160 8968
rect 4115 8928 4160 8956
rect 4154 8916 4160 8928
rect 4212 8916 4218 8968
rect 4264 8956 4292 8996
rect 4433 8993 4445 9027
rect 4479 9024 4491 9027
rect 4706 9024 4712 9036
rect 4479 8996 4712 9024
rect 4479 8993 4491 8996
rect 4433 8987 4491 8993
rect 4706 8984 4712 8996
rect 4764 8984 4770 9036
rect 5920 9033 5948 9064
rect 7282 9052 7288 9104
rect 7340 9092 7346 9104
rect 7340 9064 7420 9092
rect 7340 9052 7346 9064
rect 5905 9027 5963 9033
rect 5905 8993 5917 9027
rect 5951 8993 5963 9027
rect 5905 8987 5963 8993
rect 6457 9027 6515 9033
rect 6457 8993 6469 9027
rect 6503 9024 6515 9027
rect 6914 9024 6920 9036
rect 6503 8996 6920 9024
rect 6503 8993 6515 8996
rect 6457 8987 6515 8993
rect 6914 8984 6920 8996
rect 6972 9024 6978 9036
rect 7190 9024 7196 9036
rect 6972 8996 7196 9024
rect 6972 8984 6978 8996
rect 7190 8984 7196 8996
rect 7248 8984 7254 9036
rect 7392 9024 7420 9064
rect 10226 9052 10232 9104
rect 10284 9092 10290 9104
rect 10321 9095 10379 9101
rect 10321 9092 10333 9095
rect 10284 9064 10333 9092
rect 10284 9052 10290 9064
rect 10321 9061 10333 9064
rect 10367 9061 10379 9095
rect 10321 9055 10379 9061
rect 7392 8996 7512 9024
rect 4522 8956 4528 8968
rect 4264 8928 4528 8956
rect 4522 8916 4528 8928
rect 4580 8916 4586 8968
rect 5258 8916 5264 8968
rect 5316 8956 5322 8968
rect 5721 8959 5779 8965
rect 5721 8956 5733 8959
rect 5316 8928 5733 8956
rect 5316 8916 5322 8928
rect 5721 8925 5733 8928
rect 5767 8956 5779 8959
rect 6822 8956 6828 8968
rect 5767 8928 6828 8956
rect 5767 8925 5779 8928
rect 5721 8919 5779 8925
rect 6822 8916 6828 8928
rect 6880 8916 6886 8968
rect 7374 8956 7380 8968
rect 7335 8928 7380 8956
rect 7374 8916 7380 8928
rect 7432 8916 7438 8968
rect 7484 8956 7512 8996
rect 8386 8984 8392 9036
rect 8444 9024 8450 9036
rect 8754 9024 8760 9036
rect 8444 8996 8760 9024
rect 8444 8984 8450 8996
rect 8754 8984 8760 8996
rect 8812 8984 8818 9036
rect 7633 8959 7691 8965
rect 7633 8956 7645 8959
rect 7484 8928 7645 8956
rect 7633 8925 7645 8928
rect 7679 8925 7691 8959
rect 7633 8919 7691 8925
rect 8018 8916 8024 8968
rect 8076 8956 8082 8968
rect 8941 8959 8999 8965
rect 8941 8956 8953 8959
rect 8076 8928 8953 8956
rect 8076 8916 8082 8928
rect 8941 8925 8953 8928
rect 8987 8925 8999 8959
rect 8941 8919 8999 8925
rect 3234 8888 3240 8900
rect 3195 8860 3240 8888
rect 3234 8848 3240 8860
rect 3292 8888 3298 8900
rect 3513 8891 3571 8897
rect 3513 8888 3525 8891
rect 3292 8860 3525 8888
rect 3292 8848 3298 8860
rect 3513 8857 3525 8860
rect 3559 8857 3571 8891
rect 3513 8851 3571 8857
rect 3602 8848 3608 8900
rect 3660 8888 3666 8900
rect 4985 8891 5043 8897
rect 4985 8888 4997 8891
rect 3660 8860 4997 8888
rect 3660 8848 3666 8860
rect 4985 8857 4997 8860
rect 5031 8857 5043 8891
rect 4985 8851 5043 8857
rect 5074 8848 5080 8900
rect 5132 8888 5138 8900
rect 5629 8891 5687 8897
rect 5629 8888 5641 8891
rect 5132 8860 5641 8888
rect 5132 8848 5138 8860
rect 5629 8857 5641 8860
rect 5675 8888 5687 8891
rect 6454 8888 6460 8900
rect 5675 8860 6460 8888
rect 5675 8857 5687 8860
rect 5629 8851 5687 8857
rect 6454 8848 6460 8860
rect 6512 8848 6518 8900
rect 8478 8848 8484 8900
rect 8536 8888 8542 8900
rect 9186 8891 9244 8897
rect 9186 8888 9198 8891
rect 8536 8860 9198 8888
rect 8536 8848 8542 8860
rect 9186 8857 9198 8860
rect 9232 8857 9244 8891
rect 9186 8851 9244 8857
rect 9674 8848 9680 8900
rect 9732 8888 9738 8900
rect 9732 8860 10456 8888
rect 9732 8848 9738 8860
rect 2685 8823 2743 8829
rect 2685 8789 2697 8823
rect 2731 8820 2743 8823
rect 4154 8820 4160 8832
rect 2731 8792 4160 8820
rect 2731 8789 2743 8792
rect 2685 8783 2743 8789
rect 4154 8780 4160 8792
rect 4212 8780 4218 8832
rect 4249 8823 4307 8829
rect 4249 8789 4261 8823
rect 4295 8820 4307 8823
rect 4430 8820 4436 8832
rect 4295 8792 4436 8820
rect 4295 8789 4307 8792
rect 4249 8783 4307 8789
rect 4430 8780 4436 8792
rect 4488 8780 4494 8832
rect 4890 8820 4896 8832
rect 4851 8792 4896 8820
rect 4890 8780 4896 8792
rect 4948 8780 4954 8832
rect 5166 8780 5172 8832
rect 5224 8820 5230 8832
rect 5261 8823 5319 8829
rect 5261 8820 5273 8823
rect 5224 8792 5273 8820
rect 5224 8780 5230 8792
rect 5261 8789 5273 8792
rect 5307 8789 5319 8823
rect 5261 8783 5319 8789
rect 5902 8780 5908 8832
rect 5960 8820 5966 8832
rect 6089 8823 6147 8829
rect 6089 8820 6101 8823
rect 5960 8792 6101 8820
rect 5960 8780 5966 8792
rect 6089 8789 6101 8792
rect 6135 8820 6147 8823
rect 6549 8823 6607 8829
rect 6549 8820 6561 8823
rect 6135 8792 6561 8820
rect 6135 8789 6147 8792
rect 6089 8783 6147 8789
rect 6549 8789 6561 8792
rect 6595 8789 6607 8823
rect 6549 8783 6607 8789
rect 6638 8780 6644 8832
rect 6696 8820 6702 8832
rect 7101 8823 7159 8829
rect 7101 8820 7113 8823
rect 6696 8792 7113 8820
rect 6696 8780 6702 8792
rect 7101 8789 7113 8792
rect 7147 8820 7159 8823
rect 8386 8820 8392 8832
rect 7147 8792 8392 8820
rect 7147 8789 7159 8792
rect 7101 8783 7159 8789
rect 8386 8780 8392 8792
rect 8444 8780 8450 8832
rect 8754 8820 8760 8832
rect 8715 8792 8760 8820
rect 8754 8780 8760 8792
rect 8812 8780 8818 8832
rect 9582 8780 9588 8832
rect 9640 8820 9646 8832
rect 9858 8820 9864 8832
rect 9640 8792 9864 8820
rect 9640 8780 9646 8792
rect 9858 8780 9864 8792
rect 9916 8780 9922 8832
rect 10428 8829 10456 8860
rect 10413 8823 10471 8829
rect 10413 8789 10425 8823
rect 10459 8789 10471 8823
rect 10520 8820 10548 9132
rect 10594 9120 10600 9172
rect 10652 9160 10658 9172
rect 12158 9160 12164 9172
rect 10652 9132 12164 9160
rect 10652 9120 10658 9132
rect 12158 9120 12164 9132
rect 12216 9120 12222 9172
rect 13170 9120 13176 9172
rect 13228 9160 13234 9172
rect 13357 9163 13415 9169
rect 13357 9160 13369 9163
rect 13228 9132 13369 9160
rect 13228 9120 13234 9132
rect 13357 9129 13369 9132
rect 13403 9129 13415 9163
rect 13357 9123 13415 9129
rect 13814 9120 13820 9172
rect 13872 9160 13878 9172
rect 14826 9160 14832 9172
rect 13872 9132 14832 9160
rect 13872 9120 13878 9132
rect 14826 9120 14832 9132
rect 14884 9160 14890 9172
rect 15010 9160 15016 9172
rect 14884 9132 15016 9160
rect 14884 9120 14890 9132
rect 15010 9120 15016 9132
rect 15068 9120 15074 9172
rect 15746 9120 15752 9172
rect 15804 9160 15810 9172
rect 16298 9160 16304 9172
rect 15804 9132 16304 9160
rect 15804 9120 15810 9132
rect 16298 9120 16304 9132
rect 16356 9120 16362 9172
rect 16850 9120 16856 9172
rect 16908 9160 16914 9172
rect 16945 9163 17003 9169
rect 16945 9160 16957 9163
rect 16908 9132 16957 9160
rect 16908 9120 16914 9132
rect 16945 9129 16957 9132
rect 16991 9129 17003 9163
rect 17310 9160 17316 9172
rect 16945 9123 17003 9129
rect 17052 9132 17316 9160
rect 13630 9052 13636 9104
rect 13688 9092 13694 9104
rect 14090 9092 14096 9104
rect 13688 9064 14096 9092
rect 13688 9052 13694 9064
rect 14090 9052 14096 9064
rect 14148 9052 14154 9104
rect 11790 9024 11796 9036
rect 11751 8996 11796 9024
rect 11790 8984 11796 8996
rect 11848 9024 11854 9036
rect 11977 9027 12035 9033
rect 11977 9024 11989 9027
rect 11848 8996 11989 9024
rect 11848 8984 11854 8996
rect 11977 8993 11989 8996
rect 12023 8993 12035 9027
rect 13078 9024 13084 9036
rect 11977 8987 12035 8993
rect 13004 8996 13084 9024
rect 11238 8916 11244 8968
rect 11296 8956 11302 8968
rect 11296 8928 11652 8956
rect 11296 8916 11302 8928
rect 10778 8848 10784 8900
rect 10836 8888 10842 8900
rect 11526 8891 11584 8897
rect 11526 8888 11538 8891
rect 10836 8860 11538 8888
rect 10836 8848 10842 8860
rect 11526 8857 11538 8860
rect 11572 8857 11584 8891
rect 11624 8888 11652 8928
rect 11698 8916 11704 8968
rect 11756 8956 11762 8968
rect 11756 8928 12434 8956
rect 11756 8916 11762 8928
rect 12222 8891 12280 8897
rect 12222 8888 12234 8891
rect 11624 8860 12234 8888
rect 11526 8851 11584 8857
rect 12222 8857 12234 8860
rect 12268 8857 12280 8891
rect 12406 8888 12434 8928
rect 12618 8916 12624 8968
rect 12676 8956 12682 8968
rect 13004 8956 13032 8996
rect 13078 8984 13084 8996
rect 13136 9024 13142 9036
rect 13817 9027 13875 9033
rect 13817 9024 13829 9027
rect 13136 8996 13829 9024
rect 13136 8984 13142 8996
rect 13817 8993 13829 8996
rect 13863 8993 13875 9027
rect 13817 8987 13875 8993
rect 15194 8984 15200 9036
rect 15252 9024 15258 9036
rect 15378 9024 15384 9036
rect 15252 8996 15384 9024
rect 15252 8984 15258 8996
rect 15378 8984 15384 8996
rect 15436 8984 15442 9036
rect 17052 9033 17080 9132
rect 17310 9120 17316 9132
rect 17368 9120 17374 9172
rect 17037 9027 17095 9033
rect 17037 8993 17049 9027
rect 17083 8993 17095 9027
rect 17037 8987 17095 8993
rect 12676 8928 13032 8956
rect 12676 8916 12682 8928
rect 13538 8916 13544 8968
rect 13596 8956 13602 8968
rect 14093 8959 14151 8965
rect 14093 8956 14105 8959
rect 13596 8928 14105 8956
rect 13596 8916 13602 8928
rect 14093 8925 14105 8928
rect 14139 8956 14151 8959
rect 15562 8956 15568 8968
rect 14139 8928 15568 8956
rect 14139 8925 14151 8928
rect 14093 8919 14151 8925
rect 15562 8916 15568 8928
rect 15620 8956 15626 8968
rect 16390 8956 16396 8968
rect 15620 8928 16396 8956
rect 15620 8916 15626 8928
rect 16390 8916 16396 8928
rect 16448 8956 16454 8968
rect 17052 8956 17080 8987
rect 16448 8928 17080 8956
rect 16448 8916 16454 8928
rect 12406 8860 14136 8888
rect 12222 8851 12280 8857
rect 13170 8820 13176 8832
rect 10520 8792 13176 8820
rect 10413 8783 10471 8789
rect 13170 8780 13176 8792
rect 13228 8780 13234 8832
rect 13446 8820 13452 8832
rect 13407 8792 13452 8820
rect 13446 8780 13452 8792
rect 13504 8780 13510 8832
rect 13538 8780 13544 8832
rect 13596 8820 13602 8832
rect 13633 8823 13691 8829
rect 13633 8820 13645 8823
rect 13596 8792 13645 8820
rect 13596 8780 13602 8792
rect 13633 8789 13645 8792
rect 13679 8789 13691 8823
rect 14108 8820 14136 8860
rect 14182 8848 14188 8900
rect 14240 8888 14246 8900
rect 14338 8891 14396 8897
rect 14338 8888 14350 8891
rect 14240 8860 14350 8888
rect 14240 8848 14246 8860
rect 14338 8857 14350 8860
rect 14384 8857 14396 8891
rect 15810 8891 15868 8897
rect 15810 8888 15822 8891
rect 14338 8851 14396 8857
rect 14476 8860 15822 8888
rect 14476 8820 14504 8860
rect 15810 8857 15822 8860
rect 15856 8857 15868 8891
rect 17282 8891 17340 8897
rect 17282 8888 17294 8891
rect 15810 8851 15868 8857
rect 15948 8860 17294 8888
rect 15470 8820 15476 8832
rect 14108 8792 14504 8820
rect 15431 8792 15476 8820
rect 13633 8783 13691 8789
rect 15470 8780 15476 8792
rect 15528 8820 15534 8832
rect 15948 8820 15976 8860
rect 17282 8857 17294 8860
rect 17328 8857 17340 8891
rect 17282 8851 17340 8857
rect 15528 8792 15976 8820
rect 15528 8780 15534 8792
rect 16298 8780 16304 8832
rect 16356 8820 16362 8832
rect 17494 8820 17500 8832
rect 16356 8792 17500 8820
rect 16356 8780 16362 8792
rect 17494 8780 17500 8792
rect 17552 8780 17558 8832
rect 18417 8823 18475 8829
rect 18417 8789 18429 8823
rect 18463 8820 18475 8823
rect 18782 8820 18788 8832
rect 18463 8792 18788 8820
rect 18463 8789 18475 8792
rect 18417 8783 18475 8789
rect 18782 8780 18788 8792
rect 18840 8780 18846 8832
rect 1104 8730 18860 8752
rect 1104 8678 5398 8730
rect 5450 8678 5462 8730
rect 5514 8678 5526 8730
rect 5578 8678 5590 8730
rect 5642 8678 5654 8730
rect 5706 8678 9846 8730
rect 9898 8678 9910 8730
rect 9962 8678 9974 8730
rect 10026 8678 10038 8730
rect 10090 8678 10102 8730
rect 10154 8678 14294 8730
rect 14346 8678 14358 8730
rect 14410 8678 14422 8730
rect 14474 8678 14486 8730
rect 14538 8678 14550 8730
rect 14602 8678 18860 8730
rect 1104 8656 18860 8678
rect 2915 8619 2973 8625
rect 2915 8585 2927 8619
rect 2961 8616 2973 8619
rect 3970 8616 3976 8628
rect 2961 8588 3976 8616
rect 2961 8585 2973 8588
rect 2915 8579 2973 8585
rect 3970 8576 3976 8588
rect 4028 8576 4034 8628
rect 4430 8616 4436 8628
rect 4391 8588 4436 8616
rect 4430 8576 4436 8588
rect 4488 8576 4494 8628
rect 4522 8576 4528 8628
rect 4580 8616 4586 8628
rect 5905 8619 5963 8625
rect 5905 8616 5917 8619
rect 4580 8588 5917 8616
rect 4580 8576 4586 8588
rect 5905 8585 5917 8588
rect 5951 8585 5963 8619
rect 5905 8579 5963 8585
rect 7469 8619 7527 8625
rect 7469 8585 7481 8619
rect 7515 8616 7527 8619
rect 7929 8619 7987 8625
rect 7929 8616 7941 8619
rect 7515 8588 7941 8616
rect 7515 8585 7527 8588
rect 7469 8579 7527 8585
rect 7929 8585 7941 8588
rect 7975 8585 7987 8619
rect 7929 8579 7987 8585
rect 8018 8576 8024 8628
rect 8076 8616 8082 8628
rect 10778 8616 10784 8628
rect 8076 8588 10784 8616
rect 8076 8576 8082 8588
rect 10778 8576 10784 8588
rect 10836 8576 10842 8628
rect 11333 8619 11391 8625
rect 11333 8585 11345 8619
rect 11379 8585 11391 8619
rect 12710 8616 12716 8628
rect 12623 8588 12716 8616
rect 11333 8579 11391 8585
rect 2222 8508 2228 8560
rect 2280 8548 2286 8560
rect 6365 8551 6423 8557
rect 6365 8548 6377 8551
rect 2280 8520 6377 8548
rect 2280 8508 2286 8520
rect 6365 8517 6377 8520
rect 6411 8517 6423 8551
rect 6365 8511 6423 8517
rect 7006 8508 7012 8560
rect 7064 8508 7070 8560
rect 7282 8508 7288 8560
rect 7340 8548 7346 8560
rect 11054 8548 11060 8560
rect 7340 8520 11060 8548
rect 7340 8508 7346 8520
rect 11054 8508 11060 8520
rect 11112 8548 11118 8560
rect 11348 8548 11376 8579
rect 12710 8576 12716 8588
rect 12768 8616 12774 8628
rect 13906 8616 13912 8628
rect 12768 8588 13912 8616
rect 12768 8576 12774 8588
rect 13906 8576 13912 8588
rect 13964 8576 13970 8628
rect 14369 8619 14427 8625
rect 14369 8585 14381 8619
rect 14415 8616 14427 8619
rect 15194 8616 15200 8628
rect 14415 8588 15200 8616
rect 14415 8585 14427 8588
rect 14369 8579 14427 8585
rect 15194 8576 15200 8588
rect 15252 8576 15258 8628
rect 15378 8576 15384 8628
rect 15436 8616 15442 8628
rect 16022 8616 16028 8628
rect 15436 8588 15884 8616
rect 15983 8588 16028 8616
rect 15436 8576 15442 8588
rect 11112 8520 11376 8548
rect 11112 8508 11118 8520
rect 12894 8508 12900 8560
rect 12952 8548 12958 8560
rect 13630 8548 13636 8560
rect 12952 8520 13636 8548
rect 12952 8508 12958 8520
rect 13630 8508 13636 8520
rect 13688 8508 13694 8560
rect 15562 8548 15568 8560
rect 14108 8520 15568 8548
rect 1949 8483 2007 8489
rect 1949 8449 1961 8483
rect 1995 8480 2007 8483
rect 2038 8480 2044 8492
rect 1995 8452 2044 8480
rect 1995 8449 2007 8452
rect 1949 8443 2007 8449
rect 2038 8440 2044 8452
rect 2096 8440 2102 8492
rect 3329 8483 3387 8489
rect 3329 8449 3341 8483
rect 3375 8480 3387 8483
rect 3510 8480 3516 8492
rect 3375 8452 3516 8480
rect 3375 8449 3387 8452
rect 3329 8443 3387 8449
rect 3510 8440 3516 8452
rect 3568 8440 3574 8492
rect 4065 8483 4123 8489
rect 4065 8449 4077 8483
rect 4111 8480 4123 8483
rect 4154 8480 4160 8492
rect 4111 8452 4160 8480
rect 4111 8449 4123 8452
rect 4065 8443 4123 8449
rect 4154 8440 4160 8452
rect 4212 8480 4218 8492
rect 5074 8480 5080 8492
rect 4212 8452 5080 8480
rect 4212 8440 4218 8452
rect 5074 8440 5080 8452
rect 5132 8440 5138 8492
rect 5169 8483 5227 8489
rect 5169 8449 5181 8483
rect 5215 8480 5227 8483
rect 5258 8480 5264 8492
rect 5215 8452 5264 8480
rect 5215 8449 5227 8452
rect 5169 8443 5227 8449
rect 5258 8440 5264 8452
rect 5316 8440 5322 8492
rect 7024 8480 7052 8508
rect 5368 8452 7052 8480
rect 7101 8483 7159 8489
rect 2225 8415 2283 8421
rect 2225 8381 2237 8415
rect 2271 8412 2283 8415
rect 2774 8412 2780 8424
rect 2271 8384 2780 8412
rect 2271 8381 2283 8384
rect 2225 8375 2283 8381
rect 2746 8372 2780 8384
rect 2832 8372 2838 8424
rect 2958 8372 2964 8424
rect 3016 8412 3022 8424
rect 3145 8415 3203 8421
rect 3145 8412 3157 8415
rect 3016 8384 3157 8412
rect 3016 8372 3022 8384
rect 3145 8381 3157 8384
rect 3191 8412 3203 8415
rect 3602 8412 3608 8424
rect 3191 8384 3608 8412
rect 3191 8381 3203 8384
rect 3145 8375 3203 8381
rect 3602 8372 3608 8384
rect 3660 8372 3666 8424
rect 3694 8372 3700 8424
rect 3752 8412 3758 8424
rect 3789 8415 3847 8421
rect 3789 8412 3801 8415
rect 3752 8384 3801 8412
rect 3752 8372 3758 8384
rect 3789 8381 3801 8384
rect 3835 8381 3847 8415
rect 3789 8375 3847 8381
rect 3878 8372 3884 8424
rect 3936 8412 3942 8424
rect 5368 8421 5396 8452
rect 7101 8449 7113 8483
rect 7147 8480 7159 8483
rect 7190 8480 7196 8492
rect 7147 8452 7196 8480
rect 7147 8449 7159 8452
rect 7101 8443 7159 8449
rect 7190 8440 7196 8452
rect 7248 8480 7254 8492
rect 7742 8480 7748 8492
rect 7248 8452 7748 8480
rect 7248 8440 7254 8452
rect 7742 8440 7748 8452
rect 7800 8440 7806 8492
rect 8386 8480 8392 8492
rect 7852 8452 8392 8480
rect 3973 8415 4031 8421
rect 3973 8412 3985 8415
rect 3936 8384 3985 8412
rect 3936 8372 3942 8384
rect 3973 8381 3985 8384
rect 4019 8381 4031 8415
rect 5353 8415 5411 8421
rect 3973 8375 4031 8381
rect 4080 8384 4844 8412
rect 2746 8344 2774 8372
rect 4080 8344 4108 8384
rect 4706 8344 4712 8356
rect 2746 8316 4108 8344
rect 4667 8316 4712 8344
rect 4706 8304 4712 8316
rect 4764 8304 4770 8356
rect 4816 8344 4844 8384
rect 5353 8381 5365 8415
rect 5399 8381 5411 8415
rect 5353 8375 5411 8381
rect 5718 8372 5724 8424
rect 5776 8412 5782 8424
rect 6914 8412 6920 8424
rect 5776 8384 6224 8412
rect 6875 8384 6920 8412
rect 5776 8372 5782 8384
rect 6089 8347 6147 8353
rect 6089 8344 6101 8347
rect 4816 8316 6101 8344
rect 6089 8313 6101 8316
rect 6135 8313 6147 8347
rect 6196 8344 6224 8384
rect 6914 8372 6920 8384
rect 6972 8372 6978 8424
rect 7009 8415 7067 8421
rect 7009 8381 7021 8415
rect 7055 8412 7067 8415
rect 7852 8412 7880 8452
rect 8386 8440 8392 8452
rect 8444 8440 8450 8492
rect 9605 8483 9663 8489
rect 9605 8480 9617 8483
rect 8496 8452 9617 8480
rect 8018 8412 8024 8424
rect 7055 8384 7880 8412
rect 7979 8384 8024 8412
rect 7055 8381 7067 8384
rect 7009 8375 7067 8381
rect 8018 8372 8024 8384
rect 8076 8372 8082 8424
rect 8110 8372 8116 8424
rect 8168 8412 8174 8424
rect 8496 8412 8524 8452
rect 9605 8449 9617 8452
rect 9651 8480 9663 8483
rect 9651 8452 9812 8480
rect 9651 8449 9663 8452
rect 9605 8443 9663 8449
rect 8168 8384 8213 8412
rect 8312 8384 8524 8412
rect 9784 8412 9812 8452
rect 9858 8440 9864 8492
rect 9916 8480 9922 8492
rect 9953 8483 10011 8489
rect 9953 8480 9965 8483
rect 9916 8452 9965 8480
rect 9916 8440 9922 8452
rect 9953 8449 9965 8452
rect 9999 8449 10011 8483
rect 9953 8443 10011 8449
rect 10042 8440 10048 8492
rect 10100 8480 10106 8492
rect 10220 8483 10278 8489
rect 10220 8480 10232 8483
rect 10100 8452 10232 8480
rect 10100 8440 10106 8452
rect 10220 8449 10232 8452
rect 10266 8480 10278 8483
rect 10594 8480 10600 8492
rect 10266 8452 10600 8480
rect 10266 8449 10278 8452
rect 10220 8443 10278 8449
rect 10594 8440 10600 8452
rect 10652 8440 10658 8492
rect 11885 8483 11943 8489
rect 11885 8449 11897 8483
rect 11931 8480 11943 8483
rect 12434 8480 12440 8492
rect 11931 8452 12440 8480
rect 11931 8449 11943 8452
rect 11885 8443 11943 8449
rect 12434 8440 12440 8452
rect 12492 8440 12498 8492
rect 13814 8440 13820 8492
rect 13872 8489 13878 8492
rect 14108 8489 14136 8520
rect 13872 8480 13884 8489
rect 14093 8483 14151 8489
rect 13872 8452 13917 8480
rect 13872 8443 13884 8452
rect 14093 8449 14105 8483
rect 14139 8449 14151 8483
rect 14093 8443 14151 8449
rect 13872 8440 13878 8443
rect 14182 8440 14188 8492
rect 14240 8480 14246 8492
rect 14568 8489 14596 8520
rect 15562 8508 15568 8520
rect 15620 8508 15626 8560
rect 15856 8548 15884 8588
rect 16022 8576 16028 8588
rect 16080 8576 16086 8628
rect 17957 8619 18015 8625
rect 17957 8585 17969 8619
rect 18003 8616 18015 8619
rect 18046 8616 18052 8628
rect 18003 8588 18052 8616
rect 18003 8585 18015 8588
rect 17957 8579 18015 8585
rect 18046 8576 18052 8588
rect 18104 8576 18110 8628
rect 18414 8616 18420 8628
rect 18375 8588 18420 8616
rect 18414 8576 18420 8588
rect 18472 8576 18478 8628
rect 15856 8520 18184 8548
rect 14826 8489 14832 8492
rect 14553 8483 14611 8489
rect 14240 8452 14285 8480
rect 14240 8440 14246 8452
rect 14553 8449 14565 8483
rect 14599 8449 14611 8483
rect 14820 8480 14832 8489
rect 14787 8452 14832 8480
rect 14553 8443 14611 8449
rect 14820 8443 14832 8452
rect 14826 8440 14832 8443
rect 14884 8440 14890 8492
rect 16298 8440 16304 8492
rect 16356 8480 16362 8492
rect 16485 8483 16543 8489
rect 16485 8480 16497 8483
rect 16356 8452 16497 8480
rect 16356 8440 16362 8452
rect 16485 8449 16497 8452
rect 16531 8449 16543 8483
rect 16485 8443 16543 8449
rect 17037 8483 17095 8489
rect 17037 8449 17049 8483
rect 17083 8449 17095 8483
rect 17494 8480 17500 8492
rect 17455 8452 17500 8480
rect 17037 8443 17095 8449
rect 9784 8384 9904 8412
rect 8168 8372 8174 8384
rect 6196 8316 7420 8344
rect 6089 8307 6147 8313
rect 3421 8279 3479 8285
rect 3421 8245 3433 8279
rect 3467 8276 3479 8279
rect 4430 8276 4436 8288
rect 3467 8248 4436 8276
rect 3467 8245 3479 8248
rect 3421 8239 3479 8245
rect 4430 8236 4436 8248
rect 4488 8236 4494 8288
rect 4522 8236 4528 8288
rect 4580 8276 4586 8288
rect 4580 8248 4625 8276
rect 4580 8236 4586 8248
rect 4890 8236 4896 8288
rect 4948 8276 4954 8288
rect 5258 8276 5264 8288
rect 4948 8248 5264 8276
rect 4948 8236 4954 8248
rect 5258 8236 5264 8248
rect 5316 8276 5322 8288
rect 5537 8279 5595 8285
rect 5537 8276 5549 8279
rect 5316 8248 5549 8276
rect 5316 8236 5322 8248
rect 5537 8245 5549 8248
rect 5583 8276 5595 8279
rect 5721 8279 5779 8285
rect 5721 8276 5733 8279
rect 5583 8248 5733 8276
rect 5583 8245 5595 8248
rect 5537 8239 5595 8245
rect 5721 8245 5733 8248
rect 5767 8276 5779 8279
rect 6270 8276 6276 8288
rect 5767 8248 6276 8276
rect 5767 8245 5779 8248
rect 5721 8239 5779 8245
rect 6270 8236 6276 8248
rect 6328 8236 6334 8288
rect 7392 8276 7420 8316
rect 7466 8304 7472 8356
rect 7524 8344 7530 8356
rect 7561 8347 7619 8353
rect 7561 8344 7573 8347
rect 7524 8316 7573 8344
rect 7524 8304 7530 8316
rect 7561 8313 7573 8316
rect 7607 8313 7619 8347
rect 8312 8344 8340 8384
rect 9876 8356 9904 8384
rect 11422 8372 11428 8424
rect 11480 8412 11486 8424
rect 11974 8412 11980 8424
rect 11480 8384 11836 8412
rect 11935 8384 11980 8412
rect 11480 8372 11486 8384
rect 11808 8356 11836 8384
rect 11974 8372 11980 8384
rect 12032 8372 12038 8424
rect 12069 8415 12127 8421
rect 12069 8381 12081 8415
rect 12115 8381 12127 8415
rect 12069 8375 12127 8381
rect 12529 8415 12587 8421
rect 12529 8381 12541 8415
rect 12575 8412 12587 8415
rect 12618 8412 12624 8424
rect 12575 8384 12624 8412
rect 12575 8381 12587 8384
rect 12529 8375 12587 8381
rect 8478 8344 8484 8356
rect 7561 8307 7619 8313
rect 7668 8316 8340 8344
rect 8439 8316 8484 8344
rect 7668 8276 7696 8316
rect 8478 8304 8484 8316
rect 8536 8304 8542 8356
rect 9858 8304 9864 8356
rect 9916 8304 9922 8356
rect 11054 8304 11060 8356
rect 11112 8344 11118 8356
rect 11517 8347 11575 8353
rect 11517 8344 11529 8347
rect 11112 8316 11529 8344
rect 11112 8304 11118 8316
rect 11517 8313 11529 8316
rect 11563 8313 11575 8347
rect 11790 8344 11796 8356
rect 11703 8316 11796 8344
rect 11517 8307 11575 8313
rect 11790 8304 11796 8316
rect 11848 8344 11854 8356
rect 12084 8344 12112 8375
rect 12618 8372 12624 8384
rect 12676 8372 12682 8424
rect 15948 8384 16528 8412
rect 15948 8353 15976 8384
rect 11848 8316 12112 8344
rect 15933 8347 15991 8353
rect 11848 8304 11854 8316
rect 15933 8313 15945 8347
rect 15979 8313 15991 8347
rect 15933 8307 15991 8313
rect 16114 8304 16120 8356
rect 16172 8344 16178 8356
rect 16301 8347 16359 8353
rect 16301 8344 16313 8347
rect 16172 8316 16313 8344
rect 16172 8304 16178 8316
rect 16301 8313 16313 8316
rect 16347 8313 16359 8347
rect 16500 8344 16528 8384
rect 16853 8347 16911 8353
rect 16500 8316 16620 8344
rect 16301 8307 16359 8313
rect 7392 8248 7696 8276
rect 7742 8236 7748 8288
rect 7800 8276 7806 8288
rect 9122 8276 9128 8288
rect 7800 8248 9128 8276
rect 7800 8236 7806 8248
rect 9122 8236 9128 8248
rect 9180 8236 9186 8288
rect 11422 8236 11428 8288
rect 11480 8276 11486 8288
rect 13446 8276 13452 8288
rect 11480 8248 13452 8276
rect 11480 8236 11486 8248
rect 13446 8236 13452 8248
rect 13504 8236 13510 8288
rect 16592 8276 16620 8316
rect 16853 8313 16865 8347
rect 16899 8344 16911 8347
rect 16942 8344 16948 8356
rect 16899 8316 16948 8344
rect 16899 8313 16911 8316
rect 16853 8307 16911 8313
rect 16942 8304 16948 8316
rect 17000 8304 17006 8356
rect 17052 8344 17080 8443
rect 17494 8440 17500 8452
rect 17552 8440 17558 8492
rect 18156 8489 18184 8520
rect 18141 8483 18199 8489
rect 18141 8449 18153 8483
rect 18187 8449 18199 8483
rect 18141 8443 18199 8449
rect 18230 8440 18236 8492
rect 18288 8480 18294 8492
rect 18288 8452 18333 8480
rect 18288 8440 18294 8452
rect 17218 8412 17224 8424
rect 17179 8384 17224 8412
rect 17218 8372 17224 8384
rect 17276 8372 17282 8424
rect 17310 8372 17316 8424
rect 17368 8412 17374 8424
rect 17405 8415 17463 8421
rect 17405 8412 17417 8415
rect 17368 8384 17417 8412
rect 17368 8372 17374 8384
rect 17405 8381 17417 8384
rect 17451 8381 17463 8415
rect 17405 8375 17463 8381
rect 17052 8316 18276 8344
rect 17402 8276 17408 8288
rect 16592 8248 17408 8276
rect 17402 8236 17408 8248
rect 17460 8236 17466 8288
rect 17862 8276 17868 8288
rect 17823 8248 17868 8276
rect 17862 8236 17868 8248
rect 17920 8236 17926 8288
rect 18248 8276 18276 8316
rect 18322 8276 18328 8288
rect 18248 8248 18328 8276
rect 18322 8236 18328 8248
rect 18380 8236 18386 8288
rect 1104 8186 18860 8208
rect 1104 8134 3174 8186
rect 3226 8134 3238 8186
rect 3290 8134 3302 8186
rect 3354 8134 3366 8186
rect 3418 8134 3430 8186
rect 3482 8134 7622 8186
rect 7674 8134 7686 8186
rect 7738 8134 7750 8186
rect 7802 8134 7814 8186
rect 7866 8134 7878 8186
rect 7930 8134 12070 8186
rect 12122 8134 12134 8186
rect 12186 8134 12198 8186
rect 12250 8134 12262 8186
rect 12314 8134 12326 8186
rect 12378 8134 16518 8186
rect 16570 8134 16582 8186
rect 16634 8134 16646 8186
rect 16698 8134 16710 8186
rect 16762 8134 16774 8186
rect 16826 8134 18860 8186
rect 1104 8112 18860 8134
rect 2498 8032 2504 8084
rect 2556 8072 2562 8084
rect 3421 8075 3479 8081
rect 3421 8072 3433 8075
rect 2556 8044 3433 8072
rect 2556 8032 2562 8044
rect 3421 8041 3433 8044
rect 3467 8041 3479 8075
rect 3421 8035 3479 8041
rect 4246 8032 4252 8084
rect 4304 8072 4310 8084
rect 5074 8072 5080 8084
rect 4304 8044 5080 8072
rect 4304 8032 4310 8044
rect 5074 8032 5080 8044
rect 5132 8032 5138 8084
rect 8478 8072 8484 8084
rect 5736 8044 8484 8072
rect 2774 8004 2780 8016
rect 1964 7976 2780 8004
rect 1964 7945 1992 7976
rect 2774 7964 2780 7976
rect 2832 7964 2838 8016
rect 3053 8007 3111 8013
rect 3053 7973 3065 8007
rect 3099 8004 3111 8007
rect 3602 8004 3608 8016
rect 3099 7976 3608 8004
rect 3099 7973 3111 7976
rect 3053 7967 3111 7973
rect 3602 7964 3608 7976
rect 3660 7964 3666 8016
rect 4614 8004 4620 8016
rect 3712 7976 4620 8004
rect 1949 7939 2007 7945
rect 1949 7905 1961 7939
rect 1995 7905 2007 7939
rect 2222 7936 2228 7948
rect 2183 7908 2228 7936
rect 1949 7899 2007 7905
rect 2222 7896 2228 7908
rect 2280 7896 2286 7948
rect 2501 7939 2559 7945
rect 2501 7905 2513 7939
rect 2547 7936 2559 7939
rect 3712 7936 3740 7976
rect 4614 7964 4620 7976
rect 4672 7964 4678 8016
rect 4338 7936 4344 7948
rect 2547 7908 3740 7936
rect 4299 7908 4344 7936
rect 2547 7905 2559 7908
rect 2501 7899 2559 7905
rect 4338 7896 4344 7908
rect 4396 7896 4402 7948
rect 5166 7936 5172 7948
rect 5127 7908 5172 7936
rect 5166 7896 5172 7908
rect 5224 7896 5230 7948
rect 5258 7896 5264 7948
rect 5316 7936 5322 7948
rect 5736 7945 5764 8044
rect 8478 8032 8484 8044
rect 8536 8032 8542 8084
rect 8938 8072 8944 8084
rect 8899 8044 8944 8072
rect 8938 8032 8944 8044
rect 8996 8032 9002 8084
rect 9122 8032 9128 8084
rect 9180 8072 9186 8084
rect 10505 8075 10563 8081
rect 10505 8072 10517 8075
rect 9180 8044 10517 8072
rect 9180 8032 9186 8044
rect 10505 8041 10517 8044
rect 10551 8041 10563 8075
rect 10505 8035 10563 8041
rect 11701 8075 11759 8081
rect 11701 8041 11713 8075
rect 11747 8072 11759 8075
rect 11974 8072 11980 8084
rect 11747 8044 11980 8072
rect 11747 8041 11759 8044
rect 11701 8035 11759 8041
rect 11974 8032 11980 8044
rect 12032 8032 12038 8084
rect 12434 8032 12440 8084
rect 12492 8072 12498 8084
rect 12529 8075 12587 8081
rect 12529 8072 12541 8075
rect 12492 8044 12541 8072
rect 12492 8032 12498 8044
rect 12529 8041 12541 8044
rect 12575 8041 12587 8075
rect 18414 8072 18420 8084
rect 18375 8044 18420 8072
rect 12529 8035 12587 8041
rect 18414 8032 18420 8044
rect 18472 8032 18478 8084
rect 6178 7964 6184 8016
rect 6236 8004 6242 8016
rect 7101 8007 7159 8013
rect 6236 7976 6684 8004
rect 6236 7964 6242 7976
rect 5721 7939 5779 7945
rect 5316 7908 5361 7936
rect 5316 7896 5322 7908
rect 5721 7905 5733 7939
rect 5767 7905 5779 7939
rect 6546 7936 6552 7948
rect 6507 7908 6552 7936
rect 5721 7899 5779 7905
rect 6546 7896 6552 7908
rect 6604 7896 6610 7948
rect 6656 7936 6684 7976
rect 7101 7973 7113 8007
rect 7147 8004 7159 8007
rect 7190 8004 7196 8016
rect 7147 7976 7196 8004
rect 7147 7973 7159 7976
rect 7101 7967 7159 7973
rect 7190 7964 7196 7976
rect 7248 7964 7254 8016
rect 12360 7976 13216 8004
rect 12360 7948 12388 7976
rect 7742 7936 7748 7948
rect 6656 7908 7748 7936
rect 7742 7896 7748 7908
rect 7800 7896 7806 7948
rect 7837 7939 7895 7945
rect 7837 7905 7849 7939
rect 7883 7936 7895 7939
rect 8110 7936 8116 7948
rect 7883 7908 8116 7936
rect 7883 7905 7895 7908
rect 7837 7899 7895 7905
rect 8110 7896 8116 7908
rect 8168 7896 8174 7948
rect 8205 7939 8263 7945
rect 8205 7905 8217 7939
rect 8251 7936 8263 7939
rect 8662 7936 8668 7948
rect 8251 7908 8668 7936
rect 8251 7905 8263 7908
rect 8205 7899 8263 7905
rect 8662 7896 8668 7908
rect 8720 7896 8726 7948
rect 10502 7896 10508 7948
rect 10560 7936 10566 7948
rect 10870 7936 10876 7948
rect 10560 7908 10876 7936
rect 10560 7896 10566 7908
rect 10870 7896 10876 7908
rect 10928 7936 10934 7948
rect 11333 7939 11391 7945
rect 11333 7936 11345 7939
rect 10928 7908 11345 7936
rect 10928 7896 10934 7908
rect 11333 7905 11345 7908
rect 11379 7905 11391 7939
rect 11333 7899 11391 7905
rect 11422 7896 11428 7948
rect 11480 7936 11486 7948
rect 12161 7939 12219 7945
rect 12161 7936 12173 7939
rect 11480 7908 12173 7936
rect 11480 7896 11486 7908
rect 12161 7905 12173 7908
rect 12207 7905 12219 7939
rect 12342 7936 12348 7948
rect 12255 7908 12348 7936
rect 12161 7899 12219 7905
rect 12342 7896 12348 7908
rect 12400 7896 12406 7948
rect 13188 7945 13216 7976
rect 13446 7964 13452 8016
rect 13504 8004 13510 8016
rect 14826 8004 14832 8016
rect 13504 7976 14832 8004
rect 13504 7964 13510 7976
rect 14826 7964 14832 7976
rect 14884 8004 14890 8016
rect 15013 8007 15071 8013
rect 15013 8004 15025 8007
rect 14884 7976 15025 8004
rect 14884 7964 14890 7976
rect 15013 7973 15025 7976
rect 15059 7973 15071 8007
rect 18230 8004 18236 8016
rect 15013 7967 15071 7973
rect 17788 7976 18236 8004
rect 13173 7939 13231 7945
rect 12452 7908 13124 7936
rect 2314 7828 2320 7880
rect 2372 7868 2378 7880
rect 2685 7871 2743 7877
rect 2685 7868 2697 7871
rect 2372 7840 2697 7868
rect 2372 7828 2378 7840
rect 2685 7837 2697 7840
rect 2731 7837 2743 7871
rect 2685 7831 2743 7837
rect 3605 7871 3663 7877
rect 3605 7837 3617 7871
rect 3651 7868 3663 7871
rect 5810 7868 5816 7880
rect 3651 7840 5816 7868
rect 3651 7837 3663 7840
rect 3605 7831 3663 7837
rect 5810 7828 5816 7840
rect 5868 7828 5874 7880
rect 6641 7871 6699 7877
rect 6641 7837 6653 7871
rect 6687 7868 6699 7871
rect 9490 7868 9496 7880
rect 6687 7840 9496 7868
rect 6687 7837 6699 7840
rect 6641 7831 6699 7837
rect 9490 7828 9496 7840
rect 9548 7828 9554 7880
rect 9766 7828 9772 7880
rect 9824 7868 9830 7880
rect 10321 7871 10379 7877
rect 10321 7868 10333 7871
rect 9824 7840 10333 7868
rect 9824 7828 9830 7840
rect 10321 7837 10333 7840
rect 10367 7837 10379 7871
rect 10321 7831 10379 7837
rect 11238 7828 11244 7880
rect 11296 7868 11302 7880
rect 12452 7868 12480 7908
rect 11296 7840 12480 7868
rect 11296 7828 11302 7840
rect 12618 7828 12624 7880
rect 12676 7868 12682 7880
rect 12897 7871 12955 7877
rect 12897 7868 12909 7871
rect 12676 7840 12909 7868
rect 12676 7828 12682 7840
rect 12897 7837 12909 7840
rect 12943 7837 12955 7871
rect 12897 7831 12955 7837
rect 2406 7760 2412 7812
rect 2464 7800 2470 7812
rect 3145 7803 3203 7809
rect 3145 7800 3157 7803
rect 2464 7772 3157 7800
rect 2464 7760 2470 7772
rect 3145 7769 3157 7772
rect 3191 7769 3203 7803
rect 3145 7763 3203 7769
rect 3694 7760 3700 7812
rect 3752 7800 3758 7812
rect 4249 7803 4307 7809
rect 4249 7800 4261 7803
rect 3752 7772 4261 7800
rect 3752 7760 3758 7772
rect 4249 7769 4261 7772
rect 4295 7769 4307 7803
rect 4249 7763 4307 7769
rect 4430 7760 4436 7812
rect 4488 7800 4494 7812
rect 6733 7803 6791 7809
rect 4488 7772 5120 7800
rect 4488 7760 4494 7772
rect 2314 7692 2320 7744
rect 2372 7732 2378 7744
rect 2593 7735 2651 7741
rect 2593 7732 2605 7735
rect 2372 7704 2605 7732
rect 2372 7692 2378 7704
rect 2593 7701 2605 7704
rect 2639 7701 2651 7735
rect 2593 7695 2651 7701
rect 3510 7692 3516 7744
rect 3568 7732 3574 7744
rect 3789 7735 3847 7741
rect 3789 7732 3801 7735
rect 3568 7704 3801 7732
rect 3568 7692 3574 7704
rect 3789 7701 3801 7704
rect 3835 7701 3847 7735
rect 4154 7732 4160 7744
rect 4115 7704 4160 7732
rect 3789 7695 3847 7701
rect 4154 7692 4160 7704
rect 4212 7692 4218 7744
rect 4709 7735 4767 7741
rect 4709 7701 4721 7735
rect 4755 7732 4767 7735
rect 4890 7732 4896 7744
rect 4755 7704 4896 7732
rect 4755 7701 4767 7704
rect 4709 7695 4767 7701
rect 4890 7692 4896 7704
rect 4948 7692 4954 7744
rect 5092 7741 5120 7772
rect 6733 7769 6745 7803
rect 6779 7800 6791 7803
rect 8386 7800 8392 7812
rect 6779 7772 7236 7800
rect 8347 7772 8392 7800
rect 6779 7769 6791 7772
rect 6733 7763 6791 7769
rect 5077 7735 5135 7741
rect 5077 7701 5089 7735
rect 5123 7732 5135 7735
rect 5166 7732 5172 7744
rect 5123 7704 5172 7732
rect 5123 7701 5135 7704
rect 5077 7695 5135 7701
rect 5166 7692 5172 7704
rect 5224 7692 5230 7744
rect 5810 7732 5816 7744
rect 5771 7704 5816 7732
rect 5810 7692 5816 7704
rect 5868 7692 5874 7744
rect 5905 7735 5963 7741
rect 5905 7701 5917 7735
rect 5951 7732 5963 7735
rect 6178 7732 6184 7744
rect 5951 7704 6184 7732
rect 5951 7701 5963 7704
rect 5905 7695 5963 7701
rect 6178 7692 6184 7704
rect 6236 7692 6242 7744
rect 6270 7692 6276 7744
rect 6328 7732 6334 7744
rect 7208 7741 7236 7772
rect 8386 7760 8392 7772
rect 8444 7760 8450 7812
rect 8478 7760 8484 7812
rect 8536 7800 8542 7812
rect 8846 7800 8852 7812
rect 8536 7772 8852 7800
rect 8536 7760 8542 7772
rect 8846 7760 8852 7772
rect 8904 7760 8910 7812
rect 9674 7760 9680 7812
rect 9732 7800 9738 7812
rect 10054 7803 10112 7809
rect 10054 7800 10066 7803
rect 9732 7772 10066 7800
rect 9732 7760 9738 7772
rect 10054 7769 10066 7772
rect 10100 7769 10112 7803
rect 10594 7800 10600 7812
rect 10555 7772 10600 7800
rect 10054 7763 10112 7769
rect 10594 7760 10600 7772
rect 10652 7760 10658 7812
rect 11606 7760 11612 7812
rect 11664 7800 11670 7812
rect 11664 7772 12204 7800
rect 11664 7760 11670 7772
rect 7193 7735 7251 7741
rect 6328 7704 6373 7732
rect 6328 7692 6334 7704
rect 7193 7701 7205 7735
rect 7239 7701 7251 7735
rect 7193 7695 7251 7701
rect 7466 7692 7472 7744
rect 7524 7732 7530 7744
rect 7561 7735 7619 7741
rect 7561 7732 7573 7735
rect 7524 7704 7573 7732
rect 7524 7692 7530 7704
rect 7561 7701 7573 7704
rect 7607 7701 7619 7735
rect 7561 7695 7619 7701
rect 7653 7735 7711 7741
rect 7653 7701 7665 7735
rect 7699 7732 7711 7735
rect 8110 7732 8116 7744
rect 7699 7704 8116 7732
rect 7699 7701 7711 7704
rect 7653 7695 7711 7701
rect 8110 7692 8116 7704
rect 8168 7692 8174 7744
rect 8294 7732 8300 7744
rect 8255 7704 8300 7732
rect 8294 7692 8300 7704
rect 8352 7692 8358 7744
rect 8754 7732 8760 7744
rect 8715 7704 8760 7732
rect 8754 7692 8760 7704
rect 8812 7692 8818 7744
rect 10781 7735 10839 7741
rect 10781 7701 10793 7735
rect 10827 7732 10839 7735
rect 10962 7732 10968 7744
rect 10827 7704 10968 7732
rect 10827 7701 10839 7704
rect 10781 7695 10839 7701
rect 10962 7692 10968 7704
rect 11020 7692 11026 7744
rect 11146 7732 11152 7744
rect 11107 7704 11152 7732
rect 11146 7692 11152 7704
rect 11204 7692 11210 7744
rect 11241 7735 11299 7741
rect 11241 7701 11253 7735
rect 11287 7732 11299 7735
rect 11330 7732 11336 7744
rect 11287 7704 11336 7732
rect 11287 7701 11299 7704
rect 11241 7695 11299 7701
rect 11330 7692 11336 7704
rect 11388 7692 11394 7744
rect 11514 7692 11520 7744
rect 11572 7732 11578 7744
rect 12066 7732 12072 7744
rect 11572 7704 12072 7732
rect 11572 7692 11578 7704
rect 12066 7692 12072 7704
rect 12124 7692 12130 7744
rect 12176 7732 12204 7772
rect 12342 7760 12348 7812
rect 12400 7800 12406 7812
rect 12526 7800 12532 7812
rect 12400 7772 12532 7800
rect 12400 7760 12406 7772
rect 12526 7760 12532 7772
rect 12584 7760 12590 7812
rect 12989 7803 13047 7809
rect 12989 7769 13001 7803
rect 13035 7769 13047 7803
rect 13096 7800 13124 7908
rect 13173 7905 13185 7939
rect 13219 7936 13231 7939
rect 13262 7936 13268 7948
rect 13219 7908 13268 7936
rect 13219 7905 13231 7908
rect 13173 7899 13231 7905
rect 13262 7896 13268 7908
rect 13320 7896 13326 7948
rect 13538 7896 13544 7948
rect 13596 7936 13602 7948
rect 14277 7939 14335 7945
rect 14277 7936 14289 7939
rect 13596 7908 14289 7936
rect 13596 7896 13602 7908
rect 14277 7905 14289 7908
rect 14323 7936 14335 7939
rect 15102 7936 15108 7948
rect 14323 7908 15108 7936
rect 14323 7905 14335 7908
rect 14277 7899 14335 7905
rect 15102 7896 15108 7908
rect 15160 7896 15166 7948
rect 16390 7936 16396 7948
rect 16351 7908 16396 7936
rect 16390 7896 16396 7908
rect 16448 7896 16454 7948
rect 16669 7939 16727 7945
rect 16669 7905 16681 7939
rect 16715 7936 16727 7939
rect 17402 7936 17408 7948
rect 16715 7908 17408 7936
rect 16715 7905 16727 7908
rect 16669 7899 16727 7905
rect 17402 7896 17408 7908
rect 17460 7896 17466 7948
rect 17494 7896 17500 7948
rect 17552 7936 17558 7948
rect 17788 7945 17816 7976
rect 18230 7964 18236 7976
rect 18288 7964 18294 8016
rect 17773 7939 17831 7945
rect 17773 7936 17785 7939
rect 17552 7908 17785 7936
rect 17552 7896 17558 7908
rect 17773 7905 17785 7908
rect 17819 7905 17831 7939
rect 17773 7899 17831 7905
rect 17865 7939 17923 7945
rect 17865 7905 17877 7939
rect 17911 7936 17923 7939
rect 18138 7936 18144 7948
rect 17911 7908 18144 7936
rect 17911 7905 17923 7908
rect 17865 7899 17923 7905
rect 18138 7896 18144 7908
rect 18196 7936 18202 7948
rect 18506 7936 18512 7948
rect 18196 7908 18512 7936
rect 18196 7896 18202 7908
rect 18506 7896 18512 7908
rect 18564 7896 18570 7948
rect 13630 7828 13636 7880
rect 13688 7868 13694 7880
rect 13725 7871 13783 7877
rect 13725 7868 13737 7871
rect 13688 7840 13737 7868
rect 13688 7828 13694 7840
rect 13725 7837 13737 7840
rect 13771 7837 13783 7871
rect 13725 7831 13783 7837
rect 14369 7871 14427 7877
rect 14369 7837 14381 7871
rect 14415 7868 14427 7871
rect 16850 7868 16856 7880
rect 14415 7840 16856 7868
rect 14415 7837 14427 7840
rect 14369 7831 14427 7837
rect 16850 7828 16856 7840
rect 16908 7828 16914 7880
rect 18230 7868 18236 7880
rect 18191 7840 18236 7868
rect 18230 7828 18236 7840
rect 18288 7828 18294 7880
rect 14461 7803 14519 7809
rect 14461 7800 14473 7803
rect 13096 7772 14473 7800
rect 12989 7763 13047 7769
rect 14461 7769 14473 7772
rect 14507 7769 14519 7803
rect 14461 7763 14519 7769
rect 13004 7732 13032 7763
rect 15378 7760 15384 7812
rect 15436 7800 15442 7812
rect 15838 7800 15844 7812
rect 15436 7772 15844 7800
rect 15436 7760 15442 7772
rect 15838 7760 15844 7772
rect 15896 7800 15902 7812
rect 16126 7803 16184 7809
rect 16126 7800 16138 7803
rect 15896 7772 16138 7800
rect 15896 7760 15902 7772
rect 16126 7769 16138 7772
rect 16172 7769 16184 7803
rect 16126 7763 16184 7769
rect 16482 7760 16488 7812
rect 16540 7800 16546 7812
rect 17126 7800 17132 7812
rect 16540 7772 17132 7800
rect 16540 7760 16546 7772
rect 12176 7704 13032 7732
rect 13078 7692 13084 7744
rect 13136 7732 13142 7744
rect 13357 7735 13415 7741
rect 13357 7732 13369 7735
rect 13136 7704 13369 7732
rect 13136 7692 13142 7704
rect 13357 7701 13369 7704
rect 13403 7701 13415 7735
rect 13357 7695 13415 7701
rect 13814 7692 13820 7744
rect 13872 7732 13878 7744
rect 13909 7735 13967 7741
rect 13909 7732 13921 7735
rect 13872 7704 13921 7732
rect 13872 7692 13878 7704
rect 13909 7701 13921 7704
rect 13955 7701 13967 7735
rect 13909 7695 13967 7701
rect 14734 7692 14740 7744
rect 14792 7732 14798 7744
rect 14829 7735 14887 7741
rect 14829 7732 14841 7735
rect 14792 7704 14841 7732
rect 14792 7692 14798 7704
rect 14829 7701 14841 7704
rect 14875 7701 14887 7735
rect 14829 7695 14887 7701
rect 15930 7692 15936 7744
rect 15988 7732 15994 7744
rect 16868 7741 16896 7772
rect 17126 7760 17132 7772
rect 17184 7760 17190 7812
rect 16761 7735 16819 7741
rect 16761 7732 16773 7735
rect 15988 7704 16773 7732
rect 15988 7692 15994 7704
rect 16761 7701 16773 7704
rect 16807 7701 16819 7735
rect 16761 7695 16819 7701
rect 16853 7735 16911 7741
rect 16853 7701 16865 7735
rect 16899 7701 16911 7735
rect 17218 7732 17224 7744
rect 17179 7704 17224 7732
rect 16853 7695 16911 7701
rect 17218 7692 17224 7704
rect 17276 7692 17282 7744
rect 17310 7692 17316 7744
rect 17368 7732 17374 7744
rect 17681 7735 17739 7741
rect 17368 7704 17413 7732
rect 17368 7692 17374 7704
rect 17681 7701 17693 7735
rect 17727 7732 17739 7735
rect 18966 7732 18972 7744
rect 17727 7704 18972 7732
rect 17727 7701 17739 7704
rect 17681 7695 17739 7701
rect 18966 7692 18972 7704
rect 19024 7692 19030 7744
rect 1104 7642 18860 7664
rect 1104 7590 5398 7642
rect 5450 7590 5462 7642
rect 5514 7590 5526 7642
rect 5578 7590 5590 7642
rect 5642 7590 5654 7642
rect 5706 7590 9846 7642
rect 9898 7590 9910 7642
rect 9962 7590 9974 7642
rect 10026 7590 10038 7642
rect 10090 7590 10102 7642
rect 10154 7590 14294 7642
rect 14346 7590 14358 7642
rect 14410 7590 14422 7642
rect 14474 7590 14486 7642
rect 14538 7590 14550 7642
rect 14602 7590 18860 7642
rect 1104 7568 18860 7590
rect 1394 7528 1400 7540
rect 1355 7500 1400 7528
rect 1394 7488 1400 7500
rect 1452 7488 1458 7540
rect 2314 7528 2320 7540
rect 2275 7500 2320 7528
rect 2314 7488 2320 7500
rect 2372 7488 2378 7540
rect 2777 7531 2835 7537
rect 2777 7497 2789 7531
rect 2823 7528 2835 7531
rect 2958 7528 2964 7540
rect 2823 7500 2964 7528
rect 2823 7497 2835 7500
rect 2777 7491 2835 7497
rect 2958 7488 2964 7500
rect 3016 7488 3022 7540
rect 3418 7528 3424 7540
rect 3379 7500 3424 7528
rect 3418 7488 3424 7500
rect 3476 7488 3482 7540
rect 3786 7488 3792 7540
rect 3844 7528 3850 7540
rect 4430 7528 4436 7540
rect 3844 7500 4436 7528
rect 3844 7488 3850 7500
rect 4430 7488 4436 7500
rect 4488 7488 4494 7540
rect 4890 7528 4896 7540
rect 4851 7500 4896 7528
rect 4890 7488 4896 7500
rect 4948 7488 4954 7540
rect 4982 7488 4988 7540
rect 5040 7528 5046 7540
rect 5353 7531 5411 7537
rect 5040 7500 5085 7528
rect 5040 7488 5046 7500
rect 5353 7497 5365 7531
rect 5399 7528 5411 7531
rect 5810 7528 5816 7540
rect 5399 7500 5816 7528
rect 5399 7497 5411 7500
rect 5353 7491 5411 7497
rect 5810 7488 5816 7500
rect 5868 7488 5874 7540
rect 6178 7528 6184 7540
rect 6139 7500 6184 7528
rect 6178 7488 6184 7500
rect 6236 7488 6242 7540
rect 7282 7528 7288 7540
rect 6840 7500 7288 7528
rect 1486 7420 1492 7472
rect 1544 7460 1550 7472
rect 4246 7460 4252 7472
rect 1544 7432 3280 7460
rect 1544 7420 1550 7432
rect 1946 7392 1952 7404
rect 1907 7364 1952 7392
rect 1946 7352 1952 7364
rect 2004 7352 2010 7404
rect 3252 7401 3280 7432
rect 3896 7432 4252 7460
rect 2869 7395 2927 7401
rect 2869 7361 2881 7395
rect 2915 7392 2927 7395
rect 3237 7395 3295 7401
rect 2915 7364 3188 7392
rect 2915 7361 2927 7364
rect 2869 7355 2927 7361
rect 1670 7324 1676 7336
rect 1631 7296 1676 7324
rect 1670 7284 1676 7296
rect 1728 7284 1734 7336
rect 1854 7324 1860 7336
rect 1815 7296 1860 7324
rect 1854 7284 1860 7296
rect 1912 7284 1918 7336
rect 2958 7324 2964 7336
rect 2919 7296 2964 7324
rect 2958 7284 2964 7296
rect 3016 7284 3022 7336
rect 3160 7324 3188 7364
rect 3237 7361 3249 7395
rect 3283 7361 3295 7395
rect 3237 7355 3295 7361
rect 3697 7395 3755 7401
rect 3697 7361 3709 7395
rect 3743 7392 3755 7395
rect 3786 7392 3792 7404
rect 3743 7364 3792 7392
rect 3743 7361 3755 7364
rect 3697 7355 3755 7361
rect 3786 7352 3792 7364
rect 3844 7352 3850 7404
rect 3896 7333 3924 7432
rect 4246 7420 4252 7432
rect 4304 7420 4310 7472
rect 4338 7420 4344 7472
rect 4396 7460 4402 7472
rect 6840 7460 6868 7500
rect 7282 7488 7288 7500
rect 7340 7488 7346 7540
rect 7745 7531 7803 7537
rect 7745 7497 7757 7531
rect 7791 7528 7803 7531
rect 7926 7528 7932 7540
rect 7791 7500 7932 7528
rect 7791 7497 7803 7500
rect 7745 7491 7803 7497
rect 7926 7488 7932 7500
rect 7984 7488 7990 7540
rect 8110 7528 8116 7540
rect 8071 7500 8116 7528
rect 8110 7488 8116 7500
rect 8168 7488 8174 7540
rect 8294 7488 8300 7540
rect 8352 7528 8358 7540
rect 8941 7531 8999 7537
rect 8941 7528 8953 7531
rect 8352 7500 8953 7528
rect 8352 7488 8358 7500
rect 8941 7497 8953 7500
rect 8987 7497 8999 7531
rect 8941 7491 8999 7497
rect 9030 7488 9036 7540
rect 9088 7528 9094 7540
rect 9398 7528 9404 7540
rect 9088 7500 9404 7528
rect 9088 7488 9094 7500
rect 9398 7488 9404 7500
rect 9456 7488 9462 7540
rect 9769 7531 9827 7537
rect 9769 7497 9781 7531
rect 9815 7497 9827 7531
rect 9769 7491 9827 7497
rect 10137 7531 10195 7537
rect 10137 7497 10149 7531
rect 10183 7528 10195 7531
rect 10686 7528 10692 7540
rect 10183 7500 10692 7528
rect 10183 7497 10195 7500
rect 10137 7491 10195 7497
rect 4396 7432 6868 7460
rect 4396 7420 4402 7432
rect 6914 7420 6920 7472
rect 6972 7460 6978 7472
rect 7377 7463 7435 7469
rect 6972 7432 7144 7460
rect 6972 7420 6978 7432
rect 4157 7395 4215 7401
rect 4157 7361 4169 7395
rect 4203 7392 4215 7395
rect 5074 7392 5080 7404
rect 4203 7364 5080 7392
rect 4203 7361 4215 7364
rect 4157 7355 4215 7361
rect 5074 7352 5080 7364
rect 5132 7352 5138 7404
rect 5813 7395 5871 7401
rect 5813 7361 5825 7395
rect 5859 7392 5871 7395
rect 6822 7392 6828 7404
rect 5859 7364 6828 7392
rect 5859 7361 5871 7364
rect 5813 7355 5871 7361
rect 6822 7352 6828 7364
rect 6880 7352 6886 7404
rect 3881 7327 3939 7333
rect 3160 7296 3832 7324
rect 3513 7259 3571 7265
rect 3513 7256 3525 7259
rect 1688 7228 3525 7256
rect 1688 7200 1716 7228
rect 3513 7225 3525 7228
rect 3559 7225 3571 7259
rect 3804 7256 3832 7296
rect 3881 7293 3893 7327
rect 3927 7293 3939 7327
rect 3881 7287 3939 7293
rect 4065 7327 4123 7333
rect 4065 7293 4077 7327
rect 4111 7324 4123 7327
rect 4614 7324 4620 7336
rect 4111 7296 4620 7324
rect 4111 7293 4123 7296
rect 4065 7287 4123 7293
rect 4614 7284 4620 7296
rect 4672 7284 4678 7336
rect 4801 7327 4859 7333
rect 4801 7293 4813 7327
rect 4847 7324 4859 7327
rect 5626 7324 5632 7336
rect 4847 7296 5632 7324
rect 4847 7293 4859 7296
rect 4801 7287 4859 7293
rect 5626 7284 5632 7296
rect 5684 7284 5690 7336
rect 5721 7327 5779 7333
rect 5721 7293 5733 7327
rect 5767 7293 5779 7327
rect 6638 7324 6644 7336
rect 6599 7296 6644 7324
rect 5721 7287 5779 7293
rect 3970 7256 3976 7268
rect 3804 7228 3976 7256
rect 3513 7219 3571 7225
rect 3970 7216 3976 7228
rect 4028 7216 4034 7268
rect 4525 7259 4583 7265
rect 4525 7225 4537 7259
rect 4571 7225 4583 7259
rect 5736 7256 5764 7287
rect 6638 7284 6644 7296
rect 6696 7284 6702 7336
rect 6914 7324 6920 7336
rect 6875 7296 6920 7324
rect 6914 7284 6920 7296
rect 6972 7284 6978 7336
rect 7116 7333 7144 7432
rect 7377 7429 7389 7463
rect 7423 7460 7435 7463
rect 9306 7460 9312 7472
rect 7423 7432 9312 7460
rect 7423 7429 7435 7432
rect 7377 7423 7435 7429
rect 9306 7420 9312 7432
rect 9364 7420 9370 7472
rect 8478 7392 8484 7404
rect 7392 7364 8484 7392
rect 7392 7336 7420 7364
rect 8478 7352 8484 7364
rect 8536 7352 8542 7404
rect 8573 7395 8631 7401
rect 8573 7361 8585 7395
rect 8619 7392 8631 7395
rect 8846 7392 8852 7404
rect 8619 7364 8852 7392
rect 8619 7361 8631 7364
rect 8573 7355 8631 7361
rect 8846 7352 8852 7364
rect 8904 7352 8910 7404
rect 9784 7392 9812 7491
rect 10686 7488 10692 7500
rect 10744 7488 10750 7540
rect 10962 7528 10968 7540
rect 10923 7500 10968 7528
rect 10962 7488 10968 7500
rect 11020 7488 11026 7540
rect 11333 7531 11391 7537
rect 11333 7497 11345 7531
rect 11379 7528 11391 7531
rect 11885 7531 11943 7537
rect 11885 7528 11897 7531
rect 11379 7500 11897 7528
rect 11379 7497 11391 7500
rect 11333 7491 11391 7497
rect 11885 7497 11897 7500
rect 11931 7497 11943 7531
rect 13078 7528 13084 7540
rect 13039 7500 13084 7528
rect 11885 7491 11943 7497
rect 13078 7488 13084 7500
rect 13136 7488 13142 7540
rect 13449 7531 13507 7537
rect 13449 7497 13461 7531
rect 13495 7528 13507 7531
rect 13909 7531 13967 7537
rect 13909 7528 13921 7531
rect 13495 7500 13921 7528
rect 13495 7497 13507 7500
rect 13449 7491 13507 7497
rect 13909 7497 13921 7500
rect 13955 7497 13967 7531
rect 14734 7528 14740 7540
rect 14695 7500 14740 7528
rect 13909 7491 13967 7497
rect 14734 7488 14740 7500
rect 14792 7488 14798 7540
rect 14826 7488 14832 7540
rect 14884 7528 14890 7540
rect 15746 7528 15752 7540
rect 14884 7500 15752 7528
rect 14884 7488 14890 7500
rect 15746 7488 15752 7500
rect 15804 7488 15810 7540
rect 15930 7488 15936 7540
rect 15988 7528 15994 7540
rect 16025 7531 16083 7537
rect 16025 7528 16037 7531
rect 15988 7500 16037 7528
rect 15988 7488 15994 7500
rect 16025 7497 16037 7500
rect 16071 7497 16083 7531
rect 16390 7528 16396 7540
rect 16351 7500 16396 7528
rect 16025 7491 16083 7497
rect 16390 7488 16396 7500
rect 16448 7488 16454 7540
rect 16669 7531 16727 7537
rect 16669 7497 16681 7531
rect 16715 7497 16727 7531
rect 16669 7491 16727 7497
rect 17129 7531 17187 7537
rect 17129 7497 17141 7531
rect 17175 7528 17187 7531
rect 17310 7528 17316 7540
rect 17175 7500 17316 7528
rect 17175 7497 17187 7500
rect 17129 7491 17187 7497
rect 10226 7460 10232 7472
rect 10060 7432 10232 7460
rect 9858 7392 9864 7404
rect 9784 7364 9864 7392
rect 9858 7352 9864 7364
rect 9916 7352 9922 7404
rect 7101 7327 7159 7333
rect 7101 7293 7113 7327
rect 7147 7293 7159 7327
rect 7101 7287 7159 7293
rect 7285 7327 7343 7333
rect 7285 7293 7297 7327
rect 7331 7293 7343 7327
rect 7285 7287 7343 7293
rect 4525 7219 4583 7225
rect 4908 7228 5764 7256
rect 1670 7148 1676 7200
rect 1728 7148 1734 7200
rect 2038 7148 2044 7200
rect 2096 7188 2102 7200
rect 2409 7191 2467 7197
rect 2409 7188 2421 7191
rect 2096 7160 2421 7188
rect 2096 7148 2102 7160
rect 2409 7157 2421 7160
rect 2455 7157 2467 7191
rect 2409 7151 2467 7157
rect 2774 7148 2780 7200
rect 2832 7188 2838 7200
rect 4430 7188 4436 7200
rect 2832 7160 4436 7188
rect 2832 7148 2838 7160
rect 4430 7148 4436 7160
rect 4488 7148 4494 7200
rect 4540 7188 4568 7219
rect 4908 7188 4936 7228
rect 7006 7216 7012 7268
rect 7064 7256 7070 7268
rect 7300 7256 7328 7287
rect 7374 7284 7380 7336
rect 7432 7284 7438 7336
rect 8021 7327 8079 7333
rect 8021 7293 8033 7327
rect 8067 7324 8079 7327
rect 8294 7324 8300 7336
rect 8067 7296 8300 7324
rect 8067 7293 8079 7296
rect 8021 7287 8079 7293
rect 8294 7284 8300 7296
rect 8352 7284 8358 7336
rect 8662 7284 8668 7336
rect 8720 7324 8726 7336
rect 8757 7327 8815 7333
rect 8757 7324 8769 7327
rect 8720 7296 8769 7324
rect 8720 7284 8726 7296
rect 8757 7293 8769 7296
rect 8803 7293 8815 7327
rect 9398 7324 9404 7336
rect 9359 7296 9404 7324
rect 8757 7287 8815 7293
rect 7064 7228 7328 7256
rect 7064 7216 7070 7228
rect 7742 7216 7748 7268
rect 7800 7256 7806 7268
rect 8478 7256 8484 7268
rect 7800 7228 8484 7256
rect 7800 7216 7806 7228
rect 8478 7216 8484 7228
rect 8536 7216 8542 7268
rect 8772 7256 8800 7287
rect 9398 7284 9404 7296
rect 9456 7284 9462 7336
rect 9585 7327 9643 7333
rect 9585 7293 9597 7327
rect 9631 7324 9643 7327
rect 10060 7324 10088 7432
rect 10226 7420 10232 7432
rect 10284 7420 10290 7472
rect 11146 7420 11152 7472
rect 11204 7460 11210 7472
rect 12345 7463 12403 7469
rect 12345 7460 12357 7463
rect 11204 7432 12357 7460
rect 11204 7420 11210 7432
rect 12345 7429 12357 7432
rect 12391 7429 12403 7463
rect 12986 7460 12992 7472
rect 12947 7432 12992 7460
rect 12345 7423 12403 7429
rect 12986 7420 12992 7432
rect 13044 7420 13050 7472
rect 13262 7420 13268 7472
rect 13320 7460 13326 7472
rect 14182 7460 14188 7472
rect 13320 7432 14188 7460
rect 13320 7420 13326 7432
rect 14182 7420 14188 7432
rect 14240 7420 14246 7472
rect 14550 7420 14556 7472
rect 14608 7460 14614 7472
rect 16684 7460 16712 7491
rect 17310 7488 17316 7500
rect 17368 7488 17374 7540
rect 17862 7488 17868 7540
rect 17920 7528 17926 7540
rect 17957 7531 18015 7537
rect 17957 7528 17969 7531
rect 17920 7500 17969 7528
rect 17920 7488 17926 7500
rect 17957 7497 17969 7500
rect 18003 7497 18015 7531
rect 18322 7528 18328 7540
rect 18283 7500 18328 7528
rect 17957 7491 18015 7497
rect 18322 7488 18328 7500
rect 18380 7488 18386 7540
rect 14608 7432 16712 7460
rect 14608 7420 14614 7432
rect 17586 7420 17592 7472
rect 17644 7460 17650 7472
rect 17644 7432 18552 7460
rect 17644 7420 17650 7432
rect 10594 7392 10600 7404
rect 10244 7364 10600 7392
rect 10244 7336 10272 7364
rect 10594 7352 10600 7364
rect 10652 7352 10658 7404
rect 11698 7352 11704 7404
rect 11756 7392 11762 7404
rect 14001 7395 14059 7401
rect 11756 7364 12112 7392
rect 11756 7352 11762 7364
rect 10226 7324 10232 7336
rect 9631 7296 10088 7324
rect 10187 7296 10232 7324
rect 9631 7293 9643 7296
rect 9585 7287 9643 7293
rect 10226 7284 10232 7296
rect 10284 7284 10290 7336
rect 10318 7284 10324 7336
rect 10376 7324 10382 7336
rect 10376 7296 10421 7324
rect 10376 7284 10382 7296
rect 10502 7284 10508 7336
rect 10560 7324 10566 7336
rect 10689 7327 10747 7333
rect 10689 7324 10701 7327
rect 10560 7296 10701 7324
rect 10560 7284 10566 7296
rect 10689 7293 10701 7296
rect 10735 7293 10747 7327
rect 10689 7287 10747 7293
rect 10873 7327 10931 7333
rect 10873 7293 10885 7327
rect 10919 7324 10931 7327
rect 11422 7324 11428 7336
rect 10919 7296 11428 7324
rect 10919 7293 10931 7296
rect 10873 7287 10931 7293
rect 11422 7284 11428 7296
rect 11480 7284 11486 7336
rect 11606 7284 11612 7336
rect 11664 7324 11670 7336
rect 12084 7333 12112 7364
rect 14001 7361 14013 7395
rect 14047 7392 14059 7395
rect 15286 7392 15292 7404
rect 14047 7364 15292 7392
rect 14047 7361 14059 7364
rect 14001 7355 14059 7361
rect 15286 7352 15292 7364
rect 15344 7352 15350 7404
rect 15565 7395 15623 7401
rect 15565 7361 15577 7395
rect 15611 7392 15623 7395
rect 16206 7392 16212 7404
rect 15611 7364 16088 7392
rect 16167 7364 16212 7392
rect 15611 7361 15623 7364
rect 15565 7355 15623 7361
rect 11977 7327 12035 7333
rect 11977 7324 11989 7327
rect 11664 7296 11989 7324
rect 11664 7284 11670 7296
rect 11977 7293 11989 7296
rect 12023 7293 12035 7327
rect 11977 7287 12035 7293
rect 12069 7327 12127 7333
rect 12069 7293 12081 7327
rect 12115 7293 12127 7327
rect 12069 7287 12127 7293
rect 12434 7284 12440 7336
rect 12492 7324 12498 7336
rect 12802 7324 12808 7336
rect 12492 7296 12808 7324
rect 12492 7284 12498 7296
rect 12802 7284 12808 7296
rect 12860 7284 12866 7336
rect 12897 7327 12955 7333
rect 12897 7293 12909 7327
rect 12943 7324 12955 7327
rect 13170 7324 13176 7336
rect 12943 7296 13176 7324
rect 12943 7293 12955 7296
rect 12897 7287 12955 7293
rect 13170 7284 13176 7296
rect 13228 7324 13234 7336
rect 13538 7324 13544 7336
rect 13228 7296 13544 7324
rect 13228 7284 13234 7296
rect 13538 7284 13544 7296
rect 13596 7284 13602 7336
rect 14093 7327 14151 7333
rect 14093 7293 14105 7327
rect 14139 7293 14151 7327
rect 14093 7287 14151 7293
rect 10336 7256 10364 7284
rect 8772 7228 10364 7256
rect 10594 7216 10600 7268
rect 10652 7256 10658 7268
rect 11330 7256 11336 7268
rect 10652 7228 11336 7256
rect 10652 7216 10658 7228
rect 11330 7216 11336 7228
rect 11388 7216 11394 7268
rect 14108 7256 14136 7287
rect 14182 7284 14188 7336
rect 14240 7324 14246 7336
rect 14829 7327 14887 7333
rect 14829 7324 14841 7327
rect 14240 7296 14841 7324
rect 14240 7284 14246 7296
rect 14829 7293 14841 7296
rect 14875 7293 14887 7327
rect 14829 7287 14887 7293
rect 15013 7327 15071 7333
rect 15013 7293 15025 7327
rect 15059 7324 15071 7327
rect 15378 7324 15384 7336
rect 15059 7296 15384 7324
rect 15059 7293 15071 7296
rect 15013 7287 15071 7293
rect 15028 7256 15056 7287
rect 15378 7284 15384 7296
rect 15436 7284 15442 7336
rect 15657 7327 15715 7333
rect 15657 7293 15669 7327
rect 15703 7293 15715 7327
rect 15657 7287 15715 7293
rect 11440 7228 12434 7256
rect 14108 7228 15056 7256
rect 15672 7256 15700 7287
rect 15746 7284 15752 7336
rect 15804 7324 15810 7336
rect 16060 7324 16088 7364
rect 16206 7352 16212 7364
rect 16264 7352 16270 7404
rect 17037 7395 17095 7401
rect 17037 7361 17049 7395
rect 17083 7392 17095 7395
rect 17402 7392 17408 7404
rect 17083 7364 17408 7392
rect 17083 7361 17095 7364
rect 17037 7355 17095 7361
rect 17402 7352 17408 7364
rect 17460 7352 17466 7404
rect 17862 7392 17868 7404
rect 17823 7364 17868 7392
rect 17862 7352 17868 7364
rect 17920 7352 17926 7404
rect 18524 7401 18552 7432
rect 18509 7395 18567 7401
rect 18509 7361 18521 7395
rect 18555 7361 18567 7395
rect 18509 7355 18567 7361
rect 17126 7324 17132 7336
rect 15804 7296 15849 7324
rect 16060 7296 17132 7324
rect 15804 7284 15810 7296
rect 17126 7284 17132 7296
rect 17184 7284 17190 7336
rect 17313 7327 17371 7333
rect 17313 7293 17325 7327
rect 17359 7324 17371 7327
rect 18138 7324 18144 7336
rect 17359 7296 17632 7324
rect 18099 7296 18144 7324
rect 17359 7293 17371 7296
rect 17313 7287 17371 7293
rect 17497 7259 17555 7265
rect 17497 7256 17509 7259
rect 15672 7228 17509 7256
rect 4540 7160 4936 7188
rect 5074 7148 5080 7200
rect 5132 7188 5138 7200
rect 11440 7188 11468 7228
rect 5132 7160 11468 7188
rect 11517 7191 11575 7197
rect 5132 7148 5138 7160
rect 11517 7157 11529 7191
rect 11563 7188 11575 7191
rect 11698 7188 11704 7200
rect 11563 7160 11704 7188
rect 11563 7157 11575 7160
rect 11517 7151 11575 7157
rect 11698 7148 11704 7160
rect 11756 7148 11762 7200
rect 12406 7188 12434 7228
rect 17497 7225 17509 7228
rect 17543 7225 17555 7259
rect 17497 7219 17555 7225
rect 12986 7188 12992 7200
rect 12406 7160 12992 7188
rect 12986 7148 12992 7160
rect 13044 7148 13050 7200
rect 13538 7188 13544 7200
rect 13499 7160 13544 7188
rect 13538 7148 13544 7160
rect 13596 7148 13602 7200
rect 13630 7148 13636 7200
rect 13688 7188 13694 7200
rect 14369 7191 14427 7197
rect 14369 7188 14381 7191
rect 13688 7160 14381 7188
rect 13688 7148 13694 7160
rect 14369 7157 14381 7160
rect 14415 7157 14427 7191
rect 15194 7188 15200 7200
rect 15155 7160 15200 7188
rect 14369 7151 14427 7157
rect 15194 7148 15200 7160
rect 15252 7148 15258 7200
rect 15746 7148 15752 7200
rect 15804 7188 15810 7200
rect 17604 7188 17632 7296
rect 18138 7284 18144 7296
rect 18196 7284 18202 7336
rect 15804 7160 17632 7188
rect 15804 7148 15810 7160
rect 1104 7098 18860 7120
rect 1104 7046 3174 7098
rect 3226 7046 3238 7098
rect 3290 7046 3302 7098
rect 3354 7046 3366 7098
rect 3418 7046 3430 7098
rect 3482 7046 7622 7098
rect 7674 7046 7686 7098
rect 7738 7046 7750 7098
rect 7802 7046 7814 7098
rect 7866 7046 7878 7098
rect 7930 7046 12070 7098
rect 12122 7046 12134 7098
rect 12186 7046 12198 7098
rect 12250 7046 12262 7098
rect 12314 7046 12326 7098
rect 12378 7046 16518 7098
rect 16570 7046 16582 7098
rect 16634 7046 16646 7098
rect 16698 7046 16710 7098
rect 16762 7046 16774 7098
rect 16826 7046 18860 7098
rect 1104 7024 18860 7046
rect 2777 6987 2835 6993
rect 2777 6953 2789 6987
rect 2823 6984 2835 6987
rect 3326 6984 3332 6996
rect 2823 6956 3332 6984
rect 2823 6953 2835 6956
rect 2777 6947 2835 6953
rect 3326 6944 3332 6956
rect 3384 6944 3390 6996
rect 3605 6987 3663 6993
rect 3605 6953 3617 6987
rect 3651 6984 3663 6987
rect 3694 6984 3700 6996
rect 3651 6956 3700 6984
rect 3651 6953 3663 6956
rect 3605 6947 3663 6953
rect 3694 6944 3700 6956
rect 3752 6944 3758 6996
rect 4246 6944 4252 6996
rect 4304 6984 4310 6996
rect 4893 6987 4951 6993
rect 4304 6956 4384 6984
rect 4304 6944 4310 6956
rect 4356 6916 4384 6956
rect 4893 6953 4905 6987
rect 4939 6984 4951 6987
rect 4982 6984 4988 6996
rect 4939 6956 4988 6984
rect 4939 6953 4951 6956
rect 4893 6947 4951 6953
rect 4982 6944 4988 6956
rect 5040 6944 5046 6996
rect 5721 6987 5779 6993
rect 5721 6953 5733 6987
rect 5767 6984 5779 6987
rect 5810 6984 5816 6996
rect 5767 6956 5816 6984
rect 5767 6953 5779 6956
rect 5721 6947 5779 6953
rect 5810 6944 5816 6956
rect 5868 6944 5874 6996
rect 6454 6944 6460 6996
rect 6512 6984 6518 6996
rect 6917 6987 6975 6993
rect 6917 6984 6929 6987
rect 6512 6956 6929 6984
rect 6512 6944 6518 6956
rect 6917 6953 6929 6956
rect 6963 6953 6975 6987
rect 6917 6947 6975 6953
rect 7466 6944 7472 6996
rect 7524 6984 7530 6996
rect 7929 6987 7987 6993
rect 7929 6984 7941 6987
rect 7524 6956 7941 6984
rect 7524 6944 7530 6956
rect 7929 6953 7941 6956
rect 7975 6953 7987 6987
rect 9490 6984 9496 6996
rect 9451 6956 9496 6984
rect 7929 6947 7987 6953
rect 9490 6944 9496 6956
rect 9548 6944 9554 6996
rect 11422 6984 11428 6996
rect 11383 6956 11428 6984
rect 11422 6944 11428 6956
rect 11480 6944 11486 6996
rect 11514 6944 11520 6996
rect 11572 6984 11578 6996
rect 11698 6984 11704 6996
rect 11572 6956 11704 6984
rect 11572 6944 11578 6956
rect 11698 6944 11704 6956
rect 11756 6944 11762 6996
rect 12986 6944 12992 6996
rect 13044 6984 13050 6996
rect 15930 6984 15936 6996
rect 13044 6956 15936 6984
rect 13044 6944 13050 6956
rect 15930 6944 15936 6956
rect 15988 6944 15994 6996
rect 16669 6987 16727 6993
rect 16669 6953 16681 6987
rect 16715 6984 16727 6987
rect 16850 6984 16856 6996
rect 16715 6956 16856 6984
rect 16715 6953 16727 6956
rect 16669 6947 16727 6953
rect 16850 6944 16856 6956
rect 16908 6944 16914 6996
rect 17126 6944 17132 6996
rect 17184 6984 17190 6996
rect 17497 6987 17555 6993
rect 17497 6984 17509 6987
rect 17184 6956 17509 6984
rect 17184 6944 17190 6956
rect 17497 6953 17509 6956
rect 17543 6953 17555 6987
rect 18046 6984 18052 6996
rect 17497 6947 17555 6953
rect 17972 6956 18052 6984
rect 5258 6916 5264 6928
rect 3068 6888 4292 6916
rect 4356 6888 5264 6916
rect 3068 6857 3096 6888
rect 2225 6851 2283 6857
rect 2225 6817 2237 6851
rect 2271 6848 2283 6851
rect 3053 6851 3111 6857
rect 3053 6848 3065 6851
rect 2271 6820 3065 6848
rect 2271 6817 2283 6820
rect 2225 6811 2283 6817
rect 3053 6817 3065 6820
rect 3099 6817 3111 6851
rect 3053 6811 3111 6817
rect 3326 6808 3332 6860
rect 3384 6848 3390 6860
rect 4154 6848 4160 6860
rect 3384 6820 4160 6848
rect 3384 6808 3390 6820
rect 4154 6808 4160 6820
rect 4212 6808 4218 6860
rect 4264 6848 4292 6888
rect 5258 6876 5264 6888
rect 5316 6916 5322 6928
rect 7374 6916 7380 6928
rect 5316 6888 7380 6916
rect 5316 6876 5322 6888
rect 4709 6851 4767 6857
rect 4709 6848 4721 6851
rect 4264 6820 4721 6848
rect 4709 6817 4721 6820
rect 4755 6848 4767 6851
rect 4798 6848 4804 6860
rect 4755 6820 4804 6848
rect 4755 6817 4767 6820
rect 4709 6811 4767 6817
rect 4798 6808 4804 6820
rect 4856 6808 4862 6860
rect 4982 6808 4988 6860
rect 5040 6848 5046 6860
rect 5442 6848 5448 6860
rect 5040 6820 5448 6848
rect 5040 6808 5046 6820
rect 5442 6808 5448 6820
rect 5500 6808 5506 6860
rect 5552 6857 5580 6888
rect 7374 6876 7380 6888
rect 7432 6876 7438 6928
rect 8662 6916 8668 6928
rect 8588 6888 8668 6916
rect 5537 6851 5595 6857
rect 5537 6817 5549 6851
rect 5583 6817 5595 6851
rect 5537 6811 5595 6817
rect 5718 6808 5724 6860
rect 5776 6848 5782 6860
rect 6365 6851 6423 6857
rect 6365 6848 6377 6851
rect 5776 6820 6377 6848
rect 5776 6808 5782 6820
rect 6365 6817 6377 6820
rect 6411 6848 6423 6851
rect 7742 6848 7748 6860
rect 6411 6820 7604 6848
rect 7703 6820 7748 6848
rect 6411 6817 6423 6820
rect 6365 6811 6423 6817
rect 1673 6783 1731 6789
rect 1673 6749 1685 6783
rect 1719 6749 1731 6783
rect 1673 6743 1731 6749
rect 1949 6783 2007 6789
rect 1949 6749 1961 6783
rect 1995 6780 2007 6783
rect 2130 6780 2136 6792
rect 1995 6752 2136 6780
rect 1995 6749 2007 6752
rect 1949 6743 2007 6749
rect 1688 6712 1716 6743
rect 2130 6740 2136 6752
rect 2188 6740 2194 6792
rect 2406 6780 2412 6792
rect 2367 6752 2412 6780
rect 2406 6740 2412 6752
rect 2464 6740 2470 6792
rect 3970 6780 3976 6792
rect 2746 6752 3832 6780
rect 3931 6752 3976 6780
rect 2746 6712 2774 6752
rect 3237 6715 3295 6721
rect 3237 6712 3249 6715
rect 1688 6684 2774 6712
rect 3068 6684 3249 6712
rect 1486 6644 1492 6656
rect 1447 6616 1492 6644
rect 1486 6604 1492 6616
rect 1544 6604 1550 6656
rect 1762 6644 1768 6656
rect 1723 6616 1768 6644
rect 1762 6604 1768 6616
rect 1820 6604 1826 6656
rect 2314 6644 2320 6656
rect 2275 6616 2320 6644
rect 2314 6604 2320 6616
rect 2372 6604 2378 6656
rect 2590 6604 2596 6656
rect 2648 6644 2654 6656
rect 3068 6644 3096 6684
rect 3237 6681 3249 6684
rect 3283 6712 3295 6715
rect 3418 6712 3424 6724
rect 3283 6684 3424 6712
rect 3283 6681 3295 6684
rect 3237 6675 3295 6681
rect 3418 6672 3424 6684
rect 3476 6672 3482 6724
rect 2648 6616 3096 6644
rect 3145 6647 3203 6653
rect 2648 6604 2654 6616
rect 3145 6613 3157 6647
rect 3191 6644 3203 6647
rect 3694 6644 3700 6656
rect 3191 6616 3700 6644
rect 3191 6613 3203 6616
rect 3145 6607 3203 6613
rect 3694 6604 3700 6616
rect 3752 6604 3758 6656
rect 3804 6653 3832 6752
rect 3970 6740 3976 6752
rect 4028 6740 4034 6792
rect 4062 6740 4068 6792
rect 4120 6740 4126 6792
rect 4430 6780 4436 6792
rect 4391 6752 4436 6780
rect 4430 6740 4436 6752
rect 4488 6740 4494 6792
rect 4525 6783 4583 6789
rect 4525 6749 4537 6783
rect 4571 6780 4583 6783
rect 6730 6780 6736 6792
rect 4571 6752 6736 6780
rect 4571 6749 4583 6752
rect 4525 6743 4583 6749
rect 6730 6740 6736 6752
rect 6788 6740 6794 6792
rect 6914 6740 6920 6792
rect 6972 6780 6978 6792
rect 7469 6783 7527 6789
rect 7469 6780 7481 6783
rect 6972 6752 7481 6780
rect 6972 6740 6978 6752
rect 7469 6749 7481 6752
rect 7515 6749 7527 6783
rect 7576 6780 7604 6820
rect 7742 6808 7748 6820
rect 7800 6808 7806 6860
rect 8588 6857 8616 6888
rect 8662 6876 8668 6888
rect 8720 6876 8726 6928
rect 12710 6916 12716 6928
rect 10888 6888 12020 6916
rect 10888 6860 10916 6888
rect 8573 6851 8631 6857
rect 8573 6817 8585 6851
rect 8619 6817 8631 6851
rect 8573 6811 8631 6817
rect 8754 6808 8760 6860
rect 8812 6848 8818 6860
rect 9953 6851 10011 6857
rect 9953 6848 9965 6851
rect 8812 6820 9965 6848
rect 8812 6808 8818 6820
rect 9953 6817 9965 6820
rect 9999 6817 10011 6851
rect 10134 6848 10140 6860
rect 10095 6820 10140 6848
rect 9953 6811 10011 6817
rect 10134 6808 10140 6820
rect 10192 6808 10198 6860
rect 10870 6848 10876 6860
rect 10831 6820 10876 6848
rect 10870 6808 10876 6820
rect 10928 6808 10934 6860
rect 10980 6820 11284 6848
rect 7834 6780 7840 6792
rect 7576 6752 7840 6780
rect 7469 6743 7527 6749
rect 7834 6740 7840 6752
rect 7892 6740 7898 6792
rect 8294 6780 8300 6792
rect 8255 6752 8300 6780
rect 8294 6740 8300 6752
rect 8352 6740 8358 6792
rect 8389 6783 8447 6789
rect 8389 6749 8401 6783
rect 8435 6780 8447 6783
rect 8938 6780 8944 6792
rect 8435 6752 8944 6780
rect 8435 6749 8447 6752
rect 8389 6743 8447 6749
rect 4080 6712 4108 6740
rect 5353 6715 5411 6721
rect 5353 6712 5365 6715
rect 4080 6684 5365 6712
rect 5353 6681 5365 6684
rect 5399 6712 5411 6715
rect 5399 6684 6592 6712
rect 5399 6681 5411 6684
rect 5353 6675 5411 6681
rect 3789 6647 3847 6653
rect 3789 6613 3801 6647
rect 3835 6613 3847 6647
rect 3789 6607 3847 6613
rect 4065 6647 4123 6653
rect 4065 6613 4077 6647
rect 4111 6644 4123 6647
rect 4154 6644 4160 6656
rect 4111 6616 4160 6644
rect 4111 6613 4123 6616
rect 4065 6607 4123 6613
rect 4154 6604 4160 6616
rect 4212 6604 4218 6656
rect 5258 6644 5264 6656
rect 5219 6616 5264 6644
rect 5258 6604 5264 6616
rect 5316 6604 5322 6656
rect 5442 6604 5448 6656
rect 5500 6644 5506 6656
rect 6089 6647 6147 6653
rect 6089 6644 6101 6647
rect 5500 6616 6101 6644
rect 5500 6604 5506 6616
rect 6089 6613 6101 6616
rect 6135 6613 6147 6647
rect 6089 6607 6147 6613
rect 6181 6647 6239 6653
rect 6181 6613 6193 6647
rect 6227 6644 6239 6647
rect 6454 6644 6460 6656
rect 6227 6616 6460 6644
rect 6227 6613 6239 6616
rect 6181 6607 6239 6613
rect 6454 6604 6460 6616
rect 6512 6604 6518 6656
rect 6564 6653 6592 6684
rect 6549 6647 6607 6653
rect 6549 6613 6561 6647
rect 6595 6613 6607 6647
rect 7098 6644 7104 6656
rect 7059 6616 7104 6644
rect 6549 6607 6607 6613
rect 7098 6604 7104 6616
rect 7156 6604 7162 6656
rect 7561 6647 7619 6653
rect 7561 6613 7573 6647
rect 7607 6644 7619 6647
rect 8018 6644 8024 6656
rect 7607 6616 8024 6644
rect 7607 6613 7619 6616
rect 7561 6607 7619 6613
rect 8018 6604 8024 6616
rect 8076 6644 8082 6656
rect 8404 6644 8432 6743
rect 8938 6740 8944 6752
rect 8996 6740 9002 6792
rect 9122 6740 9128 6792
rect 9180 6780 9186 6792
rect 9309 6783 9367 6789
rect 9309 6780 9321 6783
rect 9180 6752 9321 6780
rect 9180 6740 9186 6752
rect 9309 6749 9321 6752
rect 9355 6780 9367 6783
rect 9582 6780 9588 6792
rect 9355 6752 9588 6780
rect 9355 6749 9367 6752
rect 9309 6743 9367 6749
rect 9582 6740 9588 6752
rect 9640 6740 9646 6792
rect 9858 6780 9864 6792
rect 9819 6752 9864 6780
rect 9858 6740 9864 6752
rect 9916 6740 9922 6792
rect 10502 6740 10508 6792
rect 10560 6780 10566 6792
rect 10980 6780 11008 6820
rect 11146 6780 11152 6792
rect 10560 6752 11008 6780
rect 11107 6752 11152 6780
rect 10560 6740 10566 6752
rect 11146 6740 11152 6752
rect 11204 6740 11210 6792
rect 11256 6780 11284 6820
rect 11698 6808 11704 6860
rect 11756 6848 11762 6860
rect 11882 6848 11888 6860
rect 11756 6820 11888 6848
rect 11756 6808 11762 6820
rect 11882 6808 11888 6820
rect 11940 6808 11946 6860
rect 11992 6857 12020 6888
rect 12544 6888 12716 6916
rect 11977 6851 12035 6857
rect 11977 6817 11989 6851
rect 12023 6817 12035 6851
rect 11977 6811 12035 6817
rect 12434 6808 12440 6860
rect 12492 6808 12498 6860
rect 12452 6780 12480 6808
rect 11256 6752 12480 6780
rect 8956 6712 8984 6740
rect 10781 6715 10839 6721
rect 8956 6684 9168 6712
rect 9140 6656 9168 6684
rect 10781 6681 10793 6715
rect 10827 6712 10839 6715
rect 12544 6712 12572 6888
rect 12710 6876 12716 6888
rect 12768 6876 12774 6928
rect 13446 6876 13452 6928
rect 13504 6916 13510 6928
rect 13504 6888 13676 6916
rect 13504 6876 13510 6888
rect 12802 6848 12808 6860
rect 12763 6820 12808 6848
rect 12802 6808 12808 6820
rect 12860 6808 12866 6860
rect 13648 6857 13676 6888
rect 14734 6876 14740 6928
rect 14792 6916 14798 6928
rect 17862 6916 17868 6928
rect 14792 6888 17868 6916
rect 14792 6876 14798 6888
rect 17862 6876 17868 6888
rect 17920 6876 17926 6928
rect 13633 6851 13691 6857
rect 13633 6817 13645 6851
rect 13679 6817 13691 6851
rect 13633 6811 13691 6817
rect 14369 6851 14427 6857
rect 14369 6817 14381 6851
rect 14415 6848 14427 6851
rect 14918 6848 14924 6860
rect 14415 6820 14924 6848
rect 14415 6817 14427 6820
rect 14369 6811 14427 6817
rect 14918 6808 14924 6820
rect 14976 6808 14982 6860
rect 15010 6808 15016 6860
rect 15068 6848 15074 6860
rect 15105 6851 15163 6857
rect 15105 6848 15117 6851
rect 15068 6820 15117 6848
rect 15068 6808 15074 6820
rect 15105 6817 15117 6820
rect 15151 6817 15163 6851
rect 15105 6811 15163 6817
rect 16114 6808 16120 6860
rect 16172 6848 16178 6860
rect 16301 6851 16359 6857
rect 16301 6848 16313 6851
rect 16172 6820 16313 6848
rect 16172 6808 16178 6820
rect 16301 6817 16313 6820
rect 16347 6817 16359 6851
rect 16301 6811 16359 6817
rect 16485 6851 16543 6857
rect 16485 6817 16497 6851
rect 16531 6848 16543 6851
rect 16850 6848 16856 6860
rect 16531 6820 16856 6848
rect 16531 6817 16543 6820
rect 16485 6811 16543 6817
rect 16850 6808 16856 6820
rect 16908 6848 16914 6860
rect 17034 6848 17040 6860
rect 16908 6820 17040 6848
rect 16908 6808 16914 6820
rect 17034 6808 17040 6820
rect 17092 6808 17098 6860
rect 17221 6851 17279 6857
rect 17221 6817 17233 6851
rect 17267 6817 17279 6851
rect 17221 6811 17279 6817
rect 13449 6783 13507 6789
rect 13449 6749 13461 6783
rect 13495 6780 13507 6783
rect 13538 6780 13544 6792
rect 13495 6752 13544 6780
rect 13495 6749 13507 6752
rect 13449 6743 13507 6749
rect 13538 6740 13544 6752
rect 13596 6740 13602 6792
rect 14461 6783 14519 6789
rect 14461 6749 14473 6783
rect 14507 6780 14519 6783
rect 15194 6780 15200 6792
rect 14507 6752 15200 6780
rect 14507 6749 14519 6752
rect 14461 6743 14519 6749
rect 15194 6740 15200 6752
rect 15252 6740 15258 6792
rect 15930 6740 15936 6792
rect 15988 6780 15994 6792
rect 16206 6780 16212 6792
rect 15988 6752 16212 6780
rect 15988 6740 15994 6752
rect 16206 6740 16212 6752
rect 16264 6740 16270 6792
rect 16666 6740 16672 6792
rect 16724 6780 16730 6792
rect 16942 6780 16948 6792
rect 16724 6752 16948 6780
rect 16724 6740 16730 6752
rect 16942 6740 16948 6752
rect 17000 6780 17006 6792
rect 17236 6780 17264 6811
rect 17310 6808 17316 6860
rect 17368 6848 17374 6860
rect 17972 6857 18000 6956
rect 18046 6944 18052 6956
rect 18104 6944 18110 6996
rect 18138 6944 18144 6996
rect 18196 6944 18202 6996
rect 18156 6857 18184 6944
rect 17957 6851 18015 6857
rect 17957 6848 17969 6851
rect 17368 6820 17969 6848
rect 17368 6808 17374 6820
rect 17957 6817 17969 6820
rect 18003 6817 18015 6851
rect 17957 6811 18015 6817
rect 18141 6851 18199 6857
rect 18141 6817 18153 6851
rect 18187 6817 18199 6851
rect 18141 6811 18199 6817
rect 17000 6752 17264 6780
rect 17000 6740 17006 6752
rect 17586 6740 17592 6792
rect 17644 6780 17650 6792
rect 18156 6780 18184 6811
rect 18506 6780 18512 6792
rect 17644 6752 18184 6780
rect 18467 6752 18512 6780
rect 17644 6740 17650 6752
rect 18506 6740 18512 6752
rect 18564 6740 18570 6792
rect 12621 6715 12679 6721
rect 12621 6712 12633 6715
rect 10827 6684 12296 6712
rect 12544 6684 12633 6712
rect 10827 6681 10839 6684
rect 10781 6675 10839 6681
rect 8938 6644 8944 6656
rect 8076 6616 8432 6644
rect 8899 6616 8944 6644
rect 8076 6604 8082 6616
rect 8938 6604 8944 6616
rect 8996 6604 9002 6656
rect 9122 6604 9128 6656
rect 9180 6604 9186 6656
rect 10318 6644 10324 6656
rect 10279 6616 10324 6644
rect 10318 6604 10324 6616
rect 10376 6604 10382 6656
rect 10689 6647 10747 6653
rect 10689 6613 10701 6647
rect 10735 6644 10747 6647
rect 10870 6644 10876 6656
rect 10735 6616 10876 6644
rect 10735 6613 10747 6616
rect 10689 6607 10747 6613
rect 10870 6604 10876 6616
rect 10928 6604 10934 6656
rect 11146 6604 11152 6656
rect 11204 6644 11210 6656
rect 11333 6647 11391 6653
rect 11333 6644 11345 6647
rect 11204 6616 11345 6644
rect 11204 6604 11210 6616
rect 11333 6613 11345 6616
rect 11379 6613 11391 6647
rect 11333 6607 11391 6613
rect 11793 6647 11851 6653
rect 11793 6613 11805 6647
rect 11839 6644 11851 6647
rect 11974 6644 11980 6656
rect 11839 6616 11980 6644
rect 11839 6613 11851 6616
rect 11793 6607 11851 6613
rect 11974 6604 11980 6616
rect 12032 6604 12038 6656
rect 12268 6653 12296 6684
rect 12621 6681 12633 6684
rect 12667 6681 12679 6715
rect 12621 6675 12679 6681
rect 12713 6715 12771 6721
rect 12713 6681 12725 6715
rect 12759 6712 12771 6715
rect 13814 6712 13820 6724
rect 12759 6684 13820 6712
rect 12759 6681 12771 6684
rect 12713 6675 12771 6681
rect 12253 6647 12311 6653
rect 12253 6613 12265 6647
rect 12299 6613 12311 6647
rect 12253 6607 12311 6613
rect 12434 6604 12440 6656
rect 12492 6644 12498 6656
rect 12728 6644 12756 6675
rect 13814 6672 13820 6684
rect 13872 6672 13878 6724
rect 14550 6712 14556 6724
rect 14511 6684 14556 6712
rect 14550 6672 14556 6684
rect 14608 6672 14614 6724
rect 15289 6715 15347 6721
rect 15289 6681 15301 6715
rect 15335 6712 15347 6715
rect 15335 6684 15884 6712
rect 15335 6681 15347 6684
rect 15289 6675 15347 6681
rect 12492 6616 12756 6644
rect 12492 6604 12498 6616
rect 12802 6604 12808 6656
rect 12860 6644 12866 6656
rect 13081 6647 13139 6653
rect 13081 6644 13093 6647
rect 12860 6616 13093 6644
rect 12860 6604 12866 6616
rect 13081 6613 13093 6616
rect 13127 6613 13139 6647
rect 13081 6607 13139 6613
rect 13541 6647 13599 6653
rect 13541 6613 13553 6647
rect 13587 6644 13599 6647
rect 13630 6644 13636 6656
rect 13587 6616 13636 6644
rect 13587 6613 13599 6616
rect 13541 6607 13599 6613
rect 13630 6604 13636 6616
rect 13688 6604 13694 6656
rect 13906 6604 13912 6656
rect 13964 6644 13970 6656
rect 14826 6644 14832 6656
rect 13964 6616 14832 6644
rect 13964 6604 13970 6616
rect 14826 6604 14832 6616
rect 14884 6604 14890 6656
rect 14921 6647 14979 6653
rect 14921 6613 14933 6647
rect 14967 6644 14979 6647
rect 15010 6644 15016 6656
rect 14967 6616 15016 6644
rect 14967 6613 14979 6616
rect 14921 6607 14979 6613
rect 15010 6604 15016 6616
rect 15068 6604 15074 6656
rect 15378 6644 15384 6656
rect 15339 6616 15384 6644
rect 15378 6604 15384 6616
rect 15436 6604 15442 6656
rect 15746 6644 15752 6656
rect 15707 6616 15752 6644
rect 15746 6604 15752 6616
rect 15804 6604 15810 6656
rect 15856 6653 15884 6684
rect 16114 6672 16120 6724
rect 16172 6712 16178 6724
rect 17034 6712 17040 6724
rect 16172 6684 16436 6712
rect 16995 6684 17040 6712
rect 16172 6672 16178 6684
rect 15841 6647 15899 6653
rect 15841 6613 15853 6647
rect 15887 6613 15899 6647
rect 16408 6644 16436 6684
rect 17034 6672 17040 6684
rect 17092 6712 17098 6724
rect 18598 6712 18604 6724
rect 17092 6684 18604 6712
rect 17092 6672 17098 6684
rect 18598 6672 18604 6684
rect 18656 6672 18662 6724
rect 17129 6647 17187 6653
rect 17129 6644 17141 6647
rect 16408 6616 17141 6644
rect 15841 6607 15899 6613
rect 17129 6613 17141 6616
rect 17175 6613 17187 6647
rect 17129 6607 17187 6613
rect 17678 6604 17684 6656
rect 17736 6644 17742 6656
rect 17865 6647 17923 6653
rect 17865 6644 17877 6647
rect 17736 6616 17877 6644
rect 17736 6604 17742 6616
rect 17865 6613 17877 6616
rect 17911 6613 17923 6647
rect 17865 6607 17923 6613
rect 18046 6604 18052 6656
rect 18104 6644 18110 6656
rect 18325 6647 18383 6653
rect 18325 6644 18337 6647
rect 18104 6616 18337 6644
rect 18104 6604 18110 6616
rect 18325 6613 18337 6616
rect 18371 6613 18383 6647
rect 18325 6607 18383 6613
rect 1104 6554 18860 6576
rect 1104 6502 5398 6554
rect 5450 6502 5462 6554
rect 5514 6502 5526 6554
rect 5578 6502 5590 6554
rect 5642 6502 5654 6554
rect 5706 6502 9846 6554
rect 9898 6502 9910 6554
rect 9962 6502 9974 6554
rect 10026 6502 10038 6554
rect 10090 6502 10102 6554
rect 10154 6502 14294 6554
rect 14346 6502 14358 6554
rect 14410 6502 14422 6554
rect 14474 6502 14486 6554
rect 14538 6502 14550 6554
rect 14602 6502 18860 6554
rect 1104 6480 18860 6502
rect 1946 6400 1952 6452
rect 2004 6440 2010 6452
rect 2225 6443 2283 6449
rect 2225 6440 2237 6443
rect 2004 6412 2237 6440
rect 2004 6400 2010 6412
rect 2225 6409 2237 6412
rect 2271 6409 2283 6443
rect 2406 6440 2412 6452
rect 2367 6412 2412 6440
rect 2225 6403 2283 6409
rect 2406 6400 2412 6412
rect 2464 6400 2470 6452
rect 2958 6400 2964 6452
rect 3016 6440 3022 6452
rect 3142 6440 3148 6452
rect 3016 6412 3148 6440
rect 3016 6400 3022 6412
rect 3142 6400 3148 6412
rect 3200 6400 3206 6452
rect 3237 6443 3295 6449
rect 3237 6409 3249 6443
rect 3283 6440 3295 6443
rect 3789 6443 3847 6449
rect 3789 6440 3801 6443
rect 3283 6412 3801 6440
rect 3283 6409 3295 6412
rect 3237 6403 3295 6409
rect 3789 6409 3801 6412
rect 3835 6409 3847 6443
rect 4154 6440 4160 6452
rect 4115 6412 4160 6440
rect 3789 6403 3847 6409
rect 4154 6400 4160 6412
rect 4212 6400 4218 6452
rect 4249 6443 4307 6449
rect 4249 6409 4261 6443
rect 4295 6440 4307 6443
rect 4617 6443 4675 6449
rect 4617 6440 4629 6443
rect 4295 6412 4629 6440
rect 4295 6409 4307 6412
rect 4249 6403 4307 6409
rect 4617 6409 4629 6412
rect 4663 6409 4675 6443
rect 4617 6403 4675 6409
rect 4706 6400 4712 6452
rect 4764 6440 4770 6452
rect 5077 6443 5135 6449
rect 5077 6440 5089 6443
rect 4764 6412 5089 6440
rect 4764 6400 4770 6412
rect 5077 6409 5089 6412
rect 5123 6409 5135 6443
rect 5810 6440 5816 6452
rect 5771 6412 5816 6440
rect 5077 6403 5135 6409
rect 5810 6400 5816 6412
rect 5868 6400 5874 6452
rect 6178 6440 6184 6452
rect 6139 6412 6184 6440
rect 6178 6400 6184 6412
rect 6236 6400 6242 6452
rect 6638 6400 6644 6452
rect 6696 6440 6702 6452
rect 6696 6412 6776 6440
rect 6696 6400 6702 6412
rect 1765 6375 1823 6381
rect 1765 6341 1777 6375
rect 1811 6372 1823 6375
rect 2038 6372 2044 6384
rect 1811 6344 2044 6372
rect 1811 6341 1823 6344
rect 1765 6335 1823 6341
rect 2038 6332 2044 6344
rect 2096 6332 2102 6384
rect 3329 6375 3387 6381
rect 3329 6341 3341 6375
rect 3375 6372 3387 6375
rect 3510 6372 3516 6384
rect 3375 6344 3516 6372
rect 3375 6341 3387 6344
rect 3329 6335 3387 6341
rect 3510 6332 3516 6344
rect 3568 6332 3574 6384
rect 4430 6372 4436 6384
rect 4172 6344 4436 6372
rect 1857 6307 1915 6313
rect 1857 6273 1869 6307
rect 1903 6304 1915 6307
rect 1946 6304 1952 6316
rect 1903 6276 1952 6304
rect 1903 6273 1915 6276
rect 1857 6267 1915 6273
rect 1946 6264 1952 6276
rect 2004 6264 2010 6316
rect 2593 6307 2651 6313
rect 2593 6273 2605 6307
rect 2639 6273 2651 6307
rect 2593 6267 2651 6273
rect 1673 6239 1731 6245
rect 1673 6205 1685 6239
rect 1719 6236 1731 6239
rect 2222 6236 2228 6248
rect 1719 6208 2228 6236
rect 1719 6205 1731 6208
rect 1673 6199 1731 6205
rect 2222 6196 2228 6208
rect 2280 6196 2286 6248
rect 2608 6180 2636 6267
rect 2682 6264 2688 6316
rect 2740 6304 2746 6316
rect 2740 6276 2785 6304
rect 2740 6264 2746 6276
rect 2866 6264 2872 6316
rect 2924 6304 2930 6316
rect 4172 6304 4200 6344
rect 4430 6332 4436 6344
rect 4488 6332 4494 6384
rect 4985 6375 5043 6381
rect 4985 6341 4997 6375
rect 5031 6372 5043 6375
rect 5166 6372 5172 6384
rect 5031 6344 5172 6372
rect 5031 6341 5043 6344
rect 4985 6335 5043 6341
rect 5166 6332 5172 6344
rect 5224 6372 5230 6384
rect 6748 6372 6776 6412
rect 6822 6400 6828 6452
rect 6880 6440 6886 6452
rect 8021 6443 8079 6449
rect 6880 6412 6925 6440
rect 6880 6400 6886 6412
rect 8021 6409 8033 6443
rect 8067 6440 8079 6443
rect 8938 6440 8944 6452
rect 8067 6412 8944 6440
rect 8067 6409 8079 6412
rect 8021 6403 8079 6409
rect 8938 6400 8944 6412
rect 8996 6400 9002 6452
rect 9217 6443 9275 6449
rect 9217 6409 9229 6443
rect 9263 6440 9275 6443
rect 9585 6443 9643 6449
rect 9585 6440 9597 6443
rect 9263 6412 9597 6440
rect 9263 6409 9275 6412
rect 9217 6403 9275 6409
rect 9585 6409 9597 6412
rect 9631 6409 9643 6443
rect 9585 6403 9643 6409
rect 9677 6443 9735 6449
rect 9677 6409 9689 6443
rect 9723 6440 9735 6443
rect 10318 6440 10324 6452
rect 9723 6412 10324 6440
rect 9723 6409 9735 6412
rect 9677 6403 9735 6409
rect 10318 6400 10324 6412
rect 10376 6400 10382 6452
rect 10459 6443 10517 6449
rect 10459 6409 10471 6443
rect 10505 6440 10517 6443
rect 13541 6443 13599 6449
rect 10505 6412 13492 6440
rect 10505 6409 10517 6412
rect 10459 6403 10517 6409
rect 7193 6375 7251 6381
rect 7193 6372 7205 6375
rect 5224 6344 5488 6372
rect 6748 6344 7205 6372
rect 5224 6332 5230 6344
rect 5460 6316 5488 6344
rect 7193 6341 7205 6344
rect 7239 6341 7251 6375
rect 7193 6335 7251 6341
rect 7285 6375 7343 6381
rect 7285 6341 7297 6375
rect 7331 6372 7343 6375
rect 7466 6372 7472 6384
rect 7331 6344 7472 6372
rect 7331 6341 7343 6344
rect 7285 6335 7343 6341
rect 7466 6332 7472 6344
rect 7524 6332 7530 6384
rect 9950 6332 9956 6384
rect 10008 6372 10014 6384
rect 10962 6372 10968 6384
rect 10008 6344 10968 6372
rect 10008 6332 10014 6344
rect 10962 6332 10968 6344
rect 11020 6332 11026 6384
rect 11422 6332 11428 6384
rect 11480 6372 11486 6384
rect 13464 6372 13492 6412
rect 13541 6409 13553 6443
rect 13587 6440 13599 6443
rect 14001 6443 14059 6449
rect 14001 6440 14013 6443
rect 13587 6412 14013 6440
rect 13587 6409 13599 6412
rect 13541 6403 13599 6409
rect 14001 6409 14013 6412
rect 14047 6409 14059 6443
rect 14001 6403 14059 6409
rect 14274 6400 14280 6452
rect 14332 6440 14338 6452
rect 14461 6443 14519 6449
rect 14461 6440 14473 6443
rect 14332 6412 14473 6440
rect 14332 6400 14338 6412
rect 14461 6409 14473 6412
rect 14507 6440 14519 6443
rect 14734 6440 14740 6452
rect 14507 6412 14740 6440
rect 14507 6409 14519 6412
rect 14461 6403 14519 6409
rect 14734 6400 14740 6412
rect 14792 6400 14798 6452
rect 15194 6440 15200 6452
rect 15107 6412 15200 6440
rect 15194 6400 15200 6412
rect 15252 6440 15258 6452
rect 15654 6440 15660 6452
rect 15252 6412 15660 6440
rect 15252 6400 15258 6412
rect 15654 6400 15660 6412
rect 15712 6400 15718 6452
rect 15746 6400 15752 6452
rect 15804 6440 15810 6452
rect 16025 6443 16083 6449
rect 16025 6440 16037 6443
rect 15804 6412 16037 6440
rect 15804 6400 15810 6412
rect 16025 6409 16037 6412
rect 16071 6409 16083 6443
rect 16025 6403 16083 6409
rect 17402 6400 17408 6452
rect 17460 6440 17466 6452
rect 17460 6412 17505 6440
rect 17460 6400 17466 6412
rect 11480 6344 13400 6372
rect 13464 6344 14780 6372
rect 11480 6332 11486 6344
rect 2924 6276 4200 6304
rect 2924 6264 2930 6276
rect 3528 6248 3556 6276
rect 4246 6264 4252 6316
rect 4304 6304 4310 6316
rect 5074 6304 5080 6316
rect 4304 6276 5080 6304
rect 4304 6264 4310 6276
rect 5074 6264 5080 6276
rect 5132 6264 5138 6316
rect 5442 6264 5448 6316
rect 5500 6264 5506 6316
rect 6362 6304 6368 6316
rect 5552 6276 6368 6304
rect 3145 6239 3203 6245
rect 3145 6205 3157 6239
rect 3191 6236 3203 6239
rect 3326 6236 3332 6248
rect 3191 6208 3332 6236
rect 3191 6205 3203 6208
rect 3145 6199 3203 6205
rect 3326 6196 3332 6208
rect 3384 6196 3390 6248
rect 3510 6196 3516 6248
rect 3568 6196 3574 6248
rect 3694 6196 3700 6248
rect 3752 6236 3758 6248
rect 4338 6236 4344 6248
rect 3752 6208 3924 6236
rect 4299 6208 4344 6236
rect 3752 6196 3758 6208
rect 2590 6128 2596 6180
rect 2648 6128 2654 6180
rect 3234 6128 3240 6180
rect 3292 6168 3298 6180
rect 3786 6168 3792 6180
rect 3292 6140 3792 6168
rect 3292 6128 3298 6140
rect 3786 6128 3792 6140
rect 3844 6128 3850 6180
rect 2866 6100 2872 6112
rect 2827 6072 2872 6100
rect 2866 6060 2872 6072
rect 2924 6060 2930 6112
rect 3694 6100 3700 6112
rect 3655 6072 3700 6100
rect 3694 6060 3700 6072
rect 3752 6060 3758 6112
rect 3896 6100 3924 6208
rect 4338 6196 4344 6208
rect 4396 6196 4402 6248
rect 4798 6196 4804 6248
rect 4856 6236 4862 6248
rect 5552 6245 5580 6276
rect 6362 6264 6368 6276
rect 6420 6264 6426 6316
rect 8478 6304 8484 6316
rect 6472 6276 8484 6304
rect 5169 6239 5227 6245
rect 5169 6236 5181 6239
rect 4856 6208 5181 6236
rect 4856 6196 4862 6208
rect 5169 6205 5181 6208
rect 5215 6205 5227 6239
rect 5169 6199 5227 6205
rect 5537 6239 5595 6245
rect 5537 6205 5549 6239
rect 5583 6205 5595 6239
rect 5537 6199 5595 6205
rect 5626 6196 5632 6248
rect 5684 6236 5690 6248
rect 5721 6239 5779 6245
rect 5721 6236 5733 6239
rect 5684 6208 5733 6236
rect 5684 6196 5690 6208
rect 5721 6205 5733 6208
rect 5767 6205 5779 6239
rect 5721 6199 5779 6205
rect 3970 6128 3976 6180
rect 4028 6168 4034 6180
rect 6472 6168 6500 6276
rect 8478 6264 8484 6276
rect 8536 6264 8542 6316
rect 8846 6304 8852 6316
rect 8807 6276 8852 6304
rect 8846 6264 8852 6276
rect 8904 6264 8910 6316
rect 9398 6264 9404 6316
rect 9456 6304 9462 6316
rect 10229 6307 10287 6313
rect 10229 6304 10241 6307
rect 9456 6276 10241 6304
rect 9456 6264 9462 6276
rect 10229 6273 10241 6276
rect 10275 6273 10287 6307
rect 10229 6267 10287 6273
rect 10686 6264 10692 6316
rect 10744 6304 10750 6316
rect 11330 6304 11336 6316
rect 10744 6276 11336 6304
rect 10744 6264 10750 6276
rect 11330 6264 11336 6276
rect 11388 6264 11394 6316
rect 11882 6304 11888 6316
rect 11843 6276 11888 6304
rect 11882 6264 11888 6276
rect 11940 6264 11946 6316
rect 12250 6264 12256 6316
rect 12308 6304 12314 6316
rect 12621 6307 12679 6313
rect 12621 6304 12633 6307
rect 12308 6276 12633 6304
rect 12308 6264 12314 6276
rect 12621 6273 12633 6276
rect 12667 6273 12679 6307
rect 12621 6267 12679 6273
rect 12713 6307 12771 6313
rect 12713 6273 12725 6307
rect 12759 6304 12771 6307
rect 12986 6304 12992 6316
rect 12759 6276 12992 6304
rect 12759 6273 12771 6276
rect 12713 6267 12771 6273
rect 6733 6239 6791 6245
rect 6733 6205 6745 6239
rect 6779 6205 6791 6239
rect 7374 6236 7380 6248
rect 7335 6208 7380 6236
rect 6733 6199 6791 6205
rect 4028 6140 6500 6168
rect 6549 6171 6607 6177
rect 4028 6128 4034 6140
rect 6549 6137 6561 6171
rect 6595 6168 6607 6171
rect 6638 6168 6644 6180
rect 6595 6140 6644 6168
rect 6595 6137 6607 6140
rect 6549 6131 6607 6137
rect 4706 6100 4712 6112
rect 3896 6072 4712 6100
rect 4706 6060 4712 6072
rect 4764 6060 4770 6112
rect 4798 6060 4804 6112
rect 4856 6100 4862 6112
rect 6564 6100 6592 6131
rect 6638 6128 6644 6140
rect 6696 6128 6702 6180
rect 6748 6168 6776 6199
rect 7374 6196 7380 6208
rect 7432 6196 7438 6248
rect 7834 6236 7840 6248
rect 7747 6208 7840 6236
rect 7834 6196 7840 6208
rect 7892 6196 7898 6248
rect 7929 6239 7987 6245
rect 7929 6205 7941 6239
rect 7975 6236 7987 6239
rect 8110 6236 8116 6248
rect 7975 6208 8116 6236
rect 7975 6205 7987 6208
rect 7929 6199 7987 6205
rect 8110 6196 8116 6208
rect 8168 6196 8174 6248
rect 8573 6239 8631 6245
rect 8573 6205 8585 6239
rect 8619 6205 8631 6239
rect 8754 6236 8760 6248
rect 8715 6208 8760 6236
rect 8573 6199 8631 6205
rect 7282 6168 7288 6180
rect 6748 6140 7288 6168
rect 7282 6128 7288 6140
rect 7340 6128 7346 6180
rect 7852 6168 7880 6196
rect 8588 6168 8616 6199
rect 8754 6196 8760 6208
rect 8812 6196 8818 6248
rect 9493 6239 9551 6245
rect 9493 6205 9505 6239
rect 9539 6236 9551 6239
rect 10410 6236 10416 6248
rect 9539 6208 10416 6236
rect 9539 6205 9551 6208
rect 9493 6199 9551 6205
rect 10410 6196 10416 6208
rect 10468 6196 10474 6248
rect 10520 6208 11008 6236
rect 9950 6168 9956 6180
rect 7852 6140 8524 6168
rect 8588 6140 9956 6168
rect 4856 6072 6592 6100
rect 4856 6060 4862 6072
rect 6914 6060 6920 6112
rect 6972 6100 6978 6112
rect 7374 6100 7380 6112
rect 6972 6072 7380 6100
rect 6972 6060 6978 6072
rect 7374 6060 7380 6072
rect 7432 6060 7438 6112
rect 8386 6100 8392 6112
rect 8347 6072 8392 6100
rect 8386 6060 8392 6072
rect 8444 6060 8450 6112
rect 8496 6100 8524 6140
rect 9950 6128 9956 6140
rect 10008 6128 10014 6180
rect 10045 6171 10103 6177
rect 10045 6137 10057 6171
rect 10091 6168 10103 6171
rect 10520 6168 10548 6208
rect 10091 6140 10548 6168
rect 10980 6168 11008 6208
rect 11238 6196 11244 6248
rect 11296 6236 11302 6248
rect 11977 6239 12035 6245
rect 11977 6236 11989 6239
rect 11296 6208 11989 6236
rect 11296 6196 11302 6208
rect 11977 6205 11989 6208
rect 12023 6205 12035 6239
rect 11977 6199 12035 6205
rect 12069 6239 12127 6245
rect 12069 6205 12081 6239
rect 12115 6205 12127 6239
rect 12069 6199 12127 6205
rect 12529 6239 12587 6245
rect 12529 6205 12541 6239
rect 12575 6205 12587 6239
rect 12636 6236 12664 6267
rect 12986 6264 12992 6276
rect 13044 6264 13050 6316
rect 13170 6264 13176 6316
rect 13228 6304 13234 6316
rect 13372 6304 13400 6344
rect 14752 6316 14780 6344
rect 14826 6332 14832 6384
rect 14884 6372 14890 6384
rect 17037 6375 17095 6381
rect 14884 6344 16252 6372
rect 14884 6332 14890 6344
rect 13228 6276 13308 6304
rect 13372 6276 13584 6304
rect 13228 6264 13234 6276
rect 13280 6245 13308 6276
rect 13265 6239 13323 6245
rect 12636 6208 13216 6236
rect 12529 6199 12587 6205
rect 11606 6168 11612 6180
rect 10980 6140 11612 6168
rect 10091 6137 10103 6140
rect 10045 6131 10103 6137
rect 11606 6128 11612 6140
rect 11664 6128 11670 6180
rect 11790 6128 11796 6180
rect 11848 6168 11854 6180
rect 12084 6168 12112 6199
rect 11848 6140 12112 6168
rect 12544 6168 12572 6199
rect 12894 6168 12900 6180
rect 12544 6140 12900 6168
rect 11848 6128 11854 6140
rect 12894 6128 12900 6140
rect 12952 6128 12958 6180
rect 9030 6100 9036 6112
rect 8496 6072 9036 6100
rect 9030 6060 9036 6072
rect 9088 6060 9094 6112
rect 9306 6060 9312 6112
rect 9364 6100 9370 6112
rect 9858 6100 9864 6112
rect 9364 6072 9864 6100
rect 9364 6060 9370 6072
rect 9858 6060 9864 6072
rect 9916 6100 9922 6112
rect 10686 6100 10692 6112
rect 9916 6072 10692 6100
rect 9916 6060 9922 6072
rect 10686 6060 10692 6072
rect 10744 6060 10750 6112
rect 10962 6060 10968 6112
rect 11020 6100 11026 6112
rect 11149 6103 11207 6109
rect 11149 6100 11161 6103
rect 11020 6072 11161 6100
rect 11020 6060 11026 6072
rect 11149 6069 11161 6072
rect 11195 6069 11207 6103
rect 11149 6063 11207 6069
rect 11330 6060 11336 6112
rect 11388 6100 11394 6112
rect 11517 6103 11575 6109
rect 11517 6100 11529 6103
rect 11388 6072 11529 6100
rect 11388 6060 11394 6072
rect 11517 6069 11529 6072
rect 11563 6069 11575 6103
rect 13078 6100 13084 6112
rect 13039 6072 13084 6100
rect 11517 6063 11575 6069
rect 13078 6060 13084 6072
rect 13136 6060 13142 6112
rect 13188 6100 13216 6208
rect 13265 6205 13277 6239
rect 13311 6205 13323 6239
rect 13265 6199 13323 6205
rect 13449 6239 13507 6245
rect 13449 6205 13461 6239
rect 13495 6205 13507 6239
rect 13556 6236 13584 6276
rect 14366 6264 14372 6316
rect 14424 6304 14430 6316
rect 14734 6304 14740 6316
rect 14424 6276 14469 6304
rect 14647 6276 14740 6304
rect 14424 6264 14430 6276
rect 14734 6264 14740 6276
rect 14792 6304 14798 6316
rect 15289 6307 15347 6313
rect 15289 6304 15301 6307
rect 14792 6276 15301 6304
rect 14792 6264 14798 6276
rect 15289 6273 15301 6276
rect 15335 6273 15347 6307
rect 15289 6267 15347 6273
rect 14274 6236 14280 6248
rect 13556 6208 14280 6236
rect 13449 6199 13507 6205
rect 13464 6168 13492 6199
rect 14274 6196 14280 6208
rect 14332 6196 14338 6248
rect 14645 6239 14703 6245
rect 14645 6205 14657 6239
rect 14691 6236 14703 6239
rect 15473 6239 15531 6245
rect 15473 6236 15485 6239
rect 14691 6208 15485 6236
rect 14691 6205 14703 6208
rect 14645 6199 14703 6205
rect 15473 6205 15485 6208
rect 15519 6205 15531 6239
rect 15473 6199 15531 6205
rect 14829 6171 14887 6177
rect 14829 6168 14841 6171
rect 13464 6140 14841 6168
rect 14829 6137 14841 6140
rect 14875 6137 14887 6171
rect 15488 6168 15516 6199
rect 15746 6196 15752 6248
rect 15804 6236 15810 6248
rect 16224 6245 16252 6344
rect 17037 6341 17049 6375
rect 17083 6372 17095 6375
rect 18325 6375 18383 6381
rect 18325 6372 18337 6375
rect 17083 6344 18337 6372
rect 17083 6341 17095 6344
rect 17037 6335 17095 6341
rect 18325 6341 18337 6344
rect 18371 6341 18383 6375
rect 18325 6335 18383 6341
rect 17402 6264 17408 6316
rect 17460 6304 17466 6316
rect 17865 6307 17923 6313
rect 17865 6304 17877 6307
rect 17460 6276 17877 6304
rect 17460 6264 17466 6276
rect 17865 6273 17877 6276
rect 17911 6273 17923 6307
rect 17865 6267 17923 6273
rect 16117 6239 16175 6245
rect 16117 6236 16129 6239
rect 15804 6208 16129 6236
rect 15804 6196 15810 6208
rect 16117 6205 16129 6208
rect 16163 6205 16175 6239
rect 16117 6199 16175 6205
rect 16209 6239 16267 6245
rect 16209 6205 16221 6239
rect 16255 6205 16267 6239
rect 16209 6199 16267 6205
rect 16853 6239 16911 6245
rect 16853 6205 16865 6239
rect 16899 6205 16911 6239
rect 16853 6199 16911 6205
rect 16945 6239 17003 6245
rect 16945 6205 16957 6239
rect 16991 6236 17003 6239
rect 17126 6236 17132 6248
rect 16991 6208 17132 6236
rect 16991 6205 17003 6208
rect 16945 6199 17003 6205
rect 16666 6168 16672 6180
rect 15488 6140 16672 6168
rect 14829 6131 14887 6137
rect 16666 6128 16672 6140
rect 16724 6128 16730 6180
rect 16868 6168 16896 6199
rect 17126 6196 17132 6208
rect 17184 6196 17190 6248
rect 17218 6196 17224 6248
rect 17276 6236 17282 6248
rect 17957 6239 18015 6245
rect 17957 6236 17969 6239
rect 17276 6208 17969 6236
rect 17276 6196 17282 6208
rect 17957 6205 17969 6208
rect 18003 6205 18015 6239
rect 17957 6199 18015 6205
rect 18049 6239 18107 6245
rect 18049 6205 18061 6239
rect 18095 6205 18107 6239
rect 18049 6199 18107 6205
rect 17586 6168 17592 6180
rect 16868 6140 17592 6168
rect 17586 6128 17592 6140
rect 17644 6128 17650 6180
rect 17862 6128 17868 6180
rect 17920 6168 17926 6180
rect 18064 6168 18092 6199
rect 17920 6140 18092 6168
rect 17920 6128 17926 6140
rect 13630 6100 13636 6112
rect 13188 6072 13636 6100
rect 13630 6060 13636 6072
rect 13688 6060 13694 6112
rect 13909 6103 13967 6109
rect 13909 6069 13921 6103
rect 13955 6100 13967 6103
rect 14182 6100 14188 6112
rect 13955 6072 14188 6100
rect 13955 6069 13967 6072
rect 13909 6063 13967 6069
rect 14182 6060 14188 6072
rect 14240 6060 14246 6112
rect 15286 6060 15292 6112
rect 15344 6100 15350 6112
rect 15657 6103 15715 6109
rect 15657 6100 15669 6103
rect 15344 6072 15669 6100
rect 15344 6060 15350 6072
rect 15657 6069 15669 6072
rect 15703 6069 15715 6103
rect 15657 6063 15715 6069
rect 15930 6060 15936 6112
rect 15988 6100 15994 6112
rect 17497 6103 17555 6109
rect 17497 6100 17509 6103
rect 15988 6072 17509 6100
rect 15988 6060 15994 6072
rect 17497 6069 17509 6072
rect 17543 6069 17555 6103
rect 17497 6063 17555 6069
rect 1104 6010 18860 6032
rect 1104 5958 3174 6010
rect 3226 5958 3238 6010
rect 3290 5958 3302 6010
rect 3354 5958 3366 6010
rect 3418 5958 3430 6010
rect 3482 5958 7622 6010
rect 7674 5958 7686 6010
rect 7738 5958 7750 6010
rect 7802 5958 7814 6010
rect 7866 5958 7878 6010
rect 7930 5958 12070 6010
rect 12122 5958 12134 6010
rect 12186 5958 12198 6010
rect 12250 5958 12262 6010
rect 12314 5958 12326 6010
rect 12378 5958 16518 6010
rect 16570 5958 16582 6010
rect 16634 5958 16646 6010
rect 16698 5958 16710 6010
rect 16762 5958 16774 6010
rect 16826 5958 18860 6010
rect 1104 5936 18860 5958
rect 1581 5899 1639 5905
rect 1581 5865 1593 5899
rect 1627 5896 1639 5899
rect 1854 5896 1860 5908
rect 1627 5868 1860 5896
rect 1627 5865 1639 5868
rect 1581 5859 1639 5865
rect 1854 5856 1860 5868
rect 1912 5856 1918 5908
rect 3418 5856 3424 5908
rect 3476 5896 3482 5908
rect 3973 5899 4031 5905
rect 3973 5896 3985 5899
rect 3476 5868 3985 5896
rect 3476 5856 3482 5868
rect 3973 5865 3985 5868
rect 4019 5896 4031 5899
rect 4982 5896 4988 5908
rect 4019 5868 4988 5896
rect 4019 5865 4031 5868
rect 3973 5859 4031 5865
rect 4982 5856 4988 5868
rect 5040 5856 5046 5908
rect 5626 5896 5632 5908
rect 5587 5868 5632 5896
rect 5626 5856 5632 5868
rect 5684 5856 5690 5908
rect 6454 5896 6460 5908
rect 6415 5868 6460 5896
rect 6454 5856 6460 5868
rect 6512 5856 6518 5908
rect 6733 5899 6791 5905
rect 6733 5865 6745 5899
rect 6779 5896 6791 5899
rect 8294 5896 8300 5908
rect 6779 5868 8300 5896
rect 6779 5865 6791 5868
rect 6733 5859 6791 5865
rect 8294 5856 8300 5868
rect 8352 5856 8358 5908
rect 8478 5856 8484 5908
rect 8536 5896 8542 5908
rect 8536 5868 10097 5896
rect 8536 5856 8542 5868
rect 2682 5788 2688 5840
rect 2740 5828 2746 5840
rect 4065 5831 4123 5837
rect 4065 5828 4077 5831
rect 2740 5800 4077 5828
rect 2740 5788 2746 5800
rect 4065 5797 4077 5800
rect 4111 5797 4123 5831
rect 4065 5791 4123 5797
rect 4246 5788 4252 5840
rect 4304 5788 4310 5840
rect 7929 5831 7987 5837
rect 7208 5800 7420 5828
rect 1489 5763 1547 5769
rect 1489 5729 1501 5763
rect 1535 5760 1547 5763
rect 1578 5760 1584 5772
rect 1535 5732 1584 5760
rect 1535 5729 1547 5732
rect 1489 5723 1547 5729
rect 1578 5720 1584 5732
rect 1636 5720 1642 5772
rect 2222 5760 2228 5772
rect 2183 5732 2228 5760
rect 2222 5720 2228 5732
rect 2280 5720 2286 5772
rect 2866 5760 2872 5772
rect 2827 5732 2872 5760
rect 2866 5720 2872 5732
rect 2924 5720 2930 5772
rect 3053 5763 3111 5769
rect 3053 5729 3065 5763
rect 3099 5760 3111 5763
rect 3142 5760 3148 5772
rect 3099 5732 3148 5760
rect 3099 5729 3111 5732
rect 3053 5723 3111 5729
rect 3142 5720 3148 5732
rect 3200 5720 3206 5772
rect 4264 5760 4292 5788
rect 4890 5760 4896 5772
rect 3620 5732 4292 5760
rect 4540 5732 4896 5760
rect 3237 5695 3295 5701
rect 3237 5661 3249 5695
rect 3283 5692 3295 5695
rect 3510 5692 3516 5704
rect 3283 5664 3516 5692
rect 3283 5661 3295 5664
rect 3237 5655 3295 5661
rect 3510 5652 3516 5664
rect 3568 5652 3574 5704
rect 3620 5701 3648 5732
rect 3605 5695 3663 5701
rect 3605 5661 3617 5695
rect 3651 5661 3663 5695
rect 3786 5692 3792 5704
rect 3747 5664 3792 5692
rect 3605 5655 3663 5661
rect 3786 5652 3792 5664
rect 3844 5652 3850 5704
rect 4246 5652 4252 5704
rect 4304 5701 4310 5704
rect 4540 5701 4568 5732
rect 4890 5720 4896 5732
rect 4948 5720 4954 5772
rect 5077 5763 5135 5769
rect 5077 5729 5089 5763
rect 5123 5760 5135 5763
rect 5718 5760 5724 5772
rect 5123 5732 5724 5760
rect 5123 5729 5135 5732
rect 5077 5723 5135 5729
rect 5718 5720 5724 5732
rect 5776 5720 5782 5772
rect 5905 5763 5963 5769
rect 5905 5729 5917 5763
rect 5951 5760 5963 5763
rect 5994 5760 6000 5772
rect 5951 5732 6000 5760
rect 5951 5729 5963 5732
rect 5905 5723 5963 5729
rect 5994 5720 6000 5732
rect 6052 5720 6058 5772
rect 6178 5720 6184 5772
rect 6236 5760 6242 5772
rect 7208 5769 7236 5800
rect 7193 5763 7251 5769
rect 6236 5732 6776 5760
rect 6236 5720 6242 5732
rect 4304 5692 4315 5701
rect 4525 5695 4583 5701
rect 4304 5664 4349 5692
rect 4304 5655 4315 5664
rect 4525 5661 4537 5695
rect 4571 5661 4583 5695
rect 4525 5655 4583 5661
rect 4801 5695 4859 5701
rect 4801 5661 4813 5695
rect 4847 5692 4859 5695
rect 5350 5692 5356 5704
rect 4847 5664 5356 5692
rect 4847 5661 4859 5664
rect 4801 5655 4859 5661
rect 4304 5652 4310 5655
rect 5350 5652 5356 5664
rect 5408 5692 5414 5704
rect 5408 5664 5764 5692
rect 5408 5652 5414 5664
rect 5736 5636 5764 5664
rect 6454 5652 6460 5704
rect 6512 5692 6518 5704
rect 6549 5695 6607 5701
rect 6549 5692 6561 5695
rect 6512 5664 6561 5692
rect 6512 5652 6518 5664
rect 6549 5661 6561 5664
rect 6595 5661 6607 5695
rect 6748 5692 6776 5732
rect 7193 5729 7205 5763
rect 7239 5729 7251 5763
rect 7392 5760 7420 5800
rect 7929 5797 7941 5831
rect 7975 5828 7987 5831
rect 8018 5828 8024 5840
rect 7975 5800 8024 5828
rect 7975 5797 7987 5800
rect 7929 5791 7987 5797
rect 8018 5788 8024 5800
rect 8076 5788 8082 5840
rect 8312 5828 8340 5856
rect 9674 5828 9680 5840
rect 8312 5800 9680 5828
rect 9674 5788 9680 5800
rect 9732 5828 9738 5840
rect 10069 5828 10097 5868
rect 11882 5856 11888 5908
rect 11940 5896 11946 5908
rect 12621 5899 12679 5905
rect 12621 5896 12633 5899
rect 11940 5868 12633 5896
rect 11940 5856 11946 5868
rect 12621 5865 12633 5868
rect 12667 5865 12679 5899
rect 12621 5859 12679 5865
rect 12986 5856 12992 5908
rect 13044 5896 13050 5908
rect 13446 5896 13452 5908
rect 13044 5868 13452 5896
rect 13044 5856 13050 5868
rect 13446 5856 13452 5868
rect 13504 5856 13510 5908
rect 13633 5899 13691 5905
rect 13633 5896 13645 5899
rect 13556 5868 13645 5896
rect 12066 5828 12072 5840
rect 9732 5800 9996 5828
rect 10069 5800 12072 5828
rect 9732 5788 9738 5800
rect 8202 5760 8208 5772
rect 7392 5732 8208 5760
rect 7193 5723 7251 5729
rect 8202 5720 8208 5732
rect 8260 5720 8266 5772
rect 8665 5763 8723 5769
rect 8665 5729 8677 5763
rect 8711 5760 8723 5763
rect 9030 5760 9036 5772
rect 8711 5732 9036 5760
rect 8711 5729 8723 5732
rect 8665 5723 8723 5729
rect 9030 5720 9036 5732
rect 9088 5720 9094 5772
rect 9214 5760 9220 5772
rect 9175 5732 9220 5760
rect 9214 5720 9220 5732
rect 9272 5720 9278 5772
rect 9306 5720 9312 5772
rect 9364 5760 9370 5772
rect 9968 5769 9996 5800
rect 12066 5788 12072 5800
rect 12124 5788 12130 5840
rect 12526 5788 12532 5840
rect 12584 5828 12590 5840
rect 12584 5800 13216 5828
rect 12584 5788 12590 5800
rect 9953 5763 10011 5769
rect 9364 5732 9904 5760
rect 9364 5720 9370 5732
rect 7285 5695 7343 5701
rect 7285 5692 7297 5695
rect 6748 5664 7297 5692
rect 6549 5655 6607 5661
rect 7285 5661 7297 5664
rect 7331 5661 7343 5695
rect 7285 5655 7343 5661
rect 7377 5695 7435 5701
rect 7377 5661 7389 5695
rect 7423 5688 7435 5695
rect 7834 5692 7840 5704
rect 7484 5688 7840 5692
rect 7423 5664 7840 5688
rect 7423 5661 7512 5664
rect 7377 5660 7512 5661
rect 7377 5655 7435 5660
rect 7834 5652 7840 5664
rect 7892 5652 7898 5704
rect 8478 5692 8484 5704
rect 8439 5664 8484 5692
rect 8478 5652 8484 5664
rect 8536 5652 8542 5704
rect 8570 5652 8576 5704
rect 8628 5692 8634 5704
rect 8938 5692 8944 5704
rect 8628 5664 8944 5692
rect 8628 5652 8634 5664
rect 8938 5652 8944 5664
rect 8996 5652 9002 5704
rect 9493 5695 9551 5701
rect 9493 5661 9505 5695
rect 9539 5692 9551 5695
rect 9766 5692 9772 5704
rect 9539 5664 9772 5692
rect 9539 5661 9551 5664
rect 9493 5655 9551 5661
rect 9766 5652 9772 5664
rect 9824 5652 9830 5704
rect 9876 5692 9904 5732
rect 9953 5729 9965 5763
rect 9999 5729 10011 5763
rect 9953 5723 10011 5729
rect 10229 5763 10287 5769
rect 10229 5729 10241 5763
rect 10275 5760 10287 5763
rect 11422 5760 11428 5772
rect 10275 5732 11428 5760
rect 10275 5729 10287 5732
rect 10229 5723 10287 5729
rect 11422 5720 11428 5732
rect 11480 5720 11486 5772
rect 11974 5720 11980 5772
rect 12032 5760 12038 5772
rect 12032 5732 12388 5760
rect 12032 5720 12038 5732
rect 10594 5692 10600 5704
rect 9876 5664 10600 5692
rect 10594 5652 10600 5664
rect 10652 5652 10658 5704
rect 10778 5652 10784 5704
rect 10836 5692 10842 5704
rect 10873 5695 10931 5701
rect 10873 5692 10885 5695
rect 10836 5664 10885 5692
rect 10836 5652 10842 5664
rect 10873 5661 10885 5664
rect 10919 5661 10931 5695
rect 10873 5655 10931 5661
rect 11149 5695 11207 5701
rect 11149 5661 11161 5695
rect 11195 5692 11207 5695
rect 12250 5692 12256 5704
rect 11195 5664 12256 5692
rect 11195 5661 11207 5664
rect 11149 5655 11207 5661
rect 12250 5652 12256 5664
rect 12308 5652 12314 5704
rect 12360 5692 12388 5732
rect 12434 5720 12440 5772
rect 12492 5760 12498 5772
rect 12894 5760 12900 5772
rect 12492 5732 12900 5760
rect 12492 5720 12498 5732
rect 12894 5720 12900 5732
rect 12952 5720 12958 5772
rect 13078 5760 13084 5772
rect 13039 5732 13084 5760
rect 13078 5720 13084 5732
rect 13136 5720 13142 5772
rect 13188 5769 13216 5800
rect 13262 5788 13268 5840
rect 13320 5828 13326 5840
rect 13556 5828 13584 5868
rect 13633 5865 13645 5868
rect 13679 5865 13691 5899
rect 13633 5859 13691 5865
rect 13725 5899 13783 5905
rect 13725 5865 13737 5899
rect 13771 5896 13783 5899
rect 13906 5896 13912 5908
rect 13771 5868 13912 5896
rect 13771 5865 13783 5868
rect 13725 5859 13783 5865
rect 13906 5856 13912 5868
rect 13964 5856 13970 5908
rect 15746 5896 15752 5908
rect 15707 5868 15752 5896
rect 15746 5856 15752 5868
rect 15804 5856 15810 5908
rect 16850 5856 16856 5908
rect 16908 5896 16914 5908
rect 17862 5896 17868 5908
rect 16908 5868 17868 5896
rect 16908 5856 16914 5868
rect 17862 5856 17868 5868
rect 17920 5856 17926 5908
rect 18230 5856 18236 5908
rect 18288 5896 18294 5908
rect 18325 5899 18383 5905
rect 18325 5896 18337 5899
rect 18288 5868 18337 5896
rect 18288 5856 18294 5868
rect 18325 5865 18337 5868
rect 18371 5865 18383 5899
rect 18325 5859 18383 5865
rect 13320 5800 13584 5828
rect 13648 5800 14504 5828
rect 13320 5788 13326 5800
rect 13173 5763 13231 5769
rect 13173 5729 13185 5763
rect 13219 5729 13231 5763
rect 13173 5723 13231 5729
rect 13538 5720 13544 5772
rect 13596 5760 13602 5772
rect 13648 5760 13676 5800
rect 14369 5763 14427 5769
rect 14369 5760 14381 5763
rect 13596 5732 13676 5760
rect 13823 5732 14381 5760
rect 13596 5720 13602 5732
rect 12360 5664 12940 5692
rect 12912 5636 12940 5664
rect 13262 5652 13268 5704
rect 13320 5692 13326 5704
rect 13449 5695 13507 5701
rect 13449 5692 13461 5695
rect 13320 5664 13461 5692
rect 13320 5652 13326 5664
rect 13449 5661 13461 5664
rect 13495 5692 13507 5695
rect 13722 5692 13728 5704
rect 13495 5664 13728 5692
rect 13495 5661 13507 5664
rect 13449 5655 13507 5661
rect 13722 5652 13728 5664
rect 13780 5652 13786 5704
rect 1949 5627 2007 5633
rect 1949 5593 1961 5627
rect 1995 5624 2007 5627
rect 2777 5627 2835 5633
rect 1995 5596 2452 5624
rect 1995 5593 2007 5596
rect 1949 5587 2007 5593
rect 2038 5556 2044 5568
rect 1999 5528 2044 5556
rect 2038 5516 2044 5528
rect 2096 5516 2102 5568
rect 2424 5565 2452 5596
rect 2777 5593 2789 5627
rect 2823 5624 2835 5627
rect 4062 5624 4068 5636
rect 2823 5596 4068 5624
rect 2823 5593 2835 5596
rect 2777 5587 2835 5593
rect 4062 5584 4068 5596
rect 4120 5584 4126 5636
rect 5718 5584 5724 5636
rect 5776 5584 5782 5636
rect 6822 5624 6828 5636
rect 6783 5596 6828 5624
rect 6822 5584 6828 5596
rect 6880 5584 6886 5636
rect 8294 5584 8300 5636
rect 8352 5624 8358 5636
rect 8389 5627 8447 5633
rect 8389 5624 8401 5627
rect 8352 5596 8401 5624
rect 8352 5584 8358 5596
rect 8389 5593 8401 5596
rect 8435 5593 8447 5627
rect 8389 5587 8447 5593
rect 10410 5584 10416 5636
rect 10468 5624 10474 5636
rect 10468 5596 12204 5624
rect 10468 5584 10474 5596
rect 2409 5559 2467 5565
rect 2409 5525 2421 5559
rect 2455 5525 2467 5559
rect 2409 5519 2467 5525
rect 3421 5559 3479 5565
rect 3421 5525 3433 5559
rect 3467 5556 3479 5559
rect 3878 5556 3884 5568
rect 3467 5528 3884 5556
rect 3467 5525 3479 5528
rect 3421 5519 3479 5525
rect 3878 5516 3884 5528
rect 3936 5516 3942 5568
rect 4338 5556 4344 5568
rect 4299 5528 4344 5556
rect 4338 5516 4344 5528
rect 4396 5516 4402 5568
rect 5166 5556 5172 5568
rect 5127 5528 5172 5556
rect 5166 5516 5172 5528
rect 5224 5516 5230 5568
rect 5258 5516 5264 5568
rect 5316 5556 5322 5568
rect 5316 5528 5361 5556
rect 5316 5516 5322 5528
rect 5810 5516 5816 5568
rect 5868 5556 5874 5568
rect 5997 5559 6055 5565
rect 5997 5556 6009 5559
rect 5868 5528 6009 5556
rect 5868 5516 5874 5528
rect 5997 5525 6009 5528
rect 6043 5525 6055 5559
rect 5997 5519 6055 5525
rect 6089 5559 6147 5565
rect 6089 5525 6101 5559
rect 6135 5556 6147 5559
rect 6178 5556 6184 5568
rect 6135 5528 6184 5556
rect 6135 5525 6147 5528
rect 6089 5519 6147 5525
rect 6178 5516 6184 5528
rect 6236 5516 6242 5568
rect 7466 5516 7472 5568
rect 7524 5556 7530 5568
rect 7745 5559 7803 5565
rect 7745 5556 7757 5559
rect 7524 5528 7757 5556
rect 7524 5516 7530 5528
rect 7745 5525 7757 5528
rect 7791 5525 7803 5559
rect 8018 5556 8024 5568
rect 7979 5528 8024 5556
rect 7745 5519 7803 5525
rect 8018 5516 8024 5528
rect 8076 5516 8082 5568
rect 9030 5516 9036 5568
rect 9088 5556 9094 5568
rect 9398 5556 9404 5568
rect 9088 5528 9404 5556
rect 9088 5516 9094 5528
rect 9398 5516 9404 5528
rect 9456 5516 9462 5568
rect 9766 5516 9772 5568
rect 9824 5556 9830 5568
rect 9861 5559 9919 5565
rect 9861 5556 9873 5559
rect 9824 5528 9873 5556
rect 9824 5516 9830 5528
rect 9861 5525 9873 5528
rect 9907 5525 9919 5559
rect 9861 5519 9919 5525
rect 10778 5516 10784 5568
rect 10836 5556 10842 5568
rect 12176 5565 12204 5596
rect 12894 5584 12900 5636
rect 12952 5624 12958 5636
rect 12989 5627 13047 5633
rect 12989 5624 13001 5627
rect 12952 5596 13001 5624
rect 12952 5584 12958 5596
rect 12989 5593 13001 5596
rect 13035 5593 13047 5627
rect 13823 5624 13851 5732
rect 14369 5729 14381 5732
rect 14415 5729 14427 5763
rect 14369 5723 14427 5729
rect 13909 5695 13967 5701
rect 13909 5661 13921 5695
rect 13955 5661 13967 5695
rect 13909 5655 13967 5661
rect 14093 5695 14151 5701
rect 14093 5661 14105 5695
rect 14139 5692 14151 5695
rect 14476 5692 14504 5800
rect 15378 5788 15384 5840
rect 15436 5828 15442 5840
rect 15841 5831 15899 5837
rect 15841 5828 15853 5831
rect 15436 5800 15853 5828
rect 15436 5788 15442 5800
rect 15841 5797 15853 5800
rect 15887 5797 15899 5831
rect 17497 5831 17555 5837
rect 17497 5828 17509 5831
rect 15841 5791 15899 5797
rect 16960 5800 17509 5828
rect 15102 5720 15108 5772
rect 15160 5760 15166 5772
rect 15197 5763 15255 5769
rect 15197 5760 15209 5763
rect 15160 5732 15209 5760
rect 15160 5720 15166 5732
rect 15197 5729 15209 5732
rect 15243 5729 15255 5763
rect 15197 5723 15255 5729
rect 15289 5763 15347 5769
rect 15289 5729 15301 5763
rect 15335 5760 15347 5763
rect 15930 5760 15936 5772
rect 15335 5732 15936 5760
rect 15335 5729 15347 5732
rect 15289 5723 15347 5729
rect 15930 5720 15936 5732
rect 15988 5720 15994 5772
rect 16390 5760 16396 5772
rect 16040 5732 16396 5760
rect 16040 5692 16068 5732
rect 16390 5720 16396 5732
rect 16448 5720 16454 5772
rect 16485 5763 16543 5769
rect 16485 5729 16497 5763
rect 16531 5760 16543 5763
rect 16850 5760 16856 5772
rect 16531 5732 16856 5760
rect 16531 5729 16543 5732
rect 16485 5723 16543 5729
rect 16850 5720 16856 5732
rect 16908 5720 16914 5772
rect 16206 5692 16212 5704
rect 14139 5664 16068 5692
rect 16167 5664 16212 5692
rect 14139 5661 14151 5664
rect 14093 5655 14151 5661
rect 12989 5587 13047 5593
rect 13188 5596 13851 5624
rect 13924 5624 13952 5655
rect 16206 5652 16212 5664
rect 16264 5652 16270 5704
rect 16960 5692 16988 5800
rect 17497 5797 17509 5800
rect 17543 5797 17555 5831
rect 17497 5791 17555 5797
rect 17586 5788 17592 5840
rect 17644 5828 17650 5840
rect 17644 5800 18368 5828
rect 17644 5788 17650 5800
rect 17313 5763 17371 5769
rect 17313 5729 17325 5763
rect 17359 5760 17371 5763
rect 17359 5732 17540 5760
rect 17359 5729 17371 5732
rect 17313 5723 17371 5729
rect 17512 5704 17540 5732
rect 17862 5720 17868 5772
rect 17920 5760 17926 5772
rect 18049 5763 18107 5769
rect 18049 5760 18061 5763
rect 17920 5732 18061 5760
rect 17920 5720 17926 5732
rect 18049 5729 18061 5732
rect 18095 5729 18107 5763
rect 18049 5723 18107 5729
rect 16408 5664 16988 5692
rect 15194 5624 15200 5636
rect 13924 5596 15200 5624
rect 11793 5559 11851 5565
rect 11793 5556 11805 5559
rect 10836 5528 11805 5556
rect 10836 5516 10842 5528
rect 11793 5525 11805 5528
rect 11839 5525 11851 5559
rect 11793 5519 11851 5525
rect 12161 5559 12219 5565
rect 12161 5525 12173 5559
rect 12207 5556 12219 5559
rect 13188 5556 13216 5596
rect 15194 5584 15200 5596
rect 15252 5584 15258 5636
rect 15381 5627 15439 5633
rect 15381 5593 15393 5627
rect 15427 5624 15439 5627
rect 16408 5624 16436 5664
rect 17034 5652 17040 5704
rect 17092 5652 17098 5704
rect 17494 5652 17500 5704
rect 17552 5652 17558 5704
rect 18340 5692 18368 5800
rect 18509 5695 18567 5701
rect 18509 5692 18521 5695
rect 18340 5664 18521 5692
rect 18509 5661 18521 5664
rect 18555 5661 18567 5695
rect 18509 5655 18567 5661
rect 15427 5596 16436 5624
rect 15427 5593 15439 5596
rect 15381 5587 15439 5593
rect 16758 5584 16764 5636
rect 16816 5624 16822 5636
rect 17052 5624 17080 5652
rect 17129 5627 17187 5633
rect 17129 5624 17141 5627
rect 16816 5596 17141 5624
rect 16816 5584 16822 5596
rect 17129 5593 17141 5596
rect 17175 5593 17187 5627
rect 17129 5587 17187 5593
rect 17218 5584 17224 5636
rect 17276 5624 17282 5636
rect 17276 5596 17632 5624
rect 17276 5584 17282 5596
rect 12207 5528 13216 5556
rect 12207 5525 12219 5528
rect 12161 5519 12219 5525
rect 13906 5516 13912 5568
rect 13964 5556 13970 5568
rect 14918 5556 14924 5568
rect 13964 5528 14924 5556
rect 13964 5516 13970 5528
rect 14918 5516 14924 5528
rect 14976 5556 14982 5568
rect 16301 5559 16359 5565
rect 16301 5556 16313 5559
rect 14976 5528 16313 5556
rect 14976 5516 14982 5528
rect 16301 5525 16313 5528
rect 16347 5525 16359 5559
rect 16301 5519 16359 5525
rect 16574 5516 16580 5568
rect 16632 5556 16638 5568
rect 16669 5559 16727 5565
rect 16669 5556 16681 5559
rect 16632 5528 16681 5556
rect 16632 5516 16638 5528
rect 16669 5525 16681 5528
rect 16715 5525 16727 5559
rect 17034 5556 17040 5568
rect 16995 5528 17040 5556
rect 16669 5519 16727 5525
rect 17034 5516 17040 5528
rect 17092 5516 17098 5568
rect 17604 5556 17632 5596
rect 17678 5584 17684 5636
rect 17736 5624 17742 5636
rect 17957 5627 18015 5633
rect 17957 5624 17969 5627
rect 17736 5596 17969 5624
rect 17736 5584 17742 5596
rect 17957 5593 17969 5596
rect 18003 5593 18015 5627
rect 17957 5587 18015 5593
rect 17865 5559 17923 5565
rect 17865 5556 17877 5559
rect 17604 5528 17877 5556
rect 17865 5525 17877 5528
rect 17911 5525 17923 5559
rect 17865 5519 17923 5525
rect 1104 5466 18860 5488
rect 1104 5414 5398 5466
rect 5450 5414 5462 5466
rect 5514 5414 5526 5466
rect 5578 5414 5590 5466
rect 5642 5414 5654 5466
rect 5706 5414 9846 5466
rect 9898 5414 9910 5466
rect 9962 5414 9974 5466
rect 10026 5414 10038 5466
rect 10090 5414 10102 5466
rect 10154 5414 14294 5466
rect 14346 5414 14358 5466
rect 14410 5414 14422 5466
rect 14474 5414 14486 5466
rect 14538 5414 14550 5466
rect 14602 5414 18860 5466
rect 1104 5392 18860 5414
rect 1486 5352 1492 5364
rect 1447 5324 1492 5352
rect 1486 5312 1492 5324
rect 1544 5312 1550 5364
rect 1857 5355 1915 5361
rect 1857 5321 1869 5355
rect 1903 5352 1915 5355
rect 2038 5352 2044 5364
rect 1903 5324 2044 5352
rect 1903 5321 1915 5324
rect 1857 5315 1915 5321
rect 2038 5312 2044 5324
rect 2096 5312 2102 5364
rect 2314 5352 2320 5364
rect 2275 5324 2320 5352
rect 2314 5312 2320 5324
rect 2372 5312 2378 5364
rect 2774 5312 2780 5364
rect 2832 5352 2838 5364
rect 3053 5355 3111 5361
rect 2832 5324 2877 5352
rect 2832 5312 2838 5324
rect 3053 5321 3065 5355
rect 3099 5321 3111 5355
rect 3973 5355 4031 5361
rect 3973 5352 3985 5355
rect 3053 5315 3111 5321
rect 3160 5324 3985 5352
rect 2225 5287 2283 5293
rect 2225 5253 2237 5287
rect 2271 5284 2283 5287
rect 2498 5284 2504 5296
rect 2271 5256 2504 5284
rect 2271 5253 2283 5256
rect 2225 5247 2283 5253
rect 2498 5244 2504 5256
rect 2556 5244 2562 5296
rect 2590 5244 2596 5296
rect 2648 5284 2654 5296
rect 3068 5284 3096 5315
rect 2648 5256 3096 5284
rect 2648 5244 2654 5256
rect 1673 5219 1731 5225
rect 1673 5185 1685 5219
rect 1719 5185 1731 5219
rect 1673 5179 1731 5185
rect 2961 5219 3019 5225
rect 2961 5185 2973 5219
rect 3007 5216 3019 5219
rect 3160 5216 3188 5324
rect 3973 5321 3985 5324
rect 4019 5321 4031 5355
rect 3973 5315 4031 5321
rect 4246 5312 4252 5364
rect 4304 5352 4310 5364
rect 4433 5355 4491 5361
rect 4433 5352 4445 5355
rect 4304 5324 4445 5352
rect 4304 5312 4310 5324
rect 4433 5321 4445 5324
rect 4479 5321 4491 5355
rect 4433 5315 4491 5321
rect 4801 5355 4859 5361
rect 4801 5321 4813 5355
rect 4847 5352 4859 5355
rect 5074 5352 5080 5364
rect 4847 5324 5080 5352
rect 4847 5321 4859 5324
rect 4801 5315 4859 5321
rect 5074 5312 5080 5324
rect 5132 5312 5138 5364
rect 5258 5312 5264 5364
rect 5316 5352 5322 5364
rect 5445 5355 5503 5361
rect 5445 5352 5457 5355
rect 5316 5324 5457 5352
rect 5316 5312 5322 5324
rect 5445 5321 5457 5324
rect 5491 5321 5503 5355
rect 5902 5352 5908 5364
rect 5863 5324 5908 5352
rect 5445 5315 5503 5321
rect 5902 5312 5908 5324
rect 5960 5352 5966 5364
rect 6454 5352 6460 5364
rect 5960 5324 6460 5352
rect 5960 5312 5966 5324
rect 6454 5312 6460 5324
rect 6512 5312 6518 5364
rect 6549 5355 6607 5361
rect 6549 5321 6561 5355
rect 6595 5352 6607 5355
rect 7006 5352 7012 5364
rect 6595 5324 7012 5352
rect 6595 5321 6607 5324
rect 6549 5315 6607 5321
rect 7006 5312 7012 5324
rect 7064 5312 7070 5364
rect 7282 5312 7288 5364
rect 7340 5352 7346 5364
rect 7377 5355 7435 5361
rect 7377 5352 7389 5355
rect 7340 5324 7389 5352
rect 7340 5312 7346 5324
rect 7377 5321 7389 5324
rect 7423 5321 7435 5355
rect 7834 5352 7840 5364
rect 7795 5324 7840 5352
rect 7377 5315 7435 5321
rect 7834 5312 7840 5324
rect 7892 5312 7898 5364
rect 8018 5312 8024 5364
rect 8076 5352 8082 5364
rect 8297 5355 8355 5361
rect 8297 5352 8309 5355
rect 8076 5324 8309 5352
rect 8076 5312 8082 5324
rect 8297 5321 8309 5324
rect 8343 5321 8355 5355
rect 8297 5315 8355 5321
rect 8757 5355 8815 5361
rect 8757 5321 8769 5355
rect 8803 5352 8815 5355
rect 8846 5352 8852 5364
rect 8803 5324 8852 5352
rect 8803 5321 8815 5324
rect 8757 5315 8815 5321
rect 8846 5312 8852 5324
rect 8904 5312 8910 5364
rect 9766 5312 9772 5364
rect 9824 5352 9830 5364
rect 10045 5355 10103 5361
rect 10045 5352 10057 5355
rect 9824 5324 10057 5352
rect 9824 5312 9830 5324
rect 10045 5321 10057 5324
rect 10091 5321 10103 5355
rect 10778 5352 10784 5364
rect 10739 5324 10784 5352
rect 10045 5315 10103 5321
rect 10778 5312 10784 5324
rect 10836 5312 10842 5364
rect 10873 5355 10931 5361
rect 10873 5321 10885 5355
rect 10919 5352 10931 5355
rect 11517 5355 11575 5361
rect 11517 5352 11529 5355
rect 10919 5324 11529 5352
rect 10919 5321 10931 5324
rect 10873 5315 10931 5321
rect 11517 5321 11529 5324
rect 11563 5321 11575 5355
rect 11517 5315 11575 5321
rect 12621 5355 12679 5361
rect 12621 5321 12633 5355
rect 12667 5352 12679 5355
rect 13173 5355 13231 5361
rect 13173 5352 13185 5355
rect 12667 5324 13185 5352
rect 12667 5321 12679 5324
rect 12621 5315 12679 5321
rect 13173 5321 13185 5324
rect 13219 5321 13231 5355
rect 13538 5352 13544 5364
rect 13499 5324 13544 5352
rect 13173 5315 13231 5321
rect 13538 5312 13544 5324
rect 13596 5312 13602 5364
rect 13633 5355 13691 5361
rect 13633 5321 13645 5355
rect 13679 5352 13691 5355
rect 13906 5352 13912 5364
rect 13679 5324 13912 5352
rect 13679 5321 13691 5324
rect 13633 5315 13691 5321
rect 13906 5312 13912 5324
rect 13964 5352 13970 5364
rect 15102 5352 15108 5364
rect 13964 5324 15108 5352
rect 13964 5312 13970 5324
rect 15102 5312 15108 5324
rect 15160 5312 15166 5364
rect 15841 5355 15899 5361
rect 15841 5321 15853 5355
rect 15887 5352 15899 5355
rect 15930 5352 15936 5364
rect 15887 5324 15936 5352
rect 15887 5321 15899 5324
rect 15841 5315 15899 5321
rect 15930 5312 15936 5324
rect 15988 5352 15994 5364
rect 16114 5352 16120 5364
rect 15988 5324 16120 5352
rect 15988 5312 15994 5324
rect 16114 5312 16120 5324
rect 16172 5312 16178 5364
rect 16206 5312 16212 5364
rect 16264 5352 16270 5364
rect 16301 5355 16359 5361
rect 16301 5352 16313 5355
rect 16264 5324 16313 5352
rect 16264 5312 16270 5324
rect 16301 5321 16313 5324
rect 16347 5321 16359 5355
rect 16301 5315 16359 5321
rect 17126 5312 17132 5364
rect 17184 5352 17190 5364
rect 18049 5355 18107 5361
rect 18049 5352 18061 5355
rect 17184 5324 18061 5352
rect 17184 5312 17190 5324
rect 18049 5321 18061 5324
rect 18095 5352 18107 5355
rect 18690 5352 18696 5364
rect 18095 5324 18696 5352
rect 18095 5321 18107 5324
rect 18049 5315 18107 5321
rect 18690 5312 18696 5324
rect 18748 5312 18754 5364
rect 4890 5284 4896 5296
rect 4851 5256 4896 5284
rect 4890 5244 4896 5256
rect 4948 5244 4954 5296
rect 4982 5244 4988 5296
rect 5040 5284 5046 5296
rect 5626 5284 5632 5296
rect 5040 5256 5632 5284
rect 5040 5244 5046 5256
rect 5626 5244 5632 5256
rect 5684 5284 5690 5296
rect 6733 5287 6791 5293
rect 5684 5256 6408 5284
rect 5684 5244 5690 5256
rect 3007 5188 3188 5216
rect 3007 5185 3019 5188
rect 2961 5179 3019 5185
rect 1688 5080 1716 5179
rect 3234 5176 3240 5228
rect 3292 5216 3298 5228
rect 3510 5216 3516 5228
rect 3292 5188 3337 5216
rect 3471 5188 3516 5216
rect 3292 5176 3298 5188
rect 3510 5176 3516 5188
rect 3568 5176 3574 5228
rect 4157 5219 4215 5225
rect 4157 5185 4169 5219
rect 4203 5216 4215 5219
rect 5813 5219 5871 5225
rect 4203 5188 5212 5216
rect 4203 5185 4215 5188
rect 4157 5179 4215 5185
rect 2501 5151 2559 5157
rect 2501 5117 2513 5151
rect 2547 5148 2559 5151
rect 2590 5148 2596 5160
rect 2547 5120 2596 5148
rect 2547 5117 2559 5120
rect 2501 5111 2559 5117
rect 2590 5108 2596 5120
rect 2648 5108 2654 5160
rect 3528 5148 3556 5176
rect 3528 5120 5120 5148
rect 3329 5083 3387 5089
rect 3329 5080 3341 5083
rect 1688 5052 3341 5080
rect 3329 5049 3341 5052
rect 3375 5049 3387 5083
rect 3329 5043 3387 5049
rect 3418 5040 3424 5092
rect 3476 5080 3482 5092
rect 3605 5083 3663 5089
rect 3605 5080 3617 5083
rect 3476 5052 3617 5080
rect 3476 5040 3482 5052
rect 3605 5049 3617 5052
rect 3651 5049 3663 5083
rect 3605 5043 3663 5049
rect 2590 4972 2596 5024
rect 2648 5012 2654 5024
rect 2958 5012 2964 5024
rect 2648 4984 2964 5012
rect 2648 4972 2654 4984
rect 2958 4972 2964 4984
rect 3016 5012 3022 5024
rect 3510 5012 3516 5024
rect 3016 4984 3516 5012
rect 3016 4972 3022 4984
rect 3510 4972 3516 4984
rect 3568 5012 3574 5024
rect 3789 5015 3847 5021
rect 3789 5012 3801 5015
rect 3568 4984 3801 5012
rect 3568 4972 3574 4984
rect 3789 4981 3801 4984
rect 3835 4981 3847 5015
rect 3789 4975 3847 4981
rect 4341 5015 4399 5021
rect 4341 4981 4353 5015
rect 4387 5012 4399 5015
rect 4706 5012 4712 5024
rect 4387 4984 4712 5012
rect 4387 4981 4399 4984
rect 4341 4975 4399 4981
rect 4706 4972 4712 4984
rect 4764 4972 4770 5024
rect 5092 5012 5120 5120
rect 5184 5089 5212 5188
rect 5813 5185 5825 5219
rect 5859 5216 5871 5219
rect 5902 5216 5908 5228
rect 5859 5188 5908 5216
rect 5859 5185 5871 5188
rect 5813 5179 5871 5185
rect 5902 5176 5908 5188
rect 5960 5176 5966 5228
rect 6380 5225 6408 5256
rect 6733 5253 6745 5287
rect 6779 5284 6791 5287
rect 6914 5284 6920 5296
rect 6779 5256 6920 5284
rect 6779 5253 6791 5256
rect 6733 5247 6791 5253
rect 6914 5244 6920 5256
rect 6972 5244 6978 5296
rect 7024 5284 7052 5312
rect 8205 5287 8263 5293
rect 7024 5256 8156 5284
rect 6365 5219 6423 5225
rect 6365 5185 6377 5219
rect 6411 5185 6423 5219
rect 8018 5216 8024 5228
rect 6365 5179 6423 5185
rect 7116 5188 8024 5216
rect 7116 5160 7144 5188
rect 8018 5176 8024 5188
rect 8076 5176 8082 5228
rect 8128 5216 8156 5256
rect 8205 5253 8217 5287
rect 8251 5284 8263 5287
rect 8386 5284 8392 5296
rect 8251 5256 8392 5284
rect 8251 5253 8263 5256
rect 8205 5247 8263 5253
rect 8386 5244 8392 5256
rect 8444 5244 8450 5296
rect 9674 5244 9680 5296
rect 9732 5284 9738 5296
rect 9953 5287 10011 5293
rect 9953 5284 9965 5287
rect 9732 5256 9965 5284
rect 9732 5244 9738 5256
rect 9953 5253 9965 5256
rect 9999 5253 10011 5287
rect 9953 5247 10011 5253
rect 11885 5287 11943 5293
rect 11885 5253 11897 5287
rect 11931 5284 11943 5287
rect 12986 5284 12992 5296
rect 11931 5256 12992 5284
rect 11931 5253 11943 5256
rect 11885 5247 11943 5253
rect 9030 5216 9036 5228
rect 8128 5188 9036 5216
rect 9030 5176 9036 5188
rect 9088 5176 9094 5228
rect 9125 5219 9183 5225
rect 9125 5185 9137 5219
rect 9171 5216 9183 5219
rect 11900 5216 11928 5247
rect 12986 5244 12992 5256
rect 13044 5244 13050 5296
rect 14369 5287 14427 5293
rect 14369 5253 14381 5287
rect 14415 5253 14427 5287
rect 15194 5284 15200 5296
rect 14369 5247 14427 5253
rect 15028 5256 15200 5284
rect 12526 5216 12532 5228
rect 9171 5188 11928 5216
rect 12084 5188 12532 5216
rect 9171 5185 9183 5188
rect 9125 5179 9183 5185
rect 5353 5151 5411 5157
rect 5353 5117 5365 5151
rect 5399 5148 5411 5151
rect 5994 5148 6000 5160
rect 5399 5120 6000 5148
rect 5399 5117 5411 5120
rect 5353 5111 5411 5117
rect 5994 5108 6000 5120
rect 6052 5108 6058 5160
rect 6914 5148 6920 5160
rect 6656 5120 6920 5148
rect 5169 5083 5227 5089
rect 5169 5049 5181 5083
rect 5215 5080 5227 5083
rect 6656 5080 6684 5120
rect 6914 5108 6920 5120
rect 6972 5108 6978 5160
rect 7098 5148 7104 5160
rect 7059 5120 7104 5148
rect 7098 5108 7104 5120
rect 7156 5108 7162 5160
rect 7285 5151 7343 5157
rect 7285 5117 7297 5151
rect 7331 5148 7343 5151
rect 8110 5148 8116 5160
rect 7331 5120 8116 5148
rect 7331 5117 7343 5120
rect 7285 5111 7343 5117
rect 8110 5108 8116 5120
rect 8168 5108 8174 5160
rect 8202 5108 8208 5160
rect 8260 5148 8266 5160
rect 8389 5151 8447 5157
rect 8389 5148 8401 5151
rect 8260 5120 8401 5148
rect 8260 5108 8266 5120
rect 8389 5117 8401 5120
rect 8435 5117 8447 5151
rect 8389 5111 8447 5117
rect 5215 5052 6684 5080
rect 5215 5049 5227 5052
rect 5169 5043 5227 5049
rect 6730 5040 6736 5092
rect 6788 5080 6794 5092
rect 9140 5080 9168 5179
rect 9214 5108 9220 5160
rect 9272 5148 9278 5160
rect 9401 5151 9459 5157
rect 9272 5120 9317 5148
rect 9272 5108 9278 5120
rect 9401 5117 9413 5151
rect 9447 5117 9459 5151
rect 10134 5148 10140 5160
rect 10095 5120 10140 5148
rect 9401 5111 9459 5117
rect 6788 5052 7328 5080
rect 6788 5040 6794 5052
rect 6825 5015 6883 5021
rect 6825 5012 6837 5015
rect 5092 4984 6837 5012
rect 6825 4981 6837 4984
rect 6871 5012 6883 5015
rect 7098 5012 7104 5024
rect 6871 4984 7104 5012
rect 6871 4981 6883 4984
rect 6825 4975 6883 4981
rect 7098 4972 7104 4984
rect 7156 4972 7162 5024
rect 7300 5012 7328 5052
rect 7484 5052 9168 5080
rect 9416 5080 9444 5111
rect 10134 5108 10140 5120
rect 10192 5108 10198 5160
rect 10689 5151 10747 5157
rect 10689 5117 10701 5151
rect 10735 5117 10747 5151
rect 11974 5148 11980 5160
rect 11935 5120 11980 5148
rect 10689 5111 10747 5117
rect 10502 5080 10508 5092
rect 9416 5052 10508 5080
rect 7484 5012 7512 5052
rect 10502 5040 10508 5052
rect 10560 5040 10566 5092
rect 10704 5080 10732 5111
rect 11974 5108 11980 5120
rect 12032 5108 12038 5160
rect 12084 5080 12112 5188
rect 12526 5176 12532 5188
rect 12584 5176 12590 5228
rect 12713 5219 12771 5225
rect 12713 5185 12725 5219
rect 12759 5216 12771 5219
rect 13170 5216 13176 5228
rect 12759 5188 13176 5216
rect 12759 5185 12771 5188
rect 12713 5179 12771 5185
rect 12161 5151 12219 5157
rect 12161 5117 12173 5151
rect 12207 5148 12219 5151
rect 12342 5148 12348 5160
rect 12207 5120 12348 5148
rect 12207 5117 12219 5120
rect 12161 5111 12219 5117
rect 12342 5108 12348 5120
rect 12400 5108 12406 5160
rect 12437 5151 12495 5157
rect 12437 5117 12449 5151
rect 12483 5148 12495 5151
rect 12483 5120 12572 5148
rect 12483 5117 12495 5120
rect 12437 5111 12495 5117
rect 12544 5092 12572 5120
rect 10704 5052 12112 5080
rect 12526 5040 12532 5092
rect 12584 5040 12590 5092
rect 7300 4984 7512 5012
rect 7745 5015 7803 5021
rect 7745 4981 7757 5015
rect 7791 5012 7803 5015
rect 8294 5012 8300 5024
rect 7791 4984 8300 5012
rect 7791 4981 7803 4984
rect 7745 4975 7803 4981
rect 8294 4972 8300 4984
rect 8352 4972 8358 5024
rect 9582 5012 9588 5024
rect 9543 4984 9588 5012
rect 9582 4972 9588 4984
rect 9640 4972 9646 5024
rect 11238 5012 11244 5024
rect 11199 4984 11244 5012
rect 11238 4972 11244 4984
rect 11296 4972 11302 5024
rect 11974 4972 11980 5024
rect 12032 5012 12038 5024
rect 12728 5012 12756 5179
rect 13170 5176 13176 5188
rect 13228 5176 13234 5228
rect 13262 5176 13268 5228
rect 13320 5216 13326 5228
rect 14384 5216 14412 5247
rect 15028 5225 15056 5256
rect 15194 5244 15200 5256
rect 15252 5244 15258 5296
rect 15749 5287 15807 5293
rect 15749 5253 15761 5287
rect 15795 5284 15807 5287
rect 18509 5287 18567 5293
rect 15795 5256 16712 5284
rect 15795 5253 15807 5256
rect 15749 5247 15807 5253
rect 13320 5188 14412 5216
rect 15013 5219 15071 5225
rect 13320 5176 13326 5188
rect 15013 5185 15025 5219
rect 15059 5185 15071 5219
rect 15013 5179 15071 5185
rect 15102 5176 15108 5228
rect 15160 5216 15166 5228
rect 16684 5225 16712 5256
rect 18509 5253 18521 5287
rect 18555 5284 18567 5287
rect 18966 5284 18972 5296
rect 18555 5256 18972 5284
rect 18555 5253 18567 5256
rect 18509 5247 18567 5253
rect 18966 5244 18972 5256
rect 19024 5244 19030 5296
rect 16669 5219 16727 5225
rect 15160 5188 15205 5216
rect 15160 5176 15166 5188
rect 16669 5185 16681 5219
rect 16715 5216 16727 5219
rect 17310 5216 17316 5228
rect 16715 5188 17316 5216
rect 16715 5185 16727 5188
rect 16669 5179 16727 5185
rect 17310 5176 17316 5188
rect 17368 5176 17374 5228
rect 17954 5216 17960 5228
rect 17915 5188 17960 5216
rect 17954 5176 17960 5188
rect 18012 5176 18018 5228
rect 13354 5108 13360 5160
rect 13412 5148 13418 5160
rect 13725 5151 13783 5157
rect 13725 5148 13737 5151
rect 13412 5120 13737 5148
rect 13412 5108 13418 5120
rect 13725 5117 13737 5120
rect 13771 5117 13783 5151
rect 13725 5111 13783 5117
rect 14366 5108 14372 5160
rect 14424 5148 14430 5160
rect 14461 5151 14519 5157
rect 14461 5148 14473 5151
rect 14424 5120 14473 5148
rect 14424 5108 14430 5120
rect 14461 5117 14473 5120
rect 14507 5117 14519 5151
rect 14461 5111 14519 5117
rect 14550 5108 14556 5160
rect 14608 5148 14614 5160
rect 15657 5151 15715 5157
rect 14608 5120 14653 5148
rect 14608 5108 14614 5120
rect 15657 5117 15669 5151
rect 15703 5117 15715 5151
rect 15657 5111 15715 5117
rect 12986 5040 12992 5092
rect 13044 5080 13050 5092
rect 14829 5083 14887 5089
rect 14829 5080 14841 5083
rect 13044 5052 14841 5080
rect 13044 5040 13050 5052
rect 14829 5049 14841 5052
rect 14875 5049 14887 5083
rect 14829 5043 14887 5049
rect 15378 5040 15384 5092
rect 15436 5080 15442 5092
rect 15672 5080 15700 5111
rect 16206 5108 16212 5160
rect 16264 5148 16270 5160
rect 16758 5148 16764 5160
rect 16264 5120 16764 5148
rect 16264 5108 16270 5120
rect 16758 5108 16764 5120
rect 16816 5108 16822 5160
rect 16942 5148 16948 5160
rect 16903 5120 16948 5148
rect 16942 5108 16948 5120
rect 17000 5108 17006 5160
rect 17494 5108 17500 5160
rect 17552 5148 17558 5160
rect 18141 5151 18199 5157
rect 18141 5148 18153 5151
rect 17552 5120 18153 5148
rect 17552 5108 17558 5120
rect 18141 5117 18153 5120
rect 18187 5117 18199 5151
rect 18141 5111 18199 5117
rect 17512 5080 17540 5108
rect 15436 5052 17540 5080
rect 15436 5040 15442 5052
rect 12032 4984 12756 5012
rect 13081 5015 13139 5021
rect 12032 4972 12038 4984
rect 13081 4981 13093 5015
rect 13127 5012 13139 5015
rect 13446 5012 13452 5024
rect 13127 4984 13452 5012
rect 13127 4981 13139 4984
rect 13081 4975 13139 4981
rect 13446 4972 13452 4984
rect 13504 4972 13510 5024
rect 13998 5012 14004 5024
rect 13959 4984 14004 5012
rect 13998 4972 14004 4984
rect 14056 4972 14062 5024
rect 14182 4972 14188 5024
rect 14240 5012 14246 5024
rect 14550 5012 14556 5024
rect 14240 4984 14556 5012
rect 14240 4972 14246 4984
rect 14550 4972 14556 4984
rect 14608 4972 14614 5024
rect 15286 5012 15292 5024
rect 15247 4984 15292 5012
rect 15286 4972 15292 4984
rect 15344 4972 15350 5024
rect 16114 4972 16120 5024
rect 16172 5012 16178 5024
rect 16209 5015 16267 5021
rect 16209 5012 16221 5015
rect 16172 4984 16221 5012
rect 16172 4972 16178 4984
rect 16209 4981 16221 4984
rect 16255 4981 16267 5015
rect 17586 5012 17592 5024
rect 17547 4984 17592 5012
rect 16209 4975 16267 4981
rect 17586 4972 17592 4984
rect 17644 4972 17650 5024
rect 1104 4922 18860 4944
rect 1104 4870 3174 4922
rect 3226 4870 3238 4922
rect 3290 4870 3302 4922
rect 3354 4870 3366 4922
rect 3418 4870 3430 4922
rect 3482 4870 7622 4922
rect 7674 4870 7686 4922
rect 7738 4870 7750 4922
rect 7802 4870 7814 4922
rect 7866 4870 7878 4922
rect 7930 4870 12070 4922
rect 12122 4870 12134 4922
rect 12186 4870 12198 4922
rect 12250 4870 12262 4922
rect 12314 4870 12326 4922
rect 12378 4870 16518 4922
rect 16570 4870 16582 4922
rect 16634 4870 16646 4922
rect 16698 4870 16710 4922
rect 16762 4870 16774 4922
rect 16826 4870 18860 4922
rect 1104 4848 18860 4870
rect 1394 4768 1400 4820
rect 1452 4808 1458 4820
rect 1489 4811 1547 4817
rect 1489 4808 1501 4811
rect 1452 4780 1501 4808
rect 1452 4768 1458 4780
rect 1489 4777 1501 4780
rect 1535 4777 1547 4811
rect 1854 4808 1860 4820
rect 1815 4780 1860 4808
rect 1489 4771 1547 4777
rect 1854 4768 1860 4780
rect 1912 4768 1918 4820
rect 2222 4808 2228 4820
rect 2183 4780 2228 4808
rect 2222 4768 2228 4780
rect 2280 4768 2286 4820
rect 3786 4768 3792 4820
rect 3844 4808 3850 4820
rect 4157 4811 4215 4817
rect 4157 4808 4169 4811
rect 3844 4780 4169 4808
rect 3844 4768 3850 4780
rect 4157 4777 4169 4780
rect 4203 4777 4215 4811
rect 4157 4771 4215 4777
rect 4246 4768 4252 4820
rect 4304 4808 4310 4820
rect 4341 4811 4399 4817
rect 4341 4808 4353 4811
rect 4304 4780 4353 4808
rect 4304 4768 4310 4780
rect 4341 4777 4353 4780
rect 4387 4777 4399 4811
rect 4341 4771 4399 4777
rect 4430 4768 4436 4820
rect 4488 4808 4494 4820
rect 4525 4811 4583 4817
rect 4525 4808 4537 4811
rect 4488 4780 4537 4808
rect 4488 4768 4494 4780
rect 4525 4777 4537 4780
rect 4571 4777 4583 4811
rect 4798 4808 4804 4820
rect 4759 4780 4804 4808
rect 4525 4771 4583 4777
rect 4798 4768 4804 4780
rect 4856 4768 4862 4820
rect 5166 4768 5172 4820
rect 5224 4808 5230 4820
rect 5629 4811 5687 4817
rect 5629 4808 5641 4811
rect 5224 4780 5641 4808
rect 5224 4768 5230 4780
rect 5629 4777 5641 4780
rect 5675 4777 5687 4811
rect 5629 4771 5687 4777
rect 6178 4768 6184 4820
rect 6236 4808 6242 4820
rect 6236 4780 6316 4808
rect 6236 4768 6242 4780
rect 3970 4740 3976 4752
rect 3931 4712 3976 4740
rect 3970 4700 3976 4712
rect 4028 4700 4034 4752
rect 5994 4700 6000 4752
rect 6052 4740 6058 4752
rect 6288 4740 6316 4780
rect 6362 4768 6368 4820
rect 6420 4808 6426 4820
rect 8202 4808 8208 4820
rect 6420 4780 8208 4808
rect 6420 4768 6426 4780
rect 8202 4768 8208 4780
rect 8260 4768 8266 4820
rect 8754 4768 8760 4820
rect 8812 4808 8818 4820
rect 9861 4811 9919 4817
rect 9861 4808 9873 4811
rect 8812 4780 9873 4808
rect 8812 4768 8818 4780
rect 9861 4777 9873 4780
rect 9907 4777 9919 4811
rect 11790 4808 11796 4820
rect 11751 4780 11796 4808
rect 9861 4771 9919 4777
rect 11790 4768 11796 4780
rect 11848 4768 11854 4820
rect 12342 4768 12348 4820
rect 12400 4808 12406 4820
rect 12894 4808 12900 4820
rect 12400 4780 12900 4808
rect 12400 4768 12406 4780
rect 12894 4768 12900 4780
rect 12952 4768 12958 4820
rect 13906 4768 13912 4820
rect 13964 4808 13970 4820
rect 15378 4808 15384 4820
rect 13964 4780 14412 4808
rect 13964 4768 13970 4780
rect 6457 4743 6515 4749
rect 6457 4740 6469 4743
rect 6052 4712 6224 4740
rect 6288 4712 6469 4740
rect 6052 4700 6058 4712
rect 2682 4672 2688 4684
rect 2056 4644 2688 4672
rect 1670 4604 1676 4616
rect 1631 4576 1676 4604
rect 1670 4564 1676 4576
rect 1728 4564 1734 4616
rect 2056 4613 2084 4644
rect 2682 4632 2688 4644
rect 2740 4632 2746 4684
rect 4338 4672 4344 4684
rect 2792 4644 4344 4672
rect 2041 4607 2099 4613
rect 2041 4573 2053 4607
rect 2087 4573 2099 4607
rect 2406 4604 2412 4616
rect 2367 4576 2412 4604
rect 2041 4567 2099 4573
rect 2406 4564 2412 4576
rect 2464 4564 2470 4616
rect 2792 4613 2820 4644
rect 4338 4632 4344 4644
rect 4396 4632 4402 4684
rect 5626 4632 5632 4684
rect 5684 4672 5690 4684
rect 6196 4681 6224 4712
rect 6457 4709 6469 4712
rect 6503 4709 6515 4743
rect 9674 4740 9680 4752
rect 6457 4703 6515 4709
rect 7300 4712 9680 4740
rect 7300 4681 7328 4712
rect 9674 4700 9680 4712
rect 9732 4700 9738 4752
rect 11698 4740 11704 4752
rect 11659 4712 11704 4740
rect 11698 4700 11704 4712
rect 11756 4700 11762 4752
rect 13814 4700 13820 4752
rect 13872 4740 13878 4752
rect 13872 4712 14320 4740
rect 13872 4700 13878 4712
rect 6089 4675 6147 4681
rect 6089 4672 6101 4675
rect 5684 4644 6101 4672
rect 5684 4632 5690 4644
rect 6089 4641 6101 4644
rect 6135 4641 6147 4675
rect 6089 4635 6147 4641
rect 6181 4675 6239 4681
rect 6181 4641 6193 4675
rect 6227 4641 6239 4675
rect 6181 4635 6239 4641
rect 7285 4675 7343 4681
rect 7285 4641 7297 4675
rect 7331 4641 7343 4675
rect 8018 4672 8024 4684
rect 7979 4644 8024 4672
rect 7285 4635 7343 4641
rect 8018 4632 8024 4644
rect 8076 4672 8082 4684
rect 9585 4675 9643 4681
rect 9585 4672 9597 4675
rect 8076 4644 9597 4672
rect 8076 4632 8082 4644
rect 9585 4641 9597 4644
rect 9631 4672 9643 4675
rect 10134 4672 10140 4684
rect 9631 4644 10140 4672
rect 9631 4641 9643 4644
rect 9585 4635 9643 4641
rect 10134 4632 10140 4644
rect 10192 4632 10198 4684
rect 10502 4672 10508 4684
rect 10463 4644 10508 4672
rect 10502 4632 10508 4644
rect 10560 4632 10566 4684
rect 10778 4672 10784 4684
rect 10739 4644 10784 4672
rect 10778 4632 10784 4644
rect 10836 4632 10842 4684
rect 10965 4675 11023 4681
rect 10965 4641 10977 4675
rect 11011 4672 11023 4675
rect 11330 4672 11336 4684
rect 11011 4644 11336 4672
rect 11011 4641 11023 4644
rect 10965 4635 11023 4641
rect 11330 4632 11336 4644
rect 11388 4632 11394 4684
rect 12802 4672 12808 4684
rect 12763 4644 12808 4672
rect 12802 4632 12808 4644
rect 12860 4632 12866 4684
rect 13446 4672 13452 4684
rect 13407 4644 13452 4672
rect 13446 4632 13452 4644
rect 13504 4632 13510 4684
rect 13633 4675 13691 4681
rect 13633 4641 13645 4675
rect 13679 4672 13691 4675
rect 14182 4672 14188 4684
rect 13679 4644 14188 4672
rect 13679 4641 13691 4644
rect 13633 4635 13691 4641
rect 14182 4632 14188 4644
rect 14240 4632 14246 4684
rect 2777 4607 2835 4613
rect 2777 4573 2789 4607
rect 2823 4573 2835 4607
rect 2777 4567 2835 4573
rect 3053 4607 3111 4613
rect 3053 4573 3065 4607
rect 3099 4573 3111 4607
rect 3326 4604 3332 4616
rect 3287 4576 3332 4604
rect 3053 4567 3111 4573
rect 3068 4536 3096 4567
rect 3326 4564 3332 4576
rect 3384 4564 3390 4616
rect 3602 4604 3608 4616
rect 3563 4576 3608 4604
rect 3602 4564 3608 4576
rect 3660 4564 3666 4616
rect 3786 4604 3792 4616
rect 3747 4576 3792 4604
rect 3786 4564 3792 4576
rect 3844 4564 3850 4616
rect 4982 4604 4988 4616
rect 4943 4576 4988 4604
rect 4982 4564 4988 4576
rect 5040 4564 5046 4616
rect 5074 4564 5080 4616
rect 5132 4604 5138 4616
rect 5997 4607 6055 4613
rect 5997 4604 6009 4607
rect 5132 4576 6009 4604
rect 5132 4564 5138 4576
rect 5997 4573 6009 4576
rect 6043 4604 6055 4607
rect 6454 4604 6460 4616
rect 6043 4576 6460 4604
rect 6043 4573 6055 4576
rect 5997 4567 6055 4573
rect 6454 4564 6460 4576
rect 6512 4564 6518 4616
rect 8754 4604 8760 4616
rect 6840 4576 8760 4604
rect 4154 4536 4160 4548
rect 3068 4508 4160 4536
rect 4154 4496 4160 4508
rect 4212 4496 4218 4548
rect 4522 4496 4528 4548
rect 4580 4536 4586 4548
rect 6840 4536 6868 4576
rect 8754 4564 8760 4576
rect 8812 4604 8818 4616
rect 9401 4607 9459 4613
rect 9401 4604 9413 4607
rect 8812 4576 9413 4604
rect 8812 4564 8818 4576
rect 9401 4573 9413 4576
rect 9447 4573 9459 4607
rect 9401 4567 9459 4573
rect 9493 4607 9551 4613
rect 9493 4573 9505 4607
rect 9539 4604 9551 4607
rect 10226 4604 10232 4616
rect 9539 4576 10232 4604
rect 9539 4573 9551 4576
rect 9493 4567 9551 4573
rect 10226 4564 10232 4576
rect 10284 4564 10290 4616
rect 10321 4607 10379 4613
rect 10321 4573 10333 4607
rect 10367 4604 10379 4607
rect 10686 4604 10692 4616
rect 10367 4576 10692 4604
rect 10367 4573 10379 4576
rect 10321 4567 10379 4573
rect 10686 4564 10692 4576
rect 10744 4564 10750 4616
rect 11054 4604 11060 4616
rect 11015 4576 11060 4604
rect 11054 4564 11060 4576
rect 11112 4564 11118 4616
rect 11882 4564 11888 4616
rect 11940 4604 11946 4616
rect 11977 4607 12035 4613
rect 11977 4604 11989 4607
rect 11940 4576 11989 4604
rect 11940 4564 11946 4576
rect 11977 4573 11989 4576
rect 12023 4573 12035 4607
rect 11977 4567 12035 4573
rect 12529 4607 12587 4613
rect 12529 4573 12541 4607
rect 12575 4604 12587 4607
rect 13998 4604 14004 4616
rect 12575 4576 14004 4604
rect 12575 4573 12587 4576
rect 12529 4567 12587 4573
rect 13998 4564 14004 4576
rect 14056 4564 14062 4616
rect 14090 4564 14096 4616
rect 14148 4604 14154 4616
rect 14292 4604 14320 4712
rect 14384 4672 14412 4780
rect 15028 4780 15384 4808
rect 15028 4681 15056 4780
rect 15378 4768 15384 4780
rect 15436 4768 15442 4820
rect 15470 4768 15476 4820
rect 15528 4808 15534 4820
rect 17034 4808 17040 4820
rect 15528 4780 17040 4808
rect 15528 4768 15534 4780
rect 17034 4768 17040 4780
rect 17092 4768 17098 4820
rect 17681 4811 17739 4817
rect 17681 4777 17693 4811
rect 17727 4808 17739 4811
rect 17770 4808 17776 4820
rect 17727 4780 17776 4808
rect 17727 4777 17739 4780
rect 17681 4771 17739 4777
rect 17770 4768 17776 4780
rect 17828 4768 17834 4820
rect 18049 4811 18107 4817
rect 18049 4777 18061 4811
rect 18095 4808 18107 4811
rect 18138 4808 18144 4820
rect 18095 4780 18144 4808
rect 18095 4777 18107 4780
rect 18049 4771 18107 4777
rect 18138 4768 18144 4780
rect 18196 4768 18202 4820
rect 18414 4808 18420 4820
rect 18375 4780 18420 4808
rect 18414 4768 18420 4780
rect 18472 4768 18478 4820
rect 16577 4743 16635 4749
rect 16577 4740 16589 4743
rect 15212 4712 16589 4740
rect 15212 4681 15240 4712
rect 16577 4709 16589 4712
rect 16623 4709 16635 4743
rect 16577 4703 16635 4709
rect 14645 4675 14703 4681
rect 14645 4672 14657 4675
rect 14384 4644 14657 4672
rect 14645 4641 14657 4644
rect 14691 4641 14703 4675
rect 14645 4635 14703 4641
rect 15013 4675 15071 4681
rect 15013 4641 15025 4675
rect 15059 4641 15071 4675
rect 15013 4635 15071 4641
rect 15197 4675 15255 4681
rect 15197 4641 15209 4675
rect 15243 4641 15255 4675
rect 15197 4635 15255 4641
rect 16022 4632 16028 4684
rect 16080 4672 16086 4684
rect 16301 4675 16359 4681
rect 16301 4672 16313 4675
rect 16080 4644 16313 4672
rect 16080 4632 16086 4644
rect 16301 4641 16313 4644
rect 16347 4641 16359 4675
rect 16301 4635 16359 4641
rect 17221 4675 17279 4681
rect 17221 4641 17233 4675
rect 17267 4672 17279 4675
rect 18782 4672 18788 4684
rect 17267 4644 18788 4672
rect 17267 4641 17279 4644
rect 17221 4635 17279 4641
rect 18782 4632 18788 4644
rect 18840 4632 18846 4684
rect 14461 4607 14519 4613
rect 14461 4604 14473 4607
rect 14148 4576 14228 4604
rect 14292 4576 14473 4604
rect 14148 4564 14154 4576
rect 4580 4508 6868 4536
rect 4580 4496 4586 4508
rect 6914 4496 6920 4548
rect 6972 4536 6978 4548
rect 7837 4539 7895 4545
rect 6972 4508 7604 4536
rect 6972 4496 6978 4508
rect 2593 4471 2651 4477
rect 2593 4437 2605 4471
rect 2639 4468 2651 4471
rect 2774 4468 2780 4480
rect 2639 4440 2780 4468
rect 2639 4437 2651 4440
rect 2593 4431 2651 4437
rect 2774 4428 2780 4440
rect 2832 4428 2838 4480
rect 2869 4471 2927 4477
rect 2869 4437 2881 4471
rect 2915 4468 2927 4471
rect 2958 4468 2964 4480
rect 2915 4440 2964 4468
rect 2915 4437 2927 4440
rect 2869 4431 2927 4437
rect 2958 4428 2964 4440
rect 3016 4428 3022 4480
rect 3050 4428 3056 4480
rect 3108 4468 3114 4480
rect 3145 4471 3203 4477
rect 3145 4468 3157 4471
rect 3108 4440 3157 4468
rect 3108 4428 3114 4440
rect 3145 4437 3157 4440
rect 3191 4437 3203 4471
rect 3145 4431 3203 4437
rect 3421 4471 3479 4477
rect 3421 4437 3433 4471
rect 3467 4468 3479 4471
rect 3602 4468 3608 4480
rect 3467 4440 3608 4468
rect 3467 4437 3479 4440
rect 3421 4431 3479 4437
rect 3602 4428 3608 4440
rect 3660 4428 3666 4480
rect 5166 4468 5172 4480
rect 5127 4440 5172 4468
rect 5166 4428 5172 4440
rect 5224 4428 5230 4480
rect 6638 4468 6644 4480
rect 6599 4440 6644 4468
rect 6638 4428 6644 4440
rect 6696 4428 6702 4480
rect 7006 4468 7012 4480
rect 6967 4440 7012 4468
rect 7006 4428 7012 4440
rect 7064 4428 7070 4480
rect 7098 4428 7104 4480
rect 7156 4468 7162 4480
rect 7156 4440 7201 4468
rect 7156 4428 7162 4440
rect 7374 4428 7380 4480
rect 7432 4468 7438 4480
rect 7469 4471 7527 4477
rect 7469 4468 7481 4471
rect 7432 4440 7481 4468
rect 7432 4428 7438 4440
rect 7469 4437 7481 4440
rect 7515 4437 7527 4471
rect 7576 4468 7604 4508
rect 7837 4505 7849 4539
rect 7883 4536 7895 4539
rect 8297 4539 8355 4545
rect 8297 4536 8309 4539
rect 7883 4508 8309 4536
rect 7883 4505 7895 4508
rect 7837 4499 7895 4505
rect 8297 4505 8309 4508
rect 8343 4505 8355 4539
rect 8297 4499 8355 4505
rect 13357 4539 13415 4545
rect 13357 4505 13369 4539
rect 13403 4536 13415 4539
rect 14200 4536 14228 4576
rect 14461 4573 14473 4576
rect 14507 4604 14519 4607
rect 15102 4604 15108 4616
rect 14507 4576 15108 4604
rect 14507 4573 14519 4576
rect 14461 4567 14519 4573
rect 15102 4564 15108 4576
rect 15160 4564 15166 4616
rect 16114 4604 16120 4616
rect 16075 4576 16120 4604
rect 16114 4564 16120 4576
rect 16172 4564 16178 4616
rect 16850 4564 16856 4616
rect 16908 4604 16914 4616
rect 16945 4607 17003 4613
rect 16945 4604 16957 4607
rect 16908 4576 16957 4604
rect 16908 4564 16914 4576
rect 16945 4573 16957 4576
rect 16991 4573 17003 4607
rect 16945 4567 17003 4573
rect 17034 4564 17040 4616
rect 17092 4604 17098 4616
rect 17497 4607 17555 4613
rect 17497 4604 17509 4607
rect 17092 4576 17509 4604
rect 17092 4564 17098 4576
rect 17497 4573 17509 4576
rect 17543 4573 17555 4607
rect 17497 4567 17555 4573
rect 17865 4607 17923 4613
rect 17865 4573 17877 4607
rect 17911 4573 17923 4607
rect 18230 4604 18236 4616
rect 18191 4576 18236 4604
rect 17865 4567 17923 4573
rect 14366 4536 14372 4548
rect 13403 4508 14136 4536
rect 14200 4508 14372 4536
rect 13403 4505 13415 4508
rect 13357 4499 13415 4505
rect 7929 4471 7987 4477
rect 7929 4468 7941 4471
rect 7576 4440 7941 4468
rect 7469 4431 7527 4437
rect 7929 4437 7941 4440
rect 7975 4468 7987 4471
rect 8386 4468 8392 4480
rect 7975 4440 8392 4468
rect 7975 4437 7987 4440
rect 7929 4431 7987 4437
rect 8386 4428 8392 4440
rect 8444 4468 8450 4480
rect 8570 4468 8576 4480
rect 8444 4440 8576 4468
rect 8444 4428 8450 4440
rect 8570 4428 8576 4440
rect 8628 4428 8634 4480
rect 9033 4471 9091 4477
rect 9033 4437 9045 4471
rect 9079 4468 9091 4471
rect 9306 4468 9312 4480
rect 9079 4440 9312 4468
rect 9079 4437 9091 4440
rect 9033 4431 9091 4437
rect 9306 4428 9312 4440
rect 9364 4428 9370 4480
rect 10229 4471 10287 4477
rect 10229 4437 10241 4471
rect 10275 4468 10287 4471
rect 10410 4468 10416 4480
rect 10275 4440 10416 4468
rect 10275 4437 10287 4440
rect 10229 4431 10287 4437
rect 10410 4428 10416 4440
rect 10468 4428 10474 4480
rect 11422 4468 11428 4480
rect 11383 4440 11428 4468
rect 11422 4428 11428 4440
rect 11480 4428 11486 4480
rect 11698 4428 11704 4480
rect 11756 4468 11762 4480
rect 12161 4471 12219 4477
rect 12161 4468 12173 4471
rect 11756 4440 12173 4468
rect 11756 4428 11762 4440
rect 12161 4437 12173 4440
rect 12207 4437 12219 4471
rect 12161 4431 12219 4437
rect 12621 4471 12679 4477
rect 12621 4437 12633 4471
rect 12667 4468 12679 4471
rect 12989 4471 13047 4477
rect 12989 4468 13001 4471
rect 12667 4440 13001 4468
rect 12667 4437 12679 4440
rect 12621 4431 12679 4437
rect 12989 4437 13001 4440
rect 13035 4437 13047 4471
rect 12989 4431 13047 4437
rect 13630 4428 13636 4480
rect 13688 4468 13694 4480
rect 14108 4477 14136 4508
rect 14366 4496 14372 4508
rect 14424 4496 14430 4548
rect 14553 4539 14611 4545
rect 14553 4505 14565 4539
rect 14599 4536 14611 4539
rect 15194 4536 15200 4548
rect 14599 4508 15200 4536
rect 14599 4505 14611 4508
rect 14553 4499 14611 4505
rect 15194 4496 15200 4508
rect 15252 4496 15258 4548
rect 16209 4539 16267 4545
rect 16209 4536 16221 4539
rect 15672 4508 16221 4536
rect 13817 4471 13875 4477
rect 13817 4468 13829 4471
rect 13688 4440 13829 4468
rect 13688 4428 13694 4440
rect 13817 4437 13829 4440
rect 13863 4437 13875 4471
rect 13817 4431 13875 4437
rect 14093 4471 14151 4477
rect 14093 4437 14105 4471
rect 14139 4437 14151 4471
rect 14093 4431 14151 4437
rect 14274 4428 14280 4480
rect 14332 4468 14338 4480
rect 15672 4477 15700 4508
rect 16209 4505 16221 4508
rect 16255 4505 16267 4539
rect 16209 4499 16267 4505
rect 16574 4496 16580 4548
rect 16632 4536 16638 4548
rect 17880 4536 17908 4567
rect 18230 4564 18236 4576
rect 18288 4564 18294 4616
rect 16632 4508 17908 4536
rect 16632 4496 16638 4508
rect 15289 4471 15347 4477
rect 15289 4468 15301 4471
rect 14332 4440 15301 4468
rect 14332 4428 14338 4440
rect 15289 4437 15301 4440
rect 15335 4437 15347 4471
rect 15289 4431 15347 4437
rect 15657 4471 15715 4477
rect 15657 4437 15669 4471
rect 15703 4437 15715 4471
rect 15657 4431 15715 4437
rect 15746 4428 15752 4480
rect 15804 4468 15810 4480
rect 15804 4440 15849 4468
rect 15804 4428 15810 4440
rect 16758 4428 16764 4480
rect 16816 4468 16822 4480
rect 17037 4471 17095 4477
rect 17037 4468 17049 4471
rect 16816 4440 17049 4468
rect 16816 4428 16822 4440
rect 17037 4437 17049 4440
rect 17083 4468 17095 4471
rect 17494 4468 17500 4480
rect 17083 4440 17500 4468
rect 17083 4437 17095 4440
rect 17037 4431 17095 4437
rect 17494 4428 17500 4440
rect 17552 4428 17558 4480
rect 1104 4378 18860 4400
rect 1104 4326 5398 4378
rect 5450 4326 5462 4378
rect 5514 4326 5526 4378
rect 5578 4326 5590 4378
rect 5642 4326 5654 4378
rect 5706 4326 9846 4378
rect 9898 4326 9910 4378
rect 9962 4326 9974 4378
rect 10026 4326 10038 4378
rect 10090 4326 10102 4378
rect 10154 4326 14294 4378
rect 14346 4326 14358 4378
rect 14410 4326 14422 4378
rect 14474 4326 14486 4378
rect 14538 4326 14550 4378
rect 14602 4326 18860 4378
rect 1104 4304 18860 4326
rect 1486 4264 1492 4276
rect 1447 4236 1492 4264
rect 1486 4224 1492 4236
rect 1544 4224 1550 4276
rect 1854 4264 1860 4276
rect 1815 4236 1860 4264
rect 1854 4224 1860 4236
rect 1912 4224 1918 4276
rect 3510 4224 3516 4276
rect 3568 4264 3574 4276
rect 3697 4267 3755 4273
rect 3697 4264 3709 4267
rect 3568 4236 3709 4264
rect 3568 4224 3574 4236
rect 3697 4233 3709 4236
rect 3743 4233 3755 4267
rect 3697 4227 3755 4233
rect 3786 4224 3792 4276
rect 3844 4264 3850 4276
rect 3881 4267 3939 4273
rect 3881 4264 3893 4267
rect 3844 4236 3893 4264
rect 3844 4224 3850 4236
rect 3881 4233 3893 4236
rect 3927 4233 3939 4267
rect 3881 4227 3939 4233
rect 5994 4224 6000 4276
rect 6052 4264 6058 4276
rect 6365 4267 6423 4273
rect 6365 4264 6377 4267
rect 6052 4236 6377 4264
rect 6052 4224 6058 4236
rect 6365 4233 6377 4236
rect 6411 4264 6423 4267
rect 6549 4267 6607 4273
rect 6549 4264 6561 4267
rect 6411 4236 6561 4264
rect 6411 4233 6423 4236
rect 6365 4227 6423 4233
rect 6549 4233 6561 4236
rect 6595 4233 6607 4267
rect 7006 4264 7012 4276
rect 6967 4236 7012 4264
rect 6549 4227 6607 4233
rect 7006 4224 7012 4236
rect 7064 4224 7070 4276
rect 7374 4264 7380 4276
rect 7335 4236 7380 4264
rect 7374 4224 7380 4236
rect 7432 4224 7438 4276
rect 7466 4224 7472 4276
rect 7524 4264 7530 4276
rect 8754 4264 8760 4276
rect 7524 4236 7569 4264
rect 8715 4236 8760 4264
rect 7524 4224 7530 4236
rect 8754 4224 8760 4236
rect 8812 4224 8818 4276
rect 9306 4264 9312 4276
rect 9267 4236 9312 4264
rect 9306 4224 9312 4236
rect 9364 4224 9370 4276
rect 9401 4267 9459 4273
rect 9401 4233 9413 4267
rect 9447 4264 9459 4267
rect 9582 4264 9588 4276
rect 9447 4236 9588 4264
rect 9447 4233 9459 4236
rect 9401 4227 9459 4233
rect 9582 4224 9588 4236
rect 9640 4224 9646 4276
rect 10781 4267 10839 4273
rect 10781 4233 10793 4267
rect 10827 4264 10839 4267
rect 11974 4264 11980 4276
rect 10827 4236 11980 4264
rect 10827 4233 10839 4236
rect 10781 4227 10839 4233
rect 11974 4224 11980 4236
rect 12032 4224 12038 4276
rect 12710 4264 12716 4276
rect 12452 4236 12716 4264
rect 3326 4156 3332 4208
rect 3384 4196 3390 4208
rect 6914 4196 6920 4208
rect 3384 4168 4292 4196
rect 6875 4168 6920 4196
rect 3384 4156 3390 4168
rect 1673 4131 1731 4137
rect 1673 4097 1685 4131
rect 1719 4097 1731 4131
rect 1673 4091 1731 4097
rect 2041 4131 2099 4137
rect 2041 4097 2053 4131
rect 2087 4128 2099 4131
rect 2130 4128 2136 4140
rect 2087 4100 2136 4128
rect 2087 4097 2099 4100
rect 2041 4091 2099 4097
rect 1688 4060 1716 4091
rect 2130 4088 2136 4100
rect 2188 4088 2194 4140
rect 2406 4128 2412 4140
rect 2367 4100 2412 4128
rect 2406 4088 2412 4100
rect 2464 4088 2470 4140
rect 2682 4128 2688 4140
rect 2643 4100 2688 4128
rect 2682 4088 2688 4100
rect 2740 4088 2746 4140
rect 2961 4131 3019 4137
rect 2961 4097 2973 4131
rect 3007 4097 3019 4131
rect 2961 4091 3019 4097
rect 3237 4131 3295 4137
rect 3237 4097 3249 4131
rect 3283 4097 3295 4131
rect 3418 4128 3424 4140
rect 3379 4100 3424 4128
rect 3237 4091 3295 4097
rect 1688 4032 2544 4060
rect 2516 4001 2544 4032
rect 2501 3995 2559 4001
rect 2501 3961 2513 3995
rect 2547 3961 2559 3995
rect 2501 3955 2559 3961
rect 2590 3952 2596 4004
rect 2648 3992 2654 4004
rect 2976 3992 3004 4091
rect 3252 4060 3280 4091
rect 3418 4088 3424 4100
rect 3476 4088 3482 4140
rect 3605 4131 3663 4137
rect 3605 4097 3617 4131
rect 3651 4128 3663 4131
rect 3878 4128 3884 4140
rect 3651 4100 3884 4128
rect 3651 4097 3663 4100
rect 3605 4091 3663 4097
rect 3878 4088 3884 4100
rect 3936 4088 3942 4140
rect 4154 4128 4160 4140
rect 4115 4100 4160 4128
rect 4154 4088 4160 4100
rect 4212 4088 4218 4140
rect 4264 4128 4292 4168
rect 6914 4156 6920 4168
rect 6972 4196 6978 4208
rect 7837 4199 7895 4205
rect 7837 4196 7849 4199
rect 6972 4168 7849 4196
rect 6972 4156 6978 4168
rect 7837 4165 7849 4168
rect 7883 4196 7895 4199
rect 8202 4196 8208 4208
rect 7883 4168 8208 4196
rect 7883 4165 7895 4168
rect 7837 4159 7895 4165
rect 8202 4156 8208 4168
rect 8260 4156 8266 4208
rect 10410 4196 10416 4208
rect 10371 4168 10416 4196
rect 10410 4156 10416 4168
rect 10468 4156 10474 4208
rect 10502 4156 10508 4208
rect 10560 4196 10566 4208
rect 10560 4168 10640 4196
rect 10560 4156 10566 4168
rect 4341 4131 4399 4137
rect 4341 4128 4353 4131
rect 4264 4100 4353 4128
rect 4341 4097 4353 4100
rect 4387 4128 4399 4131
rect 6178 4128 6184 4140
rect 4387 4100 6184 4128
rect 4387 4097 4399 4100
rect 4341 4091 4399 4097
rect 6178 4088 6184 4100
rect 6236 4088 6242 4140
rect 10428 4128 10456 4156
rect 10612 4137 10640 4168
rect 7484 4100 10456 4128
rect 10597 4131 10655 4137
rect 7484 4060 7512 4100
rect 10597 4097 10609 4131
rect 10643 4097 10655 4131
rect 11514 4128 11520 4140
rect 11475 4100 11520 4128
rect 10597 4091 10655 4097
rect 11514 4088 11520 4100
rect 11572 4088 11578 4140
rect 12253 4131 12311 4137
rect 12253 4097 12265 4131
rect 12299 4128 12311 4131
rect 12452 4128 12480 4236
rect 12710 4224 12716 4236
rect 12768 4224 12774 4276
rect 13262 4264 13268 4276
rect 13223 4236 13268 4264
rect 13262 4224 13268 4236
rect 13320 4224 13326 4276
rect 13722 4264 13728 4276
rect 13683 4236 13728 4264
rect 13722 4224 13728 4236
rect 13780 4224 13786 4276
rect 14090 4264 14096 4276
rect 14051 4236 14096 4264
rect 14090 4224 14096 4236
rect 14148 4224 14154 4276
rect 15105 4267 15163 4273
rect 15105 4233 15117 4267
rect 15151 4264 15163 4267
rect 15565 4267 15623 4273
rect 15565 4264 15577 4267
rect 15151 4236 15577 4264
rect 15151 4233 15163 4236
rect 15105 4227 15163 4233
rect 15565 4233 15577 4236
rect 15611 4233 15623 4267
rect 15565 4227 15623 4233
rect 15933 4267 15991 4273
rect 15933 4233 15945 4267
rect 15979 4264 15991 4267
rect 17586 4264 17592 4276
rect 15979 4236 17592 4264
rect 15979 4233 15991 4236
rect 15933 4227 15991 4233
rect 17586 4224 17592 4236
rect 17644 4224 17650 4276
rect 17678 4224 17684 4276
rect 17736 4264 17742 4276
rect 17736 4236 17781 4264
rect 17736 4224 17742 4236
rect 12526 4156 12532 4208
rect 12584 4196 12590 4208
rect 13906 4196 13912 4208
rect 12584 4168 13912 4196
rect 12584 4156 12590 4168
rect 12299 4100 12480 4128
rect 12299 4097 12311 4100
rect 12253 4091 12311 4097
rect 3252 4032 7512 4060
rect 7653 4063 7711 4069
rect 7653 4029 7665 4063
rect 7699 4060 7711 4063
rect 8294 4060 8300 4072
rect 7699 4032 8300 4060
rect 7699 4029 7711 4032
rect 7653 4023 7711 4029
rect 8294 4020 8300 4032
rect 8352 4020 8358 4072
rect 8389 4063 8447 4069
rect 8389 4029 8401 4063
rect 8435 4060 8447 4063
rect 8570 4060 8576 4072
rect 8435 4032 8576 4060
rect 8435 4029 8447 4032
rect 8389 4023 8447 4029
rect 8570 4020 8576 4032
rect 8628 4060 8634 4072
rect 8628 4032 9076 4060
rect 8628 4020 8634 4032
rect 4525 3995 4583 4001
rect 4525 3992 4537 3995
rect 2648 3964 2912 3992
rect 2976 3964 4537 3992
rect 2648 3952 2654 3964
rect 2222 3924 2228 3936
rect 2183 3896 2228 3924
rect 2222 3884 2228 3896
rect 2280 3884 2286 3936
rect 2314 3884 2320 3936
rect 2372 3924 2378 3936
rect 2777 3927 2835 3933
rect 2777 3924 2789 3927
rect 2372 3896 2789 3924
rect 2372 3884 2378 3896
rect 2777 3893 2789 3896
rect 2823 3893 2835 3927
rect 2884 3924 2912 3964
rect 4525 3961 4537 3964
rect 4571 3992 4583 3995
rect 4614 3992 4620 4004
rect 4571 3964 4620 3992
rect 4571 3961 4583 3964
rect 4525 3955 4583 3961
rect 4614 3952 4620 3964
rect 4672 3992 4678 4004
rect 4672 3964 6960 3992
rect 4672 3952 4678 3964
rect 3053 3927 3111 3933
rect 3053 3924 3065 3927
rect 2884 3896 3065 3924
rect 2777 3887 2835 3893
rect 3053 3893 3065 3896
rect 3099 3893 3111 3927
rect 6932 3924 6960 3964
rect 7098 3952 7104 4004
rect 7156 3992 7162 4004
rect 8941 3995 8999 4001
rect 8941 3992 8953 3995
rect 7156 3964 8953 3992
rect 7156 3952 7162 3964
rect 8941 3961 8953 3964
rect 8987 3961 8999 3995
rect 9048 3992 9076 4032
rect 9122 4020 9128 4072
rect 9180 4060 9186 4072
rect 9490 4060 9496 4072
rect 9180 4032 9496 4060
rect 9180 4020 9186 4032
rect 9490 4020 9496 4032
rect 9548 4020 9554 4072
rect 11974 4060 11980 4072
rect 9600 4032 11980 4060
rect 9600 3992 9628 4032
rect 11974 4020 11980 4032
rect 12032 4020 12038 4072
rect 12636 4069 12664 4168
rect 12894 4128 12900 4140
rect 12855 4100 12900 4128
rect 12894 4088 12900 4100
rect 12952 4088 12958 4140
rect 12986 4088 12992 4140
rect 13044 4088 13050 4140
rect 12621 4063 12679 4069
rect 12621 4029 12633 4063
rect 12667 4029 12679 4063
rect 12621 4023 12679 4029
rect 12805 4063 12863 4069
rect 12805 4029 12817 4063
rect 12851 4060 12863 4063
rect 13004 4060 13032 4088
rect 13556 4069 13584 4168
rect 13906 4156 13912 4168
rect 13964 4156 13970 4208
rect 13998 4156 14004 4208
rect 14056 4196 14062 4208
rect 15197 4199 15255 4205
rect 14056 4168 14780 4196
rect 14056 4156 14062 4168
rect 14182 4128 14188 4140
rect 14143 4100 14188 4128
rect 14182 4088 14188 4100
rect 14240 4088 14246 4140
rect 14476 4137 14504 4168
rect 14461 4131 14519 4137
rect 14461 4097 14473 4131
rect 14507 4097 14519 4131
rect 14461 4091 14519 4097
rect 14642 4088 14648 4140
rect 14700 4088 14706 4140
rect 14752 4128 14780 4168
rect 15197 4165 15209 4199
rect 15243 4196 15255 4199
rect 15746 4196 15752 4208
rect 15243 4168 15752 4196
rect 15243 4165 15255 4168
rect 15197 4159 15255 4165
rect 15746 4156 15752 4168
rect 15804 4156 15810 4208
rect 17402 4196 17408 4208
rect 15856 4168 17408 4196
rect 15856 4128 15884 4168
rect 17402 4156 17408 4168
rect 17460 4156 17466 4208
rect 14752 4100 15884 4128
rect 16025 4131 16083 4137
rect 16025 4097 16037 4131
rect 16071 4128 16083 4131
rect 16390 4128 16396 4140
rect 16071 4100 16396 4128
rect 16071 4097 16083 4100
rect 16025 4091 16083 4097
rect 16390 4088 16396 4100
rect 16448 4088 16454 4140
rect 16758 4128 16764 4140
rect 16719 4100 16764 4128
rect 16758 4088 16764 4100
rect 16816 4088 16822 4140
rect 17126 4128 17132 4140
rect 17087 4100 17132 4128
rect 17126 4088 17132 4100
rect 17184 4088 17190 4140
rect 17497 4131 17555 4137
rect 17497 4097 17509 4131
rect 17543 4097 17555 4131
rect 17497 4091 17555 4097
rect 17865 4131 17923 4137
rect 17865 4097 17877 4131
rect 17911 4097 17923 4131
rect 18230 4128 18236 4140
rect 18191 4100 18236 4128
rect 17865 4091 17923 4097
rect 13541 4063 13599 4069
rect 12851 4032 13492 4060
rect 12851 4029 12863 4032
rect 12805 4023 12863 4029
rect 10502 3992 10508 4004
rect 9048 3964 9628 3992
rect 10152 3964 10508 3992
rect 8941 3955 8999 3961
rect 7742 3924 7748 3936
rect 6932 3896 7748 3924
rect 3053 3887 3111 3893
rect 7742 3884 7748 3896
rect 7800 3884 7806 3936
rect 8110 3924 8116 3936
rect 8071 3896 8116 3924
rect 8110 3884 8116 3896
rect 8168 3884 8174 3936
rect 8294 3884 8300 3936
rect 8352 3924 8358 3936
rect 9122 3924 9128 3936
rect 8352 3896 9128 3924
rect 8352 3884 8358 3896
rect 9122 3884 9128 3896
rect 9180 3884 9186 3936
rect 9214 3884 9220 3936
rect 9272 3924 9278 3936
rect 10152 3924 10180 3964
rect 10502 3952 10508 3964
rect 10560 3952 10566 4004
rect 12161 3995 12219 4001
rect 12161 3961 12173 3995
rect 12207 3992 12219 3995
rect 12342 3992 12348 4004
rect 12207 3964 12348 3992
rect 12207 3961 12219 3964
rect 12161 3955 12219 3961
rect 12342 3952 12348 3964
rect 12400 3992 12406 4004
rect 12986 3992 12992 4004
rect 12400 3964 12992 3992
rect 12400 3952 12406 3964
rect 12986 3952 12992 3964
rect 13044 3952 13050 4004
rect 13464 3992 13492 4032
rect 13541 4029 13553 4063
rect 13587 4029 13599 4063
rect 13541 4023 13599 4029
rect 13633 4063 13691 4069
rect 13633 4029 13645 4063
rect 13679 4060 13691 4063
rect 14660 4060 14688 4088
rect 15289 4063 15347 4069
rect 15289 4060 15301 4063
rect 13679 4032 14044 4060
rect 14660 4032 15301 4060
rect 13679 4029 13691 4032
rect 13633 4023 13691 4029
rect 13906 3992 13912 4004
rect 13464 3964 13912 3992
rect 13906 3952 13912 3964
rect 13964 3952 13970 4004
rect 10318 3924 10324 3936
rect 9272 3896 10180 3924
rect 10279 3896 10324 3924
rect 9272 3884 9278 3896
rect 10318 3884 10324 3896
rect 10376 3884 10382 3936
rect 11698 3924 11704 3936
rect 11659 3896 11704 3924
rect 11698 3884 11704 3896
rect 11756 3884 11762 3936
rect 12434 3884 12440 3936
rect 12492 3924 12498 3936
rect 12492 3896 12537 3924
rect 12492 3884 12498 3896
rect 12802 3884 12808 3936
rect 12860 3924 12866 3936
rect 14016 3924 14044 4032
rect 15289 4029 15301 4032
rect 15335 4029 15347 4063
rect 16114 4060 16120 4072
rect 16075 4032 16120 4060
rect 15289 4023 15347 4029
rect 16114 4020 16120 4032
rect 16172 4020 16178 4072
rect 16206 4020 16212 4072
rect 16264 4060 16270 4072
rect 17512 4060 17540 4091
rect 16264 4032 17540 4060
rect 16264 4020 16270 4032
rect 14645 3995 14703 4001
rect 14645 3961 14657 3995
rect 14691 3992 14703 3995
rect 16758 3992 16764 4004
rect 14691 3964 16764 3992
rect 14691 3961 14703 3964
rect 14645 3955 14703 3961
rect 16758 3952 16764 3964
rect 16816 3952 16822 4004
rect 16942 3992 16948 4004
rect 16903 3964 16948 3992
rect 16942 3952 16948 3964
rect 17000 3952 17006 4004
rect 17310 3992 17316 4004
rect 17271 3964 17316 3992
rect 17310 3952 17316 3964
rect 17368 3952 17374 4004
rect 14182 3924 14188 3936
rect 12860 3896 14188 3924
rect 12860 3884 12866 3896
rect 14182 3884 14188 3896
rect 14240 3884 14246 3936
rect 14369 3927 14427 3933
rect 14369 3893 14381 3927
rect 14415 3924 14427 3927
rect 14550 3924 14556 3936
rect 14415 3896 14556 3924
rect 14415 3893 14427 3896
rect 14369 3887 14427 3893
rect 14550 3884 14556 3896
rect 14608 3884 14614 3936
rect 14734 3924 14740 3936
rect 14695 3896 14740 3924
rect 14734 3884 14740 3896
rect 14792 3884 14798 3936
rect 14826 3884 14832 3936
rect 14884 3924 14890 3936
rect 15102 3924 15108 3936
rect 14884 3896 15108 3924
rect 14884 3884 14890 3896
rect 15102 3884 15108 3896
rect 15160 3884 15166 3936
rect 15286 3884 15292 3936
rect 15344 3924 15350 3936
rect 15930 3924 15936 3936
rect 15344 3896 15936 3924
rect 15344 3884 15350 3896
rect 15930 3884 15936 3896
rect 15988 3924 15994 3936
rect 16393 3927 16451 3933
rect 16393 3924 16405 3927
rect 15988 3896 16405 3924
rect 15988 3884 15994 3896
rect 16393 3893 16405 3896
rect 16439 3893 16451 3927
rect 16393 3887 16451 3893
rect 16850 3884 16856 3936
rect 16908 3924 16914 3936
rect 17880 3924 17908 4091
rect 18230 4088 18236 4100
rect 18288 4088 18294 4140
rect 18046 3992 18052 4004
rect 18007 3964 18052 3992
rect 18046 3952 18052 3964
rect 18104 3952 18110 4004
rect 18417 3995 18475 4001
rect 18417 3961 18429 3995
rect 18463 3992 18475 3995
rect 18598 3992 18604 4004
rect 18463 3964 18604 3992
rect 18463 3961 18475 3964
rect 18417 3955 18475 3961
rect 18598 3952 18604 3964
rect 18656 3952 18662 4004
rect 16908 3896 17908 3924
rect 16908 3884 16914 3896
rect 1104 3834 18860 3856
rect 1104 3782 3174 3834
rect 3226 3782 3238 3834
rect 3290 3782 3302 3834
rect 3354 3782 3366 3834
rect 3418 3782 3430 3834
rect 3482 3782 7622 3834
rect 7674 3782 7686 3834
rect 7738 3782 7750 3834
rect 7802 3782 7814 3834
rect 7866 3782 7878 3834
rect 7930 3782 12070 3834
rect 12122 3782 12134 3834
rect 12186 3782 12198 3834
rect 12250 3782 12262 3834
rect 12314 3782 12326 3834
rect 12378 3782 16518 3834
rect 16570 3782 16582 3834
rect 16634 3782 16646 3834
rect 16698 3782 16710 3834
rect 16762 3782 16774 3834
rect 16826 3782 18860 3834
rect 1104 3760 18860 3782
rect 1486 3720 1492 3732
rect 1447 3692 1492 3720
rect 1486 3680 1492 3692
rect 1544 3680 1550 3732
rect 2130 3720 2136 3732
rect 2091 3692 2136 3720
rect 2130 3680 2136 3692
rect 2188 3680 2194 3732
rect 2406 3680 2412 3732
rect 2464 3720 2470 3732
rect 2685 3723 2743 3729
rect 2685 3720 2697 3723
rect 2464 3692 2697 3720
rect 2464 3680 2470 3692
rect 2685 3689 2697 3692
rect 2731 3689 2743 3723
rect 2685 3683 2743 3689
rect 2866 3680 2872 3732
rect 2924 3720 2930 3732
rect 3237 3723 3295 3729
rect 3237 3720 3249 3723
rect 2924 3692 3249 3720
rect 2924 3680 2930 3692
rect 3237 3689 3249 3692
rect 3283 3689 3295 3723
rect 3510 3720 3516 3732
rect 3471 3692 3516 3720
rect 3237 3683 3295 3689
rect 3510 3680 3516 3692
rect 3568 3680 3574 3732
rect 4157 3723 4215 3729
rect 4157 3689 4169 3723
rect 4203 3720 4215 3723
rect 8110 3720 8116 3732
rect 4203 3692 8116 3720
rect 4203 3689 4215 3692
rect 4157 3683 4215 3689
rect 2314 3652 2320 3664
rect 1688 3624 2320 3652
rect 1688 3525 1716 3624
rect 2314 3612 2320 3624
rect 2372 3612 2378 3664
rect 2498 3612 2504 3664
rect 2556 3652 2562 3664
rect 2556 3624 3188 3652
rect 2556 3612 2562 3624
rect 3160 3541 3188 3624
rect 3145 3535 3203 3541
rect 1673 3519 1731 3525
rect 1673 3485 1685 3519
rect 1719 3485 1731 3519
rect 1673 3479 1731 3485
rect 1762 3476 1768 3528
rect 1820 3516 1826 3528
rect 2314 3516 2320 3528
rect 1820 3488 1865 3516
rect 2275 3488 2320 3516
rect 1820 3476 1826 3488
rect 2314 3476 2320 3488
rect 2372 3476 2378 3528
rect 2593 3519 2651 3525
rect 2593 3485 2605 3519
rect 2639 3516 2651 3519
rect 2774 3516 2780 3528
rect 2639 3488 2780 3516
rect 2639 3485 2651 3488
rect 2593 3479 2651 3485
rect 2774 3476 2780 3488
rect 2832 3476 2838 3528
rect 2869 3519 2927 3525
rect 2869 3485 2881 3519
rect 2915 3485 2927 3519
rect 3145 3501 3157 3535
rect 3191 3501 3203 3535
rect 3145 3495 3203 3501
rect 3973 3519 4031 3525
rect 2869 3479 2927 3485
rect 3973 3485 3985 3519
rect 4019 3516 4031 3519
rect 4172 3516 4200 3683
rect 8110 3680 8116 3692
rect 8168 3680 8174 3732
rect 10778 3720 10784 3732
rect 10739 3692 10784 3720
rect 10778 3680 10784 3692
rect 10836 3680 10842 3732
rect 10870 3680 10876 3732
rect 10928 3720 10934 3732
rect 12529 3723 12587 3729
rect 12529 3720 12541 3723
rect 10928 3692 12541 3720
rect 10928 3680 10934 3692
rect 12529 3689 12541 3692
rect 12575 3720 12587 3723
rect 15473 3723 15531 3729
rect 12575 3692 14964 3720
rect 12575 3689 12587 3692
rect 12529 3683 12587 3689
rect 6825 3655 6883 3661
rect 6825 3621 6837 3655
rect 6871 3652 6883 3655
rect 8938 3652 8944 3664
rect 6871 3624 8944 3652
rect 6871 3621 6883 3624
rect 6825 3615 6883 3621
rect 8938 3612 8944 3624
rect 8996 3612 9002 3664
rect 12713 3655 12771 3661
rect 12713 3621 12725 3655
rect 12759 3652 12771 3655
rect 13078 3652 13084 3664
rect 12759 3624 13084 3652
rect 12759 3621 12771 3624
rect 12713 3615 12771 3621
rect 13078 3612 13084 3624
rect 13136 3612 13142 3664
rect 13541 3655 13599 3661
rect 13541 3621 13553 3655
rect 13587 3652 13599 3655
rect 13722 3652 13728 3664
rect 13587 3624 13728 3652
rect 13587 3621 13599 3624
rect 13541 3615 13599 3621
rect 13722 3612 13728 3624
rect 13780 3612 13786 3664
rect 13906 3652 13912 3664
rect 13867 3624 13912 3652
rect 13906 3612 13912 3624
rect 13964 3612 13970 3664
rect 14182 3652 14188 3664
rect 14143 3624 14188 3652
rect 14182 3612 14188 3624
rect 14240 3612 14246 3664
rect 14645 3655 14703 3661
rect 14645 3621 14657 3655
rect 14691 3652 14703 3655
rect 14826 3652 14832 3664
rect 14691 3624 14832 3652
rect 14691 3621 14703 3624
rect 14645 3615 14703 3621
rect 14826 3612 14832 3624
rect 14884 3612 14890 3664
rect 7466 3544 7472 3596
rect 7524 3584 7530 3596
rect 12802 3584 12808 3596
rect 7524 3556 7880 3584
rect 7524 3544 7530 3556
rect 4019 3488 4200 3516
rect 4341 3519 4399 3525
rect 4019 3485 4031 3488
rect 3973 3479 4031 3485
rect 4341 3485 4353 3519
rect 4387 3516 4399 3519
rect 4706 3516 4712 3528
rect 4387 3488 4712 3516
rect 4387 3485 4399 3488
rect 4341 3479 4399 3485
rect 2884 3448 2912 3479
rect 4706 3476 4712 3488
rect 4764 3516 4770 3528
rect 4764 3488 5856 3516
rect 4764 3476 4770 3488
rect 3510 3448 3516 3460
rect 2884 3420 3516 3448
rect 3510 3408 3516 3420
rect 3568 3448 3574 3460
rect 5828 3448 5856 3488
rect 6086 3476 6092 3528
rect 6144 3516 6150 3528
rect 6641 3519 6699 3525
rect 6641 3516 6653 3519
rect 6144 3488 6653 3516
rect 6144 3476 6150 3488
rect 6641 3485 6653 3488
rect 6687 3485 6699 3519
rect 6641 3479 6699 3485
rect 7190 3476 7196 3528
rect 7248 3516 7254 3528
rect 7852 3525 7880 3556
rect 7944 3556 12808 3584
rect 7561 3519 7619 3525
rect 7561 3516 7573 3519
rect 7248 3488 7573 3516
rect 7248 3476 7254 3488
rect 7561 3485 7573 3488
rect 7607 3485 7619 3519
rect 7561 3479 7619 3485
rect 7837 3519 7895 3525
rect 7837 3485 7849 3519
rect 7883 3485 7895 3519
rect 7837 3479 7895 3485
rect 7944 3448 7972 3556
rect 12802 3544 12808 3556
rect 12860 3544 12866 3596
rect 12894 3544 12900 3596
rect 12952 3584 12958 3596
rect 12989 3587 13047 3593
rect 12989 3584 13001 3587
rect 12952 3556 13001 3584
rect 12952 3544 12958 3556
rect 12989 3553 13001 3556
rect 13035 3553 13047 3587
rect 12989 3547 13047 3553
rect 13814 3544 13820 3596
rect 13872 3584 13878 3596
rect 14936 3584 14964 3692
rect 15473 3689 15485 3723
rect 15519 3720 15531 3723
rect 16206 3720 16212 3732
rect 15519 3692 16212 3720
rect 15519 3689 15531 3692
rect 15473 3683 15531 3689
rect 16206 3680 16212 3692
rect 16264 3680 16270 3732
rect 16298 3680 16304 3732
rect 16356 3720 16362 3732
rect 16485 3723 16543 3729
rect 16485 3720 16497 3723
rect 16356 3692 16497 3720
rect 16356 3680 16362 3692
rect 16485 3689 16497 3692
rect 16531 3689 16543 3723
rect 17678 3720 17684 3732
rect 17639 3692 17684 3720
rect 16485 3683 16543 3689
rect 17678 3680 17684 3692
rect 17736 3680 17742 3732
rect 17862 3680 17868 3732
rect 17920 3720 17926 3732
rect 18049 3723 18107 3729
rect 18049 3720 18061 3723
rect 17920 3692 18061 3720
rect 17920 3680 17926 3692
rect 18049 3689 18061 3692
rect 18095 3689 18107 3723
rect 18049 3683 18107 3689
rect 18417 3723 18475 3729
rect 18417 3689 18429 3723
rect 18463 3720 18475 3723
rect 18506 3720 18512 3732
rect 18463 3692 18512 3720
rect 18463 3689 18475 3692
rect 18417 3683 18475 3689
rect 18506 3680 18512 3692
rect 18564 3680 18570 3732
rect 15749 3655 15807 3661
rect 15749 3621 15761 3655
rect 15795 3652 15807 3655
rect 17126 3652 17132 3664
rect 15795 3624 17132 3652
rect 15795 3621 15807 3624
rect 15749 3615 15807 3621
rect 17126 3612 17132 3624
rect 17184 3612 17190 3664
rect 17310 3652 17316 3664
rect 17271 3624 17316 3652
rect 17310 3612 17316 3624
rect 17368 3612 17374 3664
rect 13872 3556 14872 3584
rect 14936 3556 16252 3584
rect 13872 3544 13878 3556
rect 8018 3476 8024 3528
rect 8076 3476 8082 3528
rect 10778 3476 10784 3528
rect 10836 3516 10842 3528
rect 10965 3519 11023 3525
rect 10965 3516 10977 3519
rect 10836 3488 10977 3516
rect 10836 3476 10842 3488
rect 10965 3485 10977 3488
rect 11011 3485 11023 3519
rect 10965 3479 11023 3485
rect 13998 3476 14004 3528
rect 14056 3516 14062 3528
rect 14737 3519 14795 3525
rect 14737 3516 14749 3519
rect 14056 3488 14749 3516
rect 14056 3476 14062 3488
rect 14737 3485 14749 3488
rect 14783 3485 14795 3519
rect 14844 3516 14872 3556
rect 15013 3519 15071 3525
rect 15013 3516 15025 3519
rect 14844 3488 15025 3516
rect 14737 3479 14795 3485
rect 15013 3485 15025 3488
rect 15059 3485 15071 3519
rect 15286 3516 15292 3528
rect 15013 3479 15071 3485
rect 15120 3488 15292 3516
rect 3568 3420 5764 3448
rect 5828 3420 7972 3448
rect 8036 3448 8064 3476
rect 8036 3420 11284 3448
rect 3568 3408 3574 3420
rect 1946 3380 1952 3392
rect 1907 3352 1952 3380
rect 1946 3340 1952 3352
rect 2004 3340 2010 3392
rect 2038 3340 2044 3392
rect 2096 3380 2102 3392
rect 2409 3383 2467 3389
rect 2409 3380 2421 3383
rect 2096 3352 2421 3380
rect 2096 3340 2102 3352
rect 2409 3349 2421 3352
rect 2455 3349 2467 3383
rect 2409 3343 2467 3349
rect 2774 3340 2780 3392
rect 2832 3380 2838 3392
rect 2961 3383 3019 3389
rect 2961 3380 2973 3383
rect 2832 3352 2973 3380
rect 2832 3340 2838 3352
rect 2961 3349 2973 3352
rect 3007 3349 3019 3383
rect 3786 3380 3792 3392
rect 3747 3352 3792 3380
rect 2961 3343 3019 3349
rect 3786 3340 3792 3352
rect 3844 3340 3850 3392
rect 5736 3380 5764 3420
rect 6822 3380 6828 3392
rect 5736 3352 6828 3380
rect 6822 3340 6828 3352
rect 6880 3340 6886 3392
rect 7745 3383 7803 3389
rect 7745 3349 7757 3383
rect 7791 3380 7803 3383
rect 7926 3380 7932 3392
rect 7791 3352 7932 3380
rect 7791 3349 7803 3352
rect 7745 3343 7803 3349
rect 7926 3340 7932 3352
rect 7984 3340 7990 3392
rect 8021 3383 8079 3389
rect 8021 3349 8033 3383
rect 8067 3380 8079 3383
rect 8202 3380 8208 3392
rect 8067 3352 8208 3380
rect 8067 3349 8079 3352
rect 8021 3343 8079 3349
rect 8202 3340 8208 3352
rect 8260 3340 8266 3392
rect 11146 3380 11152 3392
rect 11107 3352 11152 3380
rect 11146 3340 11152 3352
rect 11204 3340 11210 3392
rect 11256 3380 11284 3420
rect 12526 3408 12532 3460
rect 12584 3448 12590 3460
rect 12897 3451 12955 3457
rect 12897 3448 12909 3451
rect 12584 3420 12909 3448
rect 12584 3408 12590 3420
rect 12897 3417 12909 3420
rect 12943 3448 12955 3451
rect 13630 3448 13636 3460
rect 12943 3420 13636 3448
rect 12943 3417 12955 3420
rect 12897 3411 12955 3417
rect 13630 3408 13636 3420
rect 13688 3408 13694 3460
rect 13722 3408 13728 3460
rect 13780 3448 13786 3460
rect 14461 3451 14519 3457
rect 14461 3448 14473 3451
rect 13780 3420 14473 3448
rect 13780 3408 13786 3420
rect 14461 3417 14473 3420
rect 14507 3448 14519 3451
rect 15120 3448 15148 3488
rect 15286 3476 15292 3488
rect 15344 3476 15350 3528
rect 15562 3516 15568 3528
rect 15523 3488 15568 3516
rect 15562 3476 15568 3488
rect 15620 3476 15626 3528
rect 16224 3525 16252 3556
rect 16209 3519 16267 3525
rect 16209 3485 16221 3519
rect 16255 3485 16267 3519
rect 16666 3516 16672 3528
rect 16627 3488 16672 3516
rect 16209 3479 16267 3485
rect 16666 3476 16672 3488
rect 16724 3476 16730 3528
rect 16758 3476 16764 3528
rect 16816 3516 16822 3528
rect 17129 3519 17187 3525
rect 16816 3488 16861 3516
rect 16816 3476 16822 3488
rect 17129 3485 17141 3519
rect 17175 3485 17187 3519
rect 17494 3516 17500 3528
rect 17455 3488 17500 3516
rect 17129 3479 17187 3485
rect 17144 3448 17172 3479
rect 17494 3476 17500 3488
rect 17552 3476 17558 3528
rect 17770 3476 17776 3528
rect 17828 3516 17834 3528
rect 17865 3519 17923 3525
rect 17865 3516 17877 3519
rect 17828 3488 17877 3516
rect 17828 3476 17834 3488
rect 17865 3485 17877 3488
rect 17911 3485 17923 3519
rect 18230 3516 18236 3528
rect 18191 3488 18236 3516
rect 17865 3479 17923 3485
rect 18230 3476 18236 3488
rect 18288 3476 18294 3528
rect 14507 3420 15148 3448
rect 15212 3420 17172 3448
rect 14507 3417 14519 3420
rect 14461 3411 14519 3417
rect 13357 3383 13415 3389
rect 13357 3380 13369 3383
rect 11256 3352 13369 3380
rect 13357 3349 13369 3352
rect 13403 3380 13415 3383
rect 13538 3380 13544 3392
rect 13403 3352 13544 3380
rect 13403 3349 13415 3352
rect 13357 3343 13415 3349
rect 13538 3340 13544 3352
rect 13596 3340 13602 3392
rect 14918 3380 14924 3392
rect 14879 3352 14924 3380
rect 14918 3340 14924 3352
rect 14976 3340 14982 3392
rect 15212 3389 15240 3420
rect 15197 3383 15255 3389
rect 15197 3349 15209 3383
rect 15243 3349 15255 3383
rect 16114 3380 16120 3392
rect 16075 3352 16120 3380
rect 15197 3343 15255 3349
rect 16114 3340 16120 3352
rect 16172 3340 16178 3392
rect 16390 3380 16396 3392
rect 16351 3352 16396 3380
rect 16390 3340 16396 3352
rect 16448 3340 16454 3392
rect 16942 3380 16948 3392
rect 16903 3352 16948 3380
rect 16942 3340 16948 3352
rect 17000 3340 17006 3392
rect 1104 3290 18860 3312
rect 1104 3238 5398 3290
rect 5450 3238 5462 3290
rect 5514 3238 5526 3290
rect 5578 3238 5590 3290
rect 5642 3238 5654 3290
rect 5706 3238 9846 3290
rect 9898 3238 9910 3290
rect 9962 3238 9974 3290
rect 10026 3238 10038 3290
rect 10090 3238 10102 3290
rect 10154 3238 14294 3290
rect 14346 3238 14358 3290
rect 14410 3238 14422 3290
rect 14474 3238 14486 3290
rect 14538 3238 14550 3290
rect 14602 3238 18860 3290
rect 1104 3216 18860 3238
rect 1486 3176 1492 3188
rect 1447 3148 1492 3176
rect 1486 3136 1492 3148
rect 1544 3136 1550 3188
rect 3786 3176 3792 3188
rect 1688 3148 3792 3176
rect 1688 3049 1716 3148
rect 3786 3136 3792 3148
rect 3844 3136 3850 3188
rect 3878 3136 3884 3188
rect 3936 3176 3942 3188
rect 3936 3148 3981 3176
rect 3936 3136 3942 3148
rect 6546 3136 6552 3188
rect 6604 3176 6610 3188
rect 10318 3176 10324 3188
rect 6604 3148 10324 3176
rect 6604 3136 6610 3148
rect 10318 3136 10324 3148
rect 10376 3136 10382 3188
rect 12526 3176 12532 3188
rect 11256 3148 11928 3176
rect 12487 3148 12532 3176
rect 4062 3108 4068 3120
rect 3068 3080 4068 3108
rect 1673 3043 1731 3049
rect 1673 3009 1685 3043
rect 1719 3009 1731 3043
rect 2038 3040 2044 3052
rect 1999 3012 2044 3040
rect 1673 3003 1731 3009
rect 2038 3000 2044 3012
rect 2096 3000 2102 3052
rect 2409 3043 2467 3049
rect 2409 3009 2421 3043
rect 2455 3040 2467 3043
rect 2590 3040 2596 3052
rect 2455 3012 2596 3040
rect 2455 3009 2467 3012
rect 2409 3003 2467 3009
rect 2590 3000 2596 3012
rect 2648 3000 2654 3052
rect 3068 3049 3096 3080
rect 4062 3068 4068 3080
rect 4120 3068 4126 3120
rect 6270 3068 6276 3120
rect 6328 3108 6334 3120
rect 6328 3080 7052 3108
rect 6328 3068 6334 3080
rect 2777 3043 2835 3049
rect 2777 3009 2789 3043
rect 2823 3040 2835 3043
rect 3053 3043 3111 3049
rect 2823 3012 2912 3040
rect 2823 3009 2835 3012
rect 2777 3003 2835 3009
rect 1854 2904 1860 2916
rect 1815 2876 1860 2904
rect 1854 2864 1860 2876
rect 1912 2864 1918 2916
rect 2884 2913 2912 3012
rect 3053 3009 3065 3043
rect 3099 3009 3111 3043
rect 3053 3003 3111 3009
rect 3329 3043 3387 3049
rect 3329 3009 3341 3043
rect 3375 3040 3387 3043
rect 3694 3040 3700 3052
rect 3375 3012 3700 3040
rect 3375 3009 3387 3012
rect 3329 3003 3387 3009
rect 3694 3000 3700 3012
rect 3752 3000 3758 3052
rect 5537 3043 5595 3049
rect 5537 3009 5549 3043
rect 5583 3040 5595 3043
rect 6638 3040 6644 3052
rect 5583 3012 6644 3040
rect 5583 3009 5595 3012
rect 5537 3003 5595 3009
rect 6638 3000 6644 3012
rect 6696 3000 6702 3052
rect 7024 3049 7052 3080
rect 7009 3043 7067 3049
rect 7009 3009 7021 3043
rect 7055 3009 7067 3043
rect 7009 3003 7067 3009
rect 7282 3000 7288 3052
rect 7340 3040 7346 3052
rect 7469 3043 7527 3049
rect 7469 3040 7481 3043
rect 7340 3012 7481 3040
rect 7340 3000 7346 3012
rect 7469 3009 7481 3012
rect 7515 3009 7527 3043
rect 7469 3003 7527 3009
rect 3510 2932 3516 2984
rect 3568 2972 3574 2984
rect 3605 2975 3663 2981
rect 3605 2972 3617 2975
rect 3568 2944 3617 2972
rect 3568 2932 3574 2944
rect 3605 2941 3617 2944
rect 3651 2941 3663 2975
rect 3605 2935 3663 2941
rect 5718 2932 5724 2984
rect 5776 2972 5782 2984
rect 11256 2972 11284 3148
rect 11422 3068 11428 3120
rect 11480 3108 11486 3120
rect 11900 3108 11928 3148
rect 12526 3136 12532 3148
rect 12584 3136 12590 3188
rect 12897 3179 12955 3185
rect 12897 3145 12909 3179
rect 12943 3176 12955 3179
rect 12986 3176 12992 3188
rect 12943 3148 12992 3176
rect 12943 3145 12955 3148
rect 12897 3139 12955 3145
rect 12986 3136 12992 3148
rect 13044 3136 13050 3188
rect 13170 3176 13176 3188
rect 13131 3148 13176 3176
rect 13170 3136 13176 3148
rect 13228 3176 13234 3188
rect 15194 3176 15200 3188
rect 13228 3148 15200 3176
rect 13228 3136 13234 3148
rect 15194 3136 15200 3148
rect 15252 3136 15258 3188
rect 16206 3176 16212 3188
rect 16167 3148 16212 3176
rect 16206 3136 16212 3148
rect 16264 3136 16270 3188
rect 16485 3179 16543 3185
rect 16485 3145 16497 3179
rect 16531 3176 16543 3179
rect 16850 3176 16856 3188
rect 16531 3148 16856 3176
rect 16531 3145 16543 3148
rect 16485 3139 16543 3145
rect 16850 3136 16856 3148
rect 16908 3136 16914 3188
rect 17034 3176 17040 3188
rect 16995 3148 17040 3176
rect 17034 3136 17040 3148
rect 17092 3136 17098 3188
rect 18046 3176 18052 3188
rect 18007 3148 18052 3176
rect 18046 3136 18052 3148
rect 18104 3136 18110 3188
rect 18414 3176 18420 3188
rect 18375 3148 18420 3176
rect 18414 3136 18420 3148
rect 18472 3136 18478 3188
rect 12713 3111 12771 3117
rect 12713 3108 12725 3111
rect 11480 3080 11836 3108
rect 11900 3080 12725 3108
rect 11480 3068 11486 3080
rect 11333 3043 11391 3049
rect 11333 3009 11345 3043
rect 11379 3040 11391 3043
rect 11606 3040 11612 3052
rect 11379 3012 11612 3040
rect 11379 3009 11391 3012
rect 11333 3003 11391 3009
rect 11606 3000 11612 3012
rect 11664 3000 11670 3052
rect 11808 3049 11836 3080
rect 12713 3077 12725 3080
rect 12759 3108 12771 3111
rect 17218 3108 17224 3120
rect 12759 3080 16344 3108
rect 12759 3077 12771 3080
rect 12713 3071 12771 3077
rect 11701 3043 11759 3049
rect 11701 3009 11713 3043
rect 11747 3009 11759 3043
rect 11701 3003 11759 3009
rect 11793 3043 11851 3049
rect 11793 3009 11805 3043
rect 11839 3009 11851 3043
rect 11793 3003 11851 3009
rect 5776 2944 11284 2972
rect 11716 2972 11744 3003
rect 12618 3000 12624 3052
rect 12676 3040 12682 3052
rect 13541 3043 13599 3049
rect 13541 3040 13553 3043
rect 12676 3012 13553 3040
rect 12676 3000 12682 3012
rect 13541 3009 13553 3012
rect 13587 3009 13599 3043
rect 13814 3040 13820 3052
rect 13775 3012 13820 3040
rect 13541 3003 13599 3009
rect 13814 3000 13820 3012
rect 13872 3000 13878 3052
rect 13998 3040 14004 3052
rect 13959 3012 14004 3040
rect 13998 3000 14004 3012
rect 14056 3000 14062 3052
rect 14090 3000 14096 3052
rect 14148 3040 14154 3052
rect 14461 3043 14519 3049
rect 14148 3012 14193 3040
rect 14148 3000 14154 3012
rect 14461 3009 14473 3043
rect 14507 3040 14519 3043
rect 15010 3040 15016 3052
rect 14507 3012 14872 3040
rect 14971 3012 15016 3040
rect 14507 3009 14519 3012
rect 14461 3003 14519 3009
rect 14734 2972 14740 2984
rect 11716 2944 14740 2972
rect 5776 2932 5782 2944
rect 14734 2932 14740 2944
rect 14792 2932 14798 2984
rect 14844 2972 14872 3012
rect 15010 3000 15016 3012
rect 15068 3000 15074 3052
rect 15194 3000 15200 3052
rect 15252 3040 15258 3052
rect 15470 3040 15476 3052
rect 15252 3012 15297 3040
rect 15431 3012 15476 3040
rect 15252 3000 15258 3012
rect 15470 3000 15476 3012
rect 15528 3000 15534 3052
rect 15746 3040 15752 3052
rect 15707 3012 15752 3040
rect 15746 3000 15752 3012
rect 15804 3000 15810 3052
rect 16022 3040 16028 3052
rect 15983 3012 16028 3040
rect 16022 3000 16028 3012
rect 16080 3000 16086 3052
rect 16316 3049 16344 3080
rect 16868 3080 17224 3108
rect 16301 3043 16359 3049
rect 16301 3009 16313 3043
rect 16347 3009 16359 3043
rect 16301 3003 16359 3009
rect 16390 3000 16396 3052
rect 16448 3040 16454 3052
rect 16868 3049 16896 3080
rect 17218 3068 17224 3080
rect 17276 3068 17282 3120
rect 16853 3043 16911 3049
rect 16853 3040 16865 3043
rect 16448 3012 16865 3040
rect 16448 3000 16454 3012
rect 16853 3009 16865 3012
rect 16899 3009 16911 3043
rect 17126 3040 17132 3052
rect 17087 3012 17132 3040
rect 16853 3003 16911 3009
rect 17126 3000 17132 3012
rect 17184 3000 17190 3052
rect 17497 3043 17555 3049
rect 17497 3009 17509 3043
rect 17543 3009 17555 3043
rect 17497 3003 17555 3009
rect 15654 2972 15660 2984
rect 14844 2944 15660 2972
rect 15654 2932 15660 2944
rect 15712 2932 15718 2984
rect 17512 2972 17540 3003
rect 17586 3000 17592 3052
rect 17644 3040 17650 3052
rect 17865 3043 17923 3049
rect 17865 3040 17877 3043
rect 17644 3012 17877 3040
rect 17644 3000 17650 3012
rect 17865 3009 17877 3012
rect 17911 3009 17923 3043
rect 17865 3003 17923 3009
rect 17954 3000 17960 3052
rect 18012 3040 18018 3052
rect 18233 3043 18291 3049
rect 18233 3040 18245 3043
rect 18012 3012 18245 3040
rect 18012 3000 18018 3012
rect 18233 3009 18245 3012
rect 18279 3009 18291 3043
rect 18233 3003 18291 3009
rect 15948 2944 17540 2972
rect 2869 2907 2927 2913
rect 2869 2873 2881 2907
rect 2915 2873 2927 2907
rect 2869 2867 2927 2873
rect 7098 2864 7104 2916
rect 7156 2904 7162 2916
rect 7285 2907 7343 2913
rect 7285 2904 7297 2907
rect 7156 2876 7297 2904
rect 7156 2864 7162 2876
rect 7285 2873 7297 2876
rect 7331 2873 7343 2907
rect 7285 2867 7343 2873
rect 8754 2864 8760 2916
rect 8812 2904 8818 2916
rect 13078 2904 13084 2916
rect 8812 2876 12434 2904
rect 13039 2876 13084 2904
rect 8812 2864 8818 2876
rect 2222 2836 2228 2848
rect 2183 2808 2228 2836
rect 2222 2796 2228 2808
rect 2280 2796 2286 2848
rect 2590 2836 2596 2848
rect 2551 2808 2596 2836
rect 2590 2796 2596 2808
rect 2648 2796 2654 2848
rect 2682 2796 2688 2848
rect 2740 2836 2746 2848
rect 3145 2839 3203 2845
rect 3145 2836 3157 2839
rect 2740 2808 3157 2836
rect 2740 2796 2746 2808
rect 3145 2805 3157 2808
rect 3191 2805 3203 2839
rect 3510 2836 3516 2848
rect 3471 2808 3516 2836
rect 3145 2799 3203 2805
rect 3510 2796 3516 2808
rect 3568 2796 3574 2848
rect 4890 2796 4896 2848
rect 4948 2836 4954 2848
rect 5353 2839 5411 2845
rect 5353 2836 5365 2839
rect 4948 2808 5365 2836
rect 4948 2796 4954 2808
rect 5353 2805 5365 2808
rect 5399 2805 5411 2839
rect 7190 2836 7196 2848
rect 7151 2808 7196 2836
rect 5353 2799 5411 2805
rect 7190 2796 7196 2808
rect 7248 2796 7254 2848
rect 11146 2836 11152 2848
rect 11107 2808 11152 2836
rect 11146 2796 11152 2808
rect 11204 2796 11210 2848
rect 11514 2836 11520 2848
rect 11475 2808 11520 2836
rect 11514 2796 11520 2808
rect 11572 2796 11578 2848
rect 11974 2836 11980 2848
rect 11935 2808 11980 2836
rect 11974 2796 11980 2808
rect 12032 2796 12038 2848
rect 12406 2836 12434 2876
rect 13078 2864 13084 2876
rect 13136 2864 13142 2916
rect 13449 2907 13507 2913
rect 13449 2873 13461 2907
rect 13495 2904 13507 2907
rect 13722 2904 13728 2916
rect 13495 2876 13728 2904
rect 13495 2873 13507 2876
rect 13449 2867 13507 2873
rect 13464 2836 13492 2867
rect 13722 2864 13728 2876
rect 13780 2864 13786 2916
rect 14645 2907 14703 2913
rect 14645 2873 14657 2907
rect 14691 2904 14703 2907
rect 15102 2904 15108 2916
rect 14691 2876 15108 2904
rect 14691 2873 14703 2876
rect 14645 2867 14703 2873
rect 15102 2864 15108 2876
rect 15160 2864 15166 2916
rect 15381 2907 15439 2913
rect 15381 2873 15393 2907
rect 15427 2904 15439 2907
rect 15562 2904 15568 2916
rect 15427 2876 15568 2904
rect 15427 2873 15439 2876
rect 15381 2867 15439 2873
rect 15562 2864 15568 2876
rect 15620 2864 15626 2916
rect 15948 2913 15976 2944
rect 15933 2907 15991 2913
rect 15933 2873 15945 2907
rect 15979 2873 15991 2907
rect 15933 2867 15991 2873
rect 16574 2864 16580 2916
rect 16632 2904 16638 2916
rect 16669 2907 16727 2913
rect 16669 2904 16681 2907
rect 16632 2876 16681 2904
rect 16632 2864 16638 2876
rect 16669 2873 16681 2876
rect 16715 2873 16727 2907
rect 16669 2867 16727 2873
rect 12406 2808 13492 2836
rect 14277 2839 14335 2845
rect 14277 2805 14289 2839
rect 14323 2836 14335 2839
rect 14366 2836 14372 2848
rect 14323 2808 14372 2836
rect 14323 2805 14335 2808
rect 14277 2799 14335 2805
rect 14366 2796 14372 2808
rect 14424 2796 14430 2848
rect 14829 2839 14887 2845
rect 14829 2805 14841 2839
rect 14875 2836 14887 2839
rect 15010 2836 15016 2848
rect 14875 2808 15016 2836
rect 14875 2805 14887 2808
rect 14829 2799 14887 2805
rect 15010 2796 15016 2808
rect 15068 2796 15074 2848
rect 15654 2836 15660 2848
rect 15615 2808 15660 2836
rect 15654 2796 15660 2808
rect 15712 2796 15718 2848
rect 17310 2836 17316 2848
rect 17271 2808 17316 2836
rect 17310 2796 17316 2808
rect 17368 2796 17374 2848
rect 17678 2836 17684 2848
rect 17639 2808 17684 2836
rect 17678 2796 17684 2808
rect 17736 2796 17742 2848
rect 1104 2746 18860 2768
rect 1104 2694 3174 2746
rect 3226 2694 3238 2746
rect 3290 2694 3302 2746
rect 3354 2694 3366 2746
rect 3418 2694 3430 2746
rect 3482 2694 7622 2746
rect 7674 2694 7686 2746
rect 7738 2694 7750 2746
rect 7802 2694 7814 2746
rect 7866 2694 7878 2746
rect 7930 2694 12070 2746
rect 12122 2694 12134 2746
rect 12186 2694 12198 2746
rect 12250 2694 12262 2746
rect 12314 2694 12326 2746
rect 12378 2694 16518 2746
rect 16570 2694 16582 2746
rect 16634 2694 16646 2746
rect 16698 2694 16710 2746
rect 16762 2694 16774 2746
rect 16826 2694 18860 2746
rect 1104 2672 18860 2694
rect 1486 2632 1492 2644
rect 1447 2604 1492 2632
rect 1486 2592 1492 2604
rect 1544 2592 1550 2644
rect 2958 2632 2964 2644
rect 2056 2604 2964 2632
rect 2056 2437 2084 2604
rect 2958 2592 2964 2604
rect 3016 2592 3022 2644
rect 11882 2592 11888 2644
rect 11940 2632 11946 2644
rect 11940 2604 14320 2632
rect 11940 2592 11946 2604
rect 11238 2564 11244 2576
rect 2424 2536 11244 2564
rect 2424 2437 2452 2536
rect 11238 2524 11244 2536
rect 11296 2524 11302 2576
rect 13630 2524 13636 2576
rect 13688 2564 13694 2576
rect 14185 2567 14243 2573
rect 14185 2564 14197 2567
rect 13688 2536 14197 2564
rect 13688 2524 13694 2536
rect 14185 2533 14197 2536
rect 14231 2533 14243 2567
rect 14292 2564 14320 2604
rect 14458 2592 14464 2644
rect 14516 2632 14522 2644
rect 15013 2635 15071 2641
rect 15013 2632 15025 2635
rect 14516 2604 15025 2632
rect 14516 2592 14522 2604
rect 15013 2601 15025 2604
rect 15059 2632 15071 2635
rect 15194 2632 15200 2644
rect 15059 2604 15200 2632
rect 15059 2601 15071 2604
rect 15013 2595 15071 2601
rect 15194 2592 15200 2604
rect 15252 2592 15258 2644
rect 15289 2635 15347 2641
rect 15289 2601 15301 2635
rect 15335 2632 15347 2635
rect 15746 2632 15752 2644
rect 15335 2604 15752 2632
rect 15335 2601 15347 2604
rect 15289 2595 15347 2601
rect 15746 2592 15752 2604
rect 15804 2592 15810 2644
rect 18414 2632 18420 2644
rect 15856 2604 17724 2632
rect 18375 2604 18420 2632
rect 14292 2536 15516 2564
rect 14185 2527 14243 2533
rect 3050 2496 3056 2508
rect 2516 2468 3056 2496
rect 1673 2431 1731 2437
rect 1673 2397 1685 2431
rect 1719 2397 1731 2431
rect 1673 2391 1731 2397
rect 2041 2431 2099 2437
rect 2041 2397 2053 2431
rect 2087 2397 2099 2431
rect 2041 2391 2099 2397
rect 2409 2431 2467 2437
rect 2409 2397 2421 2431
rect 2455 2397 2467 2431
rect 2409 2391 2467 2397
rect 1688 2360 1716 2391
rect 2516 2360 2544 2468
rect 3050 2456 3056 2468
rect 3108 2456 3114 2508
rect 3602 2496 3608 2508
rect 3252 2468 3608 2496
rect 2774 2428 2780 2440
rect 2735 2400 2780 2428
rect 2774 2388 2780 2400
rect 2832 2388 2838 2440
rect 3252 2437 3280 2468
rect 3602 2456 3608 2468
rect 3660 2456 3666 2508
rect 8202 2456 8208 2508
rect 8260 2496 8266 2508
rect 8260 2468 9628 2496
rect 8260 2456 8266 2468
rect 3237 2431 3295 2437
rect 3237 2397 3249 2431
rect 3283 2397 3295 2431
rect 3237 2391 3295 2397
rect 3329 2431 3387 2437
rect 3329 2397 3341 2431
rect 3375 2397 3387 2431
rect 3329 2391 3387 2397
rect 1688 2332 2544 2360
rect 2682 2320 2688 2372
rect 2740 2360 2746 2372
rect 3344 2360 3372 2391
rect 3510 2388 3516 2440
rect 3568 2428 3574 2440
rect 3789 2431 3847 2437
rect 3789 2428 3801 2431
rect 3568 2400 3801 2428
rect 3568 2388 3574 2400
rect 3789 2397 3801 2400
rect 3835 2397 3847 2431
rect 4890 2428 4896 2440
rect 4851 2400 4896 2428
rect 3789 2391 3847 2397
rect 4890 2388 4896 2400
rect 4948 2388 4954 2440
rect 5166 2388 5172 2440
rect 5224 2428 5230 2440
rect 5445 2431 5503 2437
rect 5445 2428 5457 2431
rect 5224 2400 5457 2428
rect 5224 2388 5230 2400
rect 5445 2397 5457 2400
rect 5491 2397 5503 2431
rect 5445 2391 5503 2397
rect 6641 2431 6699 2437
rect 6641 2397 6653 2431
rect 6687 2428 6699 2431
rect 7098 2428 7104 2440
rect 6687 2400 7104 2428
rect 6687 2397 6699 2400
rect 6641 2391 6699 2397
rect 7098 2388 7104 2400
rect 7156 2388 7162 2440
rect 7190 2388 7196 2440
rect 7248 2428 7254 2440
rect 7377 2431 7435 2437
rect 7377 2428 7389 2431
rect 7248 2400 7389 2428
rect 7248 2388 7254 2400
rect 7377 2397 7389 2400
rect 7423 2397 7435 2431
rect 7377 2391 7435 2397
rect 7929 2431 7987 2437
rect 7929 2397 7941 2431
rect 7975 2428 7987 2431
rect 8018 2428 8024 2440
rect 7975 2400 8024 2428
rect 7975 2397 7987 2400
rect 7929 2391 7987 2397
rect 8018 2388 8024 2400
rect 8076 2388 8082 2440
rect 8938 2428 8944 2440
rect 8899 2400 8944 2428
rect 8938 2388 8944 2400
rect 8996 2388 9002 2440
rect 9600 2437 9628 2468
rect 11974 2456 11980 2508
rect 12032 2496 12038 2508
rect 15488 2496 15516 2536
rect 15562 2524 15568 2576
rect 15620 2564 15626 2576
rect 15856 2564 15884 2604
rect 15620 2536 15884 2564
rect 15933 2567 15991 2573
rect 15620 2524 15626 2536
rect 15933 2533 15945 2567
rect 15979 2533 15991 2567
rect 15933 2527 15991 2533
rect 16485 2567 16543 2573
rect 16485 2533 16497 2567
rect 16531 2564 16543 2567
rect 17586 2564 17592 2576
rect 16531 2536 17592 2564
rect 16531 2533 16543 2536
rect 16485 2527 16543 2533
rect 12032 2468 15424 2496
rect 15488 2468 15884 2496
rect 12032 2456 12038 2468
rect 9585 2431 9643 2437
rect 9585 2397 9597 2431
rect 9631 2397 9643 2431
rect 9585 2391 9643 2397
rect 10689 2431 10747 2437
rect 10689 2397 10701 2431
rect 10735 2428 10747 2431
rect 11146 2428 11152 2440
rect 10735 2400 11152 2428
rect 10735 2397 10747 2400
rect 10689 2391 10747 2397
rect 11146 2388 11152 2400
rect 11204 2388 11210 2440
rect 11514 2428 11520 2440
rect 11475 2400 11520 2428
rect 11514 2388 11520 2400
rect 11572 2388 11578 2440
rect 11698 2388 11704 2440
rect 11756 2428 11762 2440
rect 12069 2431 12127 2437
rect 12069 2428 12081 2431
rect 11756 2400 12081 2428
rect 11756 2388 11762 2400
rect 12069 2397 12081 2400
rect 12115 2397 12127 2431
rect 12069 2391 12127 2397
rect 12434 2388 12440 2440
rect 12492 2428 12498 2440
rect 12897 2431 12955 2437
rect 12897 2428 12909 2431
rect 12492 2400 12909 2428
rect 12492 2388 12498 2400
rect 12897 2397 12909 2400
rect 12943 2397 12955 2431
rect 12897 2391 12955 2397
rect 13357 2431 13415 2437
rect 13357 2397 13369 2431
rect 13403 2428 13415 2431
rect 13722 2428 13728 2440
rect 13403 2400 13728 2428
rect 13403 2397 13415 2400
rect 13357 2391 13415 2397
rect 13722 2388 13728 2400
rect 13780 2388 13786 2440
rect 14366 2428 14372 2440
rect 14327 2400 14372 2428
rect 14366 2388 14372 2400
rect 14424 2388 14430 2440
rect 14829 2431 14887 2437
rect 14829 2397 14841 2431
rect 14875 2428 14887 2431
rect 15010 2428 15016 2440
rect 14875 2400 15016 2428
rect 14875 2397 14887 2400
rect 14829 2391 14887 2397
rect 15010 2388 15016 2400
rect 15068 2388 15074 2440
rect 15396 2437 15424 2468
rect 15381 2431 15439 2437
rect 15381 2397 15393 2431
rect 15427 2397 15439 2431
rect 15381 2391 15439 2397
rect 15749 2431 15807 2437
rect 15749 2397 15761 2431
rect 15795 2397 15807 2431
rect 15749 2391 15807 2397
rect 4157 2363 4215 2369
rect 4157 2360 4169 2363
rect 2740 2332 4169 2360
rect 2740 2320 2746 2332
rect 4157 2329 4169 2332
rect 4203 2329 4215 2363
rect 4157 2323 4215 2329
rect 12621 2363 12679 2369
rect 12621 2329 12633 2363
rect 12667 2360 12679 2363
rect 13740 2360 13768 2388
rect 15470 2360 15476 2372
rect 12667 2332 13676 2360
rect 13740 2332 15476 2360
rect 12667 2329 12679 2332
rect 12621 2323 12679 2329
rect 1854 2292 1860 2304
rect 1815 2264 1860 2292
rect 1854 2252 1860 2264
rect 1912 2252 1918 2304
rect 2038 2252 2044 2304
rect 2096 2292 2102 2304
rect 2225 2295 2283 2301
rect 2225 2292 2237 2295
rect 2096 2264 2237 2292
rect 2096 2252 2102 2264
rect 2225 2261 2237 2264
rect 2271 2261 2283 2295
rect 2225 2255 2283 2261
rect 2593 2295 2651 2301
rect 2593 2261 2605 2295
rect 2639 2292 2651 2295
rect 2774 2292 2780 2304
rect 2639 2264 2780 2292
rect 2639 2261 2651 2264
rect 2593 2255 2651 2261
rect 2774 2252 2780 2264
rect 2832 2252 2838 2304
rect 2866 2252 2872 2304
rect 2924 2292 2930 2304
rect 3053 2295 3111 2301
rect 3053 2292 3065 2295
rect 2924 2264 3065 2292
rect 2924 2252 2930 2264
rect 3053 2261 3065 2264
rect 3099 2261 3111 2295
rect 3053 2255 3111 2261
rect 3513 2295 3571 2301
rect 3513 2261 3525 2295
rect 3559 2292 3571 2295
rect 3602 2292 3608 2304
rect 3559 2264 3608 2292
rect 3559 2261 3571 2264
rect 3513 2255 3571 2261
rect 3602 2252 3608 2264
rect 3660 2252 3666 2304
rect 3694 2252 3700 2304
rect 3752 2292 3758 2304
rect 3973 2295 4031 2301
rect 3973 2292 3985 2295
rect 3752 2264 3985 2292
rect 3752 2252 3758 2264
rect 3973 2261 3985 2264
rect 4019 2261 4031 2295
rect 3973 2255 4031 2261
rect 4522 2252 4528 2304
rect 4580 2292 4586 2304
rect 4709 2295 4767 2301
rect 4709 2292 4721 2295
rect 4580 2264 4721 2292
rect 4580 2252 4586 2264
rect 4709 2261 4721 2264
rect 4755 2261 4767 2295
rect 4709 2255 4767 2261
rect 5258 2252 5264 2304
rect 5316 2292 5322 2304
rect 5629 2295 5687 2301
rect 5629 2292 5641 2295
rect 5316 2264 5641 2292
rect 5316 2252 5322 2264
rect 5629 2261 5641 2264
rect 5675 2261 5687 2295
rect 5629 2255 5687 2261
rect 6178 2252 6184 2304
rect 6236 2292 6242 2304
rect 6457 2295 6515 2301
rect 6457 2292 6469 2295
rect 6236 2264 6469 2292
rect 6236 2252 6242 2264
rect 6457 2261 6469 2264
rect 6503 2261 6515 2295
rect 6457 2255 6515 2261
rect 7006 2252 7012 2304
rect 7064 2292 7070 2304
rect 7193 2295 7251 2301
rect 7193 2292 7205 2295
rect 7064 2264 7205 2292
rect 7064 2252 7070 2264
rect 7193 2261 7205 2264
rect 7239 2261 7251 2295
rect 7193 2255 7251 2261
rect 7834 2252 7840 2304
rect 7892 2292 7898 2304
rect 8113 2295 8171 2301
rect 8113 2292 8125 2295
rect 7892 2264 8125 2292
rect 7892 2252 7898 2264
rect 8113 2261 8125 2264
rect 8159 2261 8171 2295
rect 8113 2255 8171 2261
rect 8662 2252 8668 2304
rect 8720 2292 8726 2304
rect 9125 2295 9183 2301
rect 9125 2292 9137 2295
rect 8720 2264 9137 2292
rect 8720 2252 8726 2264
rect 9125 2261 9137 2264
rect 9171 2261 9183 2295
rect 9125 2255 9183 2261
rect 9490 2252 9496 2304
rect 9548 2292 9554 2304
rect 9769 2295 9827 2301
rect 9769 2292 9781 2295
rect 9548 2264 9781 2292
rect 9548 2252 9554 2264
rect 9769 2261 9781 2264
rect 9815 2261 9827 2295
rect 9769 2255 9827 2261
rect 10318 2252 10324 2304
rect 10376 2292 10382 2304
rect 10505 2295 10563 2301
rect 10505 2292 10517 2295
rect 10376 2264 10517 2292
rect 10376 2252 10382 2264
rect 10505 2261 10517 2264
rect 10551 2261 10563 2295
rect 10505 2255 10563 2261
rect 11146 2252 11152 2304
rect 11204 2292 11210 2304
rect 11701 2295 11759 2301
rect 11701 2292 11713 2295
rect 11204 2264 11713 2292
rect 11204 2252 11210 2264
rect 11701 2261 11713 2264
rect 11747 2261 11759 2295
rect 11701 2255 11759 2261
rect 11974 2252 11980 2304
rect 12032 2292 12038 2304
rect 12253 2295 12311 2301
rect 12253 2292 12265 2295
rect 12032 2264 12265 2292
rect 12032 2252 12038 2264
rect 12253 2261 12265 2264
rect 12299 2261 12311 2295
rect 12710 2292 12716 2304
rect 12671 2264 12716 2292
rect 12253 2255 12311 2261
rect 12710 2252 12716 2264
rect 12768 2252 12774 2304
rect 12802 2252 12808 2304
rect 12860 2292 12866 2304
rect 13081 2295 13139 2301
rect 13081 2292 13093 2295
rect 12860 2264 13093 2292
rect 12860 2252 12866 2264
rect 13081 2261 13093 2264
rect 13127 2261 13139 2295
rect 13538 2292 13544 2304
rect 13499 2264 13544 2292
rect 13081 2255 13139 2261
rect 13538 2252 13544 2264
rect 13596 2252 13602 2304
rect 13648 2292 13676 2332
rect 15470 2320 15476 2332
rect 15528 2360 15534 2372
rect 15764 2360 15792 2391
rect 15528 2332 15792 2360
rect 15528 2320 15534 2332
rect 13722 2292 13728 2304
rect 13648 2264 13728 2292
rect 13722 2252 13728 2264
rect 13780 2252 13786 2304
rect 13909 2295 13967 2301
rect 13909 2261 13921 2295
rect 13955 2292 13967 2295
rect 13998 2292 14004 2304
rect 13955 2264 14004 2292
rect 13955 2261 13967 2264
rect 13909 2255 13967 2261
rect 13998 2252 14004 2264
rect 14056 2292 14062 2304
rect 14458 2292 14464 2304
rect 14056 2264 14464 2292
rect 14056 2252 14062 2264
rect 14458 2252 14464 2264
rect 14516 2252 14522 2304
rect 14642 2292 14648 2304
rect 14603 2264 14648 2292
rect 14642 2252 14648 2264
rect 14700 2252 14706 2304
rect 15286 2252 15292 2304
rect 15344 2292 15350 2304
rect 15565 2295 15623 2301
rect 15565 2292 15577 2295
rect 15344 2264 15577 2292
rect 15344 2252 15350 2264
rect 15565 2261 15577 2264
rect 15611 2261 15623 2295
rect 15856 2292 15884 2468
rect 15948 2428 15976 2527
rect 17586 2524 17592 2536
rect 17644 2524 17650 2576
rect 16114 2456 16120 2508
rect 16172 2496 16178 2508
rect 17402 2496 17408 2508
rect 16172 2468 16252 2496
rect 16172 2456 16178 2468
rect 16224 2437 16252 2468
rect 16316 2468 17408 2496
rect 16316 2437 16344 2468
rect 17402 2456 17408 2468
rect 17460 2456 17466 2508
rect 17696 2496 17724 2604
rect 18414 2592 18420 2604
rect 18472 2592 18478 2644
rect 17696 2468 17908 2496
rect 16209 2431 16267 2437
rect 15948 2404 16068 2428
rect 15948 2400 16160 2404
rect 16040 2376 16160 2400
rect 16209 2397 16221 2431
rect 16255 2397 16267 2431
rect 16209 2391 16267 2397
rect 16301 2431 16359 2437
rect 16301 2397 16313 2431
rect 16347 2397 16359 2431
rect 16301 2391 16359 2397
rect 16390 2388 16396 2440
rect 16448 2428 16454 2440
rect 16761 2431 16819 2437
rect 16761 2428 16773 2431
rect 16448 2400 16773 2428
rect 16448 2388 16454 2400
rect 16761 2397 16773 2400
rect 16807 2397 16819 2431
rect 16761 2391 16819 2397
rect 17034 2388 17040 2440
rect 17092 2428 17098 2440
rect 17880 2437 17908 2468
rect 17497 2431 17555 2437
rect 17092 2400 17137 2428
rect 17092 2388 17098 2400
rect 17497 2397 17509 2431
rect 17543 2397 17555 2431
rect 17497 2391 17555 2397
rect 17865 2431 17923 2437
rect 17865 2397 17877 2431
rect 17911 2397 17923 2431
rect 18230 2428 18236 2440
rect 18191 2400 18236 2428
rect 17865 2391 17923 2397
rect 16132 2360 16160 2376
rect 17512 2360 17540 2391
rect 18230 2388 18236 2400
rect 18288 2388 18294 2440
rect 18598 2360 18604 2372
rect 16132 2332 17540 2360
rect 17696 2332 18604 2360
rect 16025 2295 16083 2301
rect 16025 2292 16037 2295
rect 15856 2264 16037 2292
rect 15565 2255 15623 2261
rect 16025 2261 16037 2264
rect 16071 2261 16083 2295
rect 16025 2255 16083 2261
rect 16850 2252 16856 2304
rect 16908 2292 16914 2304
rect 16945 2295 17003 2301
rect 16945 2292 16957 2295
rect 16908 2264 16957 2292
rect 16908 2252 16914 2264
rect 16945 2261 16957 2264
rect 16991 2261 17003 2295
rect 16945 2255 17003 2261
rect 17034 2252 17040 2304
rect 17092 2292 17098 2304
rect 17696 2301 17724 2332
rect 18598 2320 18604 2332
rect 18656 2320 18662 2372
rect 17221 2295 17279 2301
rect 17221 2292 17233 2295
rect 17092 2264 17233 2292
rect 17092 2252 17098 2264
rect 17221 2261 17233 2264
rect 17267 2261 17279 2295
rect 17221 2255 17279 2261
rect 17681 2295 17739 2301
rect 17681 2261 17693 2295
rect 17727 2261 17739 2295
rect 17681 2255 17739 2261
rect 17770 2252 17776 2304
rect 17828 2292 17834 2304
rect 18049 2295 18107 2301
rect 18049 2292 18061 2295
rect 17828 2264 18061 2292
rect 17828 2252 17834 2264
rect 18049 2261 18061 2264
rect 18095 2261 18107 2295
rect 18049 2255 18107 2261
rect 1104 2202 18860 2224
rect 1104 2150 5398 2202
rect 5450 2150 5462 2202
rect 5514 2150 5526 2202
rect 5578 2150 5590 2202
rect 5642 2150 5654 2202
rect 5706 2150 9846 2202
rect 9898 2150 9910 2202
rect 9962 2150 9974 2202
rect 10026 2150 10038 2202
rect 10090 2150 10102 2202
rect 10154 2150 14294 2202
rect 14346 2150 14358 2202
rect 14410 2150 14422 2202
rect 14474 2150 14486 2202
rect 14538 2150 14550 2202
rect 14602 2150 18860 2202
rect 1104 2128 18860 2150
rect 1210 2048 1216 2100
rect 1268 2088 1274 2100
rect 2682 2088 2688 2100
rect 1268 2060 2688 2088
rect 1268 2048 1274 2060
rect 2682 2048 2688 2060
rect 2740 2048 2746 2100
rect 15654 2048 15660 2100
rect 15712 2088 15718 2100
rect 18230 2088 18236 2100
rect 15712 2060 18236 2088
rect 15712 2048 15718 2060
rect 18230 2048 18236 2060
rect 18288 2048 18294 2100
rect 12710 1912 12716 1964
rect 12768 1952 12774 1964
rect 16114 1952 16120 1964
rect 12768 1924 16120 1952
rect 12768 1912 12774 1924
rect 16114 1912 16120 1924
rect 16172 1912 16178 1964
rect 16850 1912 16856 1964
rect 16908 1952 16914 1964
rect 17494 1952 17500 1964
rect 16908 1924 17500 1952
rect 16908 1912 16914 1924
rect 17494 1912 17500 1924
rect 17552 1912 17558 1964
rect 13538 1844 13544 1896
rect 13596 1884 13602 1896
rect 16022 1884 16028 1896
rect 13596 1856 16028 1884
rect 13596 1844 13602 1856
rect 16022 1844 16028 1856
rect 16080 1844 16086 1896
<< via1 >>
rect 2136 15172 2188 15224
rect 4528 15172 4580 15224
rect 11796 14900 11848 14952
rect 18328 14900 18380 14952
rect 6276 14832 6328 14884
rect 11520 14832 11572 14884
rect 12624 14832 12676 14884
rect 1860 14764 1912 14816
rect 5816 14764 5868 14816
rect 8576 14764 8628 14816
rect 13268 14764 13320 14816
rect 3174 14662 3226 14714
rect 3238 14662 3290 14714
rect 3302 14662 3354 14714
rect 3366 14662 3418 14714
rect 3430 14662 3482 14714
rect 7622 14662 7674 14714
rect 7686 14662 7738 14714
rect 7750 14662 7802 14714
rect 7814 14662 7866 14714
rect 7878 14662 7930 14714
rect 12070 14662 12122 14714
rect 12134 14662 12186 14714
rect 12198 14662 12250 14714
rect 12262 14662 12314 14714
rect 12326 14662 12378 14714
rect 16518 14662 16570 14714
rect 16582 14662 16634 14714
rect 16646 14662 16698 14714
rect 16710 14662 16762 14714
rect 16774 14662 16826 14714
rect 2044 14560 2096 14612
rect 2228 14467 2280 14476
rect 2228 14433 2237 14467
rect 2237 14433 2271 14467
rect 2271 14433 2280 14467
rect 2228 14424 2280 14433
rect 1952 14399 2004 14408
rect 1952 14365 1961 14399
rect 1961 14365 1995 14399
rect 1995 14365 2004 14399
rect 1952 14356 2004 14365
rect 3056 14492 3108 14544
rect 4804 14492 4856 14544
rect 6000 14560 6052 14612
rect 9956 14560 10008 14612
rect 4068 14424 4120 14476
rect 3056 14356 3108 14408
rect 4160 14356 4212 14408
rect 4344 14399 4396 14408
rect 4344 14365 4353 14399
rect 4353 14365 4387 14399
rect 4387 14365 4396 14399
rect 4344 14356 4396 14365
rect 8484 14424 8536 14476
rect 8760 14467 8812 14476
rect 8760 14433 8769 14467
rect 8769 14433 8803 14467
rect 8803 14433 8812 14467
rect 8760 14424 8812 14433
rect 11336 14424 11388 14476
rect 10232 14356 10284 14408
rect 15936 14560 15988 14612
rect 18328 14603 18380 14612
rect 18328 14569 18337 14603
rect 18337 14569 18371 14603
rect 18371 14569 18380 14603
rect 18328 14560 18380 14569
rect 15292 14424 15344 14476
rect 5724 14288 5776 14340
rect 12992 14356 13044 14408
rect 13360 14356 13412 14408
rect 14004 14356 14056 14408
rect 13912 14288 13964 14340
rect 2872 14220 2924 14272
rect 3792 14220 3844 14272
rect 4804 14220 4856 14272
rect 8760 14220 8812 14272
rect 9128 14220 9180 14272
rect 11520 14263 11572 14272
rect 11520 14229 11529 14263
rect 11529 14229 11563 14263
rect 11563 14229 11572 14263
rect 11520 14220 11572 14229
rect 12440 14220 12492 14272
rect 14740 14220 14792 14272
rect 14924 14263 14976 14272
rect 14924 14229 14933 14263
rect 14933 14229 14967 14263
rect 14967 14229 14976 14263
rect 14924 14220 14976 14229
rect 15660 14288 15712 14340
rect 16304 14399 16356 14408
rect 16304 14365 16313 14399
rect 16313 14365 16347 14399
rect 16347 14365 16356 14399
rect 16304 14356 16356 14365
rect 18696 14356 18748 14408
rect 16396 14263 16448 14272
rect 16396 14229 16405 14263
rect 16405 14229 16439 14263
rect 16439 14229 16448 14263
rect 16396 14220 16448 14229
rect 17592 14288 17644 14340
rect 17776 14220 17828 14272
rect 18144 14288 18196 14340
rect 18604 14288 18656 14340
rect 5398 14118 5450 14170
rect 5462 14118 5514 14170
rect 5526 14118 5578 14170
rect 5590 14118 5642 14170
rect 5654 14118 5706 14170
rect 9846 14118 9898 14170
rect 9910 14118 9962 14170
rect 9974 14118 10026 14170
rect 10038 14118 10090 14170
rect 10102 14118 10154 14170
rect 14294 14118 14346 14170
rect 14358 14118 14410 14170
rect 14422 14118 14474 14170
rect 14486 14118 14538 14170
rect 14550 14118 14602 14170
rect 3424 14016 3476 14068
rect 1952 13923 2004 13932
rect 1952 13889 1961 13923
rect 1961 13889 1995 13923
rect 1995 13889 2004 13923
rect 1952 13880 2004 13889
rect 2136 13880 2188 13932
rect 3976 13948 4028 14000
rect 3516 13923 3568 13932
rect 3516 13889 3525 13923
rect 3525 13889 3559 13923
rect 3559 13889 3568 13923
rect 3516 13880 3568 13889
rect 4252 13880 4304 13932
rect 5724 14016 5776 14068
rect 4528 13948 4580 14000
rect 4620 13923 4672 13932
rect 4620 13889 4629 13923
rect 4629 13889 4663 13923
rect 4663 13889 4672 13923
rect 4620 13880 4672 13889
rect 5080 13923 5132 13932
rect 5080 13889 5089 13923
rect 5089 13889 5123 13923
rect 5123 13889 5132 13923
rect 5080 13880 5132 13889
rect 5264 13923 5316 13932
rect 5264 13889 5273 13923
rect 5273 13889 5307 13923
rect 5307 13889 5316 13923
rect 5264 13880 5316 13889
rect 8116 14016 8168 14068
rect 9772 14016 9824 14068
rect 12440 14016 12492 14068
rect 12808 14016 12860 14068
rect 16304 14016 16356 14068
rect 7288 13948 7340 14000
rect 8576 13991 8628 14000
rect 8208 13880 8260 13932
rect 8576 13957 8610 13991
rect 8610 13957 8628 13991
rect 8576 13948 8628 13957
rect 9312 13948 9364 14000
rect 11060 13923 11112 13932
rect 2964 13812 3016 13864
rect 3332 13855 3384 13864
rect 3332 13821 3341 13855
rect 3341 13821 3375 13855
rect 3375 13821 3384 13855
rect 3332 13812 3384 13821
rect 8116 13812 8168 13864
rect 9496 13812 9548 13864
rect 4344 13676 4396 13728
rect 9588 13676 9640 13728
rect 11060 13889 11078 13923
rect 11078 13889 11112 13923
rect 11060 13880 11112 13889
rect 13728 13948 13780 14000
rect 11336 13923 11388 13932
rect 11336 13889 11345 13923
rect 11345 13889 11379 13923
rect 11379 13889 11388 13923
rect 11336 13880 11388 13889
rect 12808 13880 12860 13932
rect 13176 13880 13228 13932
rect 15200 13948 15252 14000
rect 16212 13991 16264 14000
rect 16212 13957 16230 13991
rect 16230 13957 16264 13991
rect 16212 13948 16264 13957
rect 12992 13812 13044 13864
rect 14188 13812 14240 13864
rect 14648 13855 14700 13864
rect 14648 13821 14657 13855
rect 14657 13821 14691 13855
rect 14691 13821 14700 13855
rect 14648 13812 14700 13821
rect 18420 13923 18472 13932
rect 18420 13889 18429 13923
rect 18429 13889 18463 13923
rect 18463 13889 18472 13923
rect 18420 13880 18472 13889
rect 14740 13744 14792 13796
rect 11704 13676 11756 13728
rect 12716 13676 12768 13728
rect 12900 13676 12952 13728
rect 14924 13676 14976 13728
rect 18328 13812 18380 13864
rect 18052 13719 18104 13728
rect 18052 13685 18061 13719
rect 18061 13685 18095 13719
rect 18095 13685 18104 13719
rect 18052 13676 18104 13685
rect 3174 13574 3226 13626
rect 3238 13574 3290 13626
rect 3302 13574 3354 13626
rect 3366 13574 3418 13626
rect 3430 13574 3482 13626
rect 7622 13574 7674 13626
rect 7686 13574 7738 13626
rect 7750 13574 7802 13626
rect 7814 13574 7866 13626
rect 7878 13574 7930 13626
rect 12070 13574 12122 13626
rect 12134 13574 12186 13626
rect 12198 13574 12250 13626
rect 12262 13574 12314 13626
rect 12326 13574 12378 13626
rect 16518 13574 16570 13626
rect 16582 13574 16634 13626
rect 16646 13574 16698 13626
rect 16710 13574 16762 13626
rect 16774 13574 16826 13626
rect 4988 13472 5040 13524
rect 5816 13472 5868 13524
rect 9404 13472 9456 13524
rect 2780 13404 2832 13456
rect 1952 13379 2004 13388
rect 1952 13345 1961 13379
rect 1961 13345 1995 13379
rect 1995 13345 2004 13379
rect 1952 13336 2004 13345
rect 3516 13404 3568 13456
rect 4068 13404 4120 13456
rect 14004 13472 14056 13524
rect 16396 13472 16448 13524
rect 3608 13336 3660 13388
rect 1860 13268 1912 13320
rect 3516 13268 3568 13320
rect 4252 13336 4304 13388
rect 11980 13336 12032 13388
rect 12900 13336 12952 13388
rect 17132 13379 17184 13388
rect 17132 13345 17141 13379
rect 17141 13345 17175 13379
rect 17175 13345 17184 13379
rect 17132 13336 17184 13345
rect 2964 13200 3016 13252
rect 4620 13268 4672 13320
rect 4804 13200 4856 13252
rect 5172 13311 5224 13320
rect 5172 13277 5181 13311
rect 5181 13277 5215 13311
rect 5215 13277 5224 13311
rect 5172 13268 5224 13277
rect 8116 13268 8168 13320
rect 9220 13268 9272 13320
rect 8484 13243 8536 13252
rect 8484 13209 8502 13243
rect 8502 13209 8536 13243
rect 8484 13200 8536 13209
rect 2688 13175 2740 13184
rect 2688 13141 2697 13175
rect 2697 13141 2731 13175
rect 2731 13141 2740 13175
rect 2688 13132 2740 13141
rect 3332 13132 3384 13184
rect 3884 13175 3936 13184
rect 3884 13141 3893 13175
rect 3893 13141 3927 13175
rect 3927 13141 3936 13175
rect 3884 13132 3936 13141
rect 3976 13132 4028 13184
rect 5080 13132 5132 13184
rect 5264 13175 5316 13184
rect 5264 13141 5273 13175
rect 5273 13141 5307 13175
rect 5307 13141 5316 13175
rect 5264 13132 5316 13141
rect 7380 13175 7432 13184
rect 7380 13141 7389 13175
rect 7389 13141 7423 13175
rect 7423 13141 7432 13175
rect 7380 13132 7432 13141
rect 7472 13132 7524 13184
rect 11520 13268 11572 13320
rect 13084 13268 13136 13320
rect 11796 13200 11848 13252
rect 13452 13200 13504 13252
rect 13636 13311 13688 13320
rect 13636 13277 13654 13311
rect 13654 13277 13688 13311
rect 13636 13268 13688 13277
rect 14188 13268 14240 13320
rect 15476 13311 15528 13320
rect 15476 13277 15485 13311
rect 15485 13277 15519 13311
rect 15519 13277 15528 13311
rect 15476 13268 15528 13277
rect 17868 13472 17920 13524
rect 17408 13336 17460 13388
rect 17776 13268 17828 13320
rect 10784 13132 10836 13184
rect 12072 13132 12124 13184
rect 12716 13132 12768 13184
rect 16212 13200 16264 13252
rect 16856 13243 16908 13252
rect 16856 13209 16874 13243
rect 16874 13209 16908 13243
rect 16856 13200 16908 13209
rect 14096 13175 14148 13184
rect 14096 13141 14105 13175
rect 14105 13141 14139 13175
rect 14139 13141 14148 13175
rect 14096 13132 14148 13141
rect 17776 13132 17828 13184
rect 5398 13030 5450 13082
rect 5462 13030 5514 13082
rect 5526 13030 5578 13082
rect 5590 13030 5642 13082
rect 5654 13030 5706 13082
rect 9846 13030 9898 13082
rect 9910 13030 9962 13082
rect 9974 13030 10026 13082
rect 10038 13030 10090 13082
rect 10102 13030 10154 13082
rect 14294 13030 14346 13082
rect 14358 13030 14410 13082
rect 14422 13030 14474 13082
rect 14486 13030 14538 13082
rect 14550 13030 14602 13082
rect 2320 12971 2372 12980
rect 2320 12937 2329 12971
rect 2329 12937 2363 12971
rect 2363 12937 2372 12971
rect 2320 12928 2372 12937
rect 2872 12860 2924 12912
rect 4344 12971 4396 12980
rect 4344 12937 4353 12971
rect 4353 12937 4387 12971
rect 4387 12937 4396 12971
rect 4344 12928 4396 12937
rect 4804 12971 4856 12980
rect 4804 12937 4813 12971
rect 4813 12937 4847 12971
rect 4847 12937 4856 12971
rect 4804 12928 4856 12937
rect 5080 12928 5132 12980
rect 5264 12928 5316 12980
rect 3700 12860 3752 12912
rect 3884 12860 3936 12912
rect 1768 12792 1820 12844
rect 2136 12724 2188 12776
rect 3332 12792 3384 12844
rect 4712 12792 4764 12844
rect 5264 12835 5316 12844
rect 3240 12767 3292 12776
rect 3240 12733 3249 12767
rect 3249 12733 3283 12767
rect 3283 12733 3292 12767
rect 3240 12724 3292 12733
rect 3884 12724 3936 12776
rect 4436 12767 4488 12776
rect 4436 12733 4445 12767
rect 4445 12733 4479 12767
rect 4479 12733 4488 12767
rect 4436 12724 4488 12733
rect 4620 12767 4672 12776
rect 4620 12733 4629 12767
rect 4629 12733 4663 12767
rect 4663 12733 4672 12767
rect 4620 12724 4672 12733
rect 5264 12801 5273 12835
rect 5273 12801 5307 12835
rect 5307 12801 5316 12835
rect 5264 12792 5316 12801
rect 5540 12835 5592 12844
rect 5540 12801 5549 12835
rect 5549 12801 5583 12835
rect 5583 12801 5592 12835
rect 5540 12792 5592 12801
rect 6184 12928 6236 12980
rect 8116 12860 8168 12912
rect 8852 12792 8904 12844
rect 9404 12792 9456 12844
rect 9680 12860 9732 12912
rect 11704 12860 11756 12912
rect 11428 12792 11480 12844
rect 12624 12835 12676 12844
rect 12992 12860 13044 12912
rect 12624 12801 12642 12835
rect 12642 12801 12676 12835
rect 12624 12792 12676 12801
rect 13452 12792 13504 12844
rect 15476 12860 15528 12912
rect 5172 12724 5224 12776
rect 7472 12724 7524 12776
rect 16028 12835 16080 12844
rect 16028 12801 16046 12835
rect 16046 12801 16080 12835
rect 16304 12860 16356 12912
rect 16488 12903 16540 12912
rect 16488 12869 16497 12903
rect 16497 12869 16531 12903
rect 16531 12869 16540 12903
rect 16488 12860 16540 12869
rect 17132 12860 17184 12912
rect 17408 12860 17460 12912
rect 18236 12903 18288 12912
rect 18236 12869 18245 12903
rect 18245 12869 18279 12903
rect 18279 12869 18288 12903
rect 18236 12860 18288 12869
rect 18512 12860 18564 12912
rect 16028 12792 16080 12801
rect 3056 12656 3108 12708
rect 4160 12656 4212 12708
rect 15016 12724 15068 12776
rect 17316 12792 17368 12844
rect 10600 12656 10652 12708
rect 1308 12588 1360 12640
rect 5356 12631 5408 12640
rect 5356 12597 5365 12631
rect 5365 12597 5399 12631
rect 5399 12597 5408 12631
rect 5356 12588 5408 12597
rect 6920 12588 6972 12640
rect 7380 12588 7432 12640
rect 11060 12588 11112 12640
rect 11244 12656 11296 12708
rect 11704 12656 11756 12708
rect 11888 12656 11940 12708
rect 13268 12656 13320 12708
rect 13544 12588 13596 12640
rect 15292 12656 15344 12708
rect 15108 12588 15160 12640
rect 16028 12588 16080 12640
rect 17040 12588 17092 12640
rect 3174 12486 3226 12538
rect 3238 12486 3290 12538
rect 3302 12486 3354 12538
rect 3366 12486 3418 12538
rect 3430 12486 3482 12538
rect 7622 12486 7674 12538
rect 7686 12486 7738 12538
rect 7750 12486 7802 12538
rect 7814 12486 7866 12538
rect 7878 12486 7930 12538
rect 12070 12486 12122 12538
rect 12134 12486 12186 12538
rect 12198 12486 12250 12538
rect 12262 12486 12314 12538
rect 12326 12486 12378 12538
rect 16518 12486 16570 12538
rect 16582 12486 16634 12538
rect 16646 12486 16698 12538
rect 16710 12486 16762 12538
rect 16774 12486 16826 12538
rect 3332 12384 3384 12436
rect 3516 12384 3568 12436
rect 4068 12384 4120 12436
rect 4436 12384 4488 12436
rect 4712 12384 4764 12436
rect 4804 12384 4856 12436
rect 5356 12316 5408 12368
rect 2780 12180 2832 12232
rect 3148 12223 3200 12232
rect 2412 12112 2464 12164
rect 3148 12189 3157 12223
rect 3157 12189 3191 12223
rect 3191 12189 3200 12223
rect 3148 12180 3200 12189
rect 3976 12291 4028 12300
rect 3976 12257 3985 12291
rect 3985 12257 4019 12291
rect 4019 12257 4028 12291
rect 3976 12248 4028 12257
rect 4252 12248 4304 12300
rect 3332 12180 3384 12232
rect 4804 12180 4856 12232
rect 4988 12223 5040 12232
rect 4988 12189 4997 12223
rect 4997 12189 5031 12223
rect 5031 12189 5040 12223
rect 4988 12180 5040 12189
rect 8576 12384 8628 12436
rect 13452 12427 13504 12436
rect 6000 12316 6052 12368
rect 8392 12316 8444 12368
rect 13452 12393 13461 12427
rect 13461 12393 13495 12427
rect 13495 12393 13504 12427
rect 13452 12384 13504 12393
rect 14096 12427 14148 12436
rect 14096 12393 14105 12427
rect 14105 12393 14139 12427
rect 14139 12393 14148 12427
rect 14096 12384 14148 12393
rect 14740 12384 14792 12436
rect 8208 12248 8260 12300
rect 6092 12180 6144 12232
rect 9220 12180 9272 12232
rect 11428 12291 11480 12300
rect 11428 12257 11437 12291
rect 11437 12257 11471 12291
rect 11471 12257 11480 12291
rect 11428 12248 11480 12257
rect 10692 12180 10744 12232
rect 5908 12112 5960 12164
rect 11336 12180 11388 12232
rect 11796 12223 11848 12232
rect 11796 12189 11830 12223
rect 11830 12189 11848 12223
rect 11796 12180 11848 12189
rect 12072 12180 12124 12232
rect 18052 12384 18104 12436
rect 17316 12316 17368 12368
rect 17592 12316 17644 12368
rect 17132 12291 17184 12300
rect 12808 12112 12860 12164
rect 1860 12044 1912 12096
rect 3884 12044 3936 12096
rect 4160 12044 4212 12096
rect 4804 12044 4856 12096
rect 5172 12044 5224 12096
rect 5632 12087 5684 12096
rect 5632 12053 5641 12087
rect 5641 12053 5675 12087
rect 5675 12053 5684 12087
rect 5632 12044 5684 12053
rect 5724 12044 5776 12096
rect 12900 12087 12952 12096
rect 12900 12053 12909 12087
rect 12909 12053 12943 12087
rect 12943 12053 12952 12087
rect 12900 12044 12952 12053
rect 13084 12087 13136 12096
rect 13084 12053 13093 12087
rect 13093 12053 13127 12087
rect 13127 12053 13136 12087
rect 13084 12044 13136 12053
rect 17132 12257 17141 12291
rect 17141 12257 17175 12291
rect 17175 12257 17184 12291
rect 17132 12248 17184 12257
rect 14096 12112 14148 12164
rect 14556 12112 14608 12164
rect 14648 12112 14700 12164
rect 15476 12223 15528 12232
rect 15476 12189 15485 12223
rect 15485 12189 15519 12223
rect 15519 12189 15528 12223
rect 17684 12223 17736 12232
rect 15476 12180 15528 12189
rect 17684 12189 17693 12223
rect 17693 12189 17727 12223
rect 17727 12189 17736 12223
rect 17684 12180 17736 12189
rect 18144 12248 18196 12300
rect 18236 12180 18288 12232
rect 14188 12044 14240 12096
rect 14740 12044 14792 12096
rect 16764 12112 16816 12164
rect 15476 12044 15528 12096
rect 17592 12112 17644 12164
rect 17132 12044 17184 12096
rect 5398 11942 5450 11994
rect 5462 11942 5514 11994
rect 5526 11942 5578 11994
rect 5590 11942 5642 11994
rect 5654 11942 5706 11994
rect 9846 11942 9898 11994
rect 9910 11942 9962 11994
rect 9974 11942 10026 11994
rect 10038 11942 10090 11994
rect 10102 11942 10154 11994
rect 14294 11942 14346 11994
rect 14358 11942 14410 11994
rect 14422 11942 14474 11994
rect 14486 11942 14538 11994
rect 14550 11942 14602 11994
rect 2964 11840 3016 11892
rect 3608 11840 3660 11892
rect 3976 11840 4028 11892
rect 5632 11883 5684 11892
rect 4160 11815 4212 11824
rect 4160 11781 4169 11815
rect 4169 11781 4203 11815
rect 4203 11781 4212 11815
rect 4160 11772 4212 11781
rect 2044 11704 2096 11756
rect 2964 11704 3016 11756
rect 4068 11704 4120 11756
rect 5080 11747 5132 11756
rect 4252 11713 4261 11740
rect 4261 11713 4295 11740
rect 4295 11713 4304 11740
rect 4252 11688 4304 11713
rect 5080 11713 5089 11747
rect 5089 11713 5123 11747
rect 5123 11713 5132 11747
rect 5080 11704 5132 11713
rect 1952 11679 2004 11688
rect 1952 11645 1961 11679
rect 1961 11645 1995 11679
rect 1995 11645 2004 11679
rect 1952 11636 2004 11645
rect 2228 11679 2280 11688
rect 2228 11645 2237 11679
rect 2237 11645 2271 11679
rect 2271 11645 2280 11679
rect 2228 11636 2280 11645
rect 2504 11679 2556 11688
rect 2504 11645 2513 11679
rect 2513 11645 2547 11679
rect 2547 11645 2556 11679
rect 2504 11636 2556 11645
rect 3608 11679 3660 11688
rect 3608 11645 3617 11679
rect 3617 11645 3651 11679
rect 3651 11645 3660 11679
rect 3608 11636 3660 11645
rect 3976 11679 4028 11688
rect 3976 11645 3985 11679
rect 3985 11645 4019 11679
rect 4019 11645 4028 11679
rect 3976 11636 4028 11645
rect 5172 11679 5224 11688
rect 5172 11645 5181 11679
rect 5181 11645 5215 11679
rect 5215 11645 5224 11679
rect 5172 11636 5224 11645
rect 5632 11849 5641 11883
rect 5641 11849 5675 11883
rect 5675 11849 5684 11883
rect 5632 11840 5684 11849
rect 6092 11840 6144 11892
rect 5816 11747 5868 11756
rect 5816 11713 5825 11747
rect 5825 11713 5859 11747
rect 5859 11713 5868 11747
rect 5816 11704 5868 11713
rect 8300 11840 8352 11892
rect 8576 11883 8628 11892
rect 8576 11849 8585 11883
rect 8585 11849 8619 11883
rect 8619 11849 8628 11883
rect 8576 11840 8628 11849
rect 9680 11840 9732 11892
rect 13820 11840 13872 11892
rect 15752 11840 15804 11892
rect 8116 11772 8168 11824
rect 8208 11772 8260 11824
rect 12992 11772 13044 11824
rect 7196 11747 7248 11756
rect 7196 11713 7205 11747
rect 7205 11713 7239 11747
rect 7239 11713 7248 11747
rect 7196 11704 7248 11713
rect 9220 11704 9272 11756
rect 12072 11704 12124 11756
rect 12900 11704 12952 11756
rect 14648 11747 14700 11756
rect 15384 11772 15436 11824
rect 18236 11815 18288 11824
rect 14648 11713 14666 11747
rect 14666 11713 14700 11747
rect 14648 11704 14700 11713
rect 16120 11747 16172 11756
rect 16120 11713 16138 11747
rect 16138 11713 16172 11747
rect 16120 11704 16172 11713
rect 16948 11704 17000 11756
rect 17316 11704 17368 11756
rect 17776 11747 17828 11756
rect 18236 11781 18245 11815
rect 18245 11781 18279 11815
rect 18279 11781 18288 11815
rect 18236 11772 18288 11781
rect 18420 11815 18472 11824
rect 18420 11781 18429 11815
rect 18429 11781 18463 11815
rect 18463 11781 18472 11815
rect 18420 11772 18472 11781
rect 17776 11713 17805 11747
rect 17805 11713 17828 11747
rect 17776 11704 17828 11713
rect 5908 11611 5960 11620
rect 5908 11577 5917 11611
rect 5917 11577 5951 11611
rect 5951 11577 5960 11611
rect 5908 11568 5960 11577
rect 6000 11568 6052 11620
rect 13544 11636 13596 11688
rect 13728 11636 13780 11688
rect 2412 11500 2464 11552
rect 4252 11500 4304 11552
rect 4344 11500 4396 11552
rect 4804 11500 4856 11552
rect 11612 11543 11664 11552
rect 11612 11509 11621 11543
rect 11621 11509 11655 11543
rect 11655 11509 11664 11543
rect 11612 11500 11664 11509
rect 15108 11500 15160 11552
rect 16580 11500 16632 11552
rect 17684 11500 17736 11552
rect 3174 11398 3226 11450
rect 3238 11398 3290 11450
rect 3302 11398 3354 11450
rect 3366 11398 3418 11450
rect 3430 11398 3482 11450
rect 7622 11398 7674 11450
rect 7686 11398 7738 11450
rect 7750 11398 7802 11450
rect 7814 11398 7866 11450
rect 7878 11398 7930 11450
rect 12070 11398 12122 11450
rect 12134 11398 12186 11450
rect 12198 11398 12250 11450
rect 12262 11398 12314 11450
rect 12326 11398 12378 11450
rect 16518 11398 16570 11450
rect 16582 11398 16634 11450
rect 16646 11398 16698 11450
rect 16710 11398 16762 11450
rect 16774 11398 16826 11450
rect 2872 11339 2924 11348
rect 2872 11305 2881 11339
rect 2881 11305 2915 11339
rect 2915 11305 2924 11339
rect 2872 11296 2924 11305
rect 2228 11228 2280 11280
rect 2596 11271 2648 11280
rect 2596 11237 2605 11271
rect 2605 11237 2639 11271
rect 2639 11237 2648 11271
rect 2596 11228 2648 11237
rect 2780 11271 2832 11280
rect 2780 11237 2789 11271
rect 2789 11237 2823 11271
rect 2823 11237 2832 11271
rect 2780 11228 2832 11237
rect 2964 11228 3016 11280
rect 7196 11296 7248 11348
rect 7380 11296 7432 11348
rect 8116 11296 8168 11348
rect 8944 11271 8996 11280
rect 2228 11135 2280 11144
rect 2228 11101 2237 11135
rect 2237 11101 2271 11135
rect 2271 11101 2280 11135
rect 2228 11092 2280 11101
rect 3884 11160 3936 11212
rect 4068 11160 4120 11212
rect 4160 11160 4212 11212
rect 3148 11092 3200 11144
rect 3608 11092 3660 11144
rect 4344 11135 4396 11144
rect 4344 11101 4353 11135
rect 4353 11101 4387 11135
rect 4387 11101 4396 11135
rect 4344 11092 4396 11101
rect 2872 11024 2924 11076
rect 8944 11237 8953 11271
rect 8953 11237 8987 11271
rect 8987 11237 8996 11271
rect 8944 11228 8996 11237
rect 11152 11296 11204 11348
rect 11980 11296 12032 11348
rect 12072 11296 12124 11348
rect 14004 11296 14056 11348
rect 13728 11228 13780 11280
rect 13912 11228 13964 11280
rect 16120 11228 16172 11280
rect 6644 11160 6696 11212
rect 9220 11160 9272 11212
rect 9680 11092 9732 11144
rect 13084 11092 13136 11144
rect 14740 11160 14792 11212
rect 18236 11228 18288 11280
rect 15752 11092 15804 11144
rect 16212 11092 16264 11144
rect 17684 11135 17736 11144
rect 9404 11024 9456 11076
rect 9588 11024 9640 11076
rect 11428 11024 11480 11076
rect 11796 11024 11848 11076
rect 11980 11067 12032 11076
rect 11980 11033 11998 11067
rect 11998 11033 12032 11067
rect 11980 11024 12032 11033
rect 12716 11024 12768 11076
rect 13544 11024 13596 11076
rect 3056 10956 3108 11008
rect 3884 10999 3936 11008
rect 3884 10965 3893 10999
rect 3893 10965 3927 10999
rect 3927 10965 3936 10999
rect 3884 10956 3936 10965
rect 4436 10999 4488 11008
rect 4436 10965 4445 10999
rect 4445 10965 4479 10999
rect 4479 10965 4488 10999
rect 4436 10956 4488 10965
rect 4988 10999 5040 11008
rect 4988 10965 4997 10999
rect 4997 10965 5031 10999
rect 5031 10965 5040 10999
rect 4988 10956 5040 10965
rect 5816 10956 5868 11008
rect 6092 10999 6144 11008
rect 6092 10965 6101 10999
rect 6101 10965 6135 10999
rect 6135 10965 6144 10999
rect 6092 10956 6144 10965
rect 10416 10956 10468 11008
rect 11704 10956 11756 11008
rect 15476 11024 15528 11076
rect 15568 11067 15620 11076
rect 15568 11033 15586 11067
rect 15586 11033 15620 11067
rect 15568 11024 15620 11033
rect 15936 11024 15988 11076
rect 16396 11024 16448 11076
rect 16948 11024 17000 11076
rect 17132 11024 17184 11076
rect 15660 10956 15712 11008
rect 17684 11101 17693 11135
rect 17693 11101 17727 11135
rect 17727 11101 17736 11135
rect 17684 11092 17736 11101
rect 18604 11092 18656 11144
rect 18052 11024 18104 11076
rect 18512 11024 18564 11076
rect 18972 10956 19024 11008
rect 5398 10854 5450 10906
rect 5462 10854 5514 10906
rect 5526 10854 5578 10906
rect 5590 10854 5642 10906
rect 5654 10854 5706 10906
rect 9846 10854 9898 10906
rect 9910 10854 9962 10906
rect 9974 10854 10026 10906
rect 10038 10854 10090 10906
rect 10102 10854 10154 10906
rect 14294 10854 14346 10906
rect 14358 10854 14410 10906
rect 14422 10854 14474 10906
rect 14486 10854 14538 10906
rect 14550 10854 14602 10906
rect 4436 10752 4488 10804
rect 4988 10752 5040 10804
rect 2688 10684 2740 10736
rect 3884 10684 3936 10736
rect 4068 10684 4120 10736
rect 2412 10659 2464 10668
rect 2412 10625 2421 10659
rect 2421 10625 2455 10659
rect 2455 10625 2464 10659
rect 2412 10616 2464 10625
rect 2964 10616 3016 10668
rect 3792 10616 3844 10668
rect 4160 10616 4212 10668
rect 1952 10591 2004 10600
rect 1952 10557 1961 10591
rect 1961 10557 1995 10591
rect 1995 10557 2004 10591
rect 1952 10548 2004 10557
rect 2780 10548 2832 10600
rect 3608 10548 3660 10600
rect 3884 10591 3936 10600
rect 3884 10557 3893 10591
rect 3893 10557 3927 10591
rect 3927 10557 3936 10591
rect 3884 10548 3936 10557
rect 4712 10548 4764 10600
rect 4988 10548 5040 10600
rect 5908 10684 5960 10736
rect 9404 10795 9456 10804
rect 9404 10761 9413 10795
rect 9413 10761 9447 10795
rect 9447 10761 9456 10795
rect 9404 10752 9456 10761
rect 9588 10752 9640 10804
rect 11152 10752 11204 10804
rect 12808 10752 12860 10804
rect 16028 10752 16080 10804
rect 17776 10752 17828 10804
rect 9312 10684 9364 10736
rect 9680 10684 9732 10736
rect 5724 10659 5776 10668
rect 5724 10625 5733 10659
rect 5733 10625 5767 10659
rect 5767 10625 5776 10659
rect 5724 10616 5776 10625
rect 6184 10616 6236 10668
rect 7104 10616 7156 10668
rect 5632 10591 5684 10600
rect 5632 10557 5641 10591
rect 5641 10557 5675 10591
rect 5675 10557 5684 10591
rect 5632 10548 5684 10557
rect 6276 10548 6328 10600
rect 7196 10548 7248 10600
rect 7380 10548 7432 10600
rect 5816 10480 5868 10532
rect 3516 10412 3568 10464
rect 4988 10412 5040 10464
rect 5356 10412 5408 10464
rect 6552 10412 6604 10464
rect 10600 10616 10652 10668
rect 11060 10659 11112 10668
rect 11796 10684 11848 10736
rect 11060 10625 11078 10659
rect 11078 10625 11112 10659
rect 11060 10616 11112 10625
rect 11704 10616 11756 10668
rect 15660 10684 15712 10736
rect 14556 10616 14608 10668
rect 15384 10659 15436 10668
rect 15384 10625 15393 10659
rect 15393 10625 15427 10659
rect 15427 10625 15436 10659
rect 16212 10684 16264 10736
rect 17500 10727 17552 10736
rect 17500 10693 17509 10727
rect 17509 10693 17543 10727
rect 17543 10693 17552 10727
rect 17500 10684 17552 10693
rect 15384 10616 15436 10625
rect 15936 10616 15988 10668
rect 16304 10659 16356 10668
rect 16304 10625 16313 10659
rect 16313 10625 16347 10659
rect 16347 10625 16356 10659
rect 16304 10616 16356 10625
rect 17224 10616 17276 10668
rect 18052 10616 18104 10668
rect 17592 10548 17644 10600
rect 17684 10591 17736 10600
rect 17684 10557 17693 10591
rect 17693 10557 17727 10591
rect 17727 10557 17736 10591
rect 17684 10548 17736 10557
rect 18144 10548 18196 10600
rect 9772 10480 9824 10532
rect 16948 10523 17000 10532
rect 9128 10412 9180 10464
rect 10416 10412 10468 10464
rect 12440 10412 12492 10464
rect 14188 10412 14240 10464
rect 15936 10455 15988 10464
rect 15936 10421 15945 10455
rect 15945 10421 15979 10455
rect 15979 10421 15988 10455
rect 15936 10412 15988 10421
rect 16212 10455 16264 10464
rect 16212 10421 16221 10455
rect 16221 10421 16255 10455
rect 16255 10421 16264 10455
rect 16212 10412 16264 10421
rect 16948 10489 16957 10523
rect 16957 10489 16991 10523
rect 16991 10489 17000 10523
rect 16948 10480 17000 10489
rect 17132 10412 17184 10464
rect 18696 10412 18748 10464
rect 3174 10310 3226 10362
rect 3238 10310 3290 10362
rect 3302 10310 3354 10362
rect 3366 10310 3418 10362
rect 3430 10310 3482 10362
rect 7622 10310 7674 10362
rect 7686 10310 7738 10362
rect 7750 10310 7802 10362
rect 7814 10310 7866 10362
rect 7878 10310 7930 10362
rect 12070 10310 12122 10362
rect 12134 10310 12186 10362
rect 12198 10310 12250 10362
rect 12262 10310 12314 10362
rect 12326 10310 12378 10362
rect 16518 10310 16570 10362
rect 16582 10310 16634 10362
rect 16646 10310 16698 10362
rect 16710 10310 16762 10362
rect 16774 10310 16826 10362
rect 2872 10208 2924 10260
rect 3516 10208 3568 10260
rect 4160 10251 4212 10260
rect 4160 10217 4169 10251
rect 4169 10217 4203 10251
rect 4203 10217 4212 10251
rect 4160 10208 4212 10217
rect 5632 10208 5684 10260
rect 6828 10208 6880 10260
rect 7196 10208 7248 10260
rect 13636 10208 13688 10260
rect 17684 10208 17736 10260
rect 2780 10140 2832 10192
rect 2504 10115 2556 10124
rect 2504 10081 2513 10115
rect 2513 10081 2547 10115
rect 2547 10081 2556 10115
rect 2504 10072 2556 10081
rect 3608 10072 3660 10124
rect 3792 10072 3844 10124
rect 4712 10115 4764 10124
rect 4712 10081 4721 10115
rect 4721 10081 4755 10115
rect 4755 10081 4764 10115
rect 4712 10072 4764 10081
rect 4804 10072 4856 10124
rect 6184 10140 6236 10192
rect 13452 10183 13504 10192
rect 13452 10149 13461 10183
rect 13461 10149 13495 10183
rect 13495 10149 13504 10183
rect 13452 10140 13504 10149
rect 14004 10140 14056 10192
rect 14556 10183 14608 10192
rect 14556 10149 14565 10183
rect 14565 10149 14599 10183
rect 14599 10149 14608 10183
rect 14556 10140 14608 10149
rect 16028 10183 16080 10192
rect 16028 10149 16037 10183
rect 16037 10149 16071 10183
rect 16071 10149 16080 10183
rect 16028 10140 16080 10149
rect 17592 10183 17644 10192
rect 17592 10149 17601 10183
rect 17601 10149 17635 10183
rect 17635 10149 17644 10183
rect 17592 10140 17644 10149
rect 6276 10072 6328 10124
rect 7288 10072 7340 10124
rect 8944 10072 8996 10124
rect 9956 10072 10008 10124
rect 11796 10072 11848 10124
rect 17960 10115 18012 10124
rect 17960 10081 17969 10115
rect 17969 10081 18003 10115
rect 18003 10081 18012 10115
rect 17960 10072 18012 10081
rect 1400 10047 1452 10056
rect 1400 10013 1409 10047
rect 1409 10013 1443 10047
rect 1443 10013 1452 10047
rect 1400 10004 1452 10013
rect 2872 10004 2924 10056
rect 3700 10004 3752 10056
rect 4068 10004 4120 10056
rect 6184 10004 6236 10056
rect 6552 10047 6604 10056
rect 6552 10013 6561 10047
rect 6561 10013 6595 10047
rect 6595 10013 6604 10047
rect 6552 10004 6604 10013
rect 7380 10047 7432 10056
rect 7380 10013 7389 10047
rect 7389 10013 7423 10047
rect 7423 10013 7432 10047
rect 7380 10004 7432 10013
rect 7656 10047 7708 10056
rect 7656 10013 7690 10047
rect 7690 10013 7708 10047
rect 7656 10004 7708 10013
rect 9220 10004 9272 10056
rect 9772 10004 9824 10056
rect 2780 9868 2832 9920
rect 5080 9936 5132 9988
rect 7472 9936 7524 9988
rect 9864 9936 9916 9988
rect 15292 10004 15344 10056
rect 15384 10004 15436 10056
rect 17316 10004 17368 10056
rect 10600 9936 10652 9988
rect 15200 9936 15252 9988
rect 15660 9979 15712 9988
rect 15660 9945 15678 9979
rect 15678 9945 15712 9979
rect 15660 9936 15712 9945
rect 3332 9911 3384 9920
rect 3332 9877 3341 9911
rect 3341 9877 3375 9911
rect 3375 9877 3384 9911
rect 3332 9868 3384 9877
rect 3516 9868 3568 9920
rect 4068 9868 4120 9920
rect 4620 9911 4672 9920
rect 4620 9877 4629 9911
rect 4629 9877 4663 9911
rect 4663 9877 4672 9911
rect 4620 9868 4672 9877
rect 5724 9911 5776 9920
rect 5724 9877 5733 9911
rect 5733 9877 5767 9911
rect 5767 9877 5776 9911
rect 5724 9868 5776 9877
rect 6920 9911 6972 9920
rect 6920 9877 6929 9911
rect 6929 9877 6963 9911
rect 6963 9877 6972 9911
rect 6920 9868 6972 9877
rect 8392 9868 8444 9920
rect 9404 9868 9456 9920
rect 9956 9868 10008 9920
rect 11704 9868 11756 9920
rect 13912 9911 13964 9920
rect 13912 9877 13921 9911
rect 13921 9877 13955 9911
rect 13955 9877 13964 9911
rect 13912 9868 13964 9877
rect 14648 9868 14700 9920
rect 15108 9868 15160 9920
rect 16488 9868 16540 9920
rect 17868 10004 17920 10056
rect 5398 9766 5450 9818
rect 5462 9766 5514 9818
rect 5526 9766 5578 9818
rect 5590 9766 5642 9818
rect 5654 9766 5706 9818
rect 9846 9766 9898 9818
rect 9910 9766 9962 9818
rect 9974 9766 10026 9818
rect 10038 9766 10090 9818
rect 10102 9766 10154 9818
rect 14294 9766 14346 9818
rect 14358 9766 14410 9818
rect 14422 9766 14474 9818
rect 14486 9766 14538 9818
rect 14550 9766 14602 9818
rect 2964 9664 3016 9716
rect 3332 9664 3384 9716
rect 4068 9707 4120 9716
rect 4068 9673 4077 9707
rect 4077 9673 4111 9707
rect 4111 9673 4120 9707
rect 4068 9664 4120 9673
rect 4160 9664 4212 9716
rect 4620 9664 4672 9716
rect 4896 9664 4948 9716
rect 5724 9664 5776 9716
rect 6460 9664 6512 9716
rect 7656 9664 7708 9716
rect 8392 9664 8444 9716
rect 11244 9664 11296 9716
rect 6736 9639 6788 9648
rect 6736 9605 6745 9639
rect 6745 9605 6779 9639
rect 6779 9605 6788 9639
rect 6736 9596 6788 9605
rect 2228 9571 2280 9580
rect 2228 9537 2237 9571
rect 2237 9537 2271 9571
rect 2271 9537 2280 9571
rect 2228 9528 2280 9537
rect 2780 9528 2832 9580
rect 3332 9528 3384 9580
rect 1952 9503 2004 9512
rect 1952 9469 1961 9503
rect 1961 9469 1995 9503
rect 1995 9469 2004 9503
rect 1952 9460 2004 9469
rect 2872 9503 2924 9512
rect 2872 9469 2881 9503
rect 2881 9469 2915 9503
rect 2915 9469 2924 9503
rect 2872 9460 2924 9469
rect 3608 9528 3660 9580
rect 5356 9528 5408 9580
rect 6552 9528 6604 9580
rect 7380 9528 7432 9580
rect 8024 9528 8076 9580
rect 8300 9528 8352 9580
rect 9772 9596 9824 9648
rect 9864 9596 9916 9648
rect 10784 9596 10836 9648
rect 11060 9639 11112 9648
rect 11060 9605 11078 9639
rect 11078 9605 11112 9639
rect 11060 9596 11112 9605
rect 12624 9664 12676 9716
rect 14096 9664 14148 9716
rect 14924 9664 14976 9716
rect 15292 9664 15344 9716
rect 16488 9664 16540 9716
rect 17500 9664 17552 9716
rect 17868 9664 17920 9716
rect 18052 9707 18104 9716
rect 18052 9673 18061 9707
rect 18061 9673 18095 9707
rect 18095 9673 18104 9707
rect 18052 9664 18104 9673
rect 13820 9639 13872 9648
rect 2964 9392 3016 9444
rect 3792 9460 3844 9512
rect 4344 9460 4396 9512
rect 5264 9460 5316 9512
rect 6828 9503 6880 9512
rect 6828 9469 6837 9503
rect 6837 9469 6871 9503
rect 6871 9469 6880 9503
rect 6828 9460 6880 9469
rect 6920 9460 6972 9512
rect 8116 9460 8168 9512
rect 9404 9528 9456 9580
rect 10048 9528 10100 9580
rect 11796 9528 11848 9580
rect 9680 9503 9732 9512
rect 6460 9392 6512 9444
rect 7564 9392 7616 9444
rect 8208 9392 8260 9444
rect 9680 9469 9689 9503
rect 9689 9469 9723 9503
rect 9723 9469 9732 9503
rect 9680 9460 9732 9469
rect 12624 9528 12676 9580
rect 13360 9528 13412 9580
rect 13820 9605 13854 9639
rect 13854 9605 13872 9639
rect 13820 9596 13872 9605
rect 13912 9596 13964 9648
rect 18420 9639 18472 9648
rect 18420 9605 18429 9639
rect 18429 9605 18463 9639
rect 18463 9605 18472 9639
rect 18420 9596 18472 9605
rect 14740 9528 14792 9580
rect 14924 9528 14976 9580
rect 13544 9503 13596 9512
rect 5264 9324 5316 9376
rect 6736 9324 6788 9376
rect 8576 9324 8628 9376
rect 9956 9367 10008 9376
rect 9956 9333 9965 9367
rect 9965 9333 9999 9367
rect 9999 9333 10008 9367
rect 9956 9324 10008 9333
rect 11336 9392 11388 9444
rect 11520 9435 11572 9444
rect 11520 9401 11529 9435
rect 11529 9401 11563 9435
rect 11563 9401 11572 9435
rect 11520 9392 11572 9401
rect 10600 9324 10652 9376
rect 10968 9324 11020 9376
rect 13544 9469 13553 9503
rect 13553 9469 13587 9503
rect 13587 9469 13596 9503
rect 13544 9460 13596 9469
rect 17316 9460 17368 9512
rect 13452 9367 13504 9376
rect 13452 9333 13461 9367
rect 13461 9333 13495 9367
rect 13495 9333 13504 9367
rect 15384 9392 15436 9444
rect 14924 9367 14976 9376
rect 13452 9324 13504 9333
rect 14924 9333 14933 9367
rect 14933 9333 14967 9367
rect 14967 9333 14976 9367
rect 14924 9324 14976 9333
rect 15016 9367 15068 9376
rect 15016 9333 15025 9367
rect 15025 9333 15059 9367
rect 15059 9333 15068 9367
rect 15016 9324 15068 9333
rect 15292 9324 15344 9376
rect 17592 9571 17644 9580
rect 17592 9537 17601 9571
rect 17601 9537 17635 9571
rect 17635 9537 17644 9571
rect 17592 9528 17644 9537
rect 17868 9503 17920 9512
rect 17868 9469 17877 9503
rect 17877 9469 17911 9503
rect 17911 9469 17920 9503
rect 17868 9460 17920 9469
rect 17960 9392 18012 9444
rect 16948 9367 17000 9376
rect 16948 9333 16957 9367
rect 16957 9333 16991 9367
rect 16991 9333 17000 9367
rect 16948 9324 17000 9333
rect 17500 9324 17552 9376
rect 3174 9222 3226 9274
rect 3238 9222 3290 9274
rect 3302 9222 3354 9274
rect 3366 9222 3418 9274
rect 3430 9222 3482 9274
rect 7622 9222 7674 9274
rect 7686 9222 7738 9274
rect 7750 9222 7802 9274
rect 7814 9222 7866 9274
rect 7878 9222 7930 9274
rect 12070 9222 12122 9274
rect 12134 9222 12186 9274
rect 12198 9222 12250 9274
rect 12262 9222 12314 9274
rect 12326 9222 12378 9274
rect 16518 9222 16570 9274
rect 16582 9222 16634 9274
rect 16646 9222 16698 9274
rect 16710 9222 16762 9274
rect 16774 9222 16826 9274
rect 3700 9120 3752 9172
rect 3884 9120 3936 9172
rect 4896 9120 4948 9172
rect 6276 9120 6328 9172
rect 6644 9120 6696 9172
rect 6828 9120 6880 9172
rect 2504 9027 2556 9036
rect 2504 8993 2513 9027
rect 2513 8993 2547 9027
rect 2547 8993 2556 9027
rect 2504 8984 2556 8993
rect 5172 9052 5224 9104
rect 2780 8984 2832 9036
rect 1952 8959 2004 8968
rect 1952 8925 1961 8959
rect 1961 8925 1995 8959
rect 1995 8925 2004 8959
rect 1952 8916 2004 8925
rect 3792 8916 3844 8968
rect 4160 8959 4212 8968
rect 4160 8925 4169 8959
rect 4169 8925 4203 8959
rect 4203 8925 4212 8959
rect 4160 8916 4212 8925
rect 4712 8984 4764 9036
rect 7288 9052 7340 9104
rect 6920 8984 6972 9036
rect 7196 8984 7248 9036
rect 10232 9052 10284 9104
rect 4528 8916 4580 8968
rect 5264 8916 5316 8968
rect 6828 8916 6880 8968
rect 7380 8959 7432 8968
rect 7380 8925 7389 8959
rect 7389 8925 7423 8959
rect 7423 8925 7432 8959
rect 7380 8916 7432 8925
rect 8392 8984 8444 9036
rect 8760 8984 8812 9036
rect 8024 8916 8076 8968
rect 3240 8891 3292 8900
rect 3240 8857 3249 8891
rect 3249 8857 3283 8891
rect 3283 8857 3292 8891
rect 3240 8848 3292 8857
rect 3608 8848 3660 8900
rect 5080 8848 5132 8900
rect 6460 8848 6512 8900
rect 8484 8848 8536 8900
rect 9680 8848 9732 8900
rect 4160 8780 4212 8832
rect 4436 8780 4488 8832
rect 4896 8823 4948 8832
rect 4896 8789 4905 8823
rect 4905 8789 4939 8823
rect 4939 8789 4948 8823
rect 4896 8780 4948 8789
rect 5172 8780 5224 8832
rect 5908 8780 5960 8832
rect 6644 8823 6696 8832
rect 6644 8789 6653 8823
rect 6653 8789 6687 8823
rect 6687 8789 6696 8823
rect 6644 8780 6696 8789
rect 8392 8780 8444 8832
rect 8760 8823 8812 8832
rect 8760 8789 8769 8823
rect 8769 8789 8803 8823
rect 8803 8789 8812 8823
rect 8760 8780 8812 8789
rect 9588 8780 9640 8832
rect 9864 8780 9916 8832
rect 10600 9120 10652 9172
rect 12164 9120 12216 9172
rect 13176 9120 13228 9172
rect 13820 9120 13872 9172
rect 14832 9120 14884 9172
rect 15016 9120 15068 9172
rect 15752 9120 15804 9172
rect 16304 9120 16356 9172
rect 16856 9120 16908 9172
rect 13636 9052 13688 9104
rect 14096 9052 14148 9104
rect 11796 9027 11848 9036
rect 11796 8993 11805 9027
rect 11805 8993 11839 9027
rect 11839 8993 11848 9027
rect 11796 8984 11848 8993
rect 11244 8916 11296 8968
rect 10784 8848 10836 8900
rect 11704 8916 11756 8968
rect 12624 8916 12676 8968
rect 13084 8984 13136 9036
rect 15200 8984 15252 9036
rect 15384 8984 15436 9036
rect 17316 9120 17368 9172
rect 13544 8916 13596 8968
rect 15568 8959 15620 8968
rect 15568 8925 15577 8959
rect 15577 8925 15611 8959
rect 15611 8925 15620 8959
rect 15568 8916 15620 8925
rect 16396 8916 16448 8968
rect 13176 8780 13228 8832
rect 13452 8823 13504 8832
rect 13452 8789 13461 8823
rect 13461 8789 13495 8823
rect 13495 8789 13504 8823
rect 13452 8780 13504 8789
rect 13544 8780 13596 8832
rect 14188 8848 14240 8900
rect 15476 8823 15528 8832
rect 15476 8789 15485 8823
rect 15485 8789 15519 8823
rect 15519 8789 15528 8823
rect 15476 8780 15528 8789
rect 16304 8780 16356 8832
rect 17500 8780 17552 8832
rect 18788 8780 18840 8832
rect 5398 8678 5450 8730
rect 5462 8678 5514 8730
rect 5526 8678 5578 8730
rect 5590 8678 5642 8730
rect 5654 8678 5706 8730
rect 9846 8678 9898 8730
rect 9910 8678 9962 8730
rect 9974 8678 10026 8730
rect 10038 8678 10090 8730
rect 10102 8678 10154 8730
rect 14294 8678 14346 8730
rect 14358 8678 14410 8730
rect 14422 8678 14474 8730
rect 14486 8678 14538 8730
rect 14550 8678 14602 8730
rect 3976 8576 4028 8628
rect 4436 8619 4488 8628
rect 4436 8585 4445 8619
rect 4445 8585 4479 8619
rect 4479 8585 4488 8619
rect 4436 8576 4488 8585
rect 4528 8576 4580 8628
rect 8024 8576 8076 8628
rect 10784 8576 10836 8628
rect 12716 8619 12768 8628
rect 2228 8508 2280 8560
rect 7012 8508 7064 8560
rect 7288 8508 7340 8560
rect 11060 8508 11112 8560
rect 12716 8585 12725 8619
rect 12725 8585 12759 8619
rect 12759 8585 12768 8619
rect 12716 8576 12768 8585
rect 13912 8576 13964 8628
rect 15200 8576 15252 8628
rect 15384 8576 15436 8628
rect 16028 8619 16080 8628
rect 12900 8508 12952 8560
rect 13636 8508 13688 8560
rect 2044 8440 2096 8492
rect 3516 8440 3568 8492
rect 4160 8440 4212 8492
rect 5080 8483 5132 8492
rect 5080 8449 5089 8483
rect 5089 8449 5123 8483
rect 5123 8449 5132 8483
rect 5080 8440 5132 8449
rect 5264 8440 5316 8492
rect 2780 8372 2832 8424
rect 2964 8372 3016 8424
rect 3608 8372 3660 8424
rect 3700 8372 3752 8424
rect 3884 8372 3936 8424
rect 7196 8440 7248 8492
rect 7748 8440 7800 8492
rect 4712 8347 4764 8356
rect 4712 8313 4721 8347
rect 4721 8313 4755 8347
rect 4755 8313 4764 8347
rect 4712 8304 4764 8313
rect 5724 8372 5776 8424
rect 6920 8415 6972 8424
rect 6920 8381 6929 8415
rect 6929 8381 6963 8415
rect 6963 8381 6972 8415
rect 6920 8372 6972 8381
rect 8392 8440 8444 8492
rect 8024 8415 8076 8424
rect 8024 8381 8033 8415
rect 8033 8381 8067 8415
rect 8067 8381 8076 8415
rect 8024 8372 8076 8381
rect 8116 8415 8168 8424
rect 8116 8381 8125 8415
rect 8125 8381 8159 8415
rect 8159 8381 8168 8415
rect 9864 8483 9916 8492
rect 9864 8449 9873 8483
rect 9873 8449 9907 8483
rect 9907 8449 9916 8483
rect 9864 8440 9916 8449
rect 10048 8440 10100 8492
rect 10600 8440 10652 8492
rect 12440 8440 12492 8492
rect 13820 8483 13872 8492
rect 13820 8449 13838 8483
rect 13838 8449 13872 8483
rect 13820 8440 13872 8449
rect 14188 8483 14240 8492
rect 14188 8449 14197 8483
rect 14197 8449 14231 8483
rect 14231 8449 14240 8483
rect 15568 8508 15620 8560
rect 16028 8585 16037 8619
rect 16037 8585 16071 8619
rect 16071 8585 16080 8619
rect 16028 8576 16080 8585
rect 18052 8576 18104 8628
rect 18420 8619 18472 8628
rect 18420 8585 18429 8619
rect 18429 8585 18463 8619
rect 18463 8585 18472 8619
rect 18420 8576 18472 8585
rect 14188 8440 14240 8449
rect 14832 8483 14884 8492
rect 14832 8449 14866 8483
rect 14866 8449 14884 8483
rect 14832 8440 14884 8449
rect 16304 8440 16356 8492
rect 17500 8483 17552 8492
rect 8116 8372 8168 8381
rect 4436 8236 4488 8288
rect 4528 8279 4580 8288
rect 4528 8245 4537 8279
rect 4537 8245 4571 8279
rect 4571 8245 4580 8279
rect 4528 8236 4580 8245
rect 4896 8236 4948 8288
rect 5264 8236 5316 8288
rect 6276 8236 6328 8288
rect 7472 8304 7524 8356
rect 11428 8372 11480 8424
rect 11980 8415 12032 8424
rect 11980 8381 11989 8415
rect 11989 8381 12023 8415
rect 12023 8381 12032 8415
rect 11980 8372 12032 8381
rect 8484 8347 8536 8356
rect 8484 8313 8493 8347
rect 8493 8313 8527 8347
rect 8527 8313 8536 8347
rect 8484 8304 8536 8313
rect 9864 8304 9916 8356
rect 11060 8304 11112 8356
rect 11796 8304 11848 8356
rect 12624 8372 12676 8424
rect 16120 8304 16172 8356
rect 7748 8236 7800 8288
rect 9128 8236 9180 8288
rect 11428 8236 11480 8288
rect 13452 8236 13504 8288
rect 16948 8304 17000 8356
rect 17500 8449 17509 8483
rect 17509 8449 17543 8483
rect 17543 8449 17552 8483
rect 17500 8440 17552 8449
rect 18236 8483 18288 8492
rect 18236 8449 18245 8483
rect 18245 8449 18279 8483
rect 18279 8449 18288 8483
rect 18236 8440 18288 8449
rect 17224 8415 17276 8424
rect 17224 8381 17233 8415
rect 17233 8381 17267 8415
rect 17267 8381 17276 8415
rect 17224 8372 17276 8381
rect 17316 8372 17368 8424
rect 17408 8236 17460 8288
rect 17868 8279 17920 8288
rect 17868 8245 17877 8279
rect 17877 8245 17911 8279
rect 17911 8245 17920 8279
rect 17868 8236 17920 8245
rect 18328 8236 18380 8288
rect 3174 8134 3226 8186
rect 3238 8134 3290 8186
rect 3302 8134 3354 8186
rect 3366 8134 3418 8186
rect 3430 8134 3482 8186
rect 7622 8134 7674 8186
rect 7686 8134 7738 8186
rect 7750 8134 7802 8186
rect 7814 8134 7866 8186
rect 7878 8134 7930 8186
rect 12070 8134 12122 8186
rect 12134 8134 12186 8186
rect 12198 8134 12250 8186
rect 12262 8134 12314 8186
rect 12326 8134 12378 8186
rect 16518 8134 16570 8186
rect 16582 8134 16634 8186
rect 16646 8134 16698 8186
rect 16710 8134 16762 8186
rect 16774 8134 16826 8186
rect 2504 8032 2556 8084
rect 4252 8032 4304 8084
rect 5080 8032 5132 8084
rect 2780 7964 2832 8016
rect 3608 7964 3660 8016
rect 2228 7939 2280 7948
rect 2228 7905 2237 7939
rect 2237 7905 2271 7939
rect 2271 7905 2280 7939
rect 2228 7896 2280 7905
rect 4620 7964 4672 8016
rect 4344 7939 4396 7948
rect 4344 7905 4353 7939
rect 4353 7905 4387 7939
rect 4387 7905 4396 7939
rect 4344 7896 4396 7905
rect 5172 7939 5224 7948
rect 5172 7905 5181 7939
rect 5181 7905 5215 7939
rect 5215 7905 5224 7939
rect 5172 7896 5224 7905
rect 5264 7939 5316 7948
rect 5264 7905 5273 7939
rect 5273 7905 5307 7939
rect 5307 7905 5316 7939
rect 8484 8032 8536 8084
rect 8944 8075 8996 8084
rect 8944 8041 8953 8075
rect 8953 8041 8987 8075
rect 8987 8041 8996 8075
rect 8944 8032 8996 8041
rect 9128 8032 9180 8084
rect 11980 8032 12032 8084
rect 12440 8032 12492 8084
rect 18420 8075 18472 8084
rect 18420 8041 18429 8075
rect 18429 8041 18463 8075
rect 18463 8041 18472 8075
rect 18420 8032 18472 8041
rect 6184 7964 6236 8016
rect 5264 7896 5316 7905
rect 6552 7939 6604 7948
rect 6552 7905 6561 7939
rect 6561 7905 6595 7939
rect 6595 7905 6604 7939
rect 6552 7896 6604 7905
rect 7196 7964 7248 8016
rect 7748 7896 7800 7948
rect 8116 7896 8168 7948
rect 8668 7896 8720 7948
rect 10508 7896 10560 7948
rect 10876 7896 10928 7948
rect 11428 7896 11480 7948
rect 12348 7939 12400 7948
rect 12348 7905 12357 7939
rect 12357 7905 12391 7939
rect 12391 7905 12400 7939
rect 12348 7896 12400 7905
rect 13452 7964 13504 8016
rect 14832 7964 14884 8016
rect 2320 7828 2372 7880
rect 5816 7828 5868 7880
rect 9496 7828 9548 7880
rect 9772 7828 9824 7880
rect 11244 7828 11296 7880
rect 12624 7828 12676 7880
rect 2412 7760 2464 7812
rect 3700 7760 3752 7812
rect 4436 7760 4488 7812
rect 2320 7692 2372 7744
rect 3516 7692 3568 7744
rect 4160 7735 4212 7744
rect 4160 7701 4169 7735
rect 4169 7701 4203 7735
rect 4203 7701 4212 7735
rect 4160 7692 4212 7701
rect 4896 7692 4948 7744
rect 8392 7803 8444 7812
rect 5172 7692 5224 7744
rect 5816 7735 5868 7744
rect 5816 7701 5825 7735
rect 5825 7701 5859 7735
rect 5859 7701 5868 7735
rect 5816 7692 5868 7701
rect 6184 7692 6236 7744
rect 6276 7735 6328 7744
rect 6276 7701 6285 7735
rect 6285 7701 6319 7735
rect 6319 7701 6328 7735
rect 8392 7769 8401 7803
rect 8401 7769 8435 7803
rect 8435 7769 8444 7803
rect 8392 7760 8444 7769
rect 8484 7760 8536 7812
rect 8852 7760 8904 7812
rect 9680 7760 9732 7812
rect 10600 7803 10652 7812
rect 10600 7769 10609 7803
rect 10609 7769 10643 7803
rect 10643 7769 10652 7803
rect 10600 7760 10652 7769
rect 11612 7760 11664 7812
rect 6276 7692 6328 7701
rect 7472 7692 7524 7744
rect 8116 7692 8168 7744
rect 8300 7735 8352 7744
rect 8300 7701 8309 7735
rect 8309 7701 8343 7735
rect 8343 7701 8352 7735
rect 8300 7692 8352 7701
rect 8760 7735 8812 7744
rect 8760 7701 8769 7735
rect 8769 7701 8803 7735
rect 8803 7701 8812 7735
rect 8760 7692 8812 7701
rect 10968 7692 11020 7744
rect 11152 7735 11204 7744
rect 11152 7701 11161 7735
rect 11161 7701 11195 7735
rect 11195 7701 11204 7735
rect 11152 7692 11204 7701
rect 11336 7692 11388 7744
rect 11520 7692 11572 7744
rect 12072 7735 12124 7744
rect 12072 7701 12081 7735
rect 12081 7701 12115 7735
rect 12115 7701 12124 7735
rect 12072 7692 12124 7701
rect 12348 7760 12400 7812
rect 12532 7760 12584 7812
rect 13268 7896 13320 7948
rect 13544 7896 13596 7948
rect 15108 7896 15160 7948
rect 16396 7939 16448 7948
rect 16396 7905 16405 7939
rect 16405 7905 16439 7939
rect 16439 7905 16448 7939
rect 16396 7896 16448 7905
rect 17408 7896 17460 7948
rect 17500 7896 17552 7948
rect 18236 7964 18288 8016
rect 18144 7896 18196 7948
rect 18512 7896 18564 7948
rect 13636 7828 13688 7880
rect 16856 7828 16908 7880
rect 18236 7871 18288 7880
rect 18236 7837 18245 7871
rect 18245 7837 18279 7871
rect 18279 7837 18288 7871
rect 18236 7828 18288 7837
rect 15384 7760 15436 7812
rect 15844 7760 15896 7812
rect 16488 7760 16540 7812
rect 13084 7692 13136 7744
rect 13820 7692 13872 7744
rect 14740 7692 14792 7744
rect 15936 7692 15988 7744
rect 17132 7760 17184 7812
rect 17224 7735 17276 7744
rect 17224 7701 17233 7735
rect 17233 7701 17267 7735
rect 17267 7701 17276 7735
rect 17224 7692 17276 7701
rect 17316 7735 17368 7744
rect 17316 7701 17325 7735
rect 17325 7701 17359 7735
rect 17359 7701 17368 7735
rect 17316 7692 17368 7701
rect 18972 7692 19024 7744
rect 5398 7590 5450 7642
rect 5462 7590 5514 7642
rect 5526 7590 5578 7642
rect 5590 7590 5642 7642
rect 5654 7590 5706 7642
rect 9846 7590 9898 7642
rect 9910 7590 9962 7642
rect 9974 7590 10026 7642
rect 10038 7590 10090 7642
rect 10102 7590 10154 7642
rect 14294 7590 14346 7642
rect 14358 7590 14410 7642
rect 14422 7590 14474 7642
rect 14486 7590 14538 7642
rect 14550 7590 14602 7642
rect 1400 7531 1452 7540
rect 1400 7497 1409 7531
rect 1409 7497 1443 7531
rect 1443 7497 1452 7531
rect 1400 7488 1452 7497
rect 2320 7531 2372 7540
rect 2320 7497 2329 7531
rect 2329 7497 2363 7531
rect 2363 7497 2372 7531
rect 2320 7488 2372 7497
rect 2964 7488 3016 7540
rect 3424 7531 3476 7540
rect 3424 7497 3433 7531
rect 3433 7497 3467 7531
rect 3467 7497 3476 7531
rect 3424 7488 3476 7497
rect 3792 7488 3844 7540
rect 4436 7488 4488 7540
rect 4896 7531 4948 7540
rect 4896 7497 4905 7531
rect 4905 7497 4939 7531
rect 4939 7497 4948 7531
rect 4896 7488 4948 7497
rect 4988 7531 5040 7540
rect 4988 7497 4997 7531
rect 4997 7497 5031 7531
rect 5031 7497 5040 7531
rect 4988 7488 5040 7497
rect 5816 7488 5868 7540
rect 6184 7531 6236 7540
rect 6184 7497 6193 7531
rect 6193 7497 6227 7531
rect 6227 7497 6236 7531
rect 6184 7488 6236 7497
rect 1492 7420 1544 7472
rect 1952 7395 2004 7404
rect 1952 7361 1961 7395
rect 1961 7361 1995 7395
rect 1995 7361 2004 7395
rect 1952 7352 2004 7361
rect 1676 7327 1728 7336
rect 1676 7293 1685 7327
rect 1685 7293 1719 7327
rect 1719 7293 1728 7327
rect 1676 7284 1728 7293
rect 1860 7327 1912 7336
rect 1860 7293 1869 7327
rect 1869 7293 1903 7327
rect 1903 7293 1912 7327
rect 1860 7284 1912 7293
rect 2964 7327 3016 7336
rect 2964 7293 2973 7327
rect 2973 7293 3007 7327
rect 3007 7293 3016 7327
rect 2964 7284 3016 7293
rect 3792 7352 3844 7404
rect 4252 7420 4304 7472
rect 4344 7420 4396 7472
rect 7288 7488 7340 7540
rect 7932 7488 7984 7540
rect 8116 7531 8168 7540
rect 8116 7497 8125 7531
rect 8125 7497 8159 7531
rect 8159 7497 8168 7531
rect 8116 7488 8168 7497
rect 8300 7488 8352 7540
rect 9036 7488 9088 7540
rect 9404 7488 9456 7540
rect 6920 7420 6972 7472
rect 5080 7352 5132 7404
rect 6828 7352 6880 7404
rect 4620 7284 4672 7336
rect 5632 7327 5684 7336
rect 5632 7293 5641 7327
rect 5641 7293 5675 7327
rect 5675 7293 5684 7327
rect 5632 7284 5684 7293
rect 6644 7327 6696 7336
rect 3976 7216 4028 7268
rect 6644 7293 6653 7327
rect 6653 7293 6687 7327
rect 6687 7293 6696 7327
rect 6644 7284 6696 7293
rect 6920 7327 6972 7336
rect 6920 7293 6929 7327
rect 6929 7293 6963 7327
rect 6963 7293 6972 7327
rect 6920 7284 6972 7293
rect 9312 7463 9364 7472
rect 9312 7429 9321 7463
rect 9321 7429 9355 7463
rect 9355 7429 9364 7463
rect 9312 7420 9364 7429
rect 8484 7395 8536 7404
rect 8484 7361 8493 7395
rect 8493 7361 8527 7395
rect 8527 7361 8536 7395
rect 8484 7352 8536 7361
rect 8852 7352 8904 7404
rect 10692 7488 10744 7540
rect 10968 7531 11020 7540
rect 10968 7497 10977 7531
rect 10977 7497 11011 7531
rect 11011 7497 11020 7531
rect 10968 7488 11020 7497
rect 13084 7531 13136 7540
rect 13084 7497 13093 7531
rect 13093 7497 13127 7531
rect 13127 7497 13136 7531
rect 13084 7488 13136 7497
rect 14740 7531 14792 7540
rect 14740 7497 14749 7531
rect 14749 7497 14783 7531
rect 14783 7497 14792 7531
rect 14740 7488 14792 7497
rect 14832 7488 14884 7540
rect 15752 7488 15804 7540
rect 15936 7488 15988 7540
rect 16396 7531 16448 7540
rect 16396 7497 16405 7531
rect 16405 7497 16439 7531
rect 16439 7497 16448 7531
rect 16396 7488 16448 7497
rect 9864 7352 9916 7404
rect 1676 7148 1728 7200
rect 2044 7148 2096 7200
rect 2780 7148 2832 7200
rect 4436 7148 4488 7200
rect 7012 7216 7064 7268
rect 7380 7284 7432 7336
rect 8300 7284 8352 7336
rect 8668 7284 8720 7336
rect 9404 7327 9456 7336
rect 7748 7216 7800 7268
rect 8484 7216 8536 7268
rect 9404 7293 9413 7327
rect 9413 7293 9447 7327
rect 9447 7293 9456 7327
rect 9404 7284 9456 7293
rect 10232 7420 10284 7472
rect 11152 7420 11204 7472
rect 12992 7463 13044 7472
rect 12992 7429 13001 7463
rect 13001 7429 13035 7463
rect 13035 7429 13044 7463
rect 12992 7420 13044 7429
rect 13268 7420 13320 7472
rect 14188 7420 14240 7472
rect 14556 7420 14608 7472
rect 17316 7488 17368 7540
rect 17868 7488 17920 7540
rect 18328 7531 18380 7540
rect 18328 7497 18337 7531
rect 18337 7497 18371 7531
rect 18371 7497 18380 7531
rect 18328 7488 18380 7497
rect 17592 7420 17644 7472
rect 10600 7352 10652 7404
rect 11704 7352 11756 7404
rect 10232 7327 10284 7336
rect 10232 7293 10241 7327
rect 10241 7293 10275 7327
rect 10275 7293 10284 7327
rect 10232 7284 10284 7293
rect 10324 7327 10376 7336
rect 10324 7293 10333 7327
rect 10333 7293 10367 7327
rect 10367 7293 10376 7327
rect 10324 7284 10376 7293
rect 10508 7284 10560 7336
rect 11428 7284 11480 7336
rect 11612 7284 11664 7336
rect 15292 7352 15344 7404
rect 16212 7395 16264 7404
rect 12440 7284 12492 7336
rect 12808 7284 12860 7336
rect 13176 7284 13228 7336
rect 13544 7284 13596 7336
rect 10600 7216 10652 7268
rect 11336 7216 11388 7268
rect 14188 7284 14240 7336
rect 15384 7284 15436 7336
rect 15752 7327 15804 7336
rect 15752 7293 15761 7327
rect 15761 7293 15795 7327
rect 15795 7293 15804 7327
rect 16212 7361 16221 7395
rect 16221 7361 16255 7395
rect 16255 7361 16264 7395
rect 16212 7352 16264 7361
rect 17408 7352 17460 7404
rect 17868 7395 17920 7404
rect 17868 7361 17877 7395
rect 17877 7361 17911 7395
rect 17911 7361 17920 7395
rect 17868 7352 17920 7361
rect 15752 7284 15804 7293
rect 17132 7284 17184 7336
rect 18144 7327 18196 7336
rect 5080 7148 5132 7200
rect 11704 7148 11756 7200
rect 12992 7148 13044 7200
rect 13544 7191 13596 7200
rect 13544 7157 13553 7191
rect 13553 7157 13587 7191
rect 13587 7157 13596 7191
rect 13544 7148 13596 7157
rect 13636 7148 13688 7200
rect 15200 7191 15252 7200
rect 15200 7157 15209 7191
rect 15209 7157 15243 7191
rect 15243 7157 15252 7191
rect 15200 7148 15252 7157
rect 15752 7148 15804 7200
rect 18144 7293 18153 7327
rect 18153 7293 18187 7327
rect 18187 7293 18196 7327
rect 18144 7284 18196 7293
rect 3174 7046 3226 7098
rect 3238 7046 3290 7098
rect 3302 7046 3354 7098
rect 3366 7046 3418 7098
rect 3430 7046 3482 7098
rect 7622 7046 7674 7098
rect 7686 7046 7738 7098
rect 7750 7046 7802 7098
rect 7814 7046 7866 7098
rect 7878 7046 7930 7098
rect 12070 7046 12122 7098
rect 12134 7046 12186 7098
rect 12198 7046 12250 7098
rect 12262 7046 12314 7098
rect 12326 7046 12378 7098
rect 16518 7046 16570 7098
rect 16582 7046 16634 7098
rect 16646 7046 16698 7098
rect 16710 7046 16762 7098
rect 16774 7046 16826 7098
rect 3332 6944 3384 6996
rect 3700 6944 3752 6996
rect 4252 6944 4304 6996
rect 4988 6944 5040 6996
rect 5816 6944 5868 6996
rect 6460 6944 6512 6996
rect 7472 6944 7524 6996
rect 9496 6987 9548 6996
rect 9496 6953 9505 6987
rect 9505 6953 9539 6987
rect 9539 6953 9548 6987
rect 9496 6944 9548 6953
rect 11428 6987 11480 6996
rect 11428 6953 11437 6987
rect 11437 6953 11471 6987
rect 11471 6953 11480 6987
rect 11428 6944 11480 6953
rect 11520 6944 11572 6996
rect 11704 6944 11756 6996
rect 12992 6944 13044 6996
rect 15936 6944 15988 6996
rect 16856 6944 16908 6996
rect 17132 6944 17184 6996
rect 3332 6808 3384 6860
rect 4160 6808 4212 6860
rect 5264 6876 5316 6928
rect 4804 6808 4856 6860
rect 4988 6808 5040 6860
rect 5448 6808 5500 6860
rect 7380 6876 7432 6928
rect 5724 6808 5776 6860
rect 7748 6851 7800 6860
rect 2136 6740 2188 6792
rect 2412 6783 2464 6792
rect 2412 6749 2421 6783
rect 2421 6749 2455 6783
rect 2455 6749 2464 6783
rect 2412 6740 2464 6749
rect 3976 6783 4028 6792
rect 1492 6647 1544 6656
rect 1492 6613 1501 6647
rect 1501 6613 1535 6647
rect 1535 6613 1544 6647
rect 1492 6604 1544 6613
rect 1768 6647 1820 6656
rect 1768 6613 1777 6647
rect 1777 6613 1811 6647
rect 1811 6613 1820 6647
rect 1768 6604 1820 6613
rect 2320 6647 2372 6656
rect 2320 6613 2329 6647
rect 2329 6613 2363 6647
rect 2363 6613 2372 6647
rect 2320 6604 2372 6613
rect 2596 6604 2648 6656
rect 3424 6672 3476 6724
rect 3700 6604 3752 6656
rect 3976 6749 3985 6783
rect 3985 6749 4019 6783
rect 4019 6749 4028 6783
rect 3976 6740 4028 6749
rect 4068 6740 4120 6792
rect 4436 6783 4488 6792
rect 4436 6749 4445 6783
rect 4445 6749 4479 6783
rect 4479 6749 4488 6783
rect 4436 6740 4488 6749
rect 6736 6783 6788 6792
rect 6736 6749 6745 6783
rect 6745 6749 6779 6783
rect 6779 6749 6788 6783
rect 6736 6740 6788 6749
rect 6920 6740 6972 6792
rect 7748 6817 7757 6851
rect 7757 6817 7791 6851
rect 7791 6817 7800 6851
rect 7748 6808 7800 6817
rect 8668 6876 8720 6928
rect 8760 6808 8812 6860
rect 10140 6851 10192 6860
rect 10140 6817 10149 6851
rect 10149 6817 10183 6851
rect 10183 6817 10192 6851
rect 10140 6808 10192 6817
rect 10876 6851 10928 6860
rect 10876 6817 10885 6851
rect 10885 6817 10919 6851
rect 10919 6817 10928 6851
rect 10876 6808 10928 6817
rect 7840 6740 7892 6792
rect 8300 6783 8352 6792
rect 8300 6749 8309 6783
rect 8309 6749 8343 6783
rect 8343 6749 8352 6783
rect 8300 6740 8352 6749
rect 4160 6604 4212 6656
rect 5264 6647 5316 6656
rect 5264 6613 5273 6647
rect 5273 6613 5307 6647
rect 5307 6613 5316 6647
rect 5264 6604 5316 6613
rect 5448 6604 5500 6656
rect 6460 6604 6512 6656
rect 7104 6647 7156 6656
rect 7104 6613 7113 6647
rect 7113 6613 7147 6647
rect 7147 6613 7156 6647
rect 7104 6604 7156 6613
rect 8024 6604 8076 6656
rect 8944 6740 8996 6792
rect 9128 6740 9180 6792
rect 9588 6740 9640 6792
rect 9864 6783 9916 6792
rect 9864 6749 9873 6783
rect 9873 6749 9907 6783
rect 9907 6749 9916 6783
rect 9864 6740 9916 6749
rect 10508 6740 10560 6792
rect 11152 6783 11204 6792
rect 11152 6749 11161 6783
rect 11161 6749 11195 6783
rect 11195 6749 11204 6783
rect 11152 6740 11204 6749
rect 11704 6808 11756 6860
rect 11888 6851 11940 6860
rect 11888 6817 11897 6851
rect 11897 6817 11931 6851
rect 11931 6817 11940 6851
rect 11888 6808 11940 6817
rect 12440 6808 12492 6860
rect 12716 6876 12768 6928
rect 13452 6876 13504 6928
rect 12808 6851 12860 6860
rect 12808 6817 12817 6851
rect 12817 6817 12851 6851
rect 12851 6817 12860 6851
rect 12808 6808 12860 6817
rect 14740 6876 14792 6928
rect 17868 6876 17920 6928
rect 14924 6808 14976 6860
rect 15016 6808 15068 6860
rect 16120 6808 16172 6860
rect 16856 6808 16908 6860
rect 17040 6808 17092 6860
rect 13544 6740 13596 6792
rect 15200 6740 15252 6792
rect 15936 6740 15988 6792
rect 16212 6783 16264 6792
rect 16212 6749 16221 6783
rect 16221 6749 16255 6783
rect 16255 6749 16264 6783
rect 16212 6740 16264 6749
rect 16672 6740 16724 6792
rect 16948 6740 17000 6792
rect 17316 6808 17368 6860
rect 18052 6944 18104 6996
rect 18144 6944 18196 6996
rect 17592 6740 17644 6792
rect 18512 6783 18564 6792
rect 18512 6749 18521 6783
rect 18521 6749 18555 6783
rect 18555 6749 18564 6783
rect 18512 6740 18564 6749
rect 8944 6647 8996 6656
rect 8944 6613 8953 6647
rect 8953 6613 8987 6647
rect 8987 6613 8996 6647
rect 8944 6604 8996 6613
rect 9128 6604 9180 6656
rect 10324 6647 10376 6656
rect 10324 6613 10333 6647
rect 10333 6613 10367 6647
rect 10367 6613 10376 6647
rect 10324 6604 10376 6613
rect 10876 6604 10928 6656
rect 11152 6604 11204 6656
rect 11980 6604 12032 6656
rect 12440 6604 12492 6656
rect 13820 6672 13872 6724
rect 14556 6715 14608 6724
rect 14556 6681 14565 6715
rect 14565 6681 14599 6715
rect 14599 6681 14608 6715
rect 14556 6672 14608 6681
rect 12808 6604 12860 6656
rect 13636 6604 13688 6656
rect 13912 6604 13964 6656
rect 14832 6604 14884 6656
rect 15016 6604 15068 6656
rect 15384 6647 15436 6656
rect 15384 6613 15393 6647
rect 15393 6613 15427 6647
rect 15427 6613 15436 6647
rect 15384 6604 15436 6613
rect 15752 6647 15804 6656
rect 15752 6613 15761 6647
rect 15761 6613 15795 6647
rect 15795 6613 15804 6647
rect 15752 6604 15804 6613
rect 16120 6672 16172 6724
rect 17040 6715 17092 6724
rect 17040 6681 17049 6715
rect 17049 6681 17083 6715
rect 17083 6681 17092 6715
rect 17040 6672 17092 6681
rect 18604 6672 18656 6724
rect 17684 6604 17736 6656
rect 18052 6604 18104 6656
rect 5398 6502 5450 6554
rect 5462 6502 5514 6554
rect 5526 6502 5578 6554
rect 5590 6502 5642 6554
rect 5654 6502 5706 6554
rect 9846 6502 9898 6554
rect 9910 6502 9962 6554
rect 9974 6502 10026 6554
rect 10038 6502 10090 6554
rect 10102 6502 10154 6554
rect 14294 6502 14346 6554
rect 14358 6502 14410 6554
rect 14422 6502 14474 6554
rect 14486 6502 14538 6554
rect 14550 6502 14602 6554
rect 1952 6400 2004 6452
rect 2412 6443 2464 6452
rect 2412 6409 2421 6443
rect 2421 6409 2455 6443
rect 2455 6409 2464 6443
rect 2412 6400 2464 6409
rect 2964 6400 3016 6452
rect 3148 6400 3200 6452
rect 4160 6443 4212 6452
rect 4160 6409 4169 6443
rect 4169 6409 4203 6443
rect 4203 6409 4212 6443
rect 4160 6400 4212 6409
rect 4712 6400 4764 6452
rect 5816 6443 5868 6452
rect 5816 6409 5825 6443
rect 5825 6409 5859 6443
rect 5859 6409 5868 6443
rect 5816 6400 5868 6409
rect 6184 6443 6236 6452
rect 6184 6409 6193 6443
rect 6193 6409 6227 6443
rect 6227 6409 6236 6443
rect 6184 6400 6236 6409
rect 6644 6400 6696 6452
rect 2044 6332 2096 6384
rect 3516 6332 3568 6384
rect 1952 6264 2004 6316
rect 2228 6196 2280 6248
rect 2688 6307 2740 6316
rect 2688 6273 2697 6307
rect 2697 6273 2731 6307
rect 2731 6273 2740 6307
rect 2688 6264 2740 6273
rect 2872 6264 2924 6316
rect 4436 6332 4488 6384
rect 5172 6332 5224 6384
rect 6828 6443 6880 6452
rect 6828 6409 6837 6443
rect 6837 6409 6871 6443
rect 6871 6409 6880 6443
rect 6828 6400 6880 6409
rect 8944 6400 8996 6452
rect 10324 6400 10376 6452
rect 7472 6332 7524 6384
rect 9956 6332 10008 6384
rect 10968 6332 11020 6384
rect 11428 6332 11480 6384
rect 14280 6400 14332 6452
rect 14740 6400 14792 6452
rect 15200 6443 15252 6452
rect 15200 6409 15209 6443
rect 15209 6409 15243 6443
rect 15243 6409 15252 6443
rect 15200 6400 15252 6409
rect 15660 6400 15712 6452
rect 15752 6400 15804 6452
rect 17408 6443 17460 6452
rect 17408 6409 17417 6443
rect 17417 6409 17451 6443
rect 17451 6409 17460 6443
rect 17408 6400 17460 6409
rect 4252 6264 4304 6316
rect 5080 6264 5132 6316
rect 5448 6264 5500 6316
rect 3332 6196 3384 6248
rect 3516 6196 3568 6248
rect 3700 6196 3752 6248
rect 4344 6239 4396 6248
rect 2596 6128 2648 6180
rect 3240 6128 3292 6180
rect 3792 6128 3844 6180
rect 2872 6103 2924 6112
rect 2872 6069 2881 6103
rect 2881 6069 2915 6103
rect 2915 6069 2924 6103
rect 2872 6060 2924 6069
rect 3700 6103 3752 6112
rect 3700 6069 3709 6103
rect 3709 6069 3743 6103
rect 3743 6069 3752 6103
rect 3700 6060 3752 6069
rect 4344 6205 4353 6239
rect 4353 6205 4387 6239
rect 4387 6205 4396 6239
rect 4344 6196 4396 6205
rect 4804 6196 4856 6248
rect 6368 6264 6420 6316
rect 5632 6196 5684 6248
rect 3976 6128 4028 6180
rect 8484 6264 8536 6316
rect 8852 6307 8904 6316
rect 8852 6273 8861 6307
rect 8861 6273 8895 6307
rect 8895 6273 8904 6307
rect 8852 6264 8904 6273
rect 9404 6264 9456 6316
rect 10692 6264 10744 6316
rect 11336 6307 11388 6316
rect 11336 6273 11345 6307
rect 11345 6273 11379 6307
rect 11379 6273 11388 6307
rect 11336 6264 11388 6273
rect 11888 6307 11940 6316
rect 11888 6273 11897 6307
rect 11897 6273 11931 6307
rect 11931 6273 11940 6307
rect 11888 6264 11940 6273
rect 12256 6264 12308 6316
rect 7380 6239 7432 6248
rect 4712 6060 4764 6112
rect 4804 6060 4856 6112
rect 6644 6128 6696 6180
rect 7380 6205 7389 6239
rect 7389 6205 7423 6239
rect 7423 6205 7432 6239
rect 7380 6196 7432 6205
rect 7840 6239 7892 6248
rect 7840 6205 7849 6239
rect 7849 6205 7883 6239
rect 7883 6205 7892 6239
rect 7840 6196 7892 6205
rect 8116 6196 8168 6248
rect 8760 6239 8812 6248
rect 7288 6128 7340 6180
rect 8760 6205 8769 6239
rect 8769 6205 8803 6239
rect 8803 6205 8812 6239
rect 8760 6196 8812 6205
rect 10416 6196 10468 6248
rect 6920 6060 6972 6112
rect 7380 6060 7432 6112
rect 8392 6103 8444 6112
rect 8392 6069 8401 6103
rect 8401 6069 8435 6103
rect 8435 6069 8444 6103
rect 8392 6060 8444 6069
rect 9956 6128 10008 6180
rect 11244 6196 11296 6248
rect 12992 6264 13044 6316
rect 13176 6264 13228 6316
rect 14832 6332 14884 6384
rect 11612 6128 11664 6180
rect 11796 6128 11848 6180
rect 12900 6128 12952 6180
rect 9036 6060 9088 6112
rect 9312 6060 9364 6112
rect 9864 6060 9916 6112
rect 10692 6060 10744 6112
rect 10968 6060 11020 6112
rect 11336 6060 11388 6112
rect 13084 6103 13136 6112
rect 13084 6069 13093 6103
rect 13093 6069 13127 6103
rect 13127 6069 13136 6103
rect 13084 6060 13136 6069
rect 14372 6307 14424 6316
rect 14372 6273 14381 6307
rect 14381 6273 14415 6307
rect 14415 6273 14424 6307
rect 14372 6264 14424 6273
rect 14740 6264 14792 6316
rect 14280 6196 14332 6248
rect 15752 6196 15804 6248
rect 17408 6264 17460 6316
rect 16672 6128 16724 6180
rect 17132 6196 17184 6248
rect 17224 6196 17276 6248
rect 17592 6128 17644 6180
rect 17868 6128 17920 6180
rect 13636 6060 13688 6112
rect 14188 6060 14240 6112
rect 15292 6060 15344 6112
rect 15936 6060 15988 6112
rect 3174 5958 3226 6010
rect 3238 5958 3290 6010
rect 3302 5958 3354 6010
rect 3366 5958 3418 6010
rect 3430 5958 3482 6010
rect 7622 5958 7674 6010
rect 7686 5958 7738 6010
rect 7750 5958 7802 6010
rect 7814 5958 7866 6010
rect 7878 5958 7930 6010
rect 12070 5958 12122 6010
rect 12134 5958 12186 6010
rect 12198 5958 12250 6010
rect 12262 5958 12314 6010
rect 12326 5958 12378 6010
rect 16518 5958 16570 6010
rect 16582 5958 16634 6010
rect 16646 5958 16698 6010
rect 16710 5958 16762 6010
rect 16774 5958 16826 6010
rect 1860 5856 1912 5908
rect 3424 5856 3476 5908
rect 4988 5856 5040 5908
rect 5632 5899 5684 5908
rect 5632 5865 5641 5899
rect 5641 5865 5675 5899
rect 5675 5865 5684 5899
rect 5632 5856 5684 5865
rect 6460 5899 6512 5908
rect 6460 5865 6469 5899
rect 6469 5865 6503 5899
rect 6503 5865 6512 5899
rect 6460 5856 6512 5865
rect 8300 5856 8352 5908
rect 8484 5856 8536 5908
rect 2688 5788 2740 5840
rect 4252 5788 4304 5840
rect 1584 5720 1636 5772
rect 2228 5763 2280 5772
rect 2228 5729 2237 5763
rect 2237 5729 2271 5763
rect 2271 5729 2280 5763
rect 2228 5720 2280 5729
rect 2872 5763 2924 5772
rect 2872 5729 2881 5763
rect 2881 5729 2915 5763
rect 2915 5729 2924 5763
rect 2872 5720 2924 5729
rect 3148 5720 3200 5772
rect 3516 5652 3568 5704
rect 3792 5695 3844 5704
rect 3792 5661 3801 5695
rect 3801 5661 3835 5695
rect 3835 5661 3844 5695
rect 3792 5652 3844 5661
rect 4252 5695 4304 5704
rect 4896 5720 4948 5772
rect 5724 5720 5776 5772
rect 6000 5720 6052 5772
rect 6184 5720 6236 5772
rect 4252 5661 4269 5695
rect 4269 5661 4303 5695
rect 4303 5661 4304 5695
rect 4252 5652 4304 5661
rect 5356 5652 5408 5704
rect 6460 5652 6512 5704
rect 8024 5788 8076 5840
rect 9680 5788 9732 5840
rect 11888 5856 11940 5908
rect 12992 5856 13044 5908
rect 13452 5856 13504 5908
rect 8208 5720 8260 5772
rect 9036 5720 9088 5772
rect 9220 5763 9272 5772
rect 9220 5729 9229 5763
rect 9229 5729 9263 5763
rect 9263 5729 9272 5763
rect 9220 5720 9272 5729
rect 9312 5720 9364 5772
rect 12072 5788 12124 5840
rect 12532 5788 12584 5840
rect 7840 5652 7892 5704
rect 8484 5695 8536 5704
rect 8484 5661 8493 5695
rect 8493 5661 8527 5695
rect 8527 5661 8536 5695
rect 8484 5652 8536 5661
rect 8576 5652 8628 5704
rect 8944 5695 8996 5704
rect 8944 5661 8953 5695
rect 8953 5661 8987 5695
rect 8987 5661 8996 5695
rect 8944 5652 8996 5661
rect 9772 5652 9824 5704
rect 11428 5720 11480 5772
rect 11980 5720 12032 5772
rect 10600 5652 10652 5704
rect 10784 5652 10836 5704
rect 12256 5695 12308 5704
rect 12256 5661 12265 5695
rect 12265 5661 12299 5695
rect 12299 5661 12308 5695
rect 12256 5652 12308 5661
rect 12440 5763 12492 5772
rect 12440 5729 12449 5763
rect 12449 5729 12483 5763
rect 12483 5729 12492 5763
rect 12440 5720 12492 5729
rect 12900 5720 12952 5772
rect 13084 5763 13136 5772
rect 13084 5729 13093 5763
rect 13093 5729 13127 5763
rect 13127 5729 13136 5763
rect 13084 5720 13136 5729
rect 13268 5788 13320 5840
rect 13912 5856 13964 5908
rect 15752 5899 15804 5908
rect 15752 5865 15761 5899
rect 15761 5865 15795 5899
rect 15795 5865 15804 5899
rect 15752 5856 15804 5865
rect 16856 5856 16908 5908
rect 17868 5856 17920 5908
rect 18236 5856 18288 5908
rect 13544 5720 13596 5772
rect 13268 5652 13320 5704
rect 13728 5652 13780 5704
rect 2044 5559 2096 5568
rect 2044 5525 2053 5559
rect 2053 5525 2087 5559
rect 2087 5525 2096 5559
rect 2044 5516 2096 5525
rect 4068 5584 4120 5636
rect 5724 5584 5776 5636
rect 6828 5627 6880 5636
rect 6828 5593 6837 5627
rect 6837 5593 6871 5627
rect 6871 5593 6880 5627
rect 6828 5584 6880 5593
rect 8300 5584 8352 5636
rect 10416 5584 10468 5636
rect 3884 5516 3936 5568
rect 4344 5559 4396 5568
rect 4344 5525 4353 5559
rect 4353 5525 4387 5559
rect 4387 5525 4396 5559
rect 4344 5516 4396 5525
rect 5172 5559 5224 5568
rect 5172 5525 5181 5559
rect 5181 5525 5215 5559
rect 5215 5525 5224 5559
rect 5172 5516 5224 5525
rect 5264 5559 5316 5568
rect 5264 5525 5273 5559
rect 5273 5525 5307 5559
rect 5307 5525 5316 5559
rect 5264 5516 5316 5525
rect 5816 5516 5868 5568
rect 6184 5516 6236 5568
rect 7472 5516 7524 5568
rect 8024 5559 8076 5568
rect 8024 5525 8033 5559
rect 8033 5525 8067 5559
rect 8067 5525 8076 5559
rect 8024 5516 8076 5525
rect 9036 5516 9088 5568
rect 9404 5559 9456 5568
rect 9404 5525 9413 5559
rect 9413 5525 9447 5559
rect 9447 5525 9456 5559
rect 9404 5516 9456 5525
rect 9772 5516 9824 5568
rect 10784 5516 10836 5568
rect 12900 5584 12952 5636
rect 15384 5788 15436 5840
rect 15108 5720 15160 5772
rect 15936 5720 15988 5772
rect 16396 5720 16448 5772
rect 16856 5720 16908 5772
rect 16212 5695 16264 5704
rect 16212 5661 16221 5695
rect 16221 5661 16255 5695
rect 16255 5661 16264 5695
rect 16212 5652 16264 5661
rect 17592 5788 17644 5840
rect 17868 5720 17920 5772
rect 15200 5584 15252 5636
rect 17040 5652 17092 5704
rect 17500 5652 17552 5704
rect 16764 5584 16816 5636
rect 17224 5584 17276 5636
rect 13912 5516 13964 5568
rect 14924 5516 14976 5568
rect 16580 5516 16632 5568
rect 17040 5559 17092 5568
rect 17040 5525 17049 5559
rect 17049 5525 17083 5559
rect 17083 5525 17092 5559
rect 17040 5516 17092 5525
rect 17684 5584 17736 5636
rect 5398 5414 5450 5466
rect 5462 5414 5514 5466
rect 5526 5414 5578 5466
rect 5590 5414 5642 5466
rect 5654 5414 5706 5466
rect 9846 5414 9898 5466
rect 9910 5414 9962 5466
rect 9974 5414 10026 5466
rect 10038 5414 10090 5466
rect 10102 5414 10154 5466
rect 14294 5414 14346 5466
rect 14358 5414 14410 5466
rect 14422 5414 14474 5466
rect 14486 5414 14538 5466
rect 14550 5414 14602 5466
rect 1492 5355 1544 5364
rect 1492 5321 1501 5355
rect 1501 5321 1535 5355
rect 1535 5321 1544 5355
rect 1492 5312 1544 5321
rect 2044 5312 2096 5364
rect 2320 5355 2372 5364
rect 2320 5321 2329 5355
rect 2329 5321 2363 5355
rect 2363 5321 2372 5355
rect 2320 5312 2372 5321
rect 2780 5355 2832 5364
rect 2780 5321 2789 5355
rect 2789 5321 2823 5355
rect 2823 5321 2832 5355
rect 2780 5312 2832 5321
rect 2504 5244 2556 5296
rect 2596 5244 2648 5296
rect 4252 5312 4304 5364
rect 5080 5312 5132 5364
rect 5264 5312 5316 5364
rect 5908 5355 5960 5364
rect 5908 5321 5917 5355
rect 5917 5321 5951 5355
rect 5951 5321 5960 5355
rect 5908 5312 5960 5321
rect 6460 5312 6512 5364
rect 7012 5312 7064 5364
rect 7288 5312 7340 5364
rect 7840 5355 7892 5364
rect 7840 5321 7849 5355
rect 7849 5321 7883 5355
rect 7883 5321 7892 5355
rect 7840 5312 7892 5321
rect 8024 5312 8076 5364
rect 8852 5312 8904 5364
rect 9772 5312 9824 5364
rect 10784 5355 10836 5364
rect 10784 5321 10793 5355
rect 10793 5321 10827 5355
rect 10827 5321 10836 5355
rect 10784 5312 10836 5321
rect 13544 5355 13596 5364
rect 13544 5321 13553 5355
rect 13553 5321 13587 5355
rect 13587 5321 13596 5355
rect 13544 5312 13596 5321
rect 13912 5312 13964 5364
rect 15108 5312 15160 5364
rect 15936 5312 15988 5364
rect 16120 5312 16172 5364
rect 16212 5312 16264 5364
rect 17132 5312 17184 5364
rect 18696 5312 18748 5364
rect 4896 5287 4948 5296
rect 4896 5253 4905 5287
rect 4905 5253 4939 5287
rect 4939 5253 4948 5287
rect 4896 5244 4948 5253
rect 4988 5244 5040 5296
rect 5632 5244 5684 5296
rect 3240 5219 3292 5228
rect 3240 5185 3249 5219
rect 3249 5185 3283 5219
rect 3283 5185 3292 5219
rect 3516 5219 3568 5228
rect 3240 5176 3292 5185
rect 3516 5185 3525 5219
rect 3525 5185 3559 5219
rect 3559 5185 3568 5219
rect 3516 5176 3568 5185
rect 2596 5108 2648 5160
rect 3424 5040 3476 5092
rect 2596 4972 2648 5024
rect 2964 4972 3016 5024
rect 3516 4972 3568 5024
rect 4712 4972 4764 5024
rect 5908 5176 5960 5228
rect 6920 5244 6972 5296
rect 8024 5176 8076 5228
rect 8392 5244 8444 5296
rect 9680 5244 9732 5296
rect 9036 5176 9088 5228
rect 12992 5244 13044 5296
rect 6000 5151 6052 5160
rect 6000 5117 6009 5151
rect 6009 5117 6043 5151
rect 6043 5117 6052 5151
rect 6000 5108 6052 5117
rect 6920 5108 6972 5160
rect 7104 5151 7156 5160
rect 7104 5117 7113 5151
rect 7113 5117 7147 5151
rect 7147 5117 7156 5151
rect 7104 5108 7156 5117
rect 8116 5108 8168 5160
rect 8208 5108 8260 5160
rect 6736 5040 6788 5092
rect 9220 5151 9272 5160
rect 9220 5117 9229 5151
rect 9229 5117 9263 5151
rect 9263 5117 9272 5151
rect 9220 5108 9272 5117
rect 10140 5151 10192 5160
rect 7104 4972 7156 5024
rect 10140 5117 10149 5151
rect 10149 5117 10183 5151
rect 10183 5117 10192 5151
rect 10140 5108 10192 5117
rect 11980 5151 12032 5160
rect 10508 5040 10560 5092
rect 11980 5117 11989 5151
rect 11989 5117 12023 5151
rect 12023 5117 12032 5151
rect 11980 5108 12032 5117
rect 12532 5176 12584 5228
rect 12348 5108 12400 5160
rect 12532 5040 12584 5092
rect 8300 4972 8352 5024
rect 9588 5015 9640 5024
rect 9588 4981 9597 5015
rect 9597 4981 9631 5015
rect 9631 4981 9640 5015
rect 9588 4972 9640 4981
rect 11244 5015 11296 5024
rect 11244 4981 11253 5015
rect 11253 4981 11287 5015
rect 11287 4981 11296 5015
rect 11244 4972 11296 4981
rect 11980 4972 12032 5024
rect 13176 5176 13228 5228
rect 13268 5176 13320 5228
rect 15200 5244 15252 5296
rect 15108 5219 15160 5228
rect 15108 5185 15117 5219
rect 15117 5185 15151 5219
rect 15151 5185 15160 5219
rect 18972 5244 19024 5296
rect 15108 5176 15160 5185
rect 17316 5176 17368 5228
rect 17960 5219 18012 5228
rect 17960 5185 17969 5219
rect 17969 5185 18003 5219
rect 18003 5185 18012 5219
rect 17960 5176 18012 5185
rect 13360 5108 13412 5160
rect 14372 5108 14424 5160
rect 14556 5151 14608 5160
rect 14556 5117 14565 5151
rect 14565 5117 14599 5151
rect 14599 5117 14608 5151
rect 14556 5108 14608 5117
rect 12992 5040 13044 5092
rect 15384 5040 15436 5092
rect 16212 5108 16264 5160
rect 16764 5108 16816 5160
rect 16948 5151 17000 5160
rect 16948 5117 16957 5151
rect 16957 5117 16991 5151
rect 16991 5117 17000 5151
rect 16948 5108 17000 5117
rect 17500 5108 17552 5160
rect 13452 4972 13504 5024
rect 14004 5015 14056 5024
rect 14004 4981 14013 5015
rect 14013 4981 14047 5015
rect 14047 4981 14056 5015
rect 14004 4972 14056 4981
rect 14188 4972 14240 5024
rect 14556 4972 14608 5024
rect 15292 5015 15344 5024
rect 15292 4981 15301 5015
rect 15301 4981 15335 5015
rect 15335 4981 15344 5015
rect 15292 4972 15344 4981
rect 16120 4972 16172 5024
rect 17592 5015 17644 5024
rect 17592 4981 17601 5015
rect 17601 4981 17635 5015
rect 17635 4981 17644 5015
rect 17592 4972 17644 4981
rect 3174 4870 3226 4922
rect 3238 4870 3290 4922
rect 3302 4870 3354 4922
rect 3366 4870 3418 4922
rect 3430 4870 3482 4922
rect 7622 4870 7674 4922
rect 7686 4870 7738 4922
rect 7750 4870 7802 4922
rect 7814 4870 7866 4922
rect 7878 4870 7930 4922
rect 12070 4870 12122 4922
rect 12134 4870 12186 4922
rect 12198 4870 12250 4922
rect 12262 4870 12314 4922
rect 12326 4870 12378 4922
rect 16518 4870 16570 4922
rect 16582 4870 16634 4922
rect 16646 4870 16698 4922
rect 16710 4870 16762 4922
rect 16774 4870 16826 4922
rect 1400 4768 1452 4820
rect 1860 4811 1912 4820
rect 1860 4777 1869 4811
rect 1869 4777 1903 4811
rect 1903 4777 1912 4811
rect 1860 4768 1912 4777
rect 2228 4811 2280 4820
rect 2228 4777 2237 4811
rect 2237 4777 2271 4811
rect 2271 4777 2280 4811
rect 2228 4768 2280 4777
rect 3792 4768 3844 4820
rect 4252 4768 4304 4820
rect 4436 4768 4488 4820
rect 4804 4811 4856 4820
rect 4804 4777 4813 4811
rect 4813 4777 4847 4811
rect 4847 4777 4856 4811
rect 4804 4768 4856 4777
rect 5172 4768 5224 4820
rect 6184 4768 6236 4820
rect 3976 4743 4028 4752
rect 3976 4709 3985 4743
rect 3985 4709 4019 4743
rect 4019 4709 4028 4743
rect 3976 4700 4028 4709
rect 6000 4700 6052 4752
rect 6368 4768 6420 4820
rect 8208 4768 8260 4820
rect 8760 4768 8812 4820
rect 11796 4811 11848 4820
rect 11796 4777 11805 4811
rect 11805 4777 11839 4811
rect 11839 4777 11848 4811
rect 11796 4768 11848 4777
rect 12348 4768 12400 4820
rect 12900 4768 12952 4820
rect 13912 4768 13964 4820
rect 1676 4607 1728 4616
rect 1676 4573 1685 4607
rect 1685 4573 1719 4607
rect 1719 4573 1728 4607
rect 1676 4564 1728 4573
rect 2688 4632 2740 4684
rect 2412 4607 2464 4616
rect 2412 4573 2421 4607
rect 2421 4573 2455 4607
rect 2455 4573 2464 4607
rect 2412 4564 2464 4573
rect 4344 4632 4396 4684
rect 5632 4632 5684 4684
rect 9680 4700 9732 4752
rect 11704 4743 11756 4752
rect 11704 4709 11713 4743
rect 11713 4709 11747 4743
rect 11747 4709 11756 4743
rect 11704 4700 11756 4709
rect 13820 4700 13872 4752
rect 8024 4675 8076 4684
rect 8024 4641 8033 4675
rect 8033 4641 8067 4675
rect 8067 4641 8076 4675
rect 8024 4632 8076 4641
rect 10140 4632 10192 4684
rect 10508 4675 10560 4684
rect 10508 4641 10517 4675
rect 10517 4641 10551 4675
rect 10551 4641 10560 4675
rect 10508 4632 10560 4641
rect 10784 4675 10836 4684
rect 10784 4641 10793 4675
rect 10793 4641 10827 4675
rect 10827 4641 10836 4675
rect 10784 4632 10836 4641
rect 11336 4632 11388 4684
rect 12808 4675 12860 4684
rect 12808 4641 12817 4675
rect 12817 4641 12851 4675
rect 12851 4641 12860 4675
rect 12808 4632 12860 4641
rect 13452 4675 13504 4684
rect 13452 4641 13461 4675
rect 13461 4641 13495 4675
rect 13495 4641 13504 4675
rect 13452 4632 13504 4641
rect 14188 4632 14240 4684
rect 3332 4607 3384 4616
rect 3332 4573 3341 4607
rect 3341 4573 3375 4607
rect 3375 4573 3384 4607
rect 3332 4564 3384 4573
rect 3608 4607 3660 4616
rect 3608 4573 3617 4607
rect 3617 4573 3651 4607
rect 3651 4573 3660 4607
rect 3608 4564 3660 4573
rect 3792 4607 3844 4616
rect 3792 4573 3801 4607
rect 3801 4573 3835 4607
rect 3835 4573 3844 4607
rect 3792 4564 3844 4573
rect 4988 4607 5040 4616
rect 4988 4573 4997 4607
rect 4997 4573 5031 4607
rect 5031 4573 5040 4607
rect 4988 4564 5040 4573
rect 5080 4564 5132 4616
rect 6460 4564 6512 4616
rect 4160 4496 4212 4548
rect 4528 4496 4580 4548
rect 8760 4564 8812 4616
rect 10232 4564 10284 4616
rect 10692 4564 10744 4616
rect 11060 4607 11112 4616
rect 11060 4573 11069 4607
rect 11069 4573 11103 4607
rect 11103 4573 11112 4607
rect 11060 4564 11112 4573
rect 11888 4564 11940 4616
rect 14004 4564 14056 4616
rect 14096 4564 14148 4616
rect 15384 4768 15436 4820
rect 15476 4768 15528 4820
rect 17040 4768 17092 4820
rect 17776 4768 17828 4820
rect 18144 4768 18196 4820
rect 18420 4811 18472 4820
rect 18420 4777 18429 4811
rect 18429 4777 18463 4811
rect 18463 4777 18472 4811
rect 18420 4768 18472 4777
rect 16028 4632 16080 4684
rect 18788 4632 18840 4684
rect 6920 4496 6972 4548
rect 2780 4428 2832 4480
rect 2964 4428 3016 4480
rect 3056 4428 3108 4480
rect 3608 4428 3660 4480
rect 5172 4471 5224 4480
rect 5172 4437 5181 4471
rect 5181 4437 5215 4471
rect 5215 4437 5224 4471
rect 5172 4428 5224 4437
rect 6644 4471 6696 4480
rect 6644 4437 6653 4471
rect 6653 4437 6687 4471
rect 6687 4437 6696 4471
rect 6644 4428 6696 4437
rect 7012 4471 7064 4480
rect 7012 4437 7021 4471
rect 7021 4437 7055 4471
rect 7055 4437 7064 4471
rect 7012 4428 7064 4437
rect 7104 4471 7156 4480
rect 7104 4437 7113 4471
rect 7113 4437 7147 4471
rect 7147 4437 7156 4471
rect 7104 4428 7156 4437
rect 7380 4428 7432 4480
rect 15108 4564 15160 4616
rect 16120 4607 16172 4616
rect 16120 4573 16129 4607
rect 16129 4573 16163 4607
rect 16163 4573 16172 4607
rect 16120 4564 16172 4573
rect 16856 4564 16908 4616
rect 17040 4564 17092 4616
rect 18236 4607 18288 4616
rect 8392 4428 8444 4480
rect 8576 4471 8628 4480
rect 8576 4437 8585 4471
rect 8585 4437 8619 4471
rect 8619 4437 8628 4471
rect 8576 4428 8628 4437
rect 9312 4428 9364 4480
rect 10416 4428 10468 4480
rect 11428 4471 11480 4480
rect 11428 4437 11437 4471
rect 11437 4437 11471 4471
rect 11471 4437 11480 4471
rect 11428 4428 11480 4437
rect 11704 4428 11756 4480
rect 13636 4428 13688 4480
rect 14372 4496 14424 4548
rect 15200 4496 15252 4548
rect 14280 4428 14332 4480
rect 16580 4496 16632 4548
rect 18236 4573 18245 4607
rect 18245 4573 18279 4607
rect 18279 4573 18288 4607
rect 18236 4564 18288 4573
rect 15752 4471 15804 4480
rect 15752 4437 15761 4471
rect 15761 4437 15795 4471
rect 15795 4437 15804 4471
rect 15752 4428 15804 4437
rect 16764 4428 16816 4480
rect 17500 4428 17552 4480
rect 5398 4326 5450 4378
rect 5462 4326 5514 4378
rect 5526 4326 5578 4378
rect 5590 4326 5642 4378
rect 5654 4326 5706 4378
rect 9846 4326 9898 4378
rect 9910 4326 9962 4378
rect 9974 4326 10026 4378
rect 10038 4326 10090 4378
rect 10102 4326 10154 4378
rect 14294 4326 14346 4378
rect 14358 4326 14410 4378
rect 14422 4326 14474 4378
rect 14486 4326 14538 4378
rect 14550 4326 14602 4378
rect 1492 4267 1544 4276
rect 1492 4233 1501 4267
rect 1501 4233 1535 4267
rect 1535 4233 1544 4267
rect 1492 4224 1544 4233
rect 1860 4267 1912 4276
rect 1860 4233 1869 4267
rect 1869 4233 1903 4267
rect 1903 4233 1912 4267
rect 1860 4224 1912 4233
rect 3516 4224 3568 4276
rect 3792 4224 3844 4276
rect 6000 4224 6052 4276
rect 7012 4267 7064 4276
rect 7012 4233 7021 4267
rect 7021 4233 7055 4267
rect 7055 4233 7064 4267
rect 7012 4224 7064 4233
rect 7380 4267 7432 4276
rect 7380 4233 7389 4267
rect 7389 4233 7423 4267
rect 7423 4233 7432 4267
rect 7380 4224 7432 4233
rect 7472 4267 7524 4276
rect 7472 4233 7481 4267
rect 7481 4233 7515 4267
rect 7515 4233 7524 4267
rect 8760 4267 8812 4276
rect 7472 4224 7524 4233
rect 8760 4233 8769 4267
rect 8769 4233 8803 4267
rect 8803 4233 8812 4267
rect 8760 4224 8812 4233
rect 9312 4267 9364 4276
rect 9312 4233 9321 4267
rect 9321 4233 9355 4267
rect 9355 4233 9364 4267
rect 9312 4224 9364 4233
rect 9588 4224 9640 4276
rect 11980 4224 12032 4276
rect 3332 4156 3384 4208
rect 6920 4199 6972 4208
rect 2136 4088 2188 4140
rect 2412 4131 2464 4140
rect 2412 4097 2421 4131
rect 2421 4097 2455 4131
rect 2455 4097 2464 4131
rect 2412 4088 2464 4097
rect 2688 4131 2740 4140
rect 2688 4097 2697 4131
rect 2697 4097 2731 4131
rect 2731 4097 2740 4131
rect 2688 4088 2740 4097
rect 3424 4131 3476 4140
rect 2596 3952 2648 4004
rect 3424 4097 3433 4131
rect 3433 4097 3467 4131
rect 3467 4097 3476 4131
rect 3424 4088 3476 4097
rect 3884 4088 3936 4140
rect 4160 4131 4212 4140
rect 4160 4097 4169 4131
rect 4169 4097 4203 4131
rect 4203 4097 4212 4131
rect 4160 4088 4212 4097
rect 6920 4165 6929 4199
rect 6929 4165 6963 4199
rect 6963 4165 6972 4199
rect 6920 4156 6972 4165
rect 8208 4156 8260 4208
rect 10416 4199 10468 4208
rect 10416 4165 10425 4199
rect 10425 4165 10459 4199
rect 10459 4165 10468 4199
rect 10416 4156 10468 4165
rect 10508 4156 10560 4208
rect 6184 4088 6236 4140
rect 11520 4131 11572 4140
rect 11520 4097 11529 4131
rect 11529 4097 11563 4131
rect 11563 4097 11572 4131
rect 11520 4088 11572 4097
rect 12716 4224 12768 4276
rect 13268 4267 13320 4276
rect 13268 4233 13277 4267
rect 13277 4233 13311 4267
rect 13311 4233 13320 4267
rect 13268 4224 13320 4233
rect 13728 4267 13780 4276
rect 13728 4233 13737 4267
rect 13737 4233 13771 4267
rect 13771 4233 13780 4267
rect 13728 4224 13780 4233
rect 14096 4267 14148 4276
rect 14096 4233 14105 4267
rect 14105 4233 14139 4267
rect 14139 4233 14148 4267
rect 14096 4224 14148 4233
rect 17592 4224 17644 4276
rect 17684 4267 17736 4276
rect 17684 4233 17693 4267
rect 17693 4233 17727 4267
rect 17727 4233 17736 4267
rect 17684 4224 17736 4233
rect 12532 4156 12584 4208
rect 8300 4020 8352 4072
rect 8576 4020 8628 4072
rect 2228 3927 2280 3936
rect 2228 3893 2237 3927
rect 2237 3893 2271 3927
rect 2271 3893 2280 3927
rect 2228 3884 2280 3893
rect 2320 3884 2372 3936
rect 4620 3952 4672 4004
rect 7104 3952 7156 4004
rect 9128 4020 9180 4072
rect 9496 4063 9548 4072
rect 9496 4029 9505 4063
rect 9505 4029 9539 4063
rect 9539 4029 9548 4063
rect 9496 4020 9548 4029
rect 11980 4063 12032 4072
rect 11980 4029 11989 4063
rect 11989 4029 12023 4063
rect 12023 4029 12032 4063
rect 11980 4020 12032 4029
rect 12900 4131 12952 4140
rect 12900 4097 12909 4131
rect 12909 4097 12943 4131
rect 12943 4097 12952 4131
rect 12900 4088 12952 4097
rect 12992 4088 13044 4140
rect 13912 4156 13964 4208
rect 14004 4156 14056 4208
rect 14188 4131 14240 4140
rect 14188 4097 14197 4131
rect 14197 4097 14231 4131
rect 14231 4097 14240 4131
rect 14188 4088 14240 4097
rect 14648 4088 14700 4140
rect 15752 4156 15804 4208
rect 17408 4156 17460 4208
rect 16396 4088 16448 4140
rect 16764 4131 16816 4140
rect 16764 4097 16773 4131
rect 16773 4097 16807 4131
rect 16807 4097 16816 4131
rect 16764 4088 16816 4097
rect 17132 4131 17184 4140
rect 17132 4097 17141 4131
rect 17141 4097 17175 4131
rect 17175 4097 17184 4131
rect 17132 4088 17184 4097
rect 18236 4131 18288 4140
rect 7748 3884 7800 3936
rect 8116 3927 8168 3936
rect 8116 3893 8125 3927
rect 8125 3893 8159 3927
rect 8159 3893 8168 3927
rect 8116 3884 8168 3893
rect 8300 3884 8352 3936
rect 9128 3884 9180 3936
rect 9220 3884 9272 3936
rect 10508 3952 10560 4004
rect 12348 3952 12400 4004
rect 12992 3952 13044 4004
rect 13912 3952 13964 4004
rect 10324 3927 10376 3936
rect 10324 3893 10333 3927
rect 10333 3893 10367 3927
rect 10367 3893 10376 3927
rect 10324 3884 10376 3893
rect 11704 3927 11756 3936
rect 11704 3893 11713 3927
rect 11713 3893 11747 3927
rect 11747 3893 11756 3927
rect 11704 3884 11756 3893
rect 12440 3927 12492 3936
rect 12440 3893 12449 3927
rect 12449 3893 12483 3927
rect 12483 3893 12492 3927
rect 12440 3884 12492 3893
rect 12808 3884 12860 3936
rect 16120 4063 16172 4072
rect 16120 4029 16129 4063
rect 16129 4029 16163 4063
rect 16163 4029 16172 4063
rect 16120 4020 16172 4029
rect 16212 4020 16264 4072
rect 16764 3952 16816 4004
rect 16948 3995 17000 4004
rect 16948 3961 16957 3995
rect 16957 3961 16991 3995
rect 16991 3961 17000 3995
rect 16948 3952 17000 3961
rect 17316 3995 17368 4004
rect 17316 3961 17325 3995
rect 17325 3961 17359 3995
rect 17359 3961 17368 3995
rect 17316 3952 17368 3961
rect 14188 3884 14240 3936
rect 14556 3884 14608 3936
rect 14740 3927 14792 3936
rect 14740 3893 14749 3927
rect 14749 3893 14783 3927
rect 14783 3893 14792 3927
rect 14740 3884 14792 3893
rect 14832 3884 14884 3936
rect 15108 3884 15160 3936
rect 15292 3884 15344 3936
rect 15936 3884 15988 3936
rect 16856 3884 16908 3936
rect 18236 4097 18245 4131
rect 18245 4097 18279 4131
rect 18279 4097 18288 4131
rect 18236 4088 18288 4097
rect 18052 3995 18104 4004
rect 18052 3961 18061 3995
rect 18061 3961 18095 3995
rect 18095 3961 18104 3995
rect 18052 3952 18104 3961
rect 18604 3952 18656 4004
rect 3174 3782 3226 3834
rect 3238 3782 3290 3834
rect 3302 3782 3354 3834
rect 3366 3782 3418 3834
rect 3430 3782 3482 3834
rect 7622 3782 7674 3834
rect 7686 3782 7738 3834
rect 7750 3782 7802 3834
rect 7814 3782 7866 3834
rect 7878 3782 7930 3834
rect 12070 3782 12122 3834
rect 12134 3782 12186 3834
rect 12198 3782 12250 3834
rect 12262 3782 12314 3834
rect 12326 3782 12378 3834
rect 16518 3782 16570 3834
rect 16582 3782 16634 3834
rect 16646 3782 16698 3834
rect 16710 3782 16762 3834
rect 16774 3782 16826 3834
rect 1492 3723 1544 3732
rect 1492 3689 1501 3723
rect 1501 3689 1535 3723
rect 1535 3689 1544 3723
rect 1492 3680 1544 3689
rect 2136 3723 2188 3732
rect 2136 3689 2145 3723
rect 2145 3689 2179 3723
rect 2179 3689 2188 3723
rect 2136 3680 2188 3689
rect 2412 3680 2464 3732
rect 2872 3680 2924 3732
rect 3516 3723 3568 3732
rect 3516 3689 3525 3723
rect 3525 3689 3559 3723
rect 3559 3689 3568 3723
rect 3516 3680 3568 3689
rect 2320 3612 2372 3664
rect 2504 3612 2556 3664
rect 1768 3519 1820 3528
rect 1768 3485 1777 3519
rect 1777 3485 1811 3519
rect 1811 3485 1820 3519
rect 2320 3519 2372 3528
rect 1768 3476 1820 3485
rect 2320 3485 2329 3519
rect 2329 3485 2363 3519
rect 2363 3485 2372 3519
rect 2320 3476 2372 3485
rect 2780 3476 2832 3528
rect 8116 3680 8168 3732
rect 10784 3723 10836 3732
rect 10784 3689 10793 3723
rect 10793 3689 10827 3723
rect 10827 3689 10836 3723
rect 10784 3680 10836 3689
rect 10876 3680 10928 3732
rect 8944 3612 8996 3664
rect 13084 3612 13136 3664
rect 13728 3655 13780 3664
rect 13728 3621 13737 3655
rect 13737 3621 13771 3655
rect 13771 3621 13780 3655
rect 13728 3612 13780 3621
rect 13912 3655 13964 3664
rect 13912 3621 13921 3655
rect 13921 3621 13955 3655
rect 13955 3621 13964 3655
rect 13912 3612 13964 3621
rect 14188 3655 14240 3664
rect 14188 3621 14197 3655
rect 14197 3621 14231 3655
rect 14231 3621 14240 3655
rect 14188 3612 14240 3621
rect 14832 3612 14884 3664
rect 7472 3544 7524 3596
rect 4712 3476 4764 3528
rect 3516 3408 3568 3460
rect 6092 3476 6144 3528
rect 7196 3476 7248 3528
rect 12808 3544 12860 3596
rect 12900 3544 12952 3596
rect 13820 3544 13872 3596
rect 16212 3680 16264 3732
rect 16304 3680 16356 3732
rect 17684 3723 17736 3732
rect 17684 3689 17693 3723
rect 17693 3689 17727 3723
rect 17727 3689 17736 3723
rect 17684 3680 17736 3689
rect 17868 3680 17920 3732
rect 18512 3680 18564 3732
rect 17132 3612 17184 3664
rect 17316 3655 17368 3664
rect 17316 3621 17325 3655
rect 17325 3621 17359 3655
rect 17359 3621 17368 3655
rect 17316 3612 17368 3621
rect 8024 3476 8076 3528
rect 10784 3476 10836 3528
rect 14004 3476 14056 3528
rect 15292 3519 15344 3528
rect 1952 3383 2004 3392
rect 1952 3349 1961 3383
rect 1961 3349 1995 3383
rect 1995 3349 2004 3383
rect 1952 3340 2004 3349
rect 2044 3340 2096 3392
rect 2780 3340 2832 3392
rect 3792 3383 3844 3392
rect 3792 3349 3801 3383
rect 3801 3349 3835 3383
rect 3835 3349 3844 3383
rect 3792 3340 3844 3349
rect 6828 3340 6880 3392
rect 7932 3340 7984 3392
rect 8208 3340 8260 3392
rect 11152 3383 11204 3392
rect 11152 3349 11161 3383
rect 11161 3349 11195 3383
rect 11195 3349 11204 3383
rect 11152 3340 11204 3349
rect 12532 3408 12584 3460
rect 13636 3408 13688 3460
rect 13728 3408 13780 3460
rect 15292 3485 15301 3519
rect 15301 3485 15335 3519
rect 15335 3485 15344 3519
rect 15292 3476 15344 3485
rect 15568 3519 15620 3528
rect 15568 3485 15577 3519
rect 15577 3485 15611 3519
rect 15611 3485 15620 3519
rect 15568 3476 15620 3485
rect 16672 3519 16724 3528
rect 16672 3485 16681 3519
rect 16681 3485 16715 3519
rect 16715 3485 16724 3519
rect 16672 3476 16724 3485
rect 16764 3519 16816 3528
rect 16764 3485 16773 3519
rect 16773 3485 16807 3519
rect 16807 3485 16816 3519
rect 16764 3476 16816 3485
rect 17500 3519 17552 3528
rect 17500 3485 17509 3519
rect 17509 3485 17543 3519
rect 17543 3485 17552 3519
rect 17500 3476 17552 3485
rect 17776 3476 17828 3528
rect 18236 3519 18288 3528
rect 18236 3485 18245 3519
rect 18245 3485 18279 3519
rect 18279 3485 18288 3519
rect 18236 3476 18288 3485
rect 13544 3340 13596 3392
rect 14924 3383 14976 3392
rect 14924 3349 14933 3383
rect 14933 3349 14967 3383
rect 14967 3349 14976 3383
rect 14924 3340 14976 3349
rect 16120 3383 16172 3392
rect 16120 3349 16129 3383
rect 16129 3349 16163 3383
rect 16163 3349 16172 3383
rect 16120 3340 16172 3349
rect 16396 3383 16448 3392
rect 16396 3349 16405 3383
rect 16405 3349 16439 3383
rect 16439 3349 16448 3383
rect 16396 3340 16448 3349
rect 16948 3383 17000 3392
rect 16948 3349 16957 3383
rect 16957 3349 16991 3383
rect 16991 3349 17000 3383
rect 16948 3340 17000 3349
rect 5398 3238 5450 3290
rect 5462 3238 5514 3290
rect 5526 3238 5578 3290
rect 5590 3238 5642 3290
rect 5654 3238 5706 3290
rect 9846 3238 9898 3290
rect 9910 3238 9962 3290
rect 9974 3238 10026 3290
rect 10038 3238 10090 3290
rect 10102 3238 10154 3290
rect 14294 3238 14346 3290
rect 14358 3238 14410 3290
rect 14422 3238 14474 3290
rect 14486 3238 14538 3290
rect 14550 3238 14602 3290
rect 1492 3179 1544 3188
rect 1492 3145 1501 3179
rect 1501 3145 1535 3179
rect 1535 3145 1544 3179
rect 1492 3136 1544 3145
rect 3792 3136 3844 3188
rect 3884 3179 3936 3188
rect 3884 3145 3893 3179
rect 3893 3145 3927 3179
rect 3927 3145 3936 3179
rect 3884 3136 3936 3145
rect 6552 3136 6604 3188
rect 10324 3136 10376 3188
rect 12532 3179 12584 3188
rect 2044 3043 2096 3052
rect 2044 3009 2053 3043
rect 2053 3009 2087 3043
rect 2087 3009 2096 3043
rect 2044 3000 2096 3009
rect 2596 3000 2648 3052
rect 4068 3068 4120 3120
rect 6276 3068 6328 3120
rect 1860 2907 1912 2916
rect 1860 2873 1869 2907
rect 1869 2873 1903 2907
rect 1903 2873 1912 2907
rect 1860 2864 1912 2873
rect 3700 3000 3752 3052
rect 6644 3000 6696 3052
rect 7288 3000 7340 3052
rect 3516 2932 3568 2984
rect 5724 2932 5776 2984
rect 11428 3068 11480 3120
rect 12532 3145 12541 3179
rect 12541 3145 12575 3179
rect 12575 3145 12584 3179
rect 12532 3136 12584 3145
rect 12992 3136 13044 3188
rect 13176 3179 13228 3188
rect 13176 3145 13185 3179
rect 13185 3145 13219 3179
rect 13219 3145 13228 3179
rect 13176 3136 13228 3145
rect 15200 3136 15252 3188
rect 16212 3179 16264 3188
rect 16212 3145 16221 3179
rect 16221 3145 16255 3179
rect 16255 3145 16264 3179
rect 16212 3136 16264 3145
rect 16856 3136 16908 3188
rect 17040 3179 17092 3188
rect 17040 3145 17049 3179
rect 17049 3145 17083 3179
rect 17083 3145 17092 3179
rect 17040 3136 17092 3145
rect 18052 3179 18104 3188
rect 18052 3145 18061 3179
rect 18061 3145 18095 3179
rect 18095 3145 18104 3179
rect 18052 3136 18104 3145
rect 18420 3179 18472 3188
rect 18420 3145 18429 3179
rect 18429 3145 18463 3179
rect 18463 3145 18472 3179
rect 18420 3136 18472 3145
rect 11612 3000 11664 3052
rect 12624 3000 12676 3052
rect 13820 3043 13872 3052
rect 13820 3009 13829 3043
rect 13829 3009 13863 3043
rect 13863 3009 13872 3043
rect 13820 3000 13872 3009
rect 14004 3043 14056 3052
rect 14004 3009 14013 3043
rect 14013 3009 14047 3043
rect 14047 3009 14056 3043
rect 14004 3000 14056 3009
rect 14096 3043 14148 3052
rect 14096 3009 14105 3043
rect 14105 3009 14139 3043
rect 14139 3009 14148 3043
rect 14096 3000 14148 3009
rect 15016 3043 15068 3052
rect 14740 2932 14792 2984
rect 15016 3009 15025 3043
rect 15025 3009 15059 3043
rect 15059 3009 15068 3043
rect 15016 3000 15068 3009
rect 15200 3043 15252 3052
rect 15200 3009 15209 3043
rect 15209 3009 15243 3043
rect 15243 3009 15252 3043
rect 15476 3043 15528 3052
rect 15200 3000 15252 3009
rect 15476 3009 15485 3043
rect 15485 3009 15519 3043
rect 15519 3009 15528 3043
rect 15476 3000 15528 3009
rect 15752 3043 15804 3052
rect 15752 3009 15761 3043
rect 15761 3009 15795 3043
rect 15795 3009 15804 3043
rect 15752 3000 15804 3009
rect 16028 3043 16080 3052
rect 16028 3009 16037 3043
rect 16037 3009 16071 3043
rect 16071 3009 16080 3043
rect 16028 3000 16080 3009
rect 16396 3000 16448 3052
rect 17224 3068 17276 3120
rect 17132 3043 17184 3052
rect 17132 3009 17141 3043
rect 17141 3009 17175 3043
rect 17175 3009 17184 3043
rect 17132 3000 17184 3009
rect 15660 2932 15712 2984
rect 17592 3000 17644 3052
rect 17960 3000 18012 3052
rect 7104 2864 7156 2916
rect 8760 2864 8812 2916
rect 13084 2907 13136 2916
rect 2228 2839 2280 2848
rect 2228 2805 2237 2839
rect 2237 2805 2271 2839
rect 2271 2805 2280 2839
rect 2228 2796 2280 2805
rect 2596 2839 2648 2848
rect 2596 2805 2605 2839
rect 2605 2805 2639 2839
rect 2639 2805 2648 2839
rect 2596 2796 2648 2805
rect 2688 2796 2740 2848
rect 3516 2839 3568 2848
rect 3516 2805 3525 2839
rect 3525 2805 3559 2839
rect 3559 2805 3568 2839
rect 3516 2796 3568 2805
rect 4896 2796 4948 2848
rect 7196 2839 7248 2848
rect 7196 2805 7205 2839
rect 7205 2805 7239 2839
rect 7239 2805 7248 2839
rect 7196 2796 7248 2805
rect 11152 2839 11204 2848
rect 11152 2805 11161 2839
rect 11161 2805 11195 2839
rect 11195 2805 11204 2839
rect 11152 2796 11204 2805
rect 11520 2839 11572 2848
rect 11520 2805 11529 2839
rect 11529 2805 11563 2839
rect 11563 2805 11572 2839
rect 11520 2796 11572 2805
rect 11980 2839 12032 2848
rect 11980 2805 11989 2839
rect 11989 2805 12023 2839
rect 12023 2805 12032 2839
rect 11980 2796 12032 2805
rect 13084 2873 13093 2907
rect 13093 2873 13127 2907
rect 13127 2873 13136 2907
rect 13084 2864 13136 2873
rect 13728 2864 13780 2916
rect 15108 2864 15160 2916
rect 15568 2864 15620 2916
rect 16580 2864 16632 2916
rect 14372 2796 14424 2848
rect 15016 2796 15068 2848
rect 15660 2839 15712 2848
rect 15660 2805 15669 2839
rect 15669 2805 15703 2839
rect 15703 2805 15712 2839
rect 15660 2796 15712 2805
rect 17316 2839 17368 2848
rect 17316 2805 17325 2839
rect 17325 2805 17359 2839
rect 17359 2805 17368 2839
rect 17316 2796 17368 2805
rect 17684 2839 17736 2848
rect 17684 2805 17693 2839
rect 17693 2805 17727 2839
rect 17727 2805 17736 2839
rect 17684 2796 17736 2805
rect 3174 2694 3226 2746
rect 3238 2694 3290 2746
rect 3302 2694 3354 2746
rect 3366 2694 3418 2746
rect 3430 2694 3482 2746
rect 7622 2694 7674 2746
rect 7686 2694 7738 2746
rect 7750 2694 7802 2746
rect 7814 2694 7866 2746
rect 7878 2694 7930 2746
rect 12070 2694 12122 2746
rect 12134 2694 12186 2746
rect 12198 2694 12250 2746
rect 12262 2694 12314 2746
rect 12326 2694 12378 2746
rect 16518 2694 16570 2746
rect 16582 2694 16634 2746
rect 16646 2694 16698 2746
rect 16710 2694 16762 2746
rect 16774 2694 16826 2746
rect 1492 2635 1544 2644
rect 1492 2601 1501 2635
rect 1501 2601 1535 2635
rect 1535 2601 1544 2635
rect 1492 2592 1544 2601
rect 2964 2592 3016 2644
rect 11888 2592 11940 2644
rect 11244 2524 11296 2576
rect 13636 2524 13688 2576
rect 14464 2592 14516 2644
rect 15200 2592 15252 2644
rect 15752 2592 15804 2644
rect 18420 2635 18472 2644
rect 3056 2456 3108 2508
rect 2780 2431 2832 2440
rect 2780 2397 2789 2431
rect 2789 2397 2823 2431
rect 2823 2397 2832 2431
rect 2780 2388 2832 2397
rect 3608 2456 3660 2508
rect 8208 2456 8260 2508
rect 2688 2320 2740 2372
rect 3516 2388 3568 2440
rect 4896 2431 4948 2440
rect 4896 2397 4905 2431
rect 4905 2397 4939 2431
rect 4939 2397 4948 2431
rect 4896 2388 4948 2397
rect 5172 2388 5224 2440
rect 7104 2388 7156 2440
rect 7196 2388 7248 2440
rect 8024 2388 8076 2440
rect 8944 2431 8996 2440
rect 8944 2397 8953 2431
rect 8953 2397 8987 2431
rect 8987 2397 8996 2431
rect 8944 2388 8996 2397
rect 11980 2456 12032 2508
rect 15568 2524 15620 2576
rect 11152 2388 11204 2440
rect 11520 2431 11572 2440
rect 11520 2397 11529 2431
rect 11529 2397 11563 2431
rect 11563 2397 11572 2431
rect 11520 2388 11572 2397
rect 11704 2388 11756 2440
rect 12440 2388 12492 2440
rect 13728 2431 13780 2440
rect 13728 2397 13737 2431
rect 13737 2397 13771 2431
rect 13771 2397 13780 2431
rect 13728 2388 13780 2397
rect 14372 2431 14424 2440
rect 14372 2397 14381 2431
rect 14381 2397 14415 2431
rect 14415 2397 14424 2431
rect 14372 2388 14424 2397
rect 15016 2388 15068 2440
rect 1860 2295 1912 2304
rect 1860 2261 1869 2295
rect 1869 2261 1903 2295
rect 1903 2261 1912 2295
rect 1860 2252 1912 2261
rect 2044 2252 2096 2304
rect 2780 2252 2832 2304
rect 2872 2252 2924 2304
rect 3608 2252 3660 2304
rect 3700 2252 3752 2304
rect 4528 2252 4580 2304
rect 5264 2252 5316 2304
rect 6184 2252 6236 2304
rect 7012 2252 7064 2304
rect 7840 2252 7892 2304
rect 8668 2252 8720 2304
rect 9496 2252 9548 2304
rect 10324 2252 10376 2304
rect 11152 2252 11204 2304
rect 11980 2252 12032 2304
rect 12716 2295 12768 2304
rect 12716 2261 12725 2295
rect 12725 2261 12759 2295
rect 12759 2261 12768 2295
rect 12716 2252 12768 2261
rect 12808 2252 12860 2304
rect 13544 2295 13596 2304
rect 13544 2261 13553 2295
rect 13553 2261 13587 2295
rect 13587 2261 13596 2295
rect 13544 2252 13596 2261
rect 15476 2320 15528 2372
rect 13728 2252 13780 2304
rect 14004 2252 14056 2304
rect 14464 2252 14516 2304
rect 14648 2295 14700 2304
rect 14648 2261 14657 2295
rect 14657 2261 14691 2295
rect 14691 2261 14700 2295
rect 14648 2252 14700 2261
rect 15292 2252 15344 2304
rect 17592 2524 17644 2576
rect 16120 2456 16172 2508
rect 17408 2456 17460 2508
rect 18420 2601 18429 2635
rect 18429 2601 18463 2635
rect 18463 2601 18472 2635
rect 18420 2592 18472 2601
rect 16396 2388 16448 2440
rect 17040 2431 17092 2440
rect 17040 2397 17049 2431
rect 17049 2397 17083 2431
rect 17083 2397 17092 2431
rect 17040 2388 17092 2397
rect 18236 2431 18288 2440
rect 18236 2397 18245 2431
rect 18245 2397 18279 2431
rect 18279 2397 18288 2431
rect 18236 2388 18288 2397
rect 16856 2252 16908 2304
rect 17040 2252 17092 2304
rect 18604 2320 18656 2372
rect 17776 2252 17828 2304
rect 5398 2150 5450 2202
rect 5462 2150 5514 2202
rect 5526 2150 5578 2202
rect 5590 2150 5642 2202
rect 5654 2150 5706 2202
rect 9846 2150 9898 2202
rect 9910 2150 9962 2202
rect 9974 2150 10026 2202
rect 10038 2150 10090 2202
rect 10102 2150 10154 2202
rect 14294 2150 14346 2202
rect 14358 2150 14410 2202
rect 14422 2150 14474 2202
rect 14486 2150 14538 2202
rect 14550 2150 14602 2202
rect 1216 2048 1268 2100
rect 2688 2048 2740 2100
rect 15660 2048 15712 2100
rect 18236 2048 18288 2100
rect 12716 1912 12768 1964
rect 16120 1912 16172 1964
rect 16856 1912 16908 1964
rect 17500 1912 17552 1964
rect 13544 1844 13596 1896
rect 16028 1844 16080 1896
<< metal2 >>
rect 2042 16400 2098 17200
rect 5998 16400 6054 17200
rect 9954 16400 10010 17200
rect 13910 16400 13966 17200
rect 17866 16400 17922 17200
rect 1858 14920 1914 14929
rect 1858 14855 1914 14864
rect 1872 14822 1900 14855
rect 1860 14816 1912 14822
rect 1860 14758 1912 14764
rect 1872 13326 1900 14758
rect 2056 14618 2084 16400
rect 2134 15464 2190 15473
rect 2134 15399 2190 15408
rect 2148 15230 2176 15399
rect 2136 15224 2188 15230
rect 4528 15224 4580 15230
rect 2136 15166 2188 15172
rect 3054 15192 3110 15201
rect 2044 14612 2096 14618
rect 2044 14554 2096 14560
rect 1952 14408 2004 14414
rect 1952 14350 2004 14356
rect 1964 14249 1992 14350
rect 1950 14240 2006 14249
rect 1950 14175 2006 14184
rect 1950 13968 2006 13977
rect 2148 13938 2176 15166
rect 4528 15166 4580 15172
rect 3054 15127 3110 15136
rect 2778 14920 2834 14929
rect 2778 14855 2834 14864
rect 2228 14476 2280 14482
rect 2228 14418 2280 14424
rect 2240 14113 2268 14418
rect 2226 14104 2282 14113
rect 2226 14039 2282 14048
rect 2792 13977 2820 14855
rect 2962 14648 3018 14657
rect 2962 14583 3018 14592
rect 2872 14272 2924 14278
rect 2872 14214 2924 14220
rect 2778 13968 2834 13977
rect 1950 13903 1952 13912
rect 2004 13903 2006 13912
rect 2136 13932 2188 13938
rect 1952 13874 2004 13880
rect 2778 13903 2834 13912
rect 2136 13874 2188 13880
rect 2884 13569 2912 14214
rect 2976 13870 3004 14583
rect 3068 14550 3096 15127
rect 3974 15056 4030 15065
rect 3974 14991 4030 15000
rect 3174 14716 3482 14725
rect 3174 14714 3180 14716
rect 3236 14714 3260 14716
rect 3316 14714 3340 14716
rect 3396 14714 3420 14716
rect 3476 14714 3482 14716
rect 3236 14662 3238 14714
rect 3418 14662 3420 14714
rect 3174 14660 3180 14662
rect 3236 14660 3260 14662
rect 3316 14660 3340 14662
rect 3396 14660 3420 14662
rect 3476 14660 3482 14662
rect 3174 14651 3482 14660
rect 3056 14544 3108 14550
rect 3056 14486 3108 14492
rect 3514 14512 3570 14521
rect 3514 14447 3570 14456
rect 3056 14408 3108 14414
rect 3056 14350 3108 14356
rect 3068 13977 3096 14350
rect 3528 14113 3556 14447
rect 3792 14272 3844 14278
rect 3792 14214 3844 14220
rect 3514 14104 3570 14113
rect 3424 14068 3476 14074
rect 3514 14039 3570 14048
rect 3424 14010 3476 14016
rect 3054 13968 3110 13977
rect 3054 13903 3110 13912
rect 2964 13864 3016 13870
rect 2964 13806 3016 13812
rect 3332 13864 3384 13870
rect 3436 13841 3464 14010
rect 3528 13938 3556 14039
rect 3516 13932 3568 13938
rect 3516 13874 3568 13880
rect 3332 13806 3384 13812
rect 3422 13832 3478 13841
rect 3344 13716 3372 13806
rect 3422 13767 3478 13776
rect 3344 13688 3556 13716
rect 3174 13628 3482 13637
rect 3174 13626 3180 13628
rect 3236 13626 3260 13628
rect 3316 13626 3340 13628
rect 3396 13626 3420 13628
rect 3476 13626 3482 13628
rect 3236 13574 3238 13626
rect 3418 13574 3420 13626
rect 3174 13572 3180 13574
rect 3236 13572 3260 13574
rect 3316 13572 3340 13574
rect 3396 13572 3420 13574
rect 3476 13572 3482 13574
rect 2870 13560 2926 13569
rect 3174 13563 3482 13572
rect 2870 13495 2926 13504
rect 3528 13462 3556 13688
rect 2780 13456 2832 13462
rect 1950 13424 2006 13433
rect 2780 13398 2832 13404
rect 3516 13456 3568 13462
rect 3516 13398 3568 13404
rect 1950 13359 1952 13368
rect 2004 13359 2006 13368
rect 1952 13330 2004 13336
rect 1860 13320 1912 13326
rect 1860 13262 1912 13268
rect 2688 13184 2740 13190
rect 2686 13152 2688 13161
rect 2740 13152 2742 13161
rect 2686 13087 2742 13096
rect 2320 12980 2372 12986
rect 2320 12922 2372 12928
rect 1768 12844 1820 12850
rect 1768 12786 1820 12792
rect 1308 12640 1360 12646
rect 1308 12582 1360 12588
rect 1320 4185 1348 12582
rect 1780 12434 1808 12786
rect 2136 12776 2188 12782
rect 2136 12718 2188 12724
rect 1688 12406 1808 12434
rect 1688 12345 1716 12406
rect 1674 12336 1730 12345
rect 1674 12271 1730 12280
rect 1400 10056 1452 10062
rect 1398 10024 1400 10033
rect 1452 10024 1454 10033
rect 1398 9959 1454 9968
rect 1412 7546 1440 9959
rect 1490 7848 1546 7857
rect 1490 7783 1546 7792
rect 1400 7540 1452 7546
rect 1400 7482 1452 7488
rect 1504 7478 1532 7783
rect 1688 7721 1716 12271
rect 1860 12096 1912 12102
rect 1860 12038 1912 12044
rect 1872 7970 1900 12038
rect 2044 11756 2096 11762
rect 2044 11698 2096 11704
rect 1952 11688 2004 11694
rect 1952 11630 2004 11636
rect 1964 10985 1992 11630
rect 2056 11257 2084 11698
rect 2042 11248 2098 11257
rect 2042 11183 2098 11192
rect 1950 10976 2006 10985
rect 1950 10911 2006 10920
rect 1952 10600 2004 10606
rect 1952 10542 2004 10548
rect 1964 10169 1992 10542
rect 1950 10160 2006 10169
rect 1950 10095 2006 10104
rect 1950 9616 2006 9625
rect 1950 9551 2006 9560
rect 1964 9518 1992 9551
rect 1952 9512 2004 9518
rect 1952 9454 2004 9460
rect 1964 9353 1992 9454
rect 1950 9344 2006 9353
rect 1950 9279 2006 9288
rect 1952 8968 2004 8974
rect 1952 8910 2004 8916
rect 1964 8537 1992 8910
rect 1950 8528 2006 8537
rect 2056 8498 2084 11183
rect 2148 9897 2176 12718
rect 2228 11688 2280 11694
rect 2226 11656 2228 11665
rect 2280 11656 2282 11665
rect 2226 11591 2282 11600
rect 2228 11280 2280 11286
rect 2228 11222 2280 11228
rect 2240 11150 2268 11222
rect 2228 11144 2280 11150
rect 2226 11112 2228 11121
rect 2280 11112 2282 11121
rect 2226 11047 2282 11056
rect 2134 9888 2190 9897
rect 2134 9823 2190 9832
rect 2226 9752 2282 9761
rect 2226 9687 2282 9696
rect 2240 9586 2268 9687
rect 2228 9580 2280 9586
rect 2228 9522 2280 9528
rect 2228 8560 2280 8566
rect 2228 8502 2280 8508
rect 1950 8463 2006 8472
rect 2044 8492 2096 8498
rect 2044 8434 2096 8440
rect 2240 8401 2268 8502
rect 2226 8392 2282 8401
rect 2226 8327 2282 8336
rect 1872 7942 2176 7970
rect 2240 7954 2268 8327
rect 2148 7834 2176 7942
rect 2228 7948 2280 7954
rect 2228 7890 2280 7896
rect 2332 7886 2360 12922
rect 2412 12164 2464 12170
rect 2412 12106 2464 12112
rect 2424 11558 2452 12106
rect 2504 11688 2556 11694
rect 2504 11630 2556 11636
rect 2412 11552 2464 11558
rect 2412 11494 2464 11500
rect 2412 10668 2464 10674
rect 2412 10610 2464 10616
rect 2424 10577 2452 10610
rect 2410 10568 2466 10577
rect 2410 10503 2466 10512
rect 2516 10130 2544 11630
rect 2596 11280 2648 11286
rect 2596 11222 2648 11228
rect 2504 10124 2556 10130
rect 2504 10066 2556 10072
rect 2516 9042 2544 10066
rect 2504 9036 2556 9042
rect 2504 8978 2556 8984
rect 2516 8809 2544 8978
rect 2502 8800 2558 8809
rect 2502 8735 2558 8744
rect 2608 8537 2636 11222
rect 2700 10742 2728 13087
rect 2792 12481 2820 13398
rect 3608 13388 3660 13394
rect 3608 13330 3660 13336
rect 3516 13320 3568 13326
rect 3516 13262 3568 13268
rect 2964 13252 3016 13258
rect 2964 13194 3016 13200
rect 2872 12912 2924 12918
rect 2872 12854 2924 12860
rect 2778 12472 2834 12481
rect 2778 12407 2834 12416
rect 2780 12232 2832 12238
rect 2780 12174 2832 12180
rect 2792 12073 2820 12174
rect 2778 12064 2834 12073
rect 2778 11999 2834 12008
rect 2792 11801 2820 11999
rect 2778 11792 2834 11801
rect 2778 11727 2834 11736
rect 2884 11354 2912 12854
rect 2976 11898 3004 13194
rect 3332 13184 3384 13190
rect 3332 13126 3384 13132
rect 3238 12880 3294 12889
rect 3344 12850 3372 13126
rect 3238 12815 3294 12824
rect 3332 12844 3384 12850
rect 3252 12782 3280 12815
rect 3332 12786 3384 12792
rect 3240 12776 3292 12782
rect 3240 12718 3292 12724
rect 3056 12708 3108 12714
rect 3056 12650 3108 12656
rect 3068 11937 3096 12650
rect 3174 12540 3482 12549
rect 3174 12538 3180 12540
rect 3236 12538 3260 12540
rect 3316 12538 3340 12540
rect 3396 12538 3420 12540
rect 3476 12538 3482 12540
rect 3236 12486 3238 12538
rect 3418 12486 3420 12538
rect 3174 12484 3180 12486
rect 3236 12484 3260 12486
rect 3316 12484 3340 12486
rect 3396 12484 3420 12486
rect 3476 12484 3482 12486
rect 3174 12475 3482 12484
rect 3528 12442 3556 13262
rect 3332 12436 3384 12442
rect 3332 12378 3384 12384
rect 3516 12436 3568 12442
rect 3516 12378 3568 12384
rect 3344 12238 3372 12378
rect 3148 12232 3200 12238
rect 3146 12200 3148 12209
rect 3332 12232 3384 12238
rect 3200 12200 3202 12209
rect 3332 12174 3384 12180
rect 3146 12135 3202 12144
rect 3054 11928 3110 11937
rect 2964 11892 3016 11898
rect 3620 11898 3648 13330
rect 3700 12912 3752 12918
rect 3700 12854 3752 12860
rect 3054 11863 3110 11872
rect 3608 11892 3660 11898
rect 2964 11834 3016 11840
rect 3608 11834 3660 11840
rect 3712 11778 3740 12854
rect 2964 11756 3016 11762
rect 2964 11698 3016 11704
rect 3528 11750 3740 11778
rect 2872 11348 2924 11354
rect 2872 11290 2924 11296
rect 2976 11286 3004 11698
rect 3174 11452 3482 11461
rect 3174 11450 3180 11452
rect 3236 11450 3260 11452
rect 3316 11450 3340 11452
rect 3396 11450 3420 11452
rect 3476 11450 3482 11452
rect 3236 11398 3238 11450
rect 3418 11398 3420 11450
rect 3174 11396 3180 11398
rect 3236 11396 3260 11398
rect 3316 11396 3340 11398
rect 3396 11396 3420 11398
rect 3476 11396 3482 11398
rect 3174 11387 3482 11396
rect 2780 11280 2832 11286
rect 2778 11248 2780 11257
rect 2964 11280 3016 11286
rect 2832 11248 2834 11257
rect 2964 11222 3016 11228
rect 2778 11183 2834 11192
rect 3148 11144 3200 11150
rect 3148 11086 3200 11092
rect 2872 11076 2924 11082
rect 2872 11018 2924 11024
rect 2884 10849 2912 11018
rect 3056 11008 3108 11014
rect 3056 10950 3108 10956
rect 2870 10840 2926 10849
rect 2870 10775 2926 10784
rect 2688 10736 2740 10742
rect 2688 10678 2740 10684
rect 2594 8528 2650 8537
rect 2594 8463 2650 8472
rect 2700 8344 2728 10678
rect 2964 10668 3016 10674
rect 2964 10610 3016 10616
rect 2780 10600 2832 10606
rect 2780 10542 2832 10548
rect 2792 10305 2820 10542
rect 2778 10296 2834 10305
rect 2778 10231 2834 10240
rect 2872 10260 2924 10266
rect 2792 10198 2820 10231
rect 2872 10202 2924 10208
rect 2780 10192 2832 10198
rect 2780 10134 2832 10140
rect 2884 10062 2912 10202
rect 2872 10056 2924 10062
rect 2872 9998 2924 10004
rect 2780 9920 2832 9926
rect 2780 9862 2832 9868
rect 2792 9586 2820 9862
rect 2976 9722 3004 10610
rect 2964 9716 3016 9722
rect 2964 9658 3016 9664
rect 2780 9580 2832 9586
rect 2780 9522 2832 9528
rect 2872 9512 2924 9518
rect 2778 9480 2834 9489
rect 2872 9454 2924 9460
rect 2778 9415 2834 9424
rect 2792 9042 2820 9415
rect 2884 9081 2912 9454
rect 2964 9444 3016 9450
rect 2964 9386 3016 9392
rect 2976 9217 3004 9386
rect 2962 9208 3018 9217
rect 2962 9143 3018 9152
rect 2870 9072 2926 9081
rect 2780 9036 2832 9042
rect 2870 9007 2926 9016
rect 2780 8978 2832 8984
rect 2778 8936 2834 8945
rect 2962 8936 3018 8945
rect 2778 8871 2834 8880
rect 2884 8894 2962 8922
rect 2792 8430 2820 8871
rect 2780 8424 2832 8430
rect 2780 8366 2832 8372
rect 2608 8316 2728 8344
rect 2504 8084 2556 8090
rect 2504 8026 2556 8032
rect 2320 7880 2372 7886
rect 2148 7806 2268 7834
rect 2320 7822 2372 7828
rect 1674 7712 1730 7721
rect 1674 7647 1730 7656
rect 1492 7472 1544 7478
rect 1492 7414 1544 7420
rect 1504 6882 1532 7414
rect 1688 7342 1716 7647
rect 1952 7404 2004 7410
rect 1952 7346 2004 7352
rect 1676 7336 1728 7342
rect 1676 7278 1728 7284
rect 1860 7336 1912 7342
rect 1860 7278 1912 7284
rect 1676 7200 1728 7206
rect 1676 7142 1728 7148
rect 1504 6854 1624 6882
rect 1490 6760 1546 6769
rect 1490 6695 1546 6704
rect 1504 6662 1532 6695
rect 1492 6656 1544 6662
rect 1492 6598 1544 6604
rect 1490 6216 1546 6225
rect 1490 6151 1546 6160
rect 1398 5944 1454 5953
rect 1398 5879 1454 5888
rect 1412 4826 1440 5879
rect 1504 5370 1532 6151
rect 1596 5778 1624 6854
rect 1584 5772 1636 5778
rect 1584 5714 1636 5720
rect 1492 5364 1544 5370
rect 1492 5306 1544 5312
rect 1490 5128 1546 5137
rect 1490 5063 1546 5072
rect 1400 4820 1452 4826
rect 1400 4762 1452 4768
rect 1504 4282 1532 5063
rect 1688 4622 1716 7142
rect 1768 6656 1820 6662
rect 1768 6598 1820 6604
rect 1676 4616 1728 4622
rect 1676 4558 1728 4564
rect 1492 4276 1544 4282
rect 1492 4218 1544 4224
rect 1306 4176 1362 4185
rect 1306 4111 1362 4120
rect 1490 4040 1546 4049
rect 1490 3975 1546 3984
rect 1504 3738 1532 3975
rect 1492 3732 1544 3738
rect 1492 3674 1544 3680
rect 1780 3534 1808 6598
rect 1872 5914 1900 7278
rect 1964 6458 1992 7346
rect 2044 7200 2096 7206
rect 2044 7142 2096 7148
rect 1952 6452 2004 6458
rect 1952 6394 2004 6400
rect 2056 6390 2084 7142
rect 2136 6792 2188 6798
rect 2136 6734 2188 6740
rect 2044 6384 2096 6390
rect 2044 6326 2096 6332
rect 1952 6316 2004 6322
rect 1952 6258 2004 6264
rect 1964 6225 1992 6258
rect 1950 6216 2006 6225
rect 1950 6151 2006 6160
rect 1860 5908 1912 5914
rect 1860 5850 1912 5856
rect 2148 5681 2176 6734
rect 2240 6254 2268 7806
rect 2412 7812 2464 7818
rect 2412 7754 2464 7760
rect 2320 7744 2372 7750
rect 2320 7686 2372 7692
rect 2332 7546 2360 7686
rect 2320 7540 2372 7546
rect 2320 7482 2372 7488
rect 2424 6798 2452 7754
rect 2412 6792 2464 6798
rect 2318 6760 2374 6769
rect 2412 6734 2464 6740
rect 2318 6695 2374 6704
rect 2332 6662 2360 6695
rect 2320 6656 2372 6662
rect 2320 6598 2372 6604
rect 2410 6488 2466 6497
rect 2410 6423 2412 6432
rect 2464 6423 2466 6432
rect 2412 6394 2464 6400
rect 2516 6338 2544 8026
rect 2608 6662 2636 8316
rect 2780 8016 2832 8022
rect 2780 7958 2832 7964
rect 2686 7576 2742 7585
rect 2686 7511 2742 7520
rect 2596 6656 2648 6662
rect 2596 6598 2648 6604
rect 2424 6310 2544 6338
rect 2700 6322 2728 7511
rect 2792 7206 2820 7958
rect 2884 7324 2912 8894
rect 2962 8871 3018 8880
rect 2964 8424 3016 8430
rect 2964 8366 3016 8372
rect 2976 8129 3004 8366
rect 2962 8120 3018 8129
rect 2962 8055 3018 8064
rect 2962 7576 3018 7585
rect 2962 7511 2964 7520
rect 3016 7511 3018 7520
rect 2964 7482 3016 7488
rect 2964 7336 3016 7342
rect 2884 7296 2964 7324
rect 3068 7313 3096 10950
rect 3160 10577 3188 11086
rect 3146 10568 3202 10577
rect 3146 10503 3202 10512
rect 3528 10470 3556 11750
rect 3608 11688 3660 11694
rect 3608 11630 3660 11636
rect 3620 11150 3648 11630
rect 3804 11234 3832 14214
rect 3988 14006 4016 14991
rect 4068 14476 4120 14482
rect 4068 14418 4120 14424
rect 4080 14385 4108 14418
rect 4160 14408 4212 14414
rect 4066 14376 4122 14385
rect 4160 14350 4212 14356
rect 4344 14408 4396 14414
rect 4344 14350 4396 14356
rect 4066 14311 4122 14320
rect 3976 14000 4028 14006
rect 3976 13942 4028 13948
rect 4068 13456 4120 13462
rect 4068 13398 4120 13404
rect 3974 13288 4030 13297
rect 3974 13223 4030 13232
rect 3988 13190 4016 13223
rect 3884 13184 3936 13190
rect 3884 13126 3936 13132
rect 3976 13184 4028 13190
rect 3976 13126 4028 13132
rect 3896 13025 3924 13126
rect 3882 13016 3938 13025
rect 4080 13002 4108 13398
rect 3882 12951 3938 12960
rect 3988 12974 4108 13002
rect 3884 12912 3936 12918
rect 3884 12854 3936 12860
rect 3896 12782 3924 12854
rect 3884 12776 3936 12782
rect 3884 12718 3936 12724
rect 3988 12594 4016 12974
rect 4172 12714 4200 14350
rect 4356 13977 4384 14350
rect 4540 14006 4568 15166
rect 5078 14920 5134 14929
rect 5078 14855 5134 14864
rect 4804 14544 4856 14550
rect 4804 14486 4856 14492
rect 4816 14278 4844 14486
rect 5092 14385 5120 14855
rect 5816 14816 5868 14822
rect 5816 14758 5868 14764
rect 5078 14376 5134 14385
rect 5078 14311 5134 14320
rect 5724 14340 5776 14346
rect 4804 14272 4856 14278
rect 4804 14214 4856 14220
rect 4528 14000 4580 14006
rect 4342 13968 4398 13977
rect 4252 13932 4304 13938
rect 4398 13926 4476 13954
rect 4528 13942 4580 13948
rect 5092 13938 5120 14311
rect 5724 14282 5776 14288
rect 5170 14240 5226 14249
rect 5170 14175 5226 14184
rect 4342 13903 4398 13912
rect 4252 13874 4304 13880
rect 4264 13394 4292 13874
rect 4344 13728 4396 13734
rect 4344 13670 4396 13676
rect 4252 13388 4304 13394
rect 4252 13330 4304 13336
rect 4356 12986 4384 13670
rect 4344 12980 4396 12986
rect 4344 12922 4396 12928
rect 4448 12866 4476 13926
rect 4620 13932 4672 13938
rect 4620 13874 4672 13880
rect 5080 13932 5132 13938
rect 5080 13874 5132 13880
rect 4632 13841 4660 13874
rect 4618 13832 4674 13841
rect 4618 13767 4674 13776
rect 4988 13524 5040 13530
rect 4988 13466 5040 13472
rect 4620 13320 4672 13326
rect 4620 13262 4672 13268
rect 4632 12866 4660 13262
rect 4804 13252 4856 13258
rect 4804 13194 4856 13200
rect 4816 12986 4844 13194
rect 4804 12980 4856 12986
rect 4804 12922 4856 12928
rect 4264 12838 4476 12866
rect 4540 12838 4660 12866
rect 4712 12844 4764 12850
rect 4160 12708 4212 12714
rect 4160 12650 4212 12656
rect 4264 12594 4292 12838
rect 4436 12776 4488 12782
rect 4436 12718 4488 12724
rect 3896 12566 4016 12594
rect 4080 12566 4292 12594
rect 3896 12434 3924 12566
rect 4080 12442 4108 12566
rect 4448 12442 4476 12718
rect 4068 12436 4120 12442
rect 3896 12406 4016 12434
rect 3988 12306 4016 12406
rect 4068 12378 4120 12384
rect 4436 12436 4488 12442
rect 4436 12378 4488 12384
rect 3976 12300 4028 12306
rect 3976 12242 4028 12248
rect 3884 12096 3936 12102
rect 3884 12038 3936 12044
rect 3712 11206 3832 11234
rect 3896 11218 3924 12038
rect 3988 11898 4016 12242
rect 3976 11892 4028 11898
rect 3976 11834 4028 11840
rect 4080 11762 4108 12378
rect 4252 12300 4304 12306
rect 4252 12242 4304 12248
rect 4158 12200 4214 12209
rect 4158 12135 4214 12144
rect 4172 12102 4200 12135
rect 4160 12096 4212 12102
rect 4264 12073 4292 12242
rect 4160 12038 4212 12044
rect 4250 12064 4306 12073
rect 4250 11999 4306 12008
rect 4160 11824 4212 11830
rect 4158 11792 4160 11801
rect 4212 11792 4214 11801
rect 4068 11756 4120 11762
rect 4158 11727 4214 11736
rect 4252 11740 4304 11746
rect 4068 11698 4120 11704
rect 3976 11688 4028 11694
rect 4252 11682 4304 11688
rect 3976 11630 4028 11636
rect 3988 11529 4016 11630
rect 4264 11558 4292 11682
rect 4252 11552 4304 11558
rect 3974 11520 4030 11529
rect 4252 11494 4304 11500
rect 4344 11552 4396 11558
rect 4344 11494 4396 11500
rect 3974 11455 4030 11464
rect 3974 11248 4030 11257
rect 3884 11212 3936 11218
rect 3608 11144 3660 11150
rect 3608 11086 3660 11092
rect 3606 10840 3662 10849
rect 3606 10775 3662 10784
rect 3620 10606 3648 10775
rect 3608 10600 3660 10606
rect 3608 10542 3660 10548
rect 3516 10464 3568 10470
rect 3516 10406 3568 10412
rect 3174 10364 3482 10373
rect 3174 10362 3180 10364
rect 3236 10362 3260 10364
rect 3316 10362 3340 10364
rect 3396 10362 3420 10364
rect 3476 10362 3482 10364
rect 3236 10310 3238 10362
rect 3418 10310 3420 10362
rect 3174 10308 3180 10310
rect 3236 10308 3260 10310
rect 3316 10308 3340 10310
rect 3396 10308 3420 10310
rect 3476 10308 3482 10310
rect 3174 10299 3482 10308
rect 3516 10260 3568 10266
rect 3516 10202 3568 10208
rect 3330 10024 3386 10033
rect 3330 9959 3386 9968
rect 3344 9926 3372 9959
rect 3528 9926 3556 10202
rect 3608 10124 3660 10130
rect 3608 10066 3660 10072
rect 3332 9920 3384 9926
rect 3332 9862 3384 9868
rect 3516 9920 3568 9926
rect 3516 9862 3568 9868
rect 3332 9716 3384 9722
rect 3332 9658 3384 9664
rect 3344 9586 3372 9658
rect 3620 9586 3648 10066
rect 3712 10062 3740 11206
rect 3974 11183 4030 11192
rect 4068 11212 4120 11218
rect 3884 11154 3936 11160
rect 3884 11008 3936 11014
rect 3884 10950 3936 10956
rect 3896 10742 3924 10950
rect 3884 10736 3936 10742
rect 3882 10704 3884 10713
rect 3936 10704 3938 10713
rect 3792 10668 3844 10674
rect 3882 10639 3938 10648
rect 3792 10610 3844 10616
rect 3804 10130 3832 10610
rect 3884 10600 3936 10606
rect 3884 10542 3936 10548
rect 3792 10124 3844 10130
rect 3792 10066 3844 10072
rect 3700 10056 3752 10062
rect 3700 9998 3752 10004
rect 3332 9580 3384 9586
rect 3332 9522 3384 9528
rect 3608 9580 3660 9586
rect 3608 9522 3660 9528
rect 3174 9276 3482 9285
rect 3174 9274 3180 9276
rect 3236 9274 3260 9276
rect 3316 9274 3340 9276
rect 3396 9274 3420 9276
rect 3476 9274 3482 9276
rect 3236 9222 3238 9274
rect 3418 9222 3420 9274
rect 3174 9220 3180 9222
rect 3236 9220 3260 9222
rect 3316 9220 3340 9222
rect 3396 9220 3420 9222
rect 3476 9220 3482 9222
rect 3174 9211 3482 9220
rect 3620 9024 3648 9522
rect 3792 9512 3844 9518
rect 3792 9454 3844 9460
rect 3700 9172 3752 9178
rect 3804 9160 3832 9454
rect 3896 9178 3924 10542
rect 3752 9132 3832 9160
rect 3700 9114 3752 9120
rect 3804 9058 3832 9132
rect 3884 9172 3936 9178
rect 3884 9114 3936 9120
rect 3804 9030 3924 9058
rect 3528 8996 3648 9024
rect 3240 8900 3292 8906
rect 3240 8842 3292 8848
rect 3252 8673 3280 8842
rect 3238 8664 3294 8673
rect 3238 8599 3294 8608
rect 3528 8498 3556 8996
rect 3792 8968 3844 8974
rect 3792 8910 3844 8916
rect 3608 8900 3660 8906
rect 3608 8842 3660 8848
rect 3516 8492 3568 8498
rect 3516 8434 3568 8440
rect 3174 8188 3482 8197
rect 3174 8186 3180 8188
rect 3236 8186 3260 8188
rect 3316 8186 3340 8188
rect 3396 8186 3420 8188
rect 3476 8186 3482 8188
rect 3236 8134 3238 8186
rect 3418 8134 3420 8186
rect 3174 8132 3180 8134
rect 3236 8132 3260 8134
rect 3316 8132 3340 8134
rect 3396 8132 3420 8134
rect 3476 8132 3482 8134
rect 3174 8123 3482 8132
rect 3528 8072 3556 8434
rect 3620 8430 3648 8842
rect 3698 8528 3754 8537
rect 3698 8463 3754 8472
rect 3712 8430 3740 8463
rect 3608 8424 3660 8430
rect 3608 8366 3660 8372
rect 3700 8424 3752 8430
rect 3700 8366 3752 8372
rect 3436 8044 3556 8072
rect 3436 7546 3464 8044
rect 3608 8016 3660 8022
rect 3608 7958 3660 7964
rect 3516 7744 3568 7750
rect 3516 7686 3568 7692
rect 3424 7540 3476 7546
rect 3424 7482 3476 7488
rect 2964 7278 3016 7284
rect 3054 7304 3110 7313
rect 2780 7200 2832 7206
rect 2780 7142 2832 7148
rect 2870 7168 2926 7177
rect 2976 7154 3004 7278
rect 3054 7239 3110 7248
rect 2976 7126 3096 7154
rect 2870 7103 2926 7112
rect 2884 6322 2912 7103
rect 2962 7032 3018 7041
rect 2962 6967 3018 6976
rect 2976 6458 3004 6967
rect 2964 6452 3016 6458
rect 2964 6394 3016 6400
rect 2688 6316 2740 6322
rect 2228 6248 2280 6254
rect 2228 6190 2280 6196
rect 2240 5778 2268 6190
rect 2228 5772 2280 5778
rect 2228 5714 2280 5720
rect 1858 5672 1914 5681
rect 1858 5607 1914 5616
rect 2134 5672 2190 5681
rect 2134 5607 2190 5616
rect 1872 4826 1900 5607
rect 2044 5568 2096 5574
rect 2044 5510 2096 5516
rect 2318 5536 2374 5545
rect 2056 5370 2084 5510
rect 2318 5471 2374 5480
rect 2332 5370 2360 5471
rect 2044 5364 2096 5370
rect 2044 5306 2096 5312
rect 2320 5364 2372 5370
rect 2320 5306 2372 5312
rect 2226 4856 2282 4865
rect 1860 4820 1912 4826
rect 2226 4791 2228 4800
rect 1860 4762 1912 4768
rect 2280 4791 2282 4800
rect 2228 4762 2280 4768
rect 2424 4622 2452 6310
rect 2872 6316 2924 6322
rect 2740 6276 2820 6304
rect 2688 6258 2740 6264
rect 2596 6180 2648 6186
rect 2596 6122 2648 6128
rect 2608 5302 2636 6122
rect 2688 5840 2740 5846
rect 2688 5782 2740 5788
rect 2504 5296 2556 5302
rect 2504 5238 2556 5244
rect 2596 5296 2648 5302
rect 2596 5238 2648 5244
rect 2412 4616 2464 4622
rect 1858 4584 1914 4593
rect 2516 4593 2544 5238
rect 2596 5160 2648 5166
rect 2596 5102 2648 5108
rect 2608 5030 2636 5102
rect 2596 5024 2648 5030
rect 2596 4966 2648 4972
rect 2700 4690 2728 5782
rect 2792 5522 2820 6276
rect 2872 6258 2924 6264
rect 3068 6236 3096 7126
rect 3174 7100 3482 7109
rect 3174 7098 3180 7100
rect 3236 7098 3260 7100
rect 3316 7098 3340 7100
rect 3396 7098 3420 7100
rect 3476 7098 3482 7100
rect 3236 7046 3238 7098
rect 3418 7046 3420 7098
rect 3174 7044 3180 7046
rect 3236 7044 3260 7046
rect 3316 7044 3340 7046
rect 3396 7044 3420 7046
rect 3476 7044 3482 7046
rect 3174 7035 3482 7044
rect 3332 6996 3384 7002
rect 3332 6938 3384 6944
rect 3344 6866 3372 6938
rect 3332 6860 3384 6866
rect 3332 6802 3384 6808
rect 3424 6724 3476 6730
rect 3424 6666 3476 6672
rect 3330 6488 3386 6497
rect 3148 6452 3200 6458
rect 3200 6412 3280 6440
rect 3330 6423 3386 6432
rect 3148 6394 3200 6400
rect 2870 6216 2926 6225
rect 2870 6151 2926 6160
rect 2976 6208 3096 6236
rect 2884 6118 2912 6151
rect 2872 6112 2924 6118
rect 2872 6054 2924 6060
rect 2884 5778 2912 6054
rect 2872 5772 2924 5778
rect 2872 5714 2924 5720
rect 2976 5760 3004 6208
rect 3252 6186 3280 6412
rect 3344 6254 3372 6423
rect 3436 6361 3464 6666
rect 3528 6390 3556 7686
rect 3516 6384 3568 6390
rect 3422 6352 3478 6361
rect 3516 6326 3568 6332
rect 3422 6287 3478 6296
rect 3332 6248 3384 6254
rect 3332 6190 3384 6196
rect 3516 6248 3568 6254
rect 3516 6190 3568 6196
rect 3240 6180 3292 6186
rect 3240 6122 3292 6128
rect 3174 6012 3482 6021
rect 3174 6010 3180 6012
rect 3236 6010 3260 6012
rect 3316 6010 3340 6012
rect 3396 6010 3420 6012
rect 3476 6010 3482 6012
rect 3236 5958 3238 6010
rect 3418 5958 3420 6010
rect 3174 5956 3180 5958
rect 3236 5956 3260 5958
rect 3316 5956 3340 5958
rect 3396 5956 3420 5958
rect 3476 5956 3482 5958
rect 3174 5947 3482 5956
rect 3424 5908 3476 5914
rect 3424 5850 3476 5856
rect 3148 5772 3200 5778
rect 2976 5732 3148 5760
rect 2792 5494 2912 5522
rect 2778 5400 2834 5409
rect 2778 5335 2780 5344
rect 2832 5335 2834 5344
rect 2780 5306 2832 5312
rect 2688 4684 2740 4690
rect 2688 4626 2740 4632
rect 2412 4558 2464 4564
rect 2502 4584 2558 4593
rect 1858 4519 1914 4528
rect 2502 4519 2558 4528
rect 1872 4282 1900 4519
rect 1860 4276 1912 4282
rect 1860 4218 1912 4224
rect 2136 4140 2188 4146
rect 2136 4082 2188 4088
rect 2412 4140 2464 4146
rect 2412 4082 2464 4088
rect 2148 3738 2176 4082
rect 2228 3936 2280 3942
rect 2228 3878 2280 3884
rect 2320 3936 2372 3942
rect 2320 3878 2372 3884
rect 2240 3777 2268 3878
rect 2226 3768 2282 3777
rect 2136 3732 2188 3738
rect 2226 3703 2282 3712
rect 2136 3674 2188 3680
rect 2332 3670 2360 3878
rect 2424 3738 2452 4082
rect 2412 3732 2464 3738
rect 2412 3674 2464 3680
rect 2516 3670 2544 4519
rect 2780 4480 2832 4486
rect 2780 4422 2832 4428
rect 2792 4321 2820 4422
rect 2778 4312 2834 4321
rect 2778 4247 2834 4256
rect 2688 4140 2740 4146
rect 2688 4082 2740 4088
rect 2700 4049 2728 4082
rect 2686 4040 2742 4049
rect 2596 4004 2648 4010
rect 2686 3975 2742 3984
rect 2596 3946 2648 3952
rect 2320 3664 2372 3670
rect 2320 3606 2372 3612
rect 2504 3664 2556 3670
rect 2504 3606 2556 3612
rect 1768 3528 1820 3534
rect 2320 3528 2372 3534
rect 1768 3470 1820 3476
rect 1950 3496 2006 3505
rect 2320 3470 2372 3476
rect 1950 3431 2006 3440
rect 1964 3398 1992 3431
rect 1952 3392 2004 3398
rect 1952 3334 2004 3340
rect 2044 3392 2096 3398
rect 2044 3334 2096 3340
rect 1490 3224 1546 3233
rect 1490 3159 1492 3168
rect 1544 3159 1546 3168
rect 1492 3130 1544 3136
rect 2056 3058 2084 3334
rect 2332 3233 2360 3470
rect 2318 3224 2374 3233
rect 2318 3159 2374 3168
rect 2608 3058 2636 3946
rect 2044 3052 2096 3058
rect 2044 2994 2096 3000
rect 2596 3052 2648 3058
rect 2596 2994 2648 3000
rect 1858 2952 1914 2961
rect 1858 2887 1860 2896
rect 1912 2887 1914 2896
rect 1860 2858 1912 2864
rect 2700 2854 2728 3975
rect 2884 3738 2912 5494
rect 2976 5030 3004 5732
rect 3148 5714 3200 5720
rect 3238 5672 3294 5681
rect 3238 5607 3294 5616
rect 3252 5234 3280 5607
rect 3436 5545 3464 5850
rect 3528 5710 3556 6190
rect 3516 5704 3568 5710
rect 3516 5646 3568 5652
rect 3422 5536 3478 5545
rect 3422 5471 3478 5480
rect 3514 5264 3570 5273
rect 3240 5228 3292 5234
rect 3514 5199 3516 5208
rect 3240 5170 3292 5176
rect 3568 5199 3570 5208
rect 3516 5170 3568 5176
rect 3422 5128 3478 5137
rect 3422 5063 3424 5072
rect 3476 5063 3478 5072
rect 3424 5034 3476 5040
rect 2964 5024 3016 5030
rect 2964 4966 3016 4972
rect 3516 5024 3568 5030
rect 3516 4966 3568 4972
rect 3174 4924 3482 4933
rect 3174 4922 3180 4924
rect 3236 4922 3260 4924
rect 3316 4922 3340 4924
rect 3396 4922 3420 4924
rect 3476 4922 3482 4924
rect 3236 4870 3238 4922
rect 3418 4870 3420 4922
rect 3174 4868 3180 4870
rect 3236 4868 3260 4870
rect 3316 4868 3340 4870
rect 3396 4868 3420 4870
rect 3476 4868 3482 4870
rect 3174 4859 3482 4868
rect 3330 4720 3386 4729
rect 3330 4655 3386 4664
rect 3344 4622 3372 4655
rect 3332 4616 3384 4622
rect 3332 4558 3384 4564
rect 2964 4480 3016 4486
rect 2964 4422 3016 4428
rect 3056 4480 3108 4486
rect 3056 4422 3108 4428
rect 2872 3732 2924 3738
rect 2872 3674 2924 3680
rect 2780 3528 2832 3534
rect 2778 3496 2780 3505
rect 2832 3496 2834 3505
rect 2778 3431 2834 3440
rect 2780 3392 2832 3398
rect 2780 3334 2832 3340
rect 2228 2848 2280 2854
rect 2228 2790 2280 2796
rect 2596 2848 2648 2854
rect 2596 2790 2648 2796
rect 2688 2848 2740 2854
rect 2688 2790 2740 2796
rect 1490 2680 1546 2689
rect 1490 2615 1492 2624
rect 1544 2615 1546 2624
rect 1492 2586 1544 2592
rect 1858 2408 1914 2417
rect 1858 2343 1914 2352
rect 1872 2310 1900 2343
rect 1860 2304 1912 2310
rect 1860 2246 1912 2252
rect 2044 2304 2096 2310
rect 2044 2246 2096 2252
rect 1216 2100 1268 2106
rect 1216 2042 1268 2048
rect 1228 800 1256 2042
rect 2056 800 2084 2246
rect 2240 1873 2268 2790
rect 2608 2145 2636 2790
rect 2792 2446 2820 3334
rect 2976 2650 3004 4422
rect 2964 2644 3016 2650
rect 2964 2586 3016 2592
rect 3068 2514 3096 4422
rect 3344 4214 3372 4558
rect 3528 4282 3556 4966
rect 3620 4622 3648 7958
rect 3700 7812 3752 7818
rect 3700 7754 3752 7760
rect 3712 7002 3740 7754
rect 3804 7546 3832 8910
rect 3896 8430 3924 9030
rect 3988 8945 4016 11183
rect 4068 11154 4120 11160
rect 4160 11212 4212 11218
rect 4160 11154 4212 11160
rect 4080 10742 4108 11154
rect 4172 10849 4200 11154
rect 4158 10840 4214 10849
rect 4158 10775 4214 10784
rect 4068 10736 4120 10742
rect 4068 10678 4120 10684
rect 4160 10668 4212 10674
rect 4160 10610 4212 10616
rect 4172 10266 4200 10610
rect 4160 10260 4212 10266
rect 4160 10202 4212 10208
rect 4068 10056 4120 10062
rect 4068 9998 4120 10004
rect 4080 9926 4108 9998
rect 4068 9920 4120 9926
rect 4068 9862 4120 9868
rect 4068 9716 4120 9722
rect 4068 9658 4120 9664
rect 4160 9716 4212 9722
rect 4160 9658 4212 9664
rect 3974 8936 4030 8945
rect 3974 8871 4030 8880
rect 3976 8628 4028 8634
rect 3976 8570 4028 8576
rect 3884 8424 3936 8430
rect 3884 8366 3936 8372
rect 3792 7540 3844 7546
rect 3792 7482 3844 7488
rect 3792 7404 3844 7410
rect 3792 7346 3844 7352
rect 3804 7313 3832 7346
rect 3790 7304 3846 7313
rect 3790 7239 3846 7248
rect 3700 6996 3752 7002
rect 3700 6938 3752 6944
rect 3700 6656 3752 6662
rect 3700 6598 3752 6604
rect 3712 6254 3740 6598
rect 3700 6248 3752 6254
rect 3700 6190 3752 6196
rect 3792 6180 3844 6186
rect 3792 6122 3844 6128
rect 3700 6112 3752 6118
rect 3700 6054 3752 6060
rect 3608 4616 3660 4622
rect 3608 4558 3660 4564
rect 3608 4480 3660 4486
rect 3608 4422 3660 4428
rect 3516 4276 3568 4282
rect 3516 4218 3568 4224
rect 3332 4208 3384 4214
rect 3332 4150 3384 4156
rect 3424 4140 3476 4146
rect 3424 4082 3476 4088
rect 3436 4049 3464 4082
rect 3422 4040 3478 4049
rect 3422 3975 3478 3984
rect 3174 3836 3482 3845
rect 3174 3834 3180 3836
rect 3236 3834 3260 3836
rect 3316 3834 3340 3836
rect 3396 3834 3420 3836
rect 3476 3834 3482 3836
rect 3236 3782 3238 3834
rect 3418 3782 3420 3834
rect 3174 3780 3180 3782
rect 3236 3780 3260 3782
rect 3316 3780 3340 3782
rect 3396 3780 3420 3782
rect 3476 3780 3482 3782
rect 3174 3771 3482 3780
rect 3528 3738 3556 4218
rect 3516 3732 3568 3738
rect 3516 3674 3568 3680
rect 3516 3460 3568 3466
rect 3516 3402 3568 3408
rect 3528 2990 3556 3402
rect 3516 2984 3568 2990
rect 3516 2926 3568 2932
rect 3516 2848 3568 2854
rect 3516 2790 3568 2796
rect 3174 2748 3482 2757
rect 3174 2746 3180 2748
rect 3236 2746 3260 2748
rect 3316 2746 3340 2748
rect 3396 2746 3420 2748
rect 3476 2746 3482 2748
rect 3236 2694 3238 2746
rect 3418 2694 3420 2746
rect 3174 2692 3180 2694
rect 3236 2692 3260 2694
rect 3316 2692 3340 2694
rect 3396 2692 3420 2694
rect 3476 2692 3482 2694
rect 3174 2683 3482 2692
rect 3056 2508 3108 2514
rect 3056 2450 3108 2456
rect 3528 2446 3556 2790
rect 3620 2514 3648 4422
rect 3712 3058 3740 6054
rect 3804 5710 3832 6122
rect 3792 5704 3844 5710
rect 3792 5646 3844 5652
rect 3804 4826 3832 5646
rect 3896 5574 3924 8366
rect 3988 7274 4016 8570
rect 3976 7268 4028 7274
rect 3976 7210 4028 7216
rect 3988 7041 4016 7210
rect 3974 7032 4030 7041
rect 3974 6967 4030 6976
rect 3974 6896 4030 6905
rect 3974 6831 4030 6840
rect 3988 6798 4016 6831
rect 4080 6798 4108 9658
rect 4172 8974 4200 9658
rect 4160 8968 4212 8974
rect 4160 8910 4212 8916
rect 4160 8832 4212 8838
rect 4160 8774 4212 8780
rect 4172 8498 4200 8774
rect 4160 8492 4212 8498
rect 4160 8434 4212 8440
rect 4264 8090 4292 11494
rect 4356 11150 4384 11494
rect 4344 11144 4396 11150
rect 4344 11086 4396 11092
rect 4436 11008 4488 11014
rect 4436 10950 4488 10956
rect 4448 10810 4476 10950
rect 4436 10804 4488 10810
rect 4436 10746 4488 10752
rect 4344 9512 4396 9518
rect 4344 9454 4396 9460
rect 4356 8537 4384 9454
rect 4540 9160 4568 12838
rect 4712 12786 4764 12792
rect 4620 12776 4672 12782
rect 4620 12718 4672 12724
rect 4632 12322 4660 12718
rect 4724 12442 4752 12786
rect 4712 12436 4764 12442
rect 4712 12378 4764 12384
rect 4804 12436 4856 12442
rect 4804 12378 4856 12384
rect 4816 12322 4844 12378
rect 4632 12294 4844 12322
rect 5000 12238 5028 13466
rect 5078 13424 5134 13433
rect 5078 13359 5134 13368
rect 5092 13190 5120 13359
rect 5184 13326 5212 14175
rect 5398 14172 5706 14181
rect 5398 14170 5404 14172
rect 5460 14170 5484 14172
rect 5540 14170 5564 14172
rect 5620 14170 5644 14172
rect 5700 14170 5706 14172
rect 5460 14118 5462 14170
rect 5642 14118 5644 14170
rect 5398 14116 5404 14118
rect 5460 14116 5484 14118
rect 5540 14116 5564 14118
rect 5620 14116 5644 14118
rect 5700 14116 5706 14118
rect 5398 14107 5706 14116
rect 5736 14074 5764 14282
rect 5724 14068 5776 14074
rect 5724 14010 5776 14016
rect 5264 13932 5316 13938
rect 5264 13874 5316 13880
rect 5276 13841 5304 13874
rect 5262 13832 5318 13841
rect 5262 13767 5318 13776
rect 5828 13530 5856 14758
rect 6012 14618 6040 16400
rect 6276 14884 6328 14890
rect 6276 14826 6328 14832
rect 6000 14612 6052 14618
rect 6000 14554 6052 14560
rect 5816 13524 5868 13530
rect 5816 13466 5868 13472
rect 5172 13320 5224 13326
rect 5172 13262 5224 13268
rect 5080 13184 5132 13190
rect 5080 13126 5132 13132
rect 5092 12986 5120 13126
rect 5080 12980 5132 12986
rect 5080 12922 5132 12928
rect 5184 12782 5212 13262
rect 5264 13184 5316 13190
rect 5262 13152 5264 13161
rect 5316 13152 5318 13161
rect 5262 13087 5318 13096
rect 5398 13084 5706 13093
rect 5398 13082 5404 13084
rect 5460 13082 5484 13084
rect 5540 13082 5564 13084
rect 5620 13082 5644 13084
rect 5700 13082 5706 13084
rect 5460 13030 5462 13082
rect 5642 13030 5644 13082
rect 5398 13028 5404 13030
rect 5460 13028 5484 13030
rect 5540 13028 5564 13030
rect 5620 13028 5644 13030
rect 5700 13028 5706 13030
rect 5398 13019 5706 13028
rect 5264 12980 5316 12986
rect 5264 12922 5316 12928
rect 6184 12980 6236 12986
rect 6184 12922 6236 12928
rect 5276 12850 5304 12922
rect 5264 12844 5316 12850
rect 5264 12786 5316 12792
rect 5540 12844 5592 12850
rect 5540 12786 5592 12792
rect 5172 12776 5224 12782
rect 5170 12744 5172 12753
rect 5224 12744 5226 12753
rect 5170 12679 5226 12688
rect 5356 12640 5408 12646
rect 5552 12617 5580 12786
rect 5356 12582 5408 12588
rect 5538 12608 5594 12617
rect 5368 12374 5396 12582
rect 5538 12543 5594 12552
rect 5356 12368 5408 12374
rect 5356 12310 5408 12316
rect 6000 12368 6052 12374
rect 6000 12310 6052 12316
rect 4804 12232 4856 12238
rect 4988 12232 5040 12238
rect 4856 12180 4936 12186
rect 4804 12174 4936 12180
rect 6012 12209 6040 12310
rect 6092 12232 6144 12238
rect 5998 12200 6054 12209
rect 4988 12174 5040 12180
rect 4816 12158 4936 12174
rect 4804 12096 4856 12102
rect 4804 12038 4856 12044
rect 4908 12050 4936 12158
rect 5644 12170 5948 12186
rect 5644 12164 5960 12170
rect 5644 12158 5908 12164
rect 5644 12102 5672 12158
rect 6092 12174 6144 12180
rect 5998 12135 6054 12144
rect 5908 12106 5960 12112
rect 5172 12096 5224 12102
rect 4908 12044 5172 12050
rect 4908 12038 5224 12044
rect 5632 12096 5684 12102
rect 5632 12038 5684 12044
rect 5724 12096 5776 12102
rect 5724 12038 5776 12044
rect 4816 11558 4844 12038
rect 4908 12022 5212 12038
rect 5398 11996 5706 12005
rect 5398 11994 5404 11996
rect 5460 11994 5484 11996
rect 5540 11994 5564 11996
rect 5620 11994 5644 11996
rect 5700 11994 5706 11996
rect 5460 11942 5462 11994
rect 5642 11942 5644 11994
rect 5398 11940 5404 11942
rect 5460 11940 5484 11942
rect 5540 11940 5564 11942
rect 5620 11940 5644 11942
rect 5700 11940 5706 11942
rect 5398 11931 5706 11940
rect 5632 11892 5684 11898
rect 5632 11834 5684 11840
rect 5644 11801 5672 11834
rect 5630 11792 5686 11801
rect 5080 11756 5132 11762
rect 5630 11727 5686 11736
rect 5080 11698 5132 11704
rect 4804 11552 4856 11558
rect 4710 11520 4766 11529
rect 4804 11494 4856 11500
rect 4710 11455 4766 11464
rect 4724 10606 4752 11455
rect 4894 11112 4950 11121
rect 4894 11047 4950 11056
rect 4712 10600 4764 10606
rect 4712 10542 4764 10548
rect 4724 10130 4752 10542
rect 4712 10124 4764 10130
rect 4712 10066 4764 10072
rect 4804 10124 4856 10130
rect 4804 10066 4856 10072
rect 4620 9920 4672 9926
rect 4620 9862 4672 9868
rect 4632 9722 4660 9862
rect 4620 9716 4672 9722
rect 4620 9658 4672 9664
rect 4540 9132 4660 9160
rect 4528 8968 4580 8974
rect 4528 8910 4580 8916
rect 4436 8832 4488 8838
rect 4436 8774 4488 8780
rect 4448 8634 4476 8774
rect 4540 8634 4568 8910
rect 4436 8628 4488 8634
rect 4436 8570 4488 8576
rect 4528 8628 4580 8634
rect 4528 8570 4580 8576
rect 4342 8528 4398 8537
rect 4342 8463 4398 8472
rect 4436 8288 4488 8294
rect 4436 8230 4488 8236
rect 4528 8288 4580 8294
rect 4528 8230 4580 8236
rect 4252 8084 4304 8090
rect 4252 8026 4304 8032
rect 4344 7948 4396 7954
rect 4344 7890 4396 7896
rect 4160 7744 4212 7750
rect 4160 7686 4212 7692
rect 4172 6866 4200 7686
rect 4356 7478 4384 7890
rect 4448 7818 4476 8230
rect 4436 7812 4488 7818
rect 4436 7754 4488 7760
rect 4436 7540 4488 7546
rect 4436 7482 4488 7488
rect 4252 7472 4304 7478
rect 4252 7414 4304 7420
rect 4344 7472 4396 7478
rect 4344 7414 4396 7420
rect 4264 7002 4292 7414
rect 4252 6996 4304 7002
rect 4252 6938 4304 6944
rect 4160 6860 4212 6866
rect 4160 6802 4212 6808
rect 3976 6792 4028 6798
rect 3976 6734 4028 6740
rect 4068 6792 4120 6798
rect 4068 6734 4120 6740
rect 3974 6352 4030 6361
rect 4080 6338 4108 6734
rect 4160 6656 4212 6662
rect 4160 6598 4212 6604
rect 4172 6458 4200 6598
rect 4160 6452 4212 6458
rect 4160 6394 4212 6400
rect 4080 6310 4200 6338
rect 3974 6287 4030 6296
rect 3988 6186 4016 6287
rect 3976 6180 4028 6186
rect 3976 6122 4028 6128
rect 3884 5568 3936 5574
rect 3884 5510 3936 5516
rect 3988 5352 4016 6122
rect 4068 5636 4120 5642
rect 4068 5578 4120 5584
rect 4080 5409 4108 5578
rect 3896 5324 4016 5352
rect 4066 5400 4122 5409
rect 4066 5335 4122 5344
rect 3792 4820 3844 4826
rect 3792 4762 3844 4768
rect 3790 4720 3846 4729
rect 3790 4655 3846 4664
rect 3804 4622 3832 4655
rect 3792 4616 3844 4622
rect 3792 4558 3844 4564
rect 3790 4312 3846 4321
rect 3790 4247 3792 4256
rect 3844 4247 3846 4256
rect 3792 4218 3844 4224
rect 3896 4146 3924 5324
rect 3974 5264 4030 5273
rect 3974 5199 4030 5208
rect 3988 4758 4016 5199
rect 3976 4752 4028 4758
rect 3976 4694 4028 4700
rect 3884 4140 3936 4146
rect 3884 4082 3936 4088
rect 3792 3392 3844 3398
rect 3792 3334 3844 3340
rect 3804 3194 3832 3334
rect 3882 3224 3938 3233
rect 3792 3188 3844 3194
rect 3882 3159 3884 3168
rect 3792 3130 3844 3136
rect 3936 3159 3938 3168
rect 3884 3130 3936 3136
rect 4080 3126 4108 5335
rect 4172 4554 4200 6310
rect 4252 6316 4304 6322
rect 4252 6258 4304 6264
rect 4264 5846 4292 6258
rect 4356 6254 4384 7414
rect 4448 7290 4476 7482
rect 4540 7426 4568 8230
rect 4632 8022 4660 9132
rect 4724 9042 4752 10066
rect 4816 9897 4844 10066
rect 4802 9888 4858 9897
rect 4802 9823 4858 9832
rect 4908 9722 4936 11047
rect 4988 11008 5040 11014
rect 4986 10976 4988 10985
rect 5040 10976 5042 10985
rect 4986 10911 5042 10920
rect 5000 10810 5028 10911
rect 4988 10804 5040 10810
rect 4988 10746 5040 10752
rect 4988 10600 5040 10606
rect 4988 10542 5040 10548
rect 5000 10470 5028 10542
rect 4988 10464 5040 10470
rect 4986 10432 4988 10441
rect 5040 10432 5042 10441
rect 4986 10367 5042 10376
rect 5092 9994 5120 11698
rect 5172 11688 5224 11694
rect 5172 11630 5224 11636
rect 5080 9988 5132 9994
rect 5080 9930 5132 9936
rect 4896 9716 4948 9722
rect 4896 9658 4948 9664
rect 4908 9178 4936 9658
rect 4896 9172 4948 9178
rect 4896 9114 4948 9120
rect 5184 9110 5212 11630
rect 5736 11257 5764 12038
rect 6104 11898 6132 12174
rect 6092 11892 6144 11898
rect 6092 11834 6144 11840
rect 5814 11792 5870 11801
rect 5814 11727 5816 11736
rect 5868 11727 5870 11736
rect 5816 11698 5868 11704
rect 5722 11248 5778 11257
rect 5722 11183 5778 11192
rect 5828 11121 5856 11698
rect 5906 11656 5962 11665
rect 5906 11591 5908 11600
rect 5960 11591 5962 11600
rect 6000 11620 6052 11626
rect 5908 11562 5960 11568
rect 6000 11562 6052 11568
rect 6012 11234 6040 11562
rect 5920 11206 6040 11234
rect 5814 11112 5870 11121
rect 5814 11047 5870 11056
rect 5816 11008 5868 11014
rect 5816 10950 5868 10956
rect 5398 10908 5706 10917
rect 5398 10906 5404 10908
rect 5460 10906 5484 10908
rect 5540 10906 5564 10908
rect 5620 10906 5644 10908
rect 5700 10906 5706 10908
rect 5460 10854 5462 10906
rect 5642 10854 5644 10906
rect 5398 10852 5404 10854
rect 5460 10852 5484 10854
rect 5540 10852 5564 10854
rect 5620 10852 5644 10854
rect 5700 10852 5706 10854
rect 5262 10840 5318 10849
rect 5398 10843 5706 10852
rect 5318 10784 5396 10792
rect 5262 10775 5396 10784
rect 5276 10764 5396 10775
rect 5368 10470 5396 10764
rect 5722 10704 5778 10713
rect 5722 10639 5724 10648
rect 5776 10639 5778 10648
rect 5724 10610 5776 10616
rect 5632 10600 5684 10606
rect 5632 10542 5684 10548
rect 5356 10464 5408 10470
rect 5356 10406 5408 10412
rect 5644 10266 5672 10542
rect 5632 10260 5684 10266
rect 5632 10202 5684 10208
rect 5262 10160 5318 10169
rect 5262 10095 5318 10104
rect 5276 9518 5304 10095
rect 5736 10010 5764 10610
rect 5828 10538 5856 10950
rect 5920 10742 5948 11206
rect 6196 11098 6224 12922
rect 6288 11529 6316 14826
rect 8576 14816 8628 14822
rect 8576 14758 8628 14764
rect 7622 14716 7930 14725
rect 7622 14714 7628 14716
rect 7684 14714 7708 14716
rect 7764 14714 7788 14716
rect 7844 14714 7868 14716
rect 7924 14714 7930 14716
rect 7684 14662 7686 14714
rect 7866 14662 7868 14714
rect 7622 14660 7628 14662
rect 7684 14660 7708 14662
rect 7764 14660 7788 14662
rect 7844 14660 7868 14662
rect 7924 14660 7930 14662
rect 7622 14651 7930 14660
rect 8484 14476 8536 14482
rect 8484 14418 8536 14424
rect 8116 14068 8168 14074
rect 8116 14010 8168 14016
rect 7288 14000 7340 14006
rect 7288 13942 7340 13948
rect 6920 12640 6972 12646
rect 6920 12582 6972 12588
rect 6932 12434 6960 12582
rect 6932 12406 7052 12434
rect 6458 12064 6514 12073
rect 6458 11999 6514 12008
rect 6274 11520 6330 11529
rect 6274 11455 6330 11464
rect 6472 11393 6500 11999
rect 6458 11384 6514 11393
rect 6458 11319 6514 11328
rect 6012 11070 6224 11098
rect 5908 10736 5960 10742
rect 5908 10678 5960 10684
rect 5906 10568 5962 10577
rect 5816 10532 5868 10538
rect 5906 10503 5962 10512
rect 5816 10474 5868 10480
rect 5736 9982 5856 10010
rect 5724 9920 5776 9926
rect 5724 9862 5776 9868
rect 5398 9820 5706 9829
rect 5398 9818 5404 9820
rect 5460 9818 5484 9820
rect 5540 9818 5564 9820
rect 5620 9818 5644 9820
rect 5700 9818 5706 9820
rect 5460 9766 5462 9818
rect 5642 9766 5644 9818
rect 5398 9764 5404 9766
rect 5460 9764 5484 9766
rect 5540 9764 5564 9766
rect 5620 9764 5644 9766
rect 5700 9764 5706 9766
rect 5398 9755 5706 9764
rect 5736 9722 5764 9862
rect 5724 9716 5776 9722
rect 5724 9658 5776 9664
rect 5356 9580 5408 9586
rect 5356 9522 5408 9528
rect 5264 9512 5316 9518
rect 5264 9454 5316 9460
rect 5264 9376 5316 9382
rect 5264 9318 5316 9324
rect 5172 9104 5224 9110
rect 5172 9046 5224 9052
rect 4712 9036 4764 9042
rect 4712 8978 4764 8984
rect 5276 8974 5304 9318
rect 5368 9217 5396 9522
rect 5354 9208 5410 9217
rect 5354 9143 5410 9152
rect 5264 8968 5316 8974
rect 5264 8910 5316 8916
rect 5080 8900 5132 8906
rect 5080 8842 5132 8848
rect 4896 8832 4948 8838
rect 4896 8774 4948 8780
rect 4712 8356 4764 8362
rect 4712 8298 4764 8304
rect 4620 8016 4672 8022
rect 4620 7958 4672 7964
rect 4540 7398 4660 7426
rect 4632 7342 4660 7398
rect 4620 7336 4672 7342
rect 4448 7262 4568 7290
rect 4620 7278 4672 7284
rect 4436 7200 4488 7206
rect 4436 7142 4488 7148
rect 4448 6798 4476 7142
rect 4436 6792 4488 6798
rect 4434 6760 4436 6769
rect 4488 6760 4490 6769
rect 4434 6695 4490 6704
rect 4436 6384 4488 6390
rect 4436 6326 4488 6332
rect 4344 6248 4396 6254
rect 4344 6190 4396 6196
rect 4252 5840 4304 5846
rect 4252 5782 4304 5788
rect 4252 5704 4304 5710
rect 4252 5646 4304 5652
rect 4264 5545 4292 5646
rect 4344 5568 4396 5574
rect 4250 5536 4306 5545
rect 4344 5510 4396 5516
rect 4250 5471 4306 5480
rect 4264 5370 4292 5471
rect 4252 5364 4304 5370
rect 4252 5306 4304 5312
rect 4250 4856 4306 4865
rect 4250 4791 4252 4800
rect 4304 4791 4306 4800
rect 4252 4762 4304 4768
rect 4356 4690 4384 5510
rect 4448 4826 4476 6326
rect 4436 4820 4488 4826
rect 4436 4762 4488 4768
rect 4344 4684 4396 4690
rect 4344 4626 4396 4632
rect 4540 4554 4568 7262
rect 4160 4548 4212 4554
rect 4160 4490 4212 4496
rect 4528 4548 4580 4554
rect 4528 4490 4580 4496
rect 4158 4448 4214 4457
rect 4158 4383 4214 4392
rect 4172 4146 4200 4383
rect 4160 4140 4212 4146
rect 4160 4082 4212 4088
rect 4632 4010 4660 7278
rect 4724 6458 4752 8298
rect 4908 8294 4936 8774
rect 5092 8498 5120 8842
rect 5172 8832 5224 8838
rect 5172 8774 5224 8780
rect 5080 8492 5132 8498
rect 5080 8434 5132 8440
rect 4896 8288 4948 8294
rect 4896 8230 4948 8236
rect 5080 8084 5132 8090
rect 5080 8026 5132 8032
rect 4802 7848 4858 7857
rect 4802 7783 4858 7792
rect 4816 6866 4844 7783
rect 4896 7744 4948 7750
rect 4896 7686 4948 7692
rect 4908 7546 4936 7686
rect 4896 7540 4948 7546
rect 4896 7482 4948 7488
rect 4988 7540 5040 7546
rect 4988 7482 5040 7488
rect 4894 7440 4950 7449
rect 4894 7375 4950 7384
rect 4804 6860 4856 6866
rect 4804 6802 4856 6808
rect 4712 6452 4764 6458
rect 4712 6394 4764 6400
rect 4816 6254 4844 6802
rect 4908 6497 4936 7375
rect 5000 7002 5028 7482
rect 5092 7410 5120 8026
rect 5184 7954 5212 8774
rect 5276 8498 5304 8910
rect 5398 8732 5706 8741
rect 5398 8730 5404 8732
rect 5460 8730 5484 8732
rect 5540 8730 5564 8732
rect 5620 8730 5644 8732
rect 5700 8730 5706 8732
rect 5460 8678 5462 8730
rect 5642 8678 5644 8730
rect 5398 8676 5404 8678
rect 5460 8676 5484 8678
rect 5540 8676 5564 8678
rect 5620 8676 5644 8678
rect 5700 8676 5706 8678
rect 5398 8667 5706 8676
rect 5264 8492 5316 8498
rect 5264 8434 5316 8440
rect 5724 8424 5776 8430
rect 5724 8366 5776 8372
rect 5264 8288 5316 8294
rect 5264 8230 5316 8236
rect 5276 7954 5304 8230
rect 5172 7948 5224 7954
rect 5172 7890 5224 7896
rect 5264 7948 5316 7954
rect 5264 7890 5316 7896
rect 5172 7744 5224 7750
rect 5172 7686 5224 7692
rect 5080 7404 5132 7410
rect 5080 7346 5132 7352
rect 5092 7206 5120 7346
rect 5080 7200 5132 7206
rect 5080 7142 5132 7148
rect 4988 6996 5040 7002
rect 4988 6938 5040 6944
rect 4988 6860 5040 6866
rect 4988 6802 5040 6808
rect 4894 6488 4950 6497
rect 4894 6423 4950 6432
rect 5000 6361 5028 6802
rect 4986 6352 5042 6361
rect 5092 6322 5120 7142
rect 5184 6390 5212 7686
rect 5276 6934 5304 7890
rect 5398 7644 5706 7653
rect 5398 7642 5404 7644
rect 5460 7642 5484 7644
rect 5540 7642 5564 7644
rect 5620 7642 5644 7644
rect 5700 7642 5706 7644
rect 5460 7590 5462 7642
rect 5642 7590 5644 7642
rect 5398 7588 5404 7590
rect 5460 7588 5484 7590
rect 5540 7588 5564 7590
rect 5620 7588 5644 7590
rect 5700 7588 5706 7590
rect 5398 7579 5706 7588
rect 5736 7528 5764 8366
rect 5828 7886 5856 9982
rect 5920 9897 5948 10503
rect 5906 9888 5962 9897
rect 5906 9823 5962 9832
rect 5906 9072 5962 9081
rect 5906 9007 5962 9016
rect 5920 8838 5948 9007
rect 5908 8832 5960 8838
rect 5908 8774 5960 8780
rect 5816 7880 5868 7886
rect 5816 7822 5868 7828
rect 5816 7744 5868 7750
rect 5816 7686 5868 7692
rect 5828 7546 5856 7686
rect 5644 7500 5764 7528
rect 5816 7540 5868 7546
rect 5644 7342 5672 7500
rect 5816 7482 5868 7488
rect 5632 7336 5684 7342
rect 5632 7278 5684 7284
rect 5920 7188 5948 8774
rect 5552 7160 5948 7188
rect 5264 6928 5316 6934
rect 5264 6870 5316 6876
rect 5448 6860 5500 6866
rect 5552 6848 5580 7160
rect 5906 7032 5962 7041
rect 5816 6996 5868 7002
rect 5906 6967 5962 6976
rect 5816 6938 5868 6944
rect 5500 6820 5580 6848
rect 5724 6860 5776 6866
rect 5448 6802 5500 6808
rect 5724 6802 5776 6808
rect 5460 6662 5488 6802
rect 5264 6656 5316 6662
rect 5262 6624 5264 6633
rect 5448 6656 5500 6662
rect 5316 6624 5318 6633
rect 5448 6598 5500 6604
rect 5262 6559 5318 6568
rect 5172 6384 5224 6390
rect 5172 6326 5224 6332
rect 4986 6287 5042 6296
rect 5080 6316 5132 6322
rect 5080 6258 5132 6264
rect 4804 6248 4856 6254
rect 5276 6225 5304 6559
rect 5398 6556 5706 6565
rect 5398 6554 5404 6556
rect 5460 6554 5484 6556
rect 5540 6554 5564 6556
rect 5620 6554 5644 6556
rect 5700 6554 5706 6556
rect 5460 6502 5462 6554
rect 5642 6502 5644 6554
rect 5398 6500 5404 6502
rect 5460 6500 5484 6502
rect 5540 6500 5564 6502
rect 5620 6500 5644 6502
rect 5700 6500 5706 6502
rect 5398 6491 5706 6500
rect 5354 6352 5410 6361
rect 5354 6287 5410 6296
rect 5448 6316 5500 6322
rect 5262 6216 5318 6225
rect 4804 6190 4856 6196
rect 5092 6174 5262 6202
rect 4712 6112 4764 6118
rect 4712 6054 4764 6060
rect 4804 6112 4856 6118
rect 4804 6054 4856 6060
rect 4724 5030 4752 6054
rect 4816 5681 4844 6054
rect 4988 5908 5040 5914
rect 4988 5850 5040 5856
rect 4896 5772 4948 5778
rect 4896 5714 4948 5720
rect 4802 5672 4858 5681
rect 4802 5607 4858 5616
rect 4712 5024 4764 5030
rect 4712 4966 4764 4972
rect 4620 4004 4672 4010
rect 4620 3946 4672 3952
rect 4724 3534 4752 4966
rect 4816 4826 4844 5607
rect 4908 5409 4936 5714
rect 4894 5400 4950 5409
rect 4894 5335 4950 5344
rect 4908 5302 4936 5335
rect 5000 5302 5028 5850
rect 5092 5370 5120 6174
rect 5262 6151 5318 6160
rect 5368 5710 5396 6287
rect 5448 6258 5500 6264
rect 5460 5953 5488 6258
rect 5632 6248 5684 6254
rect 5632 6190 5684 6196
rect 5446 5944 5502 5953
rect 5644 5914 5672 6190
rect 5446 5879 5502 5888
rect 5632 5908 5684 5914
rect 5632 5850 5684 5856
rect 5736 5778 5764 6802
rect 5828 6458 5856 6938
rect 5816 6452 5868 6458
rect 5816 6394 5868 6400
rect 5920 6338 5948 6967
rect 5828 6310 5948 6338
rect 5724 5772 5776 5778
rect 5724 5714 5776 5720
rect 5356 5704 5408 5710
rect 5356 5646 5408 5652
rect 5724 5636 5776 5642
rect 5724 5578 5776 5584
rect 5172 5568 5224 5574
rect 5172 5510 5224 5516
rect 5264 5568 5316 5574
rect 5264 5510 5316 5516
rect 5080 5364 5132 5370
rect 5080 5306 5132 5312
rect 4896 5296 4948 5302
rect 4896 5238 4948 5244
rect 4988 5296 5040 5302
rect 4988 5238 5040 5244
rect 5184 4826 5212 5510
rect 5276 5370 5304 5510
rect 5398 5468 5706 5477
rect 5398 5466 5404 5468
rect 5460 5466 5484 5468
rect 5540 5466 5564 5468
rect 5620 5466 5644 5468
rect 5700 5466 5706 5468
rect 5460 5414 5462 5466
rect 5642 5414 5644 5466
rect 5398 5412 5404 5414
rect 5460 5412 5484 5414
rect 5540 5412 5564 5414
rect 5620 5412 5644 5414
rect 5700 5412 5706 5414
rect 5398 5403 5706 5412
rect 5264 5364 5316 5370
rect 5264 5306 5316 5312
rect 5632 5296 5684 5302
rect 5632 5238 5684 5244
rect 4804 4820 4856 4826
rect 4804 4762 4856 4768
rect 5172 4820 5224 4826
rect 5172 4762 5224 4768
rect 5644 4690 5672 5238
rect 5632 4684 5684 4690
rect 5632 4626 5684 4632
rect 4988 4616 5040 4622
rect 5080 4616 5132 4622
rect 4988 4558 5040 4564
rect 5078 4584 5080 4593
rect 5132 4584 5134 4593
rect 5000 4185 5028 4558
rect 5078 4519 5134 4528
rect 5172 4480 5224 4486
rect 5172 4422 5224 4428
rect 4986 4176 5042 4185
rect 4986 4111 5042 4120
rect 4712 3528 4764 3534
rect 4710 3496 4712 3505
rect 4764 3496 4766 3505
rect 4710 3431 4766 3440
rect 4068 3120 4120 3126
rect 4068 3062 4120 3068
rect 3700 3052 3752 3058
rect 3700 2994 3752 3000
rect 4896 2848 4948 2854
rect 4896 2790 4948 2796
rect 3608 2508 3660 2514
rect 3608 2450 3660 2456
rect 4908 2446 4936 2790
rect 5184 2446 5212 4422
rect 5398 4380 5706 4389
rect 5398 4378 5404 4380
rect 5460 4378 5484 4380
rect 5540 4378 5564 4380
rect 5620 4378 5644 4380
rect 5700 4378 5706 4380
rect 5460 4326 5462 4378
rect 5642 4326 5644 4378
rect 5398 4324 5404 4326
rect 5460 4324 5484 4326
rect 5540 4324 5564 4326
rect 5620 4324 5644 4326
rect 5700 4324 5706 4326
rect 5398 4315 5706 4324
rect 5398 3292 5706 3301
rect 5398 3290 5404 3292
rect 5460 3290 5484 3292
rect 5540 3290 5564 3292
rect 5620 3290 5644 3292
rect 5700 3290 5706 3292
rect 5460 3238 5462 3290
rect 5642 3238 5644 3290
rect 5398 3236 5404 3238
rect 5460 3236 5484 3238
rect 5540 3236 5564 3238
rect 5620 3236 5644 3238
rect 5700 3236 5706 3238
rect 5398 3227 5706 3236
rect 5736 2990 5764 5578
rect 5828 5574 5856 6310
rect 5906 6080 5962 6089
rect 5906 6015 5962 6024
rect 5816 5568 5868 5574
rect 5816 5510 5868 5516
rect 5828 5137 5856 5510
rect 5920 5370 5948 6015
rect 6012 5778 6040 11070
rect 6092 11008 6144 11014
rect 6092 10950 6144 10956
rect 6000 5772 6052 5778
rect 6000 5714 6052 5720
rect 5908 5364 5960 5370
rect 5908 5306 5960 5312
rect 5906 5264 5962 5273
rect 5906 5199 5908 5208
rect 5960 5199 5962 5208
rect 5908 5170 5960 5176
rect 6012 5166 6040 5714
rect 6000 5160 6052 5166
rect 5814 5128 5870 5137
rect 6000 5102 6052 5108
rect 5814 5063 5870 5072
rect 6012 4758 6040 5102
rect 6000 4752 6052 4758
rect 6000 4694 6052 4700
rect 6012 4282 6040 4694
rect 6000 4276 6052 4282
rect 6000 4218 6052 4224
rect 6104 3534 6132 10950
rect 6184 10668 6236 10674
rect 6184 10610 6236 10616
rect 6196 10577 6224 10610
rect 6276 10600 6328 10606
rect 6182 10568 6238 10577
rect 6276 10542 6328 10548
rect 6182 10503 6238 10512
rect 6196 10198 6224 10503
rect 6184 10192 6236 10198
rect 6184 10134 6236 10140
rect 6288 10130 6316 10542
rect 6276 10124 6328 10130
rect 6276 10066 6328 10072
rect 6184 10056 6236 10062
rect 6184 9998 6236 10004
rect 6196 8022 6224 9998
rect 6472 9874 6500 11319
rect 6644 11212 6696 11218
rect 6644 11154 6696 11160
rect 6552 10464 6604 10470
rect 6552 10406 6604 10412
rect 6564 10062 6592 10406
rect 6552 10056 6604 10062
rect 6552 9998 6604 10004
rect 6472 9846 6592 9874
rect 6460 9716 6512 9722
rect 6380 9664 6460 9674
rect 6380 9658 6512 9664
rect 6380 9646 6500 9658
rect 6276 9172 6328 9178
rect 6276 9114 6328 9120
rect 6288 8294 6316 9114
rect 6276 8288 6328 8294
rect 6276 8230 6328 8236
rect 6184 8016 6236 8022
rect 6184 7958 6236 7964
rect 6184 7744 6236 7750
rect 6184 7686 6236 7692
rect 6276 7744 6328 7750
rect 6276 7686 6328 7692
rect 6196 7546 6224 7686
rect 6184 7540 6236 7546
rect 6184 7482 6236 7488
rect 6184 6452 6236 6458
rect 6184 6394 6236 6400
rect 6196 5778 6224 6394
rect 6184 5772 6236 5778
rect 6184 5714 6236 5720
rect 6184 5568 6236 5574
rect 6182 5536 6184 5545
rect 6236 5536 6238 5545
rect 6182 5471 6238 5480
rect 6196 4826 6224 5471
rect 6184 4820 6236 4826
rect 6184 4762 6236 4768
rect 6196 4146 6224 4762
rect 6184 4140 6236 4146
rect 6184 4082 6236 4088
rect 6092 3528 6144 3534
rect 6092 3470 6144 3476
rect 6288 3126 6316 7686
rect 6380 6322 6408 9646
rect 6564 9586 6592 9846
rect 6552 9580 6604 9586
rect 6552 9522 6604 9528
rect 6550 9480 6606 9489
rect 6460 9444 6512 9450
rect 6550 9415 6606 9424
rect 6460 9386 6512 9392
rect 6472 9081 6500 9386
rect 6458 9072 6514 9081
rect 6458 9007 6514 9016
rect 6460 8900 6512 8906
rect 6460 8842 6512 8848
rect 6472 7834 6500 8842
rect 6564 7954 6592 9415
rect 6656 9178 6684 11154
rect 6734 10296 6790 10305
rect 6734 10231 6790 10240
rect 6828 10260 6880 10266
rect 6748 9654 6776 10231
rect 6828 10202 6880 10208
rect 6736 9648 6788 9654
rect 6736 9590 6788 9596
rect 6840 9602 6868 10202
rect 6920 9920 6972 9926
rect 6920 9862 6972 9868
rect 6932 9761 6960 9862
rect 6918 9752 6974 9761
rect 6918 9687 6974 9696
rect 6748 9382 6776 9590
rect 6840 9574 6960 9602
rect 6932 9518 6960 9574
rect 6828 9512 6880 9518
rect 6828 9454 6880 9460
rect 6920 9512 6972 9518
rect 6920 9454 6972 9460
rect 6736 9376 6788 9382
rect 6736 9318 6788 9324
rect 6840 9178 6868 9454
rect 6644 9172 6696 9178
rect 6644 9114 6696 9120
rect 6828 9172 6880 9178
rect 6828 9114 6880 9120
rect 6734 9072 6790 9081
rect 6734 9007 6790 9016
rect 6920 9036 6972 9042
rect 6644 8832 6696 8838
rect 6642 8800 6644 8809
rect 6696 8800 6698 8809
rect 6642 8735 6698 8744
rect 6552 7948 6604 7954
rect 6552 7890 6604 7896
rect 6472 7806 6592 7834
rect 6458 7440 6514 7449
rect 6458 7375 6514 7384
rect 6472 7002 6500 7375
rect 6460 6996 6512 7002
rect 6460 6938 6512 6944
rect 6472 6905 6500 6938
rect 6458 6896 6514 6905
rect 6458 6831 6514 6840
rect 6460 6656 6512 6662
rect 6460 6598 6512 6604
rect 6368 6316 6420 6322
rect 6368 6258 6420 6264
rect 6380 4826 6408 6258
rect 6472 5914 6500 6598
rect 6460 5908 6512 5914
rect 6460 5850 6512 5856
rect 6460 5704 6512 5710
rect 6460 5646 6512 5652
rect 6472 5370 6500 5646
rect 6460 5364 6512 5370
rect 6460 5306 6512 5312
rect 6458 5264 6514 5273
rect 6458 5199 6514 5208
rect 6368 4820 6420 4826
rect 6368 4762 6420 4768
rect 6472 4622 6500 5199
rect 6460 4616 6512 4622
rect 6460 4558 6512 4564
rect 6564 3194 6592 7806
rect 6644 7336 6696 7342
rect 6644 7278 6696 7284
rect 6656 6458 6684 7278
rect 6748 6905 6776 9007
rect 6920 8978 6972 8984
rect 6828 8968 6880 8974
rect 6828 8910 6880 8916
rect 6840 8673 6868 8910
rect 6826 8664 6882 8673
rect 6826 8599 6882 8608
rect 6932 8430 6960 8978
rect 7024 8566 7052 12406
rect 7196 11756 7248 11762
rect 7196 11698 7248 11704
rect 7208 11354 7236 11698
rect 7196 11348 7248 11354
rect 7196 11290 7248 11296
rect 7194 10840 7250 10849
rect 7194 10775 7250 10784
rect 7104 10668 7156 10674
rect 7104 10610 7156 10616
rect 7012 8560 7064 8566
rect 7012 8502 7064 8508
rect 6920 8424 6972 8430
rect 6920 8366 6972 8372
rect 6932 7478 6960 8366
rect 6920 7472 6972 7478
rect 6920 7414 6972 7420
rect 6828 7404 6880 7410
rect 6828 7346 6880 7352
rect 6734 6896 6790 6905
rect 6734 6831 6790 6840
rect 6736 6792 6788 6798
rect 6736 6734 6788 6740
rect 6644 6452 6696 6458
rect 6644 6394 6696 6400
rect 6642 6352 6698 6361
rect 6642 6287 6698 6296
rect 6656 6186 6684 6287
rect 6644 6180 6696 6186
rect 6644 6122 6696 6128
rect 6748 5098 6776 6734
rect 6840 6458 6868 7346
rect 6920 7336 6972 7342
rect 6920 7278 6972 7284
rect 6932 6798 6960 7278
rect 7012 7268 7064 7274
rect 7012 7210 7064 7216
rect 6920 6792 6972 6798
rect 6920 6734 6972 6740
rect 6828 6452 6880 6458
rect 6828 6394 6880 6400
rect 6920 6112 6972 6118
rect 6920 6054 6972 6060
rect 6828 5636 6880 5642
rect 6828 5578 6880 5584
rect 6840 5545 6868 5578
rect 6826 5536 6882 5545
rect 6826 5471 6882 5480
rect 6736 5092 6788 5098
rect 6736 5034 6788 5040
rect 6644 4480 6696 4486
rect 6644 4422 6696 4428
rect 6552 3188 6604 3194
rect 6552 3130 6604 3136
rect 6276 3120 6328 3126
rect 6276 3062 6328 3068
rect 6656 3058 6684 4422
rect 6840 3398 6868 5471
rect 6932 5302 6960 6054
rect 7024 5370 7052 7210
rect 7116 6662 7144 10610
rect 7208 10606 7236 10775
rect 7196 10600 7248 10606
rect 7196 10542 7248 10548
rect 7196 10260 7248 10266
rect 7196 10202 7248 10208
rect 7208 9042 7236 10202
rect 7300 10130 7328 13942
rect 8128 13870 8156 14010
rect 8208 13932 8260 13938
rect 8208 13874 8260 13880
rect 8116 13864 8168 13870
rect 8116 13806 8168 13812
rect 7622 13628 7930 13637
rect 7622 13626 7628 13628
rect 7684 13626 7708 13628
rect 7764 13626 7788 13628
rect 7844 13626 7868 13628
rect 7924 13626 7930 13628
rect 7684 13574 7686 13626
rect 7866 13574 7868 13626
rect 7622 13572 7628 13574
rect 7684 13572 7708 13574
rect 7764 13572 7788 13574
rect 7844 13572 7868 13574
rect 7924 13572 7930 13574
rect 7622 13563 7930 13572
rect 8128 13326 8156 13806
rect 8220 13410 8248 13874
rect 8496 13433 8524 14418
rect 8588 14006 8616 14758
rect 9968 14618 9996 16400
rect 11796 14952 11848 14958
rect 11796 14894 11848 14900
rect 11520 14884 11572 14890
rect 11520 14826 11572 14832
rect 9956 14612 10008 14618
rect 9956 14554 10008 14560
rect 8760 14476 8812 14482
rect 8760 14418 8812 14424
rect 11336 14476 11388 14482
rect 11336 14418 11388 14424
rect 8772 14385 8800 14418
rect 10232 14408 10284 14414
rect 8758 14376 8814 14385
rect 10232 14350 10284 14356
rect 8758 14311 8814 14320
rect 8760 14272 8812 14278
rect 8680 14232 8760 14260
rect 8576 14000 8628 14006
rect 8576 13942 8628 13948
rect 8482 13424 8538 13433
rect 8220 13382 8432 13410
rect 8116 13320 8168 13326
rect 8116 13262 8168 13268
rect 7380 13184 7432 13190
rect 7380 13126 7432 13132
rect 7472 13184 7524 13190
rect 7472 13126 7524 13132
rect 7392 12646 7420 13126
rect 7484 12782 7512 13126
rect 8128 12918 8156 13262
rect 8116 12912 8168 12918
rect 8116 12854 8168 12860
rect 7472 12776 7524 12782
rect 7472 12718 7524 12724
rect 7380 12640 7432 12646
rect 7380 12582 7432 12588
rect 7380 11348 7432 11354
rect 7380 11290 7432 11296
rect 7392 10606 7420 11290
rect 7380 10600 7432 10606
rect 7380 10542 7432 10548
rect 7288 10124 7340 10130
rect 7288 10066 7340 10072
rect 7300 9110 7328 10066
rect 7392 10062 7420 10542
rect 7484 10112 7512 12718
rect 7622 12540 7930 12549
rect 7622 12538 7628 12540
rect 7684 12538 7708 12540
rect 7764 12538 7788 12540
rect 7844 12538 7868 12540
rect 7924 12538 7930 12540
rect 7684 12486 7686 12538
rect 7866 12486 7868 12538
rect 7622 12484 7628 12486
rect 7684 12484 7708 12486
rect 7764 12484 7788 12486
rect 7844 12484 7868 12486
rect 7924 12484 7930 12486
rect 7622 12475 7930 12484
rect 8128 11830 8156 12854
rect 8404 12374 8432 13382
rect 8482 13359 8538 13368
rect 8484 13252 8536 13258
rect 8484 13194 8536 13200
rect 8496 12617 8524 13194
rect 8482 12608 8538 12617
rect 8482 12543 8538 12552
rect 8576 12436 8628 12442
rect 8576 12378 8628 12384
rect 8392 12368 8444 12374
rect 8588 12345 8616 12378
rect 8392 12310 8444 12316
rect 8574 12336 8630 12345
rect 8208 12300 8260 12306
rect 8574 12271 8630 12280
rect 8208 12242 8260 12248
rect 8220 11830 8248 12242
rect 8588 11898 8616 12271
rect 8300 11892 8352 11898
rect 8300 11834 8352 11840
rect 8576 11892 8628 11898
rect 8576 11834 8628 11840
rect 8116 11824 8168 11830
rect 8116 11766 8168 11772
rect 8208 11824 8260 11830
rect 8208 11766 8260 11772
rect 7622 11452 7930 11461
rect 7622 11450 7628 11452
rect 7684 11450 7708 11452
rect 7764 11450 7788 11452
rect 7844 11450 7868 11452
rect 7924 11450 7930 11452
rect 7684 11398 7686 11450
rect 7866 11398 7868 11450
rect 7622 11396 7628 11398
rect 7684 11396 7708 11398
rect 7764 11396 7788 11398
rect 7844 11396 7868 11398
rect 7924 11396 7930 11398
rect 7622 11387 7930 11396
rect 8116 11348 8168 11354
rect 8116 11290 8168 11296
rect 7622 10364 7930 10373
rect 7622 10362 7628 10364
rect 7684 10362 7708 10364
rect 7764 10362 7788 10364
rect 7844 10362 7868 10364
rect 7924 10362 7930 10364
rect 7684 10310 7686 10362
rect 7866 10310 7868 10362
rect 7622 10308 7628 10310
rect 7684 10308 7708 10310
rect 7764 10308 7788 10310
rect 7844 10308 7868 10310
rect 7924 10308 7930 10310
rect 7622 10299 7930 10308
rect 7484 10084 7604 10112
rect 7380 10056 7432 10062
rect 7380 9998 7432 10004
rect 7392 9586 7420 9998
rect 7472 9988 7524 9994
rect 7472 9930 7524 9936
rect 7380 9580 7432 9586
rect 7380 9522 7432 9528
rect 7288 9104 7340 9110
rect 7288 9046 7340 9052
rect 7196 9036 7248 9042
rect 7196 8978 7248 8984
rect 7392 8974 7420 9522
rect 7380 8968 7432 8974
rect 7380 8910 7432 8916
rect 7288 8560 7340 8566
rect 7288 8502 7340 8508
rect 7196 8492 7248 8498
rect 7196 8434 7248 8440
rect 7208 8129 7236 8434
rect 7194 8120 7250 8129
rect 7194 8055 7250 8064
rect 7196 8016 7248 8022
rect 7196 7958 7248 7964
rect 7104 6656 7156 6662
rect 7104 6598 7156 6604
rect 7102 5400 7158 5409
rect 7012 5364 7064 5370
rect 7102 5335 7158 5344
rect 7012 5306 7064 5312
rect 6920 5296 6972 5302
rect 6920 5238 6972 5244
rect 7116 5166 7144 5335
rect 6920 5160 6972 5166
rect 6920 5102 6972 5108
rect 7104 5160 7156 5166
rect 7104 5102 7156 5108
rect 6932 4554 6960 5102
rect 7104 5024 7156 5030
rect 7104 4966 7156 4972
rect 7116 4865 7144 4966
rect 7102 4856 7158 4865
rect 7102 4791 7158 4800
rect 6920 4548 6972 4554
rect 6920 4490 6972 4496
rect 7012 4480 7064 4486
rect 7012 4422 7064 4428
rect 7104 4480 7156 4486
rect 7104 4422 7156 4428
rect 6918 4312 6974 4321
rect 7024 4282 7052 4422
rect 6918 4247 6974 4256
rect 7012 4276 7064 4282
rect 6932 4214 6960 4247
rect 7012 4218 7064 4224
rect 6920 4208 6972 4214
rect 6920 4150 6972 4156
rect 7116 4010 7144 4422
rect 7104 4004 7156 4010
rect 7104 3946 7156 3952
rect 7208 3534 7236 7958
rect 7300 7546 7328 8502
rect 7484 8362 7512 9930
rect 7576 9450 7604 10084
rect 7656 10056 7708 10062
rect 7656 9998 7708 10004
rect 7668 9722 7696 9998
rect 7656 9716 7708 9722
rect 7656 9658 7708 9664
rect 8024 9580 8076 9586
rect 8024 9522 8076 9528
rect 7564 9444 7616 9450
rect 7564 9386 7616 9392
rect 7622 9276 7930 9285
rect 7622 9274 7628 9276
rect 7684 9274 7708 9276
rect 7764 9274 7788 9276
rect 7844 9274 7868 9276
rect 7924 9274 7930 9276
rect 7684 9222 7686 9274
rect 7866 9222 7868 9274
rect 7622 9220 7628 9222
rect 7684 9220 7708 9222
rect 7764 9220 7788 9222
rect 7844 9220 7868 9222
rect 7924 9220 7930 9222
rect 7622 9211 7930 9220
rect 8036 8974 8064 9522
rect 8128 9518 8156 11290
rect 8116 9512 8168 9518
rect 8116 9454 8168 9460
rect 8024 8968 8076 8974
rect 8024 8910 8076 8916
rect 8022 8664 8078 8673
rect 8022 8599 8024 8608
rect 8076 8599 8078 8608
rect 8024 8570 8076 8576
rect 7748 8492 7800 8498
rect 7748 8434 7800 8440
rect 7472 8356 7524 8362
rect 7472 8298 7524 8304
rect 7760 8294 7788 8434
rect 8128 8430 8156 9454
rect 8220 9450 8248 11766
rect 8312 9586 8340 11834
rect 8392 9920 8444 9926
rect 8392 9862 8444 9868
rect 8404 9722 8432 9862
rect 8392 9716 8444 9722
rect 8392 9658 8444 9664
rect 8300 9580 8352 9586
rect 8300 9522 8352 9528
rect 8208 9444 8260 9450
rect 8208 9386 8260 9392
rect 8404 9160 8432 9658
rect 8576 9376 8628 9382
rect 8576 9318 8628 9324
rect 8220 9132 8432 9160
rect 8024 8424 8076 8430
rect 8116 8424 8168 8430
rect 8024 8366 8076 8372
rect 8114 8392 8116 8401
rect 8168 8392 8170 8401
rect 7748 8288 7800 8294
rect 7748 8230 7800 8236
rect 7622 8188 7930 8197
rect 7622 8186 7628 8188
rect 7684 8186 7708 8188
rect 7764 8186 7788 8188
rect 7844 8186 7868 8188
rect 7924 8186 7930 8188
rect 7684 8134 7686 8186
rect 7866 8134 7868 8186
rect 7622 8132 7628 8134
rect 7684 8132 7708 8134
rect 7764 8132 7788 8134
rect 7844 8132 7868 8134
rect 7924 8132 7930 8134
rect 7622 8123 7930 8132
rect 7748 7948 7800 7954
rect 7748 7890 7800 7896
rect 7472 7744 7524 7750
rect 7472 7686 7524 7692
rect 7288 7540 7340 7546
rect 7288 7482 7340 7488
rect 7380 7336 7432 7342
rect 7300 7296 7380 7324
rect 7300 6186 7328 7296
rect 7380 7278 7432 7284
rect 7484 7002 7512 7686
rect 7760 7274 7788 7890
rect 7932 7540 7984 7546
rect 8036 7528 8064 8366
rect 8114 8327 8170 8336
rect 8114 8256 8170 8265
rect 8114 8191 8170 8200
rect 8128 7954 8156 8191
rect 8116 7948 8168 7954
rect 8116 7890 8168 7896
rect 8116 7744 8168 7750
rect 8116 7686 8168 7692
rect 8128 7546 8156 7686
rect 7984 7500 8064 7528
rect 8116 7540 8168 7546
rect 7932 7482 7984 7488
rect 8116 7482 8168 7488
rect 7748 7268 7800 7274
rect 7748 7210 7800 7216
rect 7622 7100 7930 7109
rect 7622 7098 7628 7100
rect 7684 7098 7708 7100
rect 7764 7098 7788 7100
rect 7844 7098 7868 7100
rect 7924 7098 7930 7100
rect 7684 7046 7686 7098
rect 7866 7046 7868 7098
rect 7622 7044 7628 7046
rect 7684 7044 7708 7046
rect 7764 7044 7788 7046
rect 7844 7044 7868 7046
rect 7924 7044 7930 7046
rect 7622 7035 7930 7044
rect 7472 6996 7524 7002
rect 7472 6938 7524 6944
rect 7380 6928 7432 6934
rect 7380 6870 7432 6876
rect 7746 6896 7802 6905
rect 7392 6254 7420 6870
rect 7746 6831 7748 6840
rect 7800 6831 7802 6840
rect 7748 6802 7800 6808
rect 7840 6792 7892 6798
rect 7840 6734 7892 6740
rect 7470 6488 7526 6497
rect 7470 6423 7526 6432
rect 7484 6390 7512 6423
rect 7472 6384 7524 6390
rect 7472 6326 7524 6332
rect 7380 6248 7432 6254
rect 7380 6190 7432 6196
rect 7288 6180 7340 6186
rect 7288 6122 7340 6128
rect 7392 6118 7420 6190
rect 7380 6112 7432 6118
rect 7380 6054 7432 6060
rect 7484 5896 7512 6326
rect 7852 6254 7880 6734
rect 8024 6656 8076 6662
rect 8024 6598 8076 6604
rect 8036 6361 8064 6598
rect 8022 6352 8078 6361
rect 8022 6287 8078 6296
rect 7840 6248 7892 6254
rect 7840 6190 7892 6196
rect 7622 6012 7930 6021
rect 7622 6010 7628 6012
rect 7684 6010 7708 6012
rect 7764 6010 7788 6012
rect 7844 6010 7868 6012
rect 7924 6010 7930 6012
rect 7684 5958 7686 6010
rect 7866 5958 7868 6010
rect 7622 5956 7628 5958
rect 7684 5956 7708 5958
rect 7764 5956 7788 5958
rect 7844 5956 7868 5958
rect 7924 5956 7930 5958
rect 7622 5947 7930 5956
rect 7484 5868 7604 5896
rect 7286 5672 7342 5681
rect 7286 5607 7342 5616
rect 7300 5370 7328 5607
rect 7472 5568 7524 5574
rect 7472 5510 7524 5516
rect 7288 5364 7340 5370
rect 7288 5306 7340 5312
rect 7484 5216 7512 5510
rect 7300 5188 7512 5216
rect 7196 3528 7248 3534
rect 7196 3470 7248 3476
rect 6828 3392 6880 3398
rect 6828 3334 6880 3340
rect 7300 3058 7328 5188
rect 7576 5114 7604 5868
rect 8036 5846 8064 6287
rect 8116 6248 8168 6254
rect 8116 6190 8168 6196
rect 8024 5840 8076 5846
rect 8024 5782 8076 5788
rect 7840 5704 7892 5710
rect 7840 5646 7892 5652
rect 7852 5370 7880 5646
rect 8024 5568 8076 5574
rect 8024 5510 8076 5516
rect 8128 5522 8156 6190
rect 8220 5778 8248 9132
rect 8392 9036 8444 9042
rect 8392 8978 8444 8984
rect 8404 8838 8432 8978
rect 8484 8900 8536 8906
rect 8484 8842 8536 8848
rect 8392 8832 8444 8838
rect 8392 8774 8444 8780
rect 8392 8492 8444 8498
rect 8392 8434 8444 8440
rect 8404 7818 8432 8434
rect 8496 8362 8524 8842
rect 8484 8356 8536 8362
rect 8484 8298 8536 8304
rect 8496 8090 8524 8298
rect 8484 8084 8536 8090
rect 8484 8026 8536 8032
rect 8392 7812 8444 7818
rect 8392 7754 8444 7760
rect 8484 7812 8536 7818
rect 8484 7754 8536 7760
rect 8300 7744 8352 7750
rect 8300 7686 8352 7692
rect 8312 7546 8340 7686
rect 8300 7540 8352 7546
rect 8300 7482 8352 7488
rect 8300 7336 8352 7342
rect 8300 7278 8352 7284
rect 8312 6798 8340 7278
rect 8300 6792 8352 6798
rect 8300 6734 8352 6740
rect 8404 6202 8432 7754
rect 8496 7410 8524 7754
rect 8484 7404 8536 7410
rect 8484 7346 8536 7352
rect 8484 7268 8536 7274
rect 8484 7210 8536 7216
rect 8496 6916 8524 7210
rect 8588 7041 8616 9318
rect 8680 8265 8708 14232
rect 8760 14214 8812 14220
rect 9128 14272 9180 14278
rect 9128 14214 9180 14220
rect 8758 13288 8814 13297
rect 8758 13223 8814 13232
rect 8772 9042 8800 13223
rect 8852 12844 8904 12850
rect 8852 12786 8904 12792
rect 8864 11257 8892 12786
rect 9140 12434 9168 14214
rect 9846 14172 10154 14181
rect 9846 14170 9852 14172
rect 9908 14170 9932 14172
rect 9988 14170 10012 14172
rect 10068 14170 10092 14172
rect 10148 14170 10154 14172
rect 9908 14118 9910 14170
rect 10090 14118 10092 14170
rect 9846 14116 9852 14118
rect 9908 14116 9932 14118
rect 9988 14116 10012 14118
rect 10068 14116 10092 14118
rect 10148 14116 10154 14118
rect 9846 14107 10154 14116
rect 9772 14068 9824 14074
rect 9772 14010 9824 14016
rect 9312 14000 9364 14006
rect 9312 13942 9364 13948
rect 9220 13320 9272 13326
rect 9220 13262 9272 13268
rect 9048 12406 9168 12434
rect 8942 12336 8998 12345
rect 8942 12271 8998 12280
rect 8956 12073 8984 12271
rect 8942 12064 8998 12073
rect 8942 11999 8998 12008
rect 8944 11280 8996 11286
rect 8850 11248 8906 11257
rect 8944 11222 8996 11228
rect 8850 11183 8906 11192
rect 8956 11121 8984 11222
rect 8942 11112 8998 11121
rect 8942 11047 8998 11056
rect 8850 10568 8906 10577
rect 8850 10503 8906 10512
rect 8760 9036 8812 9042
rect 8760 8978 8812 8984
rect 8760 8832 8812 8838
rect 8760 8774 8812 8780
rect 8772 8537 8800 8774
rect 8758 8528 8814 8537
rect 8758 8463 8814 8472
rect 8666 8256 8722 8265
rect 8666 8191 8722 8200
rect 8668 7948 8720 7954
rect 8668 7890 8720 7896
rect 8680 7342 8708 7890
rect 8864 7818 8892 10503
rect 8944 10124 8996 10130
rect 8944 10066 8996 10072
rect 8956 8945 8984 10066
rect 8942 8936 8998 8945
rect 8942 8871 8998 8880
rect 8956 8090 8984 8871
rect 8944 8084 8996 8090
rect 8944 8026 8996 8032
rect 8852 7812 8904 7818
rect 8852 7754 8904 7760
rect 8760 7744 8812 7750
rect 9048 7698 9076 12406
rect 9232 12238 9260 13262
rect 9220 12232 9272 12238
rect 9220 12174 9272 12180
rect 9220 11756 9272 11762
rect 9220 11698 9272 11704
rect 9232 11218 9260 11698
rect 9220 11212 9272 11218
rect 9220 11154 9272 11160
rect 9324 10826 9352 13942
rect 9496 13864 9548 13870
rect 9496 13806 9548 13812
rect 9404 13524 9456 13530
rect 9404 13466 9456 13472
rect 9416 12850 9444 13466
rect 9404 12844 9456 12850
rect 9404 12786 9456 12792
rect 9416 12753 9444 12786
rect 9402 12744 9458 12753
rect 9402 12679 9458 12688
rect 9404 11076 9456 11082
rect 9404 11018 9456 11024
rect 9232 10798 9352 10826
rect 9416 10810 9444 11018
rect 9404 10804 9456 10810
rect 9128 10464 9180 10470
rect 9128 10406 9180 10412
rect 9140 8945 9168 10406
rect 9232 10062 9260 10798
rect 9404 10746 9456 10752
rect 9312 10736 9364 10742
rect 9312 10678 9364 10684
rect 9220 10056 9272 10062
rect 9220 9998 9272 10004
rect 9218 9888 9274 9897
rect 9218 9823 9274 9832
rect 9126 8936 9182 8945
rect 9126 8871 9182 8880
rect 9128 8288 9180 8294
rect 9128 8230 9180 8236
rect 9140 8090 9168 8230
rect 9128 8084 9180 8090
rect 9128 8026 9180 8032
rect 8760 7686 8812 7692
rect 8668 7336 8720 7342
rect 8668 7278 8720 7284
rect 8574 7032 8630 7041
rect 8574 6967 8630 6976
rect 8680 6934 8708 7278
rect 8668 6928 8720 6934
rect 8496 6888 8616 6916
rect 8484 6316 8536 6322
rect 8484 6258 8536 6264
rect 8312 6174 8432 6202
rect 8312 5914 8340 6174
rect 8392 6112 8444 6118
rect 8392 6054 8444 6060
rect 8300 5908 8352 5914
rect 8300 5850 8352 5856
rect 8208 5772 8260 5778
rect 8208 5714 8260 5720
rect 8298 5672 8354 5681
rect 8298 5607 8300 5616
rect 8352 5607 8354 5616
rect 8300 5578 8352 5584
rect 8036 5370 8064 5510
rect 8128 5494 8340 5522
rect 7840 5364 7892 5370
rect 7840 5306 7892 5312
rect 8024 5364 8076 5370
rect 8024 5306 8076 5312
rect 8024 5228 8076 5234
rect 8024 5170 8076 5176
rect 7484 5086 7604 5114
rect 7484 4865 7512 5086
rect 7622 4924 7930 4933
rect 7622 4922 7628 4924
rect 7684 4922 7708 4924
rect 7764 4922 7788 4924
rect 7844 4922 7868 4924
rect 7924 4922 7930 4924
rect 7684 4870 7686 4922
rect 7866 4870 7868 4922
rect 7622 4868 7628 4870
rect 7684 4868 7708 4870
rect 7764 4868 7788 4870
rect 7844 4868 7868 4870
rect 7924 4868 7930 4870
rect 7470 4856 7526 4865
rect 7622 4859 7930 4868
rect 7470 4791 7526 4800
rect 8036 4690 8064 5170
rect 8116 5160 8168 5166
rect 8116 5102 8168 5108
rect 8208 5160 8260 5166
rect 8208 5102 8260 5108
rect 8312 5114 8340 5494
rect 8404 5302 8432 6054
rect 8496 5914 8524 6258
rect 8484 5908 8536 5914
rect 8484 5850 8536 5856
rect 8588 5710 8616 6888
rect 8668 6870 8720 6876
rect 8772 6866 8800 7686
rect 8956 7670 9076 7698
rect 8850 7440 8906 7449
rect 8850 7375 8852 7384
rect 8904 7375 8906 7384
rect 8852 7346 8904 7352
rect 8760 6860 8812 6866
rect 8760 6802 8812 6808
rect 8956 6798 8984 7670
rect 9036 7540 9088 7546
rect 9036 7482 9088 7488
rect 8944 6792 8996 6798
rect 8944 6734 8996 6740
rect 8944 6656 8996 6662
rect 8944 6598 8996 6604
rect 8956 6458 8984 6598
rect 8944 6452 8996 6458
rect 8944 6394 8996 6400
rect 8852 6316 8904 6322
rect 8852 6258 8904 6264
rect 8760 6248 8812 6254
rect 8760 6190 8812 6196
rect 8484 5704 8536 5710
rect 8484 5646 8536 5652
rect 8576 5704 8628 5710
rect 8576 5646 8628 5652
rect 8496 5545 8524 5646
rect 8482 5536 8538 5545
rect 8482 5471 8538 5480
rect 8392 5296 8444 5302
rect 8392 5238 8444 5244
rect 8024 4684 8076 4690
rect 8024 4626 8076 4632
rect 7380 4480 7432 4486
rect 7380 4422 7432 4428
rect 7470 4448 7526 4457
rect 7392 4282 7420 4422
rect 7470 4383 7526 4392
rect 7484 4282 7512 4383
rect 7380 4276 7432 4282
rect 7380 4218 7432 4224
rect 7472 4276 7524 4282
rect 7472 4218 7524 4224
rect 7470 4176 7526 4185
rect 7470 4111 7526 4120
rect 7484 3602 7512 4111
rect 8128 3942 8156 5102
rect 8220 4826 8248 5102
rect 8312 5086 8432 5114
rect 8300 5024 8352 5030
rect 8300 4966 8352 4972
rect 8208 4820 8260 4826
rect 8208 4762 8260 4768
rect 8312 4457 8340 4966
rect 8404 4486 8432 5086
rect 8772 4826 8800 6190
rect 8864 5370 8892 6258
rect 9048 6118 9076 7482
rect 9232 7018 9260 9823
rect 9324 9674 9352 10678
rect 9416 9926 9444 10746
rect 9404 9920 9456 9926
rect 9404 9862 9456 9868
rect 9324 9646 9444 9674
rect 9416 9586 9444 9646
rect 9404 9580 9456 9586
rect 9404 9522 9456 9528
rect 9310 9344 9366 9353
rect 9310 9279 9366 9288
rect 9324 7585 9352 9279
rect 9508 7970 9536 13806
rect 9588 13728 9640 13734
rect 9588 13670 9640 13676
rect 9600 11082 9628 13670
rect 9680 12912 9732 12918
rect 9678 12880 9680 12889
rect 9732 12880 9734 12889
rect 9678 12815 9734 12824
rect 9692 11898 9720 12815
rect 9680 11892 9732 11898
rect 9680 11834 9732 11840
rect 9680 11144 9732 11150
rect 9680 11086 9732 11092
rect 9588 11076 9640 11082
rect 9588 11018 9640 11024
rect 9586 10840 9642 10849
rect 9586 10775 9588 10784
rect 9640 10775 9642 10784
rect 9588 10746 9640 10752
rect 9692 10742 9720 11086
rect 9680 10736 9732 10742
rect 9680 10678 9732 10684
rect 9692 10044 9720 10678
rect 9784 10538 9812 14010
rect 9846 13084 10154 13093
rect 9846 13082 9852 13084
rect 9908 13082 9932 13084
rect 9988 13082 10012 13084
rect 10068 13082 10092 13084
rect 10148 13082 10154 13084
rect 9908 13030 9910 13082
rect 10090 13030 10092 13082
rect 9846 13028 9852 13030
rect 9908 13028 9932 13030
rect 9988 13028 10012 13030
rect 10068 13028 10092 13030
rect 10148 13028 10154 13030
rect 9846 13019 10154 13028
rect 10244 12889 10272 14350
rect 11348 13938 11376 14418
rect 11532 14278 11560 14826
rect 11520 14272 11572 14278
rect 11520 14214 11572 14220
rect 11060 13932 11112 13938
rect 11060 13874 11112 13880
rect 11336 13932 11388 13938
rect 11336 13874 11388 13880
rect 10784 13184 10836 13190
rect 11072 13172 11100 13874
rect 11348 13308 11376 13874
rect 11704 13728 11756 13734
rect 11704 13670 11756 13676
rect 11520 13320 11572 13326
rect 11348 13280 11520 13308
rect 11072 13144 11192 13172
rect 10784 13126 10836 13132
rect 10230 12880 10286 12889
rect 10230 12815 10286 12824
rect 9846 11996 10154 12005
rect 9846 11994 9852 11996
rect 9908 11994 9932 11996
rect 9988 11994 10012 11996
rect 10068 11994 10092 11996
rect 10148 11994 10154 11996
rect 9908 11942 9910 11994
rect 10090 11942 10092 11994
rect 9846 11940 9852 11942
rect 9908 11940 9932 11942
rect 9988 11940 10012 11942
rect 10068 11940 10092 11942
rect 10148 11940 10154 11942
rect 9846 11931 10154 11940
rect 9846 10908 10154 10917
rect 9846 10906 9852 10908
rect 9908 10906 9932 10908
rect 9988 10906 10012 10908
rect 10068 10906 10092 10908
rect 10148 10906 10154 10908
rect 9908 10854 9910 10906
rect 10090 10854 10092 10906
rect 9846 10852 9852 10854
rect 9908 10852 9932 10854
rect 9988 10852 10012 10854
rect 10068 10852 10092 10854
rect 10148 10852 10154 10854
rect 9846 10843 10154 10852
rect 10244 10849 10272 12815
rect 10600 12708 10652 12714
rect 10600 12650 10652 12656
rect 10416 11008 10468 11014
rect 10416 10950 10468 10956
rect 10230 10840 10286 10849
rect 10230 10775 10286 10784
rect 10428 10554 10456 10950
rect 10612 10674 10640 12650
rect 10692 12232 10744 12238
rect 10692 12174 10744 12180
rect 10600 10668 10652 10674
rect 10600 10610 10652 10616
rect 9772 10532 9824 10538
rect 9772 10474 9824 10480
rect 9968 10526 10456 10554
rect 9784 10146 9812 10474
rect 9784 10118 9904 10146
rect 9968 10130 9996 10526
rect 10416 10464 10468 10470
rect 10046 10432 10102 10441
rect 10416 10406 10468 10412
rect 10598 10432 10654 10441
rect 10046 10367 10102 10376
rect 9772 10056 9824 10062
rect 9646 10016 9772 10044
rect 9646 9738 9674 10016
rect 9772 9998 9824 10004
rect 9876 9994 9904 10118
rect 9956 10124 10008 10130
rect 9956 10066 10008 10072
rect 9864 9988 9916 9994
rect 9864 9930 9916 9936
rect 9956 9920 10008 9926
rect 10060 9908 10088 10367
rect 10008 9880 10088 9908
rect 10230 9888 10286 9897
rect 9956 9862 10008 9868
rect 9846 9820 10154 9829
rect 10230 9823 10286 9832
rect 9846 9818 9852 9820
rect 9908 9818 9932 9820
rect 9988 9818 10012 9820
rect 10068 9818 10092 9820
rect 10148 9818 10154 9820
rect 9908 9766 9910 9818
rect 10090 9766 10092 9818
rect 9846 9764 9852 9766
rect 9908 9764 9932 9766
rect 9988 9764 10012 9766
rect 10068 9764 10092 9766
rect 10148 9764 10154 9766
rect 9846 9755 10154 9764
rect 9646 9710 9812 9738
rect 9784 9654 9812 9710
rect 9772 9648 9824 9654
rect 9678 9616 9734 9625
rect 9772 9590 9824 9596
rect 9864 9648 9916 9654
rect 9864 9590 9916 9596
rect 9678 9551 9734 9560
rect 9692 9518 9720 9551
rect 9680 9512 9732 9518
rect 9680 9454 9732 9460
rect 9680 8900 9732 8906
rect 9680 8842 9732 8848
rect 9588 8832 9640 8838
rect 9588 8774 9640 8780
rect 9416 7942 9536 7970
rect 9310 7576 9366 7585
rect 9416 7546 9444 7942
rect 9496 7880 9548 7886
rect 9496 7822 9548 7828
rect 9310 7511 9366 7520
rect 9404 7540 9456 7546
rect 9404 7482 9456 7488
rect 9312 7472 9364 7478
rect 9312 7414 9364 7420
rect 9140 6990 9260 7018
rect 9140 6798 9168 6990
rect 9218 6896 9274 6905
rect 9218 6831 9274 6840
rect 9128 6792 9180 6798
rect 9128 6734 9180 6740
rect 9128 6656 9180 6662
rect 9128 6598 9180 6604
rect 9036 6112 9088 6118
rect 9036 6054 9088 6060
rect 9048 5778 9076 6054
rect 9036 5772 9088 5778
rect 9036 5714 9088 5720
rect 8944 5704 8996 5710
rect 8942 5672 8944 5681
rect 8996 5672 8998 5681
rect 8942 5607 8998 5616
rect 9036 5568 9088 5574
rect 9036 5510 9088 5516
rect 8852 5364 8904 5370
rect 8852 5306 8904 5312
rect 9048 5234 9076 5510
rect 9036 5228 9088 5234
rect 9036 5170 9088 5176
rect 9140 5001 9168 6598
rect 9232 5778 9260 6831
rect 9324 6118 9352 7414
rect 9404 7336 9456 7342
rect 9404 7278 9456 7284
rect 9416 6322 9444 7278
rect 9508 7002 9536 7822
rect 9496 6996 9548 7002
rect 9496 6938 9548 6944
rect 9600 6882 9628 8774
rect 9692 7818 9720 8842
rect 9784 8480 9812 9590
rect 9876 8838 9904 9590
rect 10048 9580 10100 9586
rect 10048 9522 10100 9528
rect 9956 9376 10008 9382
rect 9954 9344 9956 9353
rect 10008 9344 10010 9353
rect 9954 9279 10010 9288
rect 10060 9217 10088 9522
rect 10046 9208 10102 9217
rect 10046 9143 10102 9152
rect 10244 9110 10272 9823
rect 10322 9752 10378 9761
rect 10322 9687 10378 9696
rect 10232 9104 10284 9110
rect 10232 9046 10284 9052
rect 9864 8832 9916 8838
rect 9864 8774 9916 8780
rect 9846 8732 10154 8741
rect 9846 8730 9852 8732
rect 9908 8730 9932 8732
rect 9988 8730 10012 8732
rect 10068 8730 10092 8732
rect 10148 8730 10154 8732
rect 9908 8678 9910 8730
rect 10090 8678 10092 8730
rect 9846 8676 9852 8678
rect 9908 8676 9932 8678
rect 9988 8676 10012 8678
rect 10068 8676 10092 8678
rect 10148 8676 10154 8678
rect 9846 8667 10154 8676
rect 9864 8492 9916 8498
rect 9784 8452 9864 8480
rect 9784 7886 9812 8452
rect 9864 8434 9916 8440
rect 10048 8492 10100 8498
rect 10048 8434 10100 8440
rect 9862 8392 9918 8401
rect 9862 8327 9864 8336
rect 9916 8327 9918 8336
rect 9864 8298 9916 8304
rect 9772 7880 9824 7886
rect 10060 7857 10088 8434
rect 9772 7822 9824 7828
rect 10046 7848 10102 7857
rect 9680 7812 9732 7818
rect 10046 7783 10102 7792
rect 9680 7754 9732 7760
rect 9692 7528 9720 7754
rect 9846 7644 10154 7653
rect 9846 7642 9852 7644
rect 9908 7642 9932 7644
rect 9988 7642 10012 7644
rect 10068 7642 10092 7644
rect 10148 7642 10154 7644
rect 9908 7590 9910 7642
rect 10090 7590 10092 7642
rect 9846 7588 9852 7590
rect 9908 7588 9932 7590
rect 9988 7588 10012 7590
rect 10068 7588 10092 7590
rect 10148 7588 10154 7590
rect 9846 7579 10154 7588
rect 9692 7500 9996 7528
rect 9864 7404 9916 7410
rect 9864 7346 9916 7352
rect 9508 6854 9628 6882
rect 9770 6896 9826 6905
rect 9404 6316 9456 6322
rect 9404 6258 9456 6264
rect 9312 6112 9364 6118
rect 9312 6054 9364 6060
rect 9310 5808 9366 5817
rect 9220 5772 9272 5778
rect 9310 5743 9312 5752
rect 9220 5714 9272 5720
rect 9364 5743 9366 5752
rect 9312 5714 9364 5720
rect 9416 5574 9444 6258
rect 9404 5568 9456 5574
rect 9404 5510 9456 5516
rect 9220 5160 9272 5166
rect 9220 5102 9272 5108
rect 9126 4992 9182 5001
rect 9126 4927 9182 4936
rect 8760 4820 8812 4826
rect 8760 4762 8812 4768
rect 8760 4616 8812 4622
rect 9232 4593 9260 5102
rect 8760 4558 8812 4564
rect 9218 4584 9274 4593
rect 8392 4480 8444 4486
rect 8298 4448 8354 4457
rect 8392 4422 8444 4428
rect 8576 4480 8628 4486
rect 8576 4422 8628 4428
rect 8298 4383 8354 4392
rect 8208 4208 8260 4214
rect 8208 4150 8260 4156
rect 7748 3936 7800 3942
rect 8116 3936 8168 3942
rect 7800 3896 8064 3924
rect 7748 3878 7800 3884
rect 7622 3836 7930 3845
rect 7622 3834 7628 3836
rect 7684 3834 7708 3836
rect 7764 3834 7788 3836
rect 7844 3834 7868 3836
rect 7924 3834 7930 3836
rect 7684 3782 7686 3834
rect 7866 3782 7868 3834
rect 7622 3780 7628 3782
rect 7684 3780 7708 3782
rect 7764 3780 7788 3782
rect 7844 3780 7868 3782
rect 7924 3780 7930 3782
rect 7622 3771 7930 3780
rect 7472 3596 7524 3602
rect 7472 3538 7524 3544
rect 8036 3534 8064 3896
rect 8116 3878 8168 3884
rect 8128 3738 8156 3878
rect 8116 3732 8168 3738
rect 8116 3674 8168 3680
rect 8024 3528 8076 3534
rect 8024 3470 8076 3476
rect 7932 3392 7984 3398
rect 7932 3334 7984 3340
rect 7944 3074 7972 3334
rect 6644 3052 6696 3058
rect 6644 2994 6696 3000
rect 7288 3052 7340 3058
rect 7944 3046 8064 3074
rect 7288 2994 7340 3000
rect 5724 2984 5776 2990
rect 5724 2926 5776 2932
rect 7104 2916 7156 2922
rect 7104 2858 7156 2864
rect 7116 2446 7144 2858
rect 7196 2848 7248 2854
rect 7196 2790 7248 2796
rect 7208 2446 7236 2790
rect 7622 2748 7930 2757
rect 7622 2746 7628 2748
rect 7684 2746 7708 2748
rect 7764 2746 7788 2748
rect 7844 2746 7868 2748
rect 7924 2746 7930 2748
rect 7684 2694 7686 2746
rect 7866 2694 7868 2746
rect 7622 2692 7628 2694
rect 7684 2692 7708 2694
rect 7764 2692 7788 2694
rect 7844 2692 7868 2694
rect 7924 2692 7930 2694
rect 7622 2683 7930 2692
rect 8036 2446 8064 3046
rect 2780 2440 2832 2446
rect 2780 2382 2832 2388
rect 3516 2440 3568 2446
rect 4896 2440 4948 2446
rect 3516 2382 3568 2388
rect 3606 2408 3662 2417
rect 2688 2372 2740 2378
rect 4896 2382 4948 2388
rect 5172 2440 5224 2446
rect 5172 2382 5224 2388
rect 7104 2440 7156 2446
rect 7104 2382 7156 2388
rect 7196 2440 7248 2446
rect 7196 2382 7248 2388
rect 8024 2440 8076 2446
rect 8024 2382 8076 2388
rect 3606 2343 3662 2352
rect 2688 2314 2740 2320
rect 2594 2136 2650 2145
rect 2700 2106 2728 2314
rect 3620 2310 3648 2343
rect 2780 2304 2832 2310
rect 2780 2246 2832 2252
rect 2872 2304 2924 2310
rect 2872 2246 2924 2252
rect 3608 2304 3660 2310
rect 3608 2246 3660 2252
rect 3700 2304 3752 2310
rect 3700 2246 3752 2252
rect 4528 2304 4580 2310
rect 4528 2246 4580 2252
rect 5264 2304 5316 2310
rect 5264 2246 5316 2252
rect 6184 2304 6236 2310
rect 6184 2246 6236 2252
rect 7012 2304 7064 2310
rect 7012 2246 7064 2252
rect 7840 2304 7892 2310
rect 7840 2246 7892 2252
rect 2594 2071 2650 2080
rect 2688 2100 2740 2106
rect 2688 2042 2740 2048
rect 2226 1864 2282 1873
rect 2226 1799 2282 1808
rect 2792 1601 2820 2246
rect 2778 1592 2834 1601
rect 2778 1527 2834 1536
rect 2884 800 2912 2246
rect 3712 800 3740 2246
rect 4540 800 4568 2246
rect 5276 1170 5304 2246
rect 5398 2204 5706 2213
rect 5398 2202 5404 2204
rect 5460 2202 5484 2204
rect 5540 2202 5564 2204
rect 5620 2202 5644 2204
rect 5700 2202 5706 2204
rect 5460 2150 5462 2202
rect 5642 2150 5644 2202
rect 5398 2148 5404 2150
rect 5460 2148 5484 2150
rect 5540 2148 5564 2150
rect 5620 2148 5644 2150
rect 5700 2148 5706 2150
rect 5398 2139 5706 2148
rect 5276 1142 5396 1170
rect 5368 800 5396 1142
rect 6196 800 6224 2246
rect 7024 800 7052 2246
rect 7852 800 7880 2246
rect 8128 2009 8156 3674
rect 8220 3641 8248 4150
rect 8588 4078 8616 4422
rect 8772 4282 8800 4558
rect 9218 4519 9274 4528
rect 8760 4276 8812 4282
rect 8760 4218 8812 4224
rect 8300 4072 8352 4078
rect 8300 4014 8352 4020
rect 8576 4072 8628 4078
rect 8576 4014 8628 4020
rect 8312 3942 8340 4014
rect 8300 3936 8352 3942
rect 8300 3878 8352 3884
rect 8206 3632 8262 3641
rect 8206 3567 8262 3576
rect 8208 3392 8260 3398
rect 8208 3334 8260 3340
rect 8220 2514 8248 3334
rect 8772 2922 8800 4218
rect 9128 4072 9180 4078
rect 9128 4014 9180 4020
rect 9140 3942 9168 4014
rect 9232 3942 9260 4519
rect 9312 4480 9364 4486
rect 9312 4422 9364 4428
rect 9324 4282 9352 4422
rect 9312 4276 9364 4282
rect 9312 4218 9364 4224
rect 9508 4078 9536 6854
rect 9770 6831 9826 6840
rect 9588 6792 9640 6798
rect 9784 6780 9812 6831
rect 9876 6798 9904 7346
rect 9640 6752 9812 6780
rect 9864 6792 9916 6798
rect 9588 6734 9640 6740
rect 9864 6734 9916 6740
rect 9968 6644 9996 7500
rect 10244 7478 10272 9046
rect 10232 7472 10284 7478
rect 10232 7414 10284 7420
rect 10336 7342 10364 9687
rect 10428 7426 10456 10406
rect 10598 10367 10654 10376
rect 10612 9994 10640 10367
rect 10600 9988 10652 9994
rect 10600 9930 10652 9936
rect 10704 9738 10732 12174
rect 10612 9710 10732 9738
rect 10612 9674 10640 9710
rect 10520 9646 10640 9674
rect 10796 9654 10824 13126
rect 11060 12640 11112 12646
rect 11060 12582 11112 12588
rect 10874 11656 10930 11665
rect 10874 11591 10930 11600
rect 10784 9648 10836 9654
rect 10520 7954 10548 9646
rect 10690 9616 10746 9625
rect 10784 9590 10836 9596
rect 10690 9551 10746 9560
rect 10600 9376 10652 9382
rect 10600 9318 10652 9324
rect 10612 9178 10640 9318
rect 10600 9172 10652 9178
rect 10600 9114 10652 9120
rect 10598 8936 10654 8945
rect 10598 8871 10654 8880
rect 10612 8498 10640 8871
rect 10704 8809 10732 9551
rect 10796 8906 10824 9590
rect 10888 9353 10916 11591
rect 11072 10674 11100 12582
rect 11164 11354 11192 13144
rect 11440 12850 11468 13280
rect 11520 13262 11572 13268
rect 11716 12918 11744 13670
rect 11808 13258 11836 14894
rect 12624 14884 12676 14890
rect 12624 14826 12676 14832
rect 12070 14716 12378 14725
rect 12070 14714 12076 14716
rect 12132 14714 12156 14716
rect 12212 14714 12236 14716
rect 12292 14714 12316 14716
rect 12372 14714 12378 14716
rect 12132 14662 12134 14714
rect 12314 14662 12316 14714
rect 12070 14660 12076 14662
rect 12132 14660 12156 14662
rect 12212 14660 12236 14662
rect 12292 14660 12316 14662
rect 12372 14660 12378 14662
rect 12070 14651 12378 14660
rect 11978 14512 12034 14521
rect 11978 14447 12034 14456
rect 11992 13394 12020 14447
rect 12440 14272 12492 14278
rect 12440 14214 12492 14220
rect 12452 14074 12480 14214
rect 12440 14068 12492 14074
rect 12440 14010 12492 14016
rect 12070 13628 12378 13637
rect 12070 13626 12076 13628
rect 12132 13626 12156 13628
rect 12212 13626 12236 13628
rect 12292 13626 12316 13628
rect 12372 13626 12378 13628
rect 12132 13574 12134 13626
rect 12314 13574 12316 13626
rect 12070 13572 12076 13574
rect 12132 13572 12156 13574
rect 12212 13572 12236 13574
rect 12292 13572 12316 13574
rect 12372 13572 12378 13574
rect 12070 13563 12378 13572
rect 11980 13388 12032 13394
rect 11900 13348 11980 13376
rect 11796 13252 11848 13258
rect 11796 13194 11848 13200
rect 11704 12912 11756 12918
rect 11704 12854 11756 12860
rect 11428 12844 11480 12850
rect 11428 12786 11480 12792
rect 11244 12708 11296 12714
rect 11244 12650 11296 12656
rect 11256 11937 11284 12650
rect 11440 12306 11468 12786
rect 11704 12708 11756 12714
rect 11704 12650 11756 12656
rect 11428 12300 11480 12306
rect 11428 12242 11480 12248
rect 11336 12232 11388 12238
rect 11336 12174 11388 12180
rect 11242 11928 11298 11937
rect 11242 11863 11298 11872
rect 11348 11778 11376 12174
rect 11256 11750 11376 11778
rect 11152 11348 11204 11354
rect 11152 11290 11204 11296
rect 11164 10810 11192 11290
rect 11152 10804 11204 10810
rect 11152 10746 11204 10752
rect 11060 10668 11112 10674
rect 11060 10610 11112 10616
rect 11256 9874 11284 11750
rect 11612 11552 11664 11558
rect 11610 11520 11612 11529
rect 11664 11520 11666 11529
rect 11610 11455 11666 11464
rect 11716 11370 11744 12650
rect 11808 12434 11836 13194
rect 11900 12714 11928 13348
rect 11980 13330 12032 13336
rect 12072 13184 12124 13190
rect 11992 13144 12072 13172
rect 11888 12708 11940 12714
rect 11888 12650 11940 12656
rect 11808 12406 11928 12434
rect 11796 12232 11848 12238
rect 11796 12174 11848 12180
rect 11808 11529 11836 12174
rect 11794 11520 11850 11529
rect 11794 11455 11850 11464
rect 11624 11342 11744 11370
rect 11428 11076 11480 11082
rect 11428 11018 11480 11024
rect 11164 9846 11284 9874
rect 11060 9648 11112 9654
rect 11164 9625 11192 9846
rect 11244 9716 11296 9722
rect 11244 9658 11296 9664
rect 11060 9590 11112 9596
rect 11150 9616 11206 9625
rect 10968 9376 11020 9382
rect 10874 9344 10930 9353
rect 10968 9318 11020 9324
rect 10874 9279 10930 9288
rect 10784 8900 10836 8906
rect 10784 8842 10836 8848
rect 10690 8800 10746 8809
rect 10690 8735 10746 8744
rect 10600 8492 10652 8498
rect 10600 8434 10652 8440
rect 10508 7948 10560 7954
rect 10508 7890 10560 7896
rect 10600 7812 10652 7818
rect 10600 7754 10652 7760
rect 10428 7398 10548 7426
rect 10612 7410 10640 7754
rect 10704 7546 10732 8735
rect 10784 8628 10836 8634
rect 10784 8570 10836 8576
rect 10692 7540 10744 7546
rect 10692 7482 10744 7488
rect 10232 7336 10284 7342
rect 10232 7278 10284 7284
rect 10324 7336 10376 7342
rect 10324 7278 10376 7284
rect 10138 7168 10194 7177
rect 10138 7103 10194 7112
rect 10152 6866 10180 7103
rect 10140 6860 10192 6866
rect 10140 6802 10192 6808
rect 9692 6616 9996 6644
rect 9692 5930 9720 6616
rect 9846 6556 10154 6565
rect 9846 6554 9852 6556
rect 9908 6554 9932 6556
rect 9988 6554 10012 6556
rect 10068 6554 10092 6556
rect 10148 6554 10154 6556
rect 9908 6502 9910 6554
rect 10090 6502 10092 6554
rect 9846 6500 9852 6502
rect 9908 6500 9932 6502
rect 9988 6500 10012 6502
rect 10068 6500 10092 6502
rect 10148 6500 10154 6502
rect 9846 6491 10154 6500
rect 9956 6384 10008 6390
rect 10244 6361 10272 7278
rect 10324 6656 10376 6662
rect 10324 6598 10376 6604
rect 10336 6458 10364 6598
rect 10324 6452 10376 6458
rect 10324 6394 10376 6400
rect 9956 6326 10008 6332
rect 10046 6352 10102 6361
rect 9968 6186 9996 6326
rect 10046 6287 10102 6296
rect 10230 6352 10286 6361
rect 10230 6287 10286 6296
rect 9956 6180 10008 6186
rect 9956 6122 10008 6128
rect 9864 6112 9916 6118
rect 10060 6089 10088 6287
rect 9864 6054 9916 6060
rect 10046 6080 10102 6089
rect 9600 5902 9720 5930
rect 9600 5114 9628 5902
rect 9680 5840 9732 5846
rect 9680 5782 9732 5788
rect 9692 5302 9720 5782
rect 9772 5704 9824 5710
rect 9876 5692 9904 6054
rect 10046 6015 10102 6024
rect 9824 5664 9904 5692
rect 9772 5646 9824 5652
rect 9772 5568 9824 5574
rect 9772 5510 9824 5516
rect 9784 5370 9812 5510
rect 9846 5468 10154 5477
rect 9846 5466 9852 5468
rect 9908 5466 9932 5468
rect 9988 5466 10012 5468
rect 10068 5466 10092 5468
rect 10148 5466 10154 5468
rect 9908 5414 9910 5466
rect 10090 5414 10092 5466
rect 9846 5412 9852 5414
rect 9908 5412 9932 5414
rect 9988 5412 10012 5414
rect 10068 5412 10092 5414
rect 10148 5412 10154 5414
rect 9846 5403 10154 5412
rect 9772 5364 9824 5370
rect 9772 5306 9824 5312
rect 9680 5296 9732 5302
rect 9680 5238 9732 5244
rect 10140 5160 10192 5166
rect 9600 5086 9720 5114
rect 10140 5102 10192 5108
rect 9588 5024 9640 5030
rect 9588 4966 9640 4972
rect 9600 4282 9628 4966
rect 9692 4758 9720 5086
rect 9680 4752 9732 4758
rect 9680 4694 9732 4700
rect 10152 4690 10180 5102
rect 10140 4684 10192 4690
rect 10140 4626 10192 4632
rect 10244 4622 10272 6287
rect 10428 6254 10456 7398
rect 10520 7342 10548 7398
rect 10600 7404 10652 7410
rect 10600 7346 10652 7352
rect 10508 7336 10560 7342
rect 10508 7278 10560 7284
rect 10600 7268 10652 7274
rect 10600 7210 10652 7216
rect 10508 6792 10560 6798
rect 10508 6734 10560 6740
rect 10416 6248 10468 6254
rect 10416 6190 10468 6196
rect 10416 5636 10468 5642
rect 10416 5578 10468 5584
rect 10232 4616 10284 4622
rect 10232 4558 10284 4564
rect 10428 4486 10456 5578
rect 10520 5098 10548 6734
rect 10612 5710 10640 7210
rect 10692 6316 10744 6322
rect 10692 6258 10744 6264
rect 10704 6118 10732 6258
rect 10692 6112 10744 6118
rect 10692 6054 10744 6060
rect 10796 5710 10824 8570
rect 10980 8265 11008 9318
rect 11072 8566 11100 9590
rect 11150 9551 11206 9560
rect 11256 8974 11284 9658
rect 11336 9444 11388 9450
rect 11336 9386 11388 9392
rect 11348 9217 11376 9386
rect 11334 9208 11390 9217
rect 11334 9143 11390 9152
rect 11244 8968 11296 8974
rect 11348 8945 11376 9143
rect 11244 8910 11296 8916
rect 11334 8936 11390 8945
rect 11334 8871 11390 8880
rect 11060 8560 11112 8566
rect 11060 8502 11112 8508
rect 11440 8430 11468 11018
rect 11518 9616 11574 9625
rect 11518 9551 11574 9560
rect 11532 9450 11560 9551
rect 11520 9444 11572 9450
rect 11520 9386 11572 9392
rect 11428 8424 11480 8430
rect 11428 8366 11480 8372
rect 11060 8356 11112 8362
rect 11060 8298 11112 8304
rect 10966 8256 11022 8265
rect 10966 8191 11022 8200
rect 10876 7948 10928 7954
rect 10876 7890 10928 7896
rect 10888 6866 10916 7890
rect 10968 7744 11020 7750
rect 10968 7686 11020 7692
rect 10980 7546 11008 7686
rect 10968 7540 11020 7546
rect 10968 7482 11020 7488
rect 10876 6860 10928 6866
rect 10928 6820 11008 6848
rect 10876 6802 10928 6808
rect 10876 6656 10928 6662
rect 10876 6598 10928 6604
rect 10600 5704 10652 5710
rect 10784 5704 10836 5710
rect 10600 5646 10652 5652
rect 10704 5664 10784 5692
rect 10508 5092 10560 5098
rect 10508 5034 10560 5040
rect 10520 4690 10548 5034
rect 10508 4684 10560 4690
rect 10508 4626 10560 4632
rect 10704 4622 10732 5664
rect 10888 5681 10916 6598
rect 10980 6390 11008 6820
rect 10968 6384 11020 6390
rect 10968 6326 11020 6332
rect 10968 6112 11020 6118
rect 10968 6054 11020 6060
rect 10784 5646 10836 5652
rect 10874 5672 10930 5681
rect 10874 5607 10930 5616
rect 10784 5568 10836 5574
rect 10784 5510 10836 5516
rect 10796 5370 10824 5510
rect 10784 5364 10836 5370
rect 10784 5306 10836 5312
rect 10782 4720 10838 4729
rect 10782 4655 10784 4664
rect 10836 4655 10838 4664
rect 10784 4626 10836 4632
rect 10692 4616 10744 4622
rect 10692 4558 10744 4564
rect 10416 4480 10468 4486
rect 10416 4422 10468 4428
rect 9846 4380 10154 4389
rect 9846 4378 9852 4380
rect 9908 4378 9932 4380
rect 9988 4378 10012 4380
rect 10068 4378 10092 4380
rect 10148 4378 10154 4380
rect 9908 4326 9910 4378
rect 10090 4326 10092 4378
rect 9846 4324 9852 4326
rect 9908 4324 9932 4326
rect 9988 4324 10012 4326
rect 10068 4324 10092 4326
rect 10148 4324 10154 4326
rect 9846 4315 10154 4324
rect 9588 4276 9640 4282
rect 9588 4218 9640 4224
rect 10428 4214 10456 4422
rect 10416 4208 10468 4214
rect 10416 4150 10468 4156
rect 10508 4208 10560 4214
rect 10508 4150 10560 4156
rect 9496 4072 9548 4078
rect 9496 4014 9548 4020
rect 10520 4010 10548 4150
rect 10782 4040 10838 4049
rect 10508 4004 10560 4010
rect 10782 3975 10838 3984
rect 10508 3946 10560 3952
rect 9128 3936 9180 3942
rect 9128 3878 9180 3884
rect 9220 3936 9272 3942
rect 9220 3878 9272 3884
rect 10324 3936 10376 3942
rect 10324 3878 10376 3884
rect 8944 3664 8996 3670
rect 8944 3606 8996 3612
rect 8760 2916 8812 2922
rect 8760 2858 8812 2864
rect 8208 2508 8260 2514
rect 8208 2450 8260 2456
rect 8956 2446 8984 3606
rect 9846 3292 10154 3301
rect 9846 3290 9852 3292
rect 9908 3290 9932 3292
rect 9988 3290 10012 3292
rect 10068 3290 10092 3292
rect 10148 3290 10154 3292
rect 9908 3238 9910 3290
rect 10090 3238 10092 3290
rect 9846 3236 9852 3238
rect 9908 3236 9932 3238
rect 9988 3236 10012 3238
rect 10068 3236 10092 3238
rect 10148 3236 10154 3238
rect 9846 3227 10154 3236
rect 10336 3194 10364 3878
rect 10796 3738 10824 3975
rect 10888 3738 10916 5607
rect 10980 5273 11008 6054
rect 10966 5264 11022 5273
rect 10966 5199 11022 5208
rect 11072 4622 11100 8298
rect 11428 8288 11480 8294
rect 11428 8230 11480 8236
rect 11440 7954 11468 8230
rect 11428 7948 11480 7954
rect 11348 7908 11428 7936
rect 11244 7880 11296 7886
rect 11244 7822 11296 7828
rect 11152 7744 11204 7750
rect 11152 7686 11204 7692
rect 11164 7478 11192 7686
rect 11152 7472 11204 7478
rect 11152 7414 11204 7420
rect 11150 7032 11206 7041
rect 11256 7018 11284 7822
rect 11348 7750 11376 7908
rect 11428 7890 11480 7896
rect 11532 7750 11560 9386
rect 11624 7818 11652 11342
rect 11796 11076 11848 11082
rect 11796 11018 11848 11024
rect 11704 11008 11756 11014
rect 11704 10950 11756 10956
rect 11716 10674 11744 10950
rect 11808 10742 11836 11018
rect 11796 10736 11848 10742
rect 11796 10678 11848 10684
rect 11704 10668 11756 10674
rect 11704 10610 11756 10616
rect 11808 10130 11836 10678
rect 11796 10124 11848 10130
rect 11796 10066 11848 10072
rect 11704 9920 11756 9926
rect 11704 9862 11756 9868
rect 11716 8974 11744 9862
rect 11808 9586 11836 10066
rect 11796 9580 11848 9586
rect 11796 9522 11848 9528
rect 11808 9042 11836 9522
rect 11796 9036 11848 9042
rect 11796 8978 11848 8984
rect 11704 8968 11756 8974
rect 11704 8910 11756 8916
rect 11612 7812 11664 7818
rect 11612 7754 11664 7760
rect 11336 7744 11388 7750
rect 11336 7686 11388 7692
rect 11520 7744 11572 7750
rect 11520 7686 11572 7692
rect 11348 7274 11376 7686
rect 11716 7410 11744 8910
rect 11796 8356 11848 8362
rect 11796 8298 11848 8304
rect 11704 7404 11756 7410
rect 11704 7346 11756 7352
rect 11428 7336 11480 7342
rect 11428 7278 11480 7284
rect 11612 7336 11664 7342
rect 11612 7278 11664 7284
rect 11336 7268 11388 7274
rect 11336 7210 11388 7216
rect 11206 6990 11284 7018
rect 11440 7002 11468 7278
rect 11428 6996 11480 7002
rect 11150 6967 11206 6976
rect 11164 6798 11192 6967
rect 11428 6938 11480 6944
rect 11520 6996 11572 7002
rect 11520 6938 11572 6944
rect 11152 6792 11204 6798
rect 11152 6734 11204 6740
rect 11152 6656 11204 6662
rect 11152 6598 11204 6604
rect 11060 4616 11112 4622
rect 11164 4593 11192 6598
rect 11426 6488 11482 6497
rect 11348 6446 11426 6474
rect 11348 6322 11376 6446
rect 11426 6423 11482 6432
rect 11428 6384 11480 6390
rect 11428 6326 11480 6332
rect 11336 6316 11388 6322
rect 11336 6258 11388 6264
rect 11244 6248 11296 6254
rect 11244 6190 11296 6196
rect 11256 5030 11284 6190
rect 11336 6112 11388 6118
rect 11336 6054 11388 6060
rect 11244 5024 11296 5030
rect 11244 4966 11296 4972
rect 11242 4720 11298 4729
rect 11348 4690 11376 6054
rect 11440 5778 11468 6326
rect 11428 5772 11480 5778
rect 11428 5714 11480 5720
rect 11426 5264 11482 5273
rect 11426 5199 11482 5208
rect 11440 5001 11468 5199
rect 11426 4992 11482 5001
rect 11426 4927 11482 4936
rect 11242 4655 11298 4664
rect 11336 4684 11388 4690
rect 11060 4558 11112 4564
rect 11150 4584 11206 4593
rect 11150 4519 11206 4528
rect 10784 3732 10836 3738
rect 10784 3674 10836 3680
rect 10876 3732 10928 3738
rect 10876 3674 10928 3680
rect 10796 3534 10824 3674
rect 10784 3528 10836 3534
rect 10784 3470 10836 3476
rect 11152 3392 11204 3398
rect 11152 3334 11204 3340
rect 10324 3188 10376 3194
rect 10324 3130 10376 3136
rect 11164 3097 11192 3334
rect 11150 3088 11206 3097
rect 11150 3023 11206 3032
rect 11152 2848 11204 2854
rect 11152 2790 11204 2796
rect 11164 2446 11192 2790
rect 11256 2582 11284 4655
rect 11336 4626 11388 4632
rect 11428 4480 11480 4486
rect 11428 4422 11480 4428
rect 11440 3126 11468 4422
rect 11532 4146 11560 6938
rect 11624 6186 11652 7278
rect 11704 7200 11756 7206
rect 11704 7142 11756 7148
rect 11716 7002 11744 7142
rect 11704 6996 11756 7002
rect 11704 6938 11756 6944
rect 11704 6860 11756 6866
rect 11704 6802 11756 6808
rect 11612 6180 11664 6186
rect 11612 6122 11664 6128
rect 11716 4758 11744 6802
rect 11808 6186 11836 8298
rect 11900 6866 11928 12406
rect 11992 11354 12020 13144
rect 12072 13126 12124 13132
rect 12636 12850 12664 14826
rect 13268 14816 13320 14822
rect 13268 14758 13320 14764
rect 12992 14408 13044 14414
rect 12992 14350 13044 14356
rect 12808 14068 12860 14074
rect 12808 14010 12860 14016
rect 12820 13938 12848 14010
rect 12808 13932 12860 13938
rect 12808 13874 12860 13880
rect 13004 13870 13032 14350
rect 13176 13932 13228 13938
rect 13176 13874 13228 13880
rect 12992 13864 13044 13870
rect 12992 13806 13044 13812
rect 12716 13728 12768 13734
rect 12716 13670 12768 13676
rect 12900 13728 12952 13734
rect 12900 13670 12952 13676
rect 12728 13190 12756 13670
rect 12912 13394 12940 13670
rect 12900 13388 12952 13394
rect 12900 13330 12952 13336
rect 13004 13308 13032 13806
rect 13084 13320 13136 13326
rect 13004 13280 13084 13308
rect 12716 13184 12768 13190
rect 12716 13126 12768 13132
rect 13004 12918 13032 13280
rect 13084 13262 13136 13268
rect 12992 12912 13044 12918
rect 12992 12854 13044 12860
rect 12624 12844 12676 12850
rect 12624 12786 12676 12792
rect 12070 12540 12378 12549
rect 12070 12538 12076 12540
rect 12132 12538 12156 12540
rect 12212 12538 12236 12540
rect 12292 12538 12316 12540
rect 12372 12538 12378 12540
rect 12132 12486 12134 12538
rect 12314 12486 12316 12538
rect 12070 12484 12076 12486
rect 12132 12484 12156 12486
rect 12212 12484 12236 12486
rect 12292 12484 12316 12486
rect 12372 12484 12378 12486
rect 12070 12475 12378 12484
rect 12072 12232 12124 12238
rect 12072 12174 12124 12180
rect 12084 11762 12112 12174
rect 12808 12164 12860 12170
rect 12808 12106 12860 12112
rect 12072 11756 12124 11762
rect 12072 11698 12124 11704
rect 12070 11452 12378 11461
rect 12070 11450 12076 11452
rect 12132 11450 12156 11452
rect 12212 11450 12236 11452
rect 12292 11450 12316 11452
rect 12372 11450 12378 11452
rect 12132 11398 12134 11450
rect 12314 11398 12316 11450
rect 12070 11396 12076 11398
rect 12132 11396 12156 11398
rect 12212 11396 12236 11398
rect 12292 11396 12316 11398
rect 12372 11396 12378 11398
rect 12070 11387 12378 11396
rect 11980 11348 12032 11354
rect 11980 11290 12032 11296
rect 12072 11348 12124 11354
rect 12072 11290 12124 11296
rect 11992 11082 12020 11290
rect 11980 11076 12032 11082
rect 11980 11018 12032 11024
rect 12084 10452 12112 11290
rect 12716 11076 12768 11082
rect 12716 11018 12768 11024
rect 11992 10424 12112 10452
rect 12440 10464 12492 10470
rect 11992 8514 12020 10424
rect 12440 10406 12492 10412
rect 12070 10364 12378 10373
rect 12070 10362 12076 10364
rect 12132 10362 12156 10364
rect 12212 10362 12236 10364
rect 12292 10362 12316 10364
rect 12372 10362 12378 10364
rect 12132 10310 12134 10362
rect 12314 10310 12316 10362
rect 12070 10308 12076 10310
rect 12132 10308 12156 10310
rect 12212 10308 12236 10310
rect 12292 10308 12316 10310
rect 12372 10308 12378 10310
rect 12070 10299 12378 10308
rect 12070 9276 12378 9285
rect 12070 9274 12076 9276
rect 12132 9274 12156 9276
rect 12212 9274 12236 9276
rect 12292 9274 12316 9276
rect 12372 9274 12378 9276
rect 12132 9222 12134 9274
rect 12314 9222 12316 9274
rect 12070 9220 12076 9222
rect 12132 9220 12156 9222
rect 12212 9220 12236 9222
rect 12292 9220 12316 9222
rect 12372 9220 12378 9222
rect 12070 9211 12378 9220
rect 12164 9172 12216 9178
rect 12452 9160 12480 10406
rect 12622 10296 12678 10305
rect 12622 10231 12678 10240
rect 12636 10033 12664 10231
rect 12622 10024 12678 10033
rect 12622 9959 12678 9968
rect 12624 9716 12676 9722
rect 12624 9658 12676 9664
rect 12636 9586 12664 9658
rect 12624 9580 12676 9586
rect 12624 9522 12676 9528
rect 12216 9132 12480 9160
rect 12164 9114 12216 9120
rect 12624 8968 12676 8974
rect 12624 8910 12676 8916
rect 12636 8514 12664 8910
rect 12728 8634 12756 11018
rect 12820 10810 12848 12106
rect 12900 12096 12952 12102
rect 12900 12038 12952 12044
rect 12912 11762 12940 12038
rect 13004 11830 13032 12854
rect 13084 12096 13136 12102
rect 13084 12038 13136 12044
rect 12992 11824 13044 11830
rect 13096 11801 13124 12038
rect 12992 11766 13044 11772
rect 13082 11792 13138 11801
rect 12900 11756 12952 11762
rect 13082 11727 13138 11736
rect 12900 11698 12952 11704
rect 13084 11144 13136 11150
rect 13084 11086 13136 11092
rect 12808 10804 12860 10810
rect 12808 10746 12860 10752
rect 12716 8628 12768 8634
rect 12716 8570 12768 8576
rect 11992 8486 12112 8514
rect 11980 8424 12032 8430
rect 12084 8401 12112 8486
rect 12440 8492 12492 8498
rect 12636 8486 12756 8514
rect 12440 8434 12492 8440
rect 11980 8366 12032 8372
rect 12070 8392 12126 8401
rect 11992 8090 12020 8366
rect 12070 8327 12126 8336
rect 12070 8188 12378 8197
rect 12070 8186 12076 8188
rect 12132 8186 12156 8188
rect 12212 8186 12236 8188
rect 12292 8186 12316 8188
rect 12372 8186 12378 8188
rect 12132 8134 12134 8186
rect 12314 8134 12316 8186
rect 12070 8132 12076 8134
rect 12132 8132 12156 8134
rect 12212 8132 12236 8134
rect 12292 8132 12316 8134
rect 12372 8132 12378 8134
rect 12070 8123 12378 8132
rect 12452 8090 12480 8434
rect 12624 8424 12676 8430
rect 12624 8366 12676 8372
rect 11980 8084 12032 8090
rect 11980 8026 12032 8032
rect 12440 8084 12492 8090
rect 12440 8026 12492 8032
rect 12348 7948 12400 7954
rect 12348 7890 12400 7896
rect 12070 7848 12126 7857
rect 12360 7818 12388 7890
rect 12636 7886 12664 8366
rect 12624 7880 12676 7886
rect 12624 7822 12676 7828
rect 12070 7783 12126 7792
rect 12348 7812 12400 7818
rect 12084 7750 12112 7783
rect 12348 7754 12400 7760
rect 12532 7812 12584 7818
rect 12532 7754 12584 7760
rect 12072 7744 12124 7750
rect 12072 7686 12124 7692
rect 12440 7336 12492 7342
rect 12440 7278 12492 7284
rect 12070 7100 12378 7109
rect 12070 7098 12076 7100
rect 12132 7098 12156 7100
rect 12212 7098 12236 7100
rect 12292 7098 12316 7100
rect 12372 7098 12378 7100
rect 12132 7046 12134 7098
rect 12314 7046 12316 7098
rect 12070 7044 12076 7046
rect 12132 7044 12156 7046
rect 12212 7044 12236 7046
rect 12292 7044 12316 7046
rect 12372 7044 12378 7046
rect 12070 7035 12378 7044
rect 11978 6896 12034 6905
rect 11888 6860 11940 6866
rect 12452 6866 12480 7278
rect 11978 6831 12034 6840
rect 12440 6860 12492 6866
rect 11888 6802 11940 6808
rect 11992 6662 12020 6831
rect 12440 6802 12492 6808
rect 12438 6760 12494 6769
rect 12438 6695 12494 6704
rect 12452 6662 12480 6695
rect 11980 6656 12032 6662
rect 11980 6598 12032 6604
rect 12440 6656 12492 6662
rect 12440 6598 12492 6604
rect 11888 6316 11940 6322
rect 11888 6258 11940 6264
rect 11796 6180 11848 6186
rect 11796 6122 11848 6128
rect 11900 5914 11928 6258
rect 11888 5908 11940 5914
rect 11888 5850 11940 5856
rect 11992 5778 12020 6598
rect 12256 6316 12308 6322
rect 12256 6258 12308 6264
rect 12268 6225 12296 6258
rect 12254 6216 12310 6225
rect 12254 6151 12310 6160
rect 12070 6012 12378 6021
rect 12070 6010 12076 6012
rect 12132 6010 12156 6012
rect 12212 6010 12236 6012
rect 12292 6010 12316 6012
rect 12372 6010 12378 6012
rect 12132 5958 12134 6010
rect 12314 5958 12316 6010
rect 12070 5956 12076 5958
rect 12132 5956 12156 5958
rect 12212 5956 12236 5958
rect 12292 5956 12316 5958
rect 12372 5956 12378 5958
rect 12070 5947 12378 5956
rect 12544 5846 12572 7754
rect 12622 7712 12678 7721
rect 12622 7647 12678 7656
rect 12072 5840 12124 5846
rect 12072 5782 12124 5788
rect 12532 5840 12584 5846
rect 12532 5782 12584 5788
rect 11980 5772 12032 5778
rect 11980 5714 12032 5720
rect 12084 5681 12112 5782
rect 12440 5772 12492 5778
rect 12440 5714 12492 5720
rect 12256 5704 12308 5710
rect 12070 5672 12126 5681
rect 12256 5646 12308 5652
rect 12070 5607 12126 5616
rect 12268 5409 12296 5646
rect 12452 5556 12480 5714
rect 12360 5528 12480 5556
rect 12254 5400 12310 5409
rect 12254 5335 12310 5344
rect 12360 5166 12388 5528
rect 12544 5234 12572 5782
rect 12532 5228 12584 5234
rect 12532 5170 12584 5176
rect 11980 5160 12032 5166
rect 11980 5102 12032 5108
rect 12348 5160 12400 5166
rect 12348 5102 12400 5108
rect 11992 5030 12020 5102
rect 12532 5092 12584 5098
rect 12532 5034 12584 5040
rect 11980 5024 12032 5030
rect 11980 4966 12032 4972
rect 11794 4856 11850 4865
rect 11794 4791 11796 4800
rect 11848 4791 11850 4800
rect 11796 4762 11848 4768
rect 11704 4752 11756 4758
rect 11704 4694 11756 4700
rect 11888 4616 11940 4622
rect 11888 4558 11940 4564
rect 11704 4480 11756 4486
rect 11704 4422 11756 4428
rect 11520 4140 11572 4146
rect 11520 4082 11572 4088
rect 11716 4026 11744 4422
rect 11624 3998 11744 4026
rect 11428 3120 11480 3126
rect 11428 3062 11480 3068
rect 11624 3058 11652 3998
rect 11704 3936 11756 3942
rect 11704 3878 11756 3884
rect 11612 3052 11664 3058
rect 11612 2994 11664 3000
rect 11520 2848 11572 2854
rect 11520 2790 11572 2796
rect 11244 2576 11296 2582
rect 11244 2518 11296 2524
rect 11532 2446 11560 2790
rect 11716 2446 11744 3878
rect 11900 2650 11928 4558
rect 11992 4282 12020 4966
rect 12070 4924 12378 4933
rect 12070 4922 12076 4924
rect 12132 4922 12156 4924
rect 12212 4922 12236 4924
rect 12292 4922 12316 4924
rect 12372 4922 12378 4924
rect 12132 4870 12134 4922
rect 12314 4870 12316 4922
rect 12070 4868 12076 4870
rect 12132 4868 12156 4870
rect 12212 4868 12236 4870
rect 12292 4868 12316 4870
rect 12372 4868 12378 4870
rect 12070 4859 12378 4868
rect 12348 4820 12400 4826
rect 12348 4762 12400 4768
rect 11980 4276 12032 4282
rect 11980 4218 12032 4224
rect 11980 4072 12032 4078
rect 11978 4040 11980 4049
rect 12032 4040 12034 4049
rect 12360 4010 12388 4762
rect 12544 4214 12572 5034
rect 12532 4208 12584 4214
rect 12532 4150 12584 4156
rect 11978 3975 12034 3984
rect 12348 4004 12400 4010
rect 12348 3946 12400 3952
rect 12440 3936 12492 3942
rect 12440 3878 12492 3884
rect 12070 3836 12378 3845
rect 12070 3834 12076 3836
rect 12132 3834 12156 3836
rect 12212 3834 12236 3836
rect 12292 3834 12316 3836
rect 12372 3834 12378 3836
rect 12132 3782 12134 3834
rect 12314 3782 12316 3834
rect 12070 3780 12076 3782
rect 12132 3780 12156 3782
rect 12212 3780 12236 3782
rect 12292 3780 12316 3782
rect 12372 3780 12378 3782
rect 12070 3771 12378 3780
rect 11980 2848 12032 2854
rect 11980 2790 12032 2796
rect 11888 2644 11940 2650
rect 11888 2586 11940 2592
rect 11992 2514 12020 2790
rect 12070 2748 12378 2757
rect 12070 2746 12076 2748
rect 12132 2746 12156 2748
rect 12212 2746 12236 2748
rect 12292 2746 12316 2748
rect 12372 2746 12378 2748
rect 12132 2694 12134 2746
rect 12314 2694 12316 2746
rect 12070 2692 12076 2694
rect 12132 2692 12156 2694
rect 12212 2692 12236 2694
rect 12292 2692 12316 2694
rect 12372 2692 12378 2694
rect 12070 2683 12378 2692
rect 11980 2508 12032 2514
rect 11980 2450 12032 2456
rect 12452 2446 12480 3878
rect 12532 3460 12584 3466
rect 12532 3402 12584 3408
rect 12544 3194 12572 3402
rect 12532 3188 12584 3194
rect 12532 3130 12584 3136
rect 12636 3058 12664 7647
rect 12728 6934 12756 8486
rect 12820 7342 12848 10746
rect 12990 10024 13046 10033
rect 12990 9959 13046 9968
rect 12900 8560 12952 8566
rect 12900 8502 12952 8508
rect 12808 7336 12860 7342
rect 12808 7278 12860 7284
rect 12716 6928 12768 6934
rect 12714 6896 12716 6905
rect 12768 6896 12770 6905
rect 12820 6866 12848 7278
rect 12714 6831 12770 6840
rect 12808 6860 12860 6866
rect 12808 6802 12860 6808
rect 12808 6656 12860 6662
rect 12728 6616 12808 6644
rect 12728 4282 12756 6616
rect 12808 6598 12860 6604
rect 12912 6186 12940 8502
rect 13004 7478 13032 9959
rect 13096 9042 13124 11086
rect 13188 9178 13216 13874
rect 13280 12714 13308 14758
rect 13450 14512 13506 14521
rect 13924 14498 13952 16400
rect 16518 14716 16826 14725
rect 16518 14714 16524 14716
rect 16580 14714 16604 14716
rect 16660 14714 16684 14716
rect 16740 14714 16764 14716
rect 16820 14714 16826 14716
rect 16580 14662 16582 14714
rect 16762 14662 16764 14714
rect 16518 14660 16524 14662
rect 16580 14660 16604 14662
rect 16660 14660 16684 14662
rect 16740 14660 16764 14662
rect 16820 14660 16826 14662
rect 16518 14651 16826 14660
rect 15936 14612 15988 14618
rect 15936 14554 15988 14560
rect 13924 14470 14044 14498
rect 13450 14447 13506 14456
rect 13360 14408 13412 14414
rect 13360 14350 13412 14356
rect 13268 12708 13320 12714
rect 13268 12650 13320 12656
rect 13176 9172 13228 9178
rect 13176 9114 13228 9120
rect 13084 9036 13136 9042
rect 13084 8978 13136 8984
rect 13188 8838 13216 9114
rect 13176 8832 13228 8838
rect 13176 8774 13228 8780
rect 13280 7954 13308 12650
rect 13372 9586 13400 14350
rect 13464 13258 13492 14447
rect 14016 14414 14044 14470
rect 15292 14476 15344 14482
rect 15292 14418 15344 14424
rect 14004 14408 14056 14414
rect 14004 14350 14056 14356
rect 13912 14340 13964 14346
rect 13912 14282 13964 14288
rect 13728 14000 13780 14006
rect 13728 13942 13780 13948
rect 13636 13320 13688 13326
rect 13636 13262 13688 13268
rect 13452 13252 13504 13258
rect 13452 13194 13504 13200
rect 13452 12844 13504 12850
rect 13452 12786 13504 12792
rect 13464 12594 13492 12786
rect 13544 12640 13596 12646
rect 13464 12588 13544 12594
rect 13464 12582 13596 12588
rect 13464 12566 13584 12582
rect 13464 12442 13492 12566
rect 13452 12436 13504 12442
rect 13452 12378 13504 12384
rect 13544 11688 13596 11694
rect 13544 11630 13596 11636
rect 13556 11082 13584 11630
rect 13544 11076 13596 11082
rect 13544 11018 13596 11024
rect 13450 10568 13506 10577
rect 13450 10503 13506 10512
rect 13464 10198 13492 10503
rect 13452 10192 13504 10198
rect 13452 10134 13504 10140
rect 13556 10146 13584 11018
rect 13648 10266 13676 13262
rect 13740 11694 13768 13942
rect 13820 11892 13872 11898
rect 13820 11834 13872 11840
rect 13728 11688 13780 11694
rect 13728 11630 13780 11636
rect 13728 11280 13780 11286
rect 13728 11222 13780 11228
rect 13636 10260 13688 10266
rect 13636 10202 13688 10208
rect 13740 10169 13768 11222
rect 13726 10160 13782 10169
rect 13556 10118 13676 10146
rect 13360 9580 13412 9586
rect 13360 9522 13412 9528
rect 13372 8820 13400 9522
rect 13544 9512 13596 9518
rect 13450 9480 13506 9489
rect 13648 9489 13676 10118
rect 13726 10095 13782 10104
rect 13832 9654 13860 11834
rect 13924 11286 13952 14282
rect 14016 13530 14044 14350
rect 14740 14272 14792 14278
rect 14740 14214 14792 14220
rect 14924 14272 14976 14278
rect 14924 14214 14976 14220
rect 14294 14172 14602 14181
rect 14294 14170 14300 14172
rect 14356 14170 14380 14172
rect 14436 14170 14460 14172
rect 14516 14170 14540 14172
rect 14596 14170 14602 14172
rect 14356 14118 14358 14170
rect 14538 14118 14540 14170
rect 14294 14116 14300 14118
rect 14356 14116 14380 14118
rect 14436 14116 14460 14118
rect 14516 14116 14540 14118
rect 14596 14116 14602 14118
rect 14294 14107 14602 14116
rect 14188 13864 14240 13870
rect 14188 13806 14240 13812
rect 14648 13864 14700 13870
rect 14648 13806 14700 13812
rect 14004 13524 14056 13530
rect 14004 13466 14056 13472
rect 14200 13326 14228 13806
rect 14188 13320 14240 13326
rect 14188 13262 14240 13268
rect 14096 13184 14148 13190
rect 14016 13144 14096 13172
rect 14016 11354 14044 13144
rect 14096 13126 14148 13132
rect 14094 12744 14150 12753
rect 14094 12679 14150 12688
rect 14108 12442 14136 12679
rect 14096 12436 14148 12442
rect 14096 12378 14148 12384
rect 14096 12164 14148 12170
rect 14096 12106 14148 12112
rect 14108 12073 14136 12106
rect 14200 12102 14228 13262
rect 14294 13084 14602 13093
rect 14294 13082 14300 13084
rect 14356 13082 14380 13084
rect 14436 13082 14460 13084
rect 14516 13082 14540 13084
rect 14596 13082 14602 13084
rect 14356 13030 14358 13082
rect 14538 13030 14540 13082
rect 14294 13028 14300 13030
rect 14356 13028 14380 13030
rect 14436 13028 14460 13030
rect 14516 13028 14540 13030
rect 14596 13028 14602 13030
rect 14294 13019 14602 13028
rect 14660 12434 14688 13806
rect 14752 13802 14780 14214
rect 14740 13796 14792 13802
rect 14740 13738 14792 13744
rect 14936 13734 14964 14214
rect 15200 14000 15252 14006
rect 15200 13942 15252 13948
rect 14924 13728 14976 13734
rect 14924 13670 14976 13676
rect 15212 12889 15240 13942
rect 15304 13433 15332 14418
rect 15660 14340 15712 14346
rect 15660 14282 15712 14288
rect 15382 13968 15438 13977
rect 15382 13903 15438 13912
rect 15290 13424 15346 13433
rect 15290 13359 15346 13368
rect 14738 12880 14794 12889
rect 15198 12880 15254 12889
rect 14738 12815 14794 12824
rect 14936 12838 15148 12866
rect 14752 12442 14780 12815
rect 14568 12406 14688 12434
rect 14740 12436 14792 12442
rect 14568 12170 14596 12406
rect 14936 12434 14964 12838
rect 15016 12776 15068 12782
rect 15016 12718 15068 12724
rect 14740 12378 14792 12384
rect 14844 12406 14964 12434
rect 14556 12164 14608 12170
rect 14556 12106 14608 12112
rect 14648 12164 14700 12170
rect 14648 12106 14700 12112
rect 14188 12096 14240 12102
rect 14094 12064 14150 12073
rect 14188 12038 14240 12044
rect 14094 11999 14150 12008
rect 14294 11996 14602 12005
rect 14294 11994 14300 11996
rect 14356 11994 14380 11996
rect 14436 11994 14460 11996
rect 14516 11994 14540 11996
rect 14596 11994 14602 11996
rect 14356 11942 14358 11994
rect 14538 11942 14540 11994
rect 14294 11940 14300 11942
rect 14356 11940 14380 11942
rect 14436 11940 14460 11942
rect 14516 11940 14540 11942
rect 14596 11940 14602 11942
rect 14294 11931 14602 11940
rect 14660 11762 14688 12106
rect 14740 12096 14792 12102
rect 14740 12038 14792 12044
rect 14648 11756 14700 11762
rect 14648 11698 14700 11704
rect 14094 11656 14150 11665
rect 14094 11591 14150 11600
rect 14004 11348 14056 11354
rect 14004 11290 14056 11296
rect 13912 11280 13964 11286
rect 13912 11222 13964 11228
rect 14004 10192 14056 10198
rect 14004 10134 14056 10140
rect 13912 9920 13964 9926
rect 13912 9862 13964 9868
rect 13924 9654 13952 9862
rect 13820 9648 13872 9654
rect 13820 9590 13872 9596
rect 13912 9648 13964 9654
rect 13912 9590 13964 9596
rect 13544 9454 13596 9460
rect 13634 9480 13690 9489
rect 13450 9415 13506 9424
rect 13464 9382 13492 9415
rect 13452 9376 13504 9382
rect 13452 9318 13504 9324
rect 13556 8974 13584 9454
rect 13634 9415 13690 9424
rect 13820 9172 13872 9178
rect 13820 9114 13872 9120
rect 13636 9104 13688 9110
rect 13636 9046 13688 9052
rect 13544 8968 13596 8974
rect 13544 8910 13596 8916
rect 13452 8832 13504 8838
rect 13372 8792 13452 8820
rect 13544 8832 13596 8838
rect 13452 8774 13504 8780
rect 13542 8800 13544 8809
rect 13596 8800 13598 8809
rect 13358 8528 13414 8537
rect 13358 8463 13414 8472
rect 13268 7948 13320 7954
rect 13268 7890 13320 7896
rect 13084 7744 13136 7750
rect 13084 7686 13136 7692
rect 13096 7546 13124 7686
rect 13084 7540 13136 7546
rect 13084 7482 13136 7488
rect 12992 7472 13044 7478
rect 12992 7414 13044 7420
rect 13268 7472 13320 7478
rect 13268 7414 13320 7420
rect 13004 7313 13032 7414
rect 13176 7336 13228 7342
rect 12990 7304 13046 7313
rect 13176 7278 13228 7284
rect 12990 7239 13046 7248
rect 12992 7200 13044 7206
rect 12992 7142 13044 7148
rect 13004 7002 13032 7142
rect 12992 6996 13044 7002
rect 12992 6938 13044 6944
rect 13004 6474 13032 6938
rect 13004 6446 13124 6474
rect 12992 6316 13044 6322
rect 12992 6258 13044 6264
rect 12900 6180 12952 6186
rect 12900 6122 12952 6128
rect 12806 6080 12862 6089
rect 12806 6015 12862 6024
rect 12820 4690 12848 6015
rect 12912 5778 12940 6122
rect 13004 5914 13032 6258
rect 13096 6202 13124 6446
rect 13188 6322 13216 7278
rect 13176 6316 13228 6322
rect 13176 6258 13228 6264
rect 13096 6174 13216 6202
rect 13084 6112 13136 6118
rect 13084 6054 13136 6060
rect 12992 5908 13044 5914
rect 12992 5850 13044 5856
rect 13096 5778 13124 6054
rect 12900 5772 12952 5778
rect 12900 5714 12952 5720
rect 13084 5772 13136 5778
rect 13084 5714 13136 5720
rect 13188 5658 13216 6174
rect 13280 5846 13308 7414
rect 13268 5840 13320 5846
rect 13268 5782 13320 5788
rect 13268 5704 13320 5710
rect 12900 5636 12952 5642
rect 12900 5578 12952 5584
rect 13096 5630 13216 5658
rect 13266 5672 13268 5681
rect 13320 5672 13322 5681
rect 12912 4826 12940 5578
rect 12992 5296 13044 5302
rect 12992 5238 13044 5244
rect 13004 5098 13032 5238
rect 12992 5092 13044 5098
rect 12992 5034 13044 5040
rect 12900 4820 12952 4826
rect 12900 4762 12952 4768
rect 12808 4684 12860 4690
rect 12808 4626 12860 4632
rect 12806 4448 12862 4457
rect 12806 4383 12862 4392
rect 12990 4448 13046 4457
rect 12990 4383 13046 4392
rect 12716 4276 12768 4282
rect 12716 4218 12768 4224
rect 12820 3942 12848 4383
rect 13004 4146 13032 4383
rect 12900 4140 12952 4146
rect 12900 4082 12952 4088
rect 12992 4140 13044 4146
rect 12992 4082 13044 4088
rect 12808 3936 12860 3942
rect 12808 3878 12860 3884
rect 12820 3602 12848 3878
rect 12912 3602 12940 4082
rect 12992 4004 13044 4010
rect 12992 3946 13044 3952
rect 13004 3641 13032 3946
rect 13096 3670 13124 5630
rect 13266 5607 13322 5616
rect 13176 5228 13228 5234
rect 13176 5170 13228 5176
rect 13268 5228 13320 5234
rect 13268 5170 13320 5176
rect 13188 4457 13216 5170
rect 13174 4448 13230 4457
rect 13174 4383 13230 4392
rect 13280 4282 13308 5170
rect 13372 5166 13400 8463
rect 13464 8294 13492 8774
rect 13542 8735 13598 8744
rect 13556 8378 13584 8735
rect 13648 8566 13676 9046
rect 13636 8560 13688 8566
rect 13636 8502 13688 8508
rect 13832 8498 13860 9114
rect 13912 8628 13964 8634
rect 13912 8570 13964 8576
rect 13820 8492 13872 8498
rect 13820 8434 13872 8440
rect 13556 8350 13676 8378
rect 13452 8288 13504 8294
rect 13452 8230 13504 8236
rect 13452 8016 13504 8022
rect 13648 7993 13676 8350
rect 13452 7958 13504 7964
rect 13634 7984 13690 7993
rect 13464 6934 13492 7958
rect 13544 7948 13596 7954
rect 13634 7919 13690 7928
rect 13544 7890 13596 7896
rect 13556 7342 13584 7890
rect 13648 7886 13676 7919
rect 13636 7880 13688 7886
rect 13636 7822 13688 7828
rect 13820 7744 13872 7750
rect 13820 7686 13872 7692
rect 13544 7336 13596 7342
rect 13832 7313 13860 7686
rect 13544 7278 13596 7284
rect 13818 7304 13874 7313
rect 13818 7239 13874 7248
rect 13544 7200 13596 7206
rect 13544 7142 13596 7148
rect 13636 7200 13688 7206
rect 13636 7142 13688 7148
rect 13452 6928 13504 6934
rect 13452 6870 13504 6876
rect 13556 6798 13584 7142
rect 13544 6792 13596 6798
rect 13544 6734 13596 6740
rect 13648 6662 13676 7142
rect 13820 6724 13872 6730
rect 13820 6666 13872 6672
rect 13636 6656 13688 6662
rect 13636 6598 13688 6604
rect 13636 6112 13688 6118
rect 13636 6054 13688 6060
rect 13452 5908 13504 5914
rect 13452 5850 13504 5856
rect 13464 5250 13492 5850
rect 13544 5772 13596 5778
rect 13544 5714 13596 5720
rect 13556 5370 13584 5714
rect 13544 5364 13596 5370
rect 13544 5306 13596 5312
rect 13464 5222 13584 5250
rect 13360 5160 13412 5166
rect 13360 5102 13412 5108
rect 13452 5024 13504 5030
rect 13452 4966 13504 4972
rect 13464 4690 13492 4966
rect 13452 4684 13504 4690
rect 13452 4626 13504 4632
rect 13268 4276 13320 4282
rect 13268 4218 13320 4224
rect 13084 3664 13136 3670
rect 12990 3632 13046 3641
rect 12808 3596 12860 3602
rect 12808 3538 12860 3544
rect 12900 3596 12952 3602
rect 13084 3606 13136 3612
rect 12990 3567 13046 3576
rect 12900 3538 12952 3544
rect 13004 3194 13032 3567
rect 13082 3496 13138 3505
rect 13082 3431 13138 3440
rect 12992 3188 13044 3194
rect 12992 3130 13044 3136
rect 12624 3052 12676 3058
rect 12624 2994 12676 3000
rect 13096 2961 13124 3431
rect 13556 3398 13584 5222
rect 13648 4486 13676 6054
rect 13728 5704 13780 5710
rect 13728 5646 13780 5652
rect 13636 4480 13688 4486
rect 13636 4422 13688 4428
rect 13648 3505 13676 4422
rect 13740 4282 13768 5646
rect 13832 4758 13860 6666
rect 13924 6662 13952 8570
rect 13912 6656 13964 6662
rect 13912 6598 13964 6604
rect 13910 6488 13966 6497
rect 13910 6423 13966 6432
rect 13924 5914 13952 6423
rect 13912 5908 13964 5914
rect 13912 5850 13964 5856
rect 13912 5568 13964 5574
rect 13910 5536 13912 5545
rect 13964 5536 13966 5545
rect 13910 5471 13966 5480
rect 13910 5400 13966 5409
rect 13910 5335 13912 5344
rect 13964 5335 13966 5344
rect 13912 5306 13964 5312
rect 14016 5114 14044 10134
rect 14108 9897 14136 11591
rect 14752 11218 14780 12038
rect 14740 11212 14792 11218
rect 14740 11154 14792 11160
rect 14294 10908 14602 10917
rect 14294 10906 14300 10908
rect 14356 10906 14380 10908
rect 14436 10906 14460 10908
rect 14516 10906 14540 10908
rect 14596 10906 14602 10908
rect 14356 10854 14358 10906
rect 14538 10854 14540 10906
rect 14294 10852 14300 10854
rect 14356 10852 14380 10854
rect 14436 10852 14460 10854
rect 14516 10852 14540 10854
rect 14596 10852 14602 10854
rect 14294 10843 14602 10852
rect 14556 10668 14608 10674
rect 14556 10610 14608 10616
rect 14188 10464 14240 10470
rect 14188 10406 14240 10412
rect 14094 9888 14150 9897
rect 14094 9823 14150 9832
rect 14096 9716 14148 9722
rect 14096 9658 14148 9664
rect 14108 9110 14136 9658
rect 14096 9104 14148 9110
rect 14096 9046 14148 9052
rect 14200 8906 14228 10406
rect 14568 10198 14596 10610
rect 14556 10192 14608 10198
rect 14556 10134 14608 10140
rect 14648 9920 14700 9926
rect 14648 9862 14700 9868
rect 14294 9820 14602 9829
rect 14294 9818 14300 9820
rect 14356 9818 14380 9820
rect 14436 9818 14460 9820
rect 14516 9818 14540 9820
rect 14596 9818 14602 9820
rect 14356 9766 14358 9818
rect 14538 9766 14540 9818
rect 14294 9764 14300 9766
rect 14356 9764 14380 9766
rect 14436 9764 14460 9766
rect 14516 9764 14540 9766
rect 14596 9764 14602 9766
rect 14294 9755 14602 9764
rect 14188 8900 14240 8906
rect 14108 8860 14188 8888
rect 14108 5148 14136 8860
rect 14188 8842 14240 8848
rect 14294 8732 14602 8741
rect 14294 8730 14300 8732
rect 14356 8730 14380 8732
rect 14436 8730 14460 8732
rect 14516 8730 14540 8732
rect 14596 8730 14602 8732
rect 14356 8678 14358 8730
rect 14538 8678 14540 8730
rect 14294 8676 14300 8678
rect 14356 8676 14380 8678
rect 14436 8676 14460 8678
rect 14516 8676 14540 8678
rect 14596 8676 14602 8678
rect 14294 8667 14602 8676
rect 14188 8492 14240 8498
rect 14188 8434 14240 8440
rect 14200 7478 14228 8434
rect 14294 7644 14602 7653
rect 14294 7642 14300 7644
rect 14356 7642 14380 7644
rect 14436 7642 14460 7644
rect 14516 7642 14540 7644
rect 14596 7642 14602 7644
rect 14356 7590 14358 7642
rect 14538 7590 14540 7642
rect 14294 7588 14300 7590
rect 14356 7588 14380 7590
rect 14436 7588 14460 7590
rect 14516 7588 14540 7590
rect 14596 7588 14602 7590
rect 14294 7579 14602 7588
rect 14188 7472 14240 7478
rect 14188 7414 14240 7420
rect 14556 7472 14608 7478
rect 14556 7414 14608 7420
rect 14188 7336 14240 7342
rect 14188 7278 14240 7284
rect 14200 6118 14228 7278
rect 14568 6730 14596 7414
rect 14556 6724 14608 6730
rect 14556 6666 14608 6672
rect 14294 6556 14602 6565
rect 14294 6554 14300 6556
rect 14356 6554 14380 6556
rect 14436 6554 14460 6556
rect 14516 6554 14540 6556
rect 14596 6554 14602 6556
rect 14356 6502 14358 6554
rect 14538 6502 14540 6554
rect 14294 6500 14300 6502
rect 14356 6500 14380 6502
rect 14436 6500 14460 6502
rect 14516 6500 14540 6502
rect 14596 6500 14602 6502
rect 14294 6491 14602 6500
rect 14280 6452 14332 6458
rect 14280 6394 14332 6400
rect 14292 6254 14320 6394
rect 14372 6316 14424 6322
rect 14372 6258 14424 6264
rect 14280 6248 14332 6254
rect 14384 6225 14412 6258
rect 14280 6190 14332 6196
rect 14370 6216 14426 6225
rect 14188 6112 14240 6118
rect 14188 6054 14240 6060
rect 14292 5556 14320 6190
rect 14370 6151 14426 6160
rect 14200 5528 14320 5556
rect 14200 5250 14228 5528
rect 14294 5468 14602 5477
rect 14294 5466 14300 5468
rect 14356 5466 14380 5468
rect 14436 5466 14460 5468
rect 14516 5466 14540 5468
rect 14596 5466 14602 5468
rect 14356 5414 14358 5466
rect 14538 5414 14540 5466
rect 14294 5412 14300 5414
rect 14356 5412 14380 5414
rect 14436 5412 14460 5414
rect 14516 5412 14540 5414
rect 14596 5412 14602 5414
rect 14294 5403 14602 5412
rect 14200 5222 14320 5250
rect 14108 5120 14228 5148
rect 13924 5086 14044 5114
rect 13924 4826 13952 5086
rect 14200 5030 14228 5120
rect 14004 5024 14056 5030
rect 14004 4966 14056 4972
rect 14188 5024 14240 5030
rect 14188 4966 14240 4972
rect 13912 4820 13964 4826
rect 13912 4762 13964 4768
rect 13820 4752 13872 4758
rect 13820 4694 13872 4700
rect 13728 4276 13780 4282
rect 13728 4218 13780 4224
rect 13740 3670 13768 4218
rect 13924 4214 13952 4762
rect 14016 4622 14044 4966
rect 14200 4690 14228 4966
rect 14188 4684 14240 4690
rect 14188 4626 14240 4632
rect 14004 4616 14056 4622
rect 14004 4558 14056 4564
rect 14096 4616 14148 4622
rect 14292 4570 14320 5222
rect 14372 5160 14424 5166
rect 14372 5102 14424 5108
rect 14556 5160 14608 5166
rect 14556 5102 14608 5108
rect 14096 4558 14148 4564
rect 14002 4448 14058 4457
rect 14002 4383 14058 4392
rect 14016 4214 14044 4383
rect 14108 4282 14136 4558
rect 14200 4542 14320 4570
rect 14384 4554 14412 5102
rect 14568 5030 14596 5102
rect 14556 5024 14608 5030
rect 14556 4966 14608 4972
rect 14096 4276 14148 4282
rect 14096 4218 14148 4224
rect 13912 4208 13964 4214
rect 13912 4150 13964 4156
rect 14004 4208 14056 4214
rect 14004 4150 14056 4156
rect 14200 4146 14228 4542
rect 14292 4486 14320 4542
rect 14372 4548 14424 4554
rect 14372 4490 14424 4496
rect 14280 4480 14332 4486
rect 14280 4422 14332 4428
rect 14294 4380 14602 4389
rect 14294 4378 14300 4380
rect 14356 4378 14380 4380
rect 14436 4378 14460 4380
rect 14516 4378 14540 4380
rect 14596 4378 14602 4380
rect 14356 4326 14358 4378
rect 14538 4326 14540 4378
rect 14294 4324 14300 4326
rect 14356 4324 14380 4326
rect 14436 4324 14460 4326
rect 14516 4324 14540 4326
rect 14596 4324 14602 4326
rect 14294 4315 14602 4324
rect 14660 4146 14688 9862
rect 14740 9580 14792 9586
rect 14740 9522 14792 9528
rect 14752 7834 14780 9522
rect 14844 9178 14872 12406
rect 15028 11642 15056 12718
rect 15120 12646 15148 12838
rect 15198 12815 15254 12824
rect 15396 12730 15424 13903
rect 15476 13320 15528 13326
rect 15476 13262 15528 13268
rect 15488 12918 15516 13262
rect 15476 12912 15528 12918
rect 15476 12854 15528 12860
rect 15304 12714 15424 12730
rect 15292 12708 15424 12714
rect 15344 12702 15424 12708
rect 15292 12650 15344 12656
rect 15108 12640 15160 12646
rect 15108 12582 15160 12588
rect 15488 12238 15516 12854
rect 15476 12232 15528 12238
rect 15396 12192 15476 12220
rect 15396 11830 15424 12192
rect 15476 12174 15528 12180
rect 15476 12096 15528 12102
rect 15476 12038 15528 12044
rect 15384 11824 15436 11830
rect 15384 11766 15436 11772
rect 14936 11614 15056 11642
rect 14936 9738 14964 11614
rect 15108 11552 15160 11558
rect 15108 11494 15160 11500
rect 15120 9926 15148 11494
rect 15488 11082 15516 12038
rect 15672 11801 15700 14282
rect 15948 14249 15976 14554
rect 16304 14408 16356 14414
rect 16304 14350 16356 14356
rect 15934 14240 15990 14249
rect 15934 14175 15990 14184
rect 16316 14074 16344 14350
rect 17592 14340 17644 14346
rect 17592 14282 17644 14288
rect 16396 14272 16448 14278
rect 16396 14214 16448 14220
rect 16304 14068 16356 14074
rect 16304 14010 16356 14016
rect 16212 14000 16264 14006
rect 16212 13942 16264 13948
rect 16224 13258 16252 13942
rect 16212 13252 16264 13258
rect 16212 13194 16264 13200
rect 16316 12918 16344 14010
rect 16408 13530 16436 14214
rect 17222 13696 17278 13705
rect 16518 13628 16826 13637
rect 17222 13631 17278 13640
rect 16518 13626 16524 13628
rect 16580 13626 16604 13628
rect 16660 13626 16684 13628
rect 16740 13626 16764 13628
rect 16820 13626 16826 13628
rect 16580 13574 16582 13626
rect 16762 13574 16764 13626
rect 16518 13572 16524 13574
rect 16580 13572 16604 13574
rect 16660 13572 16684 13574
rect 16740 13572 16764 13574
rect 16820 13572 16826 13574
rect 16518 13563 16826 13572
rect 16396 13524 16448 13530
rect 16396 13466 16448 13472
rect 17132 13388 17184 13394
rect 17132 13330 17184 13336
rect 16856 13252 16908 13258
rect 16856 13194 16908 13200
rect 16304 12912 16356 12918
rect 16488 12912 16540 12918
rect 16304 12854 16356 12860
rect 16486 12880 16488 12889
rect 16540 12880 16542 12889
rect 16028 12844 16080 12850
rect 16486 12815 16542 12824
rect 16028 12786 16080 12792
rect 16040 12646 16068 12786
rect 16028 12640 16080 12646
rect 16028 12582 16080 12588
rect 16518 12540 16826 12549
rect 16518 12538 16524 12540
rect 16580 12538 16604 12540
rect 16660 12538 16684 12540
rect 16740 12538 16764 12540
rect 16820 12538 16826 12540
rect 16580 12486 16582 12538
rect 16762 12486 16764 12538
rect 16518 12484 16524 12486
rect 16580 12484 16604 12486
rect 16660 12484 16684 12486
rect 16740 12484 16764 12486
rect 16820 12484 16826 12486
rect 16518 12475 16826 12484
rect 16764 12164 16816 12170
rect 16764 12106 16816 12112
rect 15752 11892 15804 11898
rect 15752 11834 15804 11840
rect 15658 11792 15714 11801
rect 15658 11727 15714 11736
rect 15764 11150 15792 11834
rect 16120 11756 16172 11762
rect 16120 11698 16172 11704
rect 16132 11286 16160 11698
rect 16776 11665 16804 12106
rect 16762 11656 16818 11665
rect 16408 11614 16620 11642
rect 16120 11280 16172 11286
rect 16120 11222 16172 11228
rect 15752 11144 15804 11150
rect 15752 11086 15804 11092
rect 15476 11076 15528 11082
rect 15476 11018 15528 11024
rect 15568 11076 15620 11082
rect 15936 11076 15988 11082
rect 15568 11018 15620 11024
rect 15856 11036 15936 11064
rect 15384 10668 15436 10674
rect 15384 10610 15436 10616
rect 15396 10062 15424 10610
rect 15292 10056 15344 10062
rect 15292 9998 15344 10004
rect 15384 10056 15436 10062
rect 15384 9998 15436 10004
rect 15200 9988 15252 9994
rect 15200 9930 15252 9936
rect 15108 9920 15160 9926
rect 15212 9897 15240 9930
rect 15108 9862 15160 9868
rect 15198 9888 15254 9897
rect 15198 9823 15254 9832
rect 15106 9752 15162 9761
rect 14936 9722 15056 9738
rect 14924 9716 15056 9722
rect 14976 9710 15056 9716
rect 14924 9658 14976 9664
rect 14924 9580 14976 9586
rect 14924 9522 14976 9528
rect 14936 9382 14964 9522
rect 15028 9382 15056 9710
rect 15106 9687 15162 9696
rect 14924 9376 14976 9382
rect 14924 9318 14976 9324
rect 15016 9376 15068 9382
rect 15016 9318 15068 9324
rect 14832 9172 14884 9178
rect 14832 9114 14884 9120
rect 14832 8492 14884 8498
rect 14832 8434 14884 8440
rect 14844 8022 14872 8434
rect 14832 8016 14884 8022
rect 14832 7958 14884 7964
rect 14752 7806 14872 7834
rect 14740 7744 14792 7750
rect 14740 7686 14792 7692
rect 14752 7546 14780 7686
rect 14844 7546 14872 7806
rect 14740 7540 14792 7546
rect 14740 7482 14792 7488
rect 14832 7540 14884 7546
rect 14832 7482 14884 7488
rect 14740 6928 14792 6934
rect 14740 6870 14792 6876
rect 14752 6458 14780 6870
rect 14936 6866 14964 9318
rect 15016 9172 15068 9178
rect 15016 9114 15068 9120
rect 15028 6866 15056 9114
rect 15120 9081 15148 9687
rect 15106 9072 15162 9081
rect 15212 9042 15240 9823
rect 15304 9722 15332 9998
rect 15292 9716 15344 9722
rect 15292 9658 15344 9664
rect 15384 9444 15436 9450
rect 15580 9432 15608 11018
rect 15660 11008 15712 11014
rect 15660 10950 15712 10956
rect 15672 10742 15700 10950
rect 15660 10736 15712 10742
rect 15660 10678 15712 10684
rect 15672 10441 15700 10678
rect 15658 10432 15714 10441
rect 15658 10367 15714 10376
rect 15660 9988 15712 9994
rect 15660 9930 15712 9936
rect 15436 9404 15608 9432
rect 15384 9386 15436 9392
rect 15292 9376 15344 9382
rect 15292 9318 15344 9324
rect 15106 9007 15162 9016
rect 15200 9036 15252 9042
rect 15200 8978 15252 8984
rect 15200 8628 15252 8634
rect 15200 8570 15252 8576
rect 15106 8392 15162 8401
rect 15106 8327 15162 8336
rect 15120 7954 15148 8327
rect 15108 7948 15160 7954
rect 15108 7890 15160 7896
rect 15212 7449 15240 8570
rect 15198 7440 15254 7449
rect 15304 7410 15332 9318
rect 15384 9036 15436 9042
rect 15384 8978 15436 8984
rect 15396 8634 15424 8978
rect 15568 8968 15620 8974
rect 15568 8910 15620 8916
rect 15476 8832 15528 8838
rect 15476 8774 15528 8780
rect 15384 8628 15436 8634
rect 15384 8570 15436 8576
rect 15384 7812 15436 7818
rect 15384 7754 15436 7760
rect 15198 7375 15254 7384
rect 15292 7404 15344 7410
rect 15292 7346 15344 7352
rect 15396 7342 15424 7754
rect 15384 7336 15436 7342
rect 15384 7278 15436 7284
rect 15200 7200 15252 7206
rect 15200 7142 15252 7148
rect 14924 6860 14976 6866
rect 14924 6802 14976 6808
rect 15016 6860 15068 6866
rect 15068 6820 15148 6848
rect 15016 6802 15068 6808
rect 14832 6656 14884 6662
rect 14832 6598 14884 6604
rect 15016 6656 15068 6662
rect 15016 6598 15068 6604
rect 14740 6452 14792 6458
rect 14740 6394 14792 6400
rect 14844 6390 14872 6598
rect 14832 6384 14884 6390
rect 14832 6326 14884 6332
rect 14740 6316 14792 6322
rect 14740 6258 14792 6264
rect 14752 4729 14780 6258
rect 14830 5672 14886 5681
rect 14830 5607 14886 5616
rect 14844 5273 14872 5607
rect 14924 5568 14976 5574
rect 14924 5510 14976 5516
rect 14830 5264 14886 5273
rect 14830 5199 14886 5208
rect 14738 4720 14794 4729
rect 14738 4655 14794 4664
rect 14188 4140 14240 4146
rect 14188 4082 14240 4088
rect 14648 4140 14700 4146
rect 14648 4082 14700 4088
rect 13912 4004 13964 4010
rect 13912 3946 13964 3952
rect 13924 3670 13952 3946
rect 14844 3942 14872 5199
rect 14188 3936 14240 3942
rect 14188 3878 14240 3884
rect 14556 3936 14608 3942
rect 14556 3878 14608 3884
rect 14740 3936 14792 3942
rect 14740 3878 14792 3884
rect 14832 3936 14884 3942
rect 14832 3878 14884 3884
rect 14094 3768 14150 3777
rect 14094 3703 14150 3712
rect 13728 3664 13780 3670
rect 13728 3606 13780 3612
rect 13912 3664 13964 3670
rect 13912 3606 13964 3612
rect 13820 3596 13872 3602
rect 13820 3538 13872 3544
rect 13634 3496 13690 3505
rect 13634 3431 13636 3440
rect 13688 3431 13690 3440
rect 13728 3460 13780 3466
rect 13636 3402 13688 3408
rect 13728 3402 13780 3408
rect 13544 3392 13596 3398
rect 13648 3371 13676 3402
rect 13544 3334 13596 3340
rect 13174 3224 13230 3233
rect 13174 3159 13176 3168
rect 13228 3159 13230 3168
rect 13176 3130 13228 3136
rect 13082 2952 13138 2961
rect 13082 2887 13084 2896
rect 13136 2887 13138 2896
rect 13084 2858 13136 2864
rect 13556 2825 13584 3334
rect 13740 2922 13768 3402
rect 13832 3233 13860 3538
rect 14004 3528 14056 3534
rect 14004 3470 14056 3476
rect 14016 3233 14044 3470
rect 13818 3224 13874 3233
rect 13818 3159 13874 3168
rect 14002 3224 14058 3233
rect 14002 3159 14058 3168
rect 13832 3058 13860 3159
rect 14016 3058 14044 3159
rect 14108 3058 14136 3703
rect 14200 3670 14228 3878
rect 14188 3664 14240 3670
rect 14188 3606 14240 3612
rect 14568 3380 14596 3878
rect 14568 3352 14688 3380
rect 14294 3292 14602 3301
rect 14294 3290 14300 3292
rect 14356 3290 14380 3292
rect 14436 3290 14460 3292
rect 14516 3290 14540 3292
rect 14596 3290 14602 3292
rect 14356 3238 14358 3290
rect 14538 3238 14540 3290
rect 14294 3236 14300 3238
rect 14356 3236 14380 3238
rect 14436 3236 14460 3238
rect 14516 3236 14540 3238
rect 14596 3236 14602 3238
rect 14294 3227 14602 3236
rect 13820 3052 13872 3058
rect 13820 2994 13872 3000
rect 14004 3052 14056 3058
rect 14004 2994 14056 3000
rect 14096 3052 14148 3058
rect 14096 2994 14148 3000
rect 13728 2916 13780 2922
rect 13728 2858 13780 2864
rect 14372 2848 14424 2854
rect 13542 2816 13598 2825
rect 14372 2790 14424 2796
rect 13542 2751 13598 2760
rect 13542 2680 13598 2689
rect 13542 2615 13598 2624
rect 8944 2440 8996 2446
rect 8944 2382 8996 2388
rect 11152 2440 11204 2446
rect 11152 2382 11204 2388
rect 11520 2440 11572 2446
rect 11520 2382 11572 2388
rect 11704 2440 11756 2446
rect 11704 2382 11756 2388
rect 12440 2440 12492 2446
rect 12440 2382 12492 2388
rect 13556 2310 13584 2615
rect 13636 2576 13688 2582
rect 13636 2518 13688 2524
rect 13726 2544 13782 2553
rect 8668 2304 8720 2310
rect 8668 2246 8720 2252
rect 9496 2304 9548 2310
rect 9496 2246 9548 2252
rect 10324 2304 10376 2310
rect 10324 2246 10376 2252
rect 11152 2304 11204 2310
rect 11152 2246 11204 2252
rect 11980 2304 12032 2310
rect 11980 2246 12032 2252
rect 12716 2304 12768 2310
rect 12716 2246 12768 2252
rect 12808 2304 12860 2310
rect 12808 2246 12860 2252
rect 13544 2304 13596 2310
rect 13544 2246 13596 2252
rect 8114 2000 8170 2009
rect 8114 1935 8170 1944
rect 8680 800 8708 2246
rect 9508 800 9536 2246
rect 9846 2204 10154 2213
rect 9846 2202 9852 2204
rect 9908 2202 9932 2204
rect 9988 2202 10012 2204
rect 10068 2202 10092 2204
rect 10148 2202 10154 2204
rect 9908 2150 9910 2202
rect 10090 2150 10092 2202
rect 9846 2148 9852 2150
rect 9908 2148 9932 2150
rect 9988 2148 10012 2150
rect 10068 2148 10092 2150
rect 10148 2148 10154 2150
rect 9846 2139 10154 2148
rect 10336 800 10364 2246
rect 11164 800 11192 2246
rect 11992 800 12020 2246
rect 12728 1970 12756 2246
rect 12716 1964 12768 1970
rect 12716 1906 12768 1912
rect 12820 800 12848 2246
rect 13556 1902 13584 2246
rect 13544 1896 13596 1902
rect 13544 1838 13596 1844
rect 13648 800 13676 2518
rect 13726 2479 13782 2488
rect 13910 2544 13966 2553
rect 13910 2479 13966 2488
rect 13740 2446 13768 2479
rect 13728 2440 13780 2446
rect 13728 2382 13780 2388
rect 13728 2304 13780 2310
rect 13924 2292 13952 2479
rect 14384 2446 14412 2790
rect 14464 2644 14516 2650
rect 14464 2586 14516 2592
rect 14372 2440 14424 2446
rect 14372 2382 14424 2388
rect 14476 2310 14504 2586
rect 14660 2417 14688 3352
rect 14752 2990 14780 3878
rect 14832 3664 14884 3670
rect 14936 3652 14964 5510
rect 14884 3624 14964 3652
rect 14832 3606 14884 3612
rect 14924 3392 14976 3398
rect 14922 3360 14924 3369
rect 14976 3360 14978 3369
rect 14922 3295 14978 3304
rect 15028 3058 15056 6598
rect 15120 5778 15148 6820
rect 15212 6798 15240 7142
rect 15200 6792 15252 6798
rect 15200 6734 15252 6740
rect 15384 6656 15436 6662
rect 15384 6598 15436 6604
rect 15200 6452 15252 6458
rect 15200 6394 15252 6400
rect 15108 5772 15160 5778
rect 15108 5714 15160 5720
rect 15212 5642 15240 6394
rect 15292 6112 15344 6118
rect 15292 6054 15344 6060
rect 15200 5636 15252 5642
rect 15200 5578 15252 5584
rect 15106 5536 15162 5545
rect 15106 5471 15162 5480
rect 15120 5370 15148 5471
rect 15198 5400 15254 5409
rect 15108 5364 15160 5370
rect 15198 5335 15254 5344
rect 15108 5306 15160 5312
rect 15212 5302 15240 5335
rect 15200 5296 15252 5302
rect 15200 5238 15252 5244
rect 15304 5250 15332 6054
rect 15396 5846 15424 6598
rect 15488 6089 15516 8774
rect 15580 8566 15608 8910
rect 15568 8560 15620 8566
rect 15672 8537 15700 9930
rect 15752 9172 15804 9178
rect 15752 9114 15804 9120
rect 15568 8502 15620 8508
rect 15658 8528 15714 8537
rect 15658 8463 15714 8472
rect 15566 7984 15622 7993
rect 15566 7919 15622 7928
rect 15580 6633 15608 7919
rect 15764 7698 15792 9114
rect 15856 7818 15884 11036
rect 15936 11018 15988 11024
rect 16028 10804 16080 10810
rect 16028 10746 16080 10752
rect 15936 10668 15988 10674
rect 15936 10610 15988 10616
rect 15948 10470 15976 10610
rect 15936 10464 15988 10470
rect 15936 10406 15988 10412
rect 15948 10169 15976 10406
rect 16040 10198 16068 10746
rect 16028 10192 16080 10198
rect 15934 10160 15990 10169
rect 16028 10134 16080 10140
rect 15934 10095 15990 10104
rect 16026 8936 16082 8945
rect 16026 8871 16082 8880
rect 16040 8634 16068 8871
rect 16028 8628 16080 8634
rect 16028 8570 16080 8576
rect 16132 8514 16160 11222
rect 16212 11144 16264 11150
rect 16212 11086 16264 11092
rect 16224 10742 16252 11086
rect 16408 11082 16436 11614
rect 16592 11558 16620 11614
rect 16762 11591 16818 11600
rect 16580 11552 16632 11558
rect 16580 11494 16632 11500
rect 16518 11452 16826 11461
rect 16518 11450 16524 11452
rect 16580 11450 16604 11452
rect 16660 11450 16684 11452
rect 16740 11450 16764 11452
rect 16820 11450 16826 11452
rect 16580 11398 16582 11450
rect 16762 11398 16764 11450
rect 16518 11396 16524 11398
rect 16580 11396 16604 11398
rect 16660 11396 16684 11398
rect 16740 11396 16764 11398
rect 16820 11396 16826 11398
rect 16518 11387 16826 11396
rect 16396 11076 16448 11082
rect 16396 11018 16448 11024
rect 16212 10736 16264 10742
rect 16212 10678 16264 10684
rect 16304 10668 16356 10674
rect 16304 10610 16356 10616
rect 16212 10464 16264 10470
rect 16212 10406 16264 10412
rect 16040 8486 16160 8514
rect 15844 7812 15896 7818
rect 15844 7754 15896 7760
rect 15936 7744 15988 7750
rect 15672 7670 15792 7698
rect 15934 7712 15936 7721
rect 15988 7712 15990 7721
rect 15566 6624 15622 6633
rect 15566 6559 15622 6568
rect 15474 6080 15530 6089
rect 15474 6015 15530 6024
rect 15384 5840 15436 5846
rect 15384 5782 15436 5788
rect 15580 5794 15608 6559
rect 15672 6458 15700 7670
rect 15934 7647 15990 7656
rect 15752 7540 15804 7546
rect 15752 7482 15804 7488
rect 15936 7540 15988 7546
rect 15936 7482 15988 7488
rect 15764 7342 15792 7482
rect 15752 7336 15804 7342
rect 15752 7278 15804 7284
rect 15764 7206 15792 7278
rect 15752 7200 15804 7206
rect 15752 7142 15804 7148
rect 15948 7002 15976 7482
rect 15936 6996 15988 7002
rect 15936 6938 15988 6944
rect 15948 6798 15976 6938
rect 15936 6792 15988 6798
rect 15936 6734 15988 6740
rect 15752 6656 15804 6662
rect 15752 6598 15804 6604
rect 15764 6458 15792 6598
rect 15660 6452 15712 6458
rect 15660 6394 15712 6400
rect 15752 6452 15804 6458
rect 15752 6394 15804 6400
rect 15672 6338 15700 6394
rect 15672 6310 15884 6338
rect 15752 6248 15804 6254
rect 15752 6190 15804 6196
rect 15764 5914 15792 6190
rect 15752 5908 15804 5914
rect 15752 5850 15804 5856
rect 15580 5766 15792 5794
rect 15108 5228 15160 5234
rect 15108 5170 15160 5176
rect 15120 4622 15148 5170
rect 15108 4616 15160 4622
rect 15108 4558 15160 4564
rect 15212 4554 15240 5238
rect 15304 5222 15700 5250
rect 15566 5128 15622 5137
rect 15384 5092 15436 5098
rect 15566 5063 15622 5072
rect 15384 5034 15436 5040
rect 15292 5024 15344 5030
rect 15292 4966 15344 4972
rect 15200 4548 15252 4554
rect 15200 4490 15252 4496
rect 15304 4049 15332 4966
rect 15396 4826 15424 5034
rect 15384 4820 15436 4826
rect 15384 4762 15436 4768
rect 15476 4820 15528 4826
rect 15476 4762 15528 4768
rect 15382 4448 15438 4457
rect 15382 4383 15438 4392
rect 15290 4040 15346 4049
rect 15290 3975 15346 3984
rect 15108 3936 15160 3942
rect 15108 3878 15160 3884
rect 15292 3936 15344 3942
rect 15292 3878 15344 3884
rect 15016 3052 15068 3058
rect 15016 2994 15068 3000
rect 14740 2984 14792 2990
rect 14740 2926 14792 2932
rect 15120 2922 15148 3878
rect 15304 3534 15332 3878
rect 15292 3528 15344 3534
rect 15292 3470 15344 3476
rect 15200 3188 15252 3194
rect 15200 3130 15252 3136
rect 15212 3058 15240 3130
rect 15200 3052 15252 3058
rect 15200 2994 15252 3000
rect 15108 2916 15160 2922
rect 15108 2858 15160 2864
rect 15016 2848 15068 2854
rect 15016 2790 15068 2796
rect 15028 2446 15056 2790
rect 15200 2644 15252 2650
rect 15396 2632 15424 4383
rect 15488 3777 15516 4762
rect 15474 3768 15530 3777
rect 15474 3703 15530 3712
rect 15580 3534 15608 5063
rect 15568 3528 15620 3534
rect 15568 3470 15620 3476
rect 15476 3052 15528 3058
rect 15476 2994 15528 3000
rect 15252 2604 15424 2632
rect 15200 2586 15252 2592
rect 15016 2440 15068 2446
rect 14646 2408 14702 2417
rect 15016 2382 15068 2388
rect 15488 2378 15516 2994
rect 15672 2990 15700 5222
rect 15764 5012 15792 5766
rect 15856 5137 15884 6310
rect 15936 6112 15988 6118
rect 15936 6054 15988 6060
rect 15948 5778 15976 6054
rect 15936 5772 15988 5778
rect 15936 5714 15988 5720
rect 15936 5364 15988 5370
rect 15936 5306 15988 5312
rect 15842 5128 15898 5137
rect 15842 5063 15898 5072
rect 15764 4984 15884 5012
rect 15752 4480 15804 4486
rect 15752 4422 15804 4428
rect 15764 4214 15792 4422
rect 15752 4208 15804 4214
rect 15752 4150 15804 4156
rect 15752 3052 15804 3058
rect 15752 2994 15804 3000
rect 15660 2984 15712 2990
rect 15764 2961 15792 2994
rect 15660 2926 15712 2932
rect 15750 2952 15806 2961
rect 15568 2916 15620 2922
rect 15750 2887 15806 2896
rect 15568 2858 15620 2864
rect 15580 2582 15608 2858
rect 15660 2848 15712 2854
rect 15660 2790 15712 2796
rect 15568 2576 15620 2582
rect 15568 2518 15620 2524
rect 14646 2343 14702 2352
rect 15476 2372 15528 2378
rect 15476 2314 15528 2320
rect 13780 2264 13952 2292
rect 14004 2304 14056 2310
rect 13728 2246 13780 2252
rect 14004 2246 14056 2252
rect 14464 2304 14516 2310
rect 14464 2246 14516 2252
rect 14648 2304 14700 2310
rect 14648 2246 14700 2252
rect 15292 2304 15344 2310
rect 15292 2246 15344 2252
rect 14016 2009 14044 2246
rect 14294 2204 14602 2213
rect 14294 2202 14300 2204
rect 14356 2202 14380 2204
rect 14436 2202 14460 2204
rect 14516 2202 14540 2204
rect 14596 2202 14602 2204
rect 14356 2150 14358 2202
rect 14538 2150 14540 2202
rect 14294 2148 14300 2150
rect 14356 2148 14380 2150
rect 14436 2148 14460 2150
rect 14516 2148 14540 2150
rect 14596 2148 14602 2150
rect 14294 2139 14602 2148
rect 14002 2000 14058 2009
rect 14002 1935 14058 1944
rect 14660 1170 14688 2246
rect 14476 1142 14688 1170
rect 14476 800 14504 1142
rect 15304 800 15332 2246
rect 15672 2106 15700 2790
rect 15856 2774 15884 4984
rect 15948 3942 15976 5306
rect 16040 4690 16068 8486
rect 16120 8356 16172 8362
rect 16120 8298 16172 8304
rect 16132 7993 16160 8298
rect 16118 7984 16174 7993
rect 16118 7919 16174 7928
rect 16118 7712 16174 7721
rect 16118 7647 16174 7656
rect 16132 6866 16160 7647
rect 16224 7410 16252 10406
rect 16316 9625 16344 10610
rect 16518 10364 16826 10373
rect 16518 10362 16524 10364
rect 16580 10362 16604 10364
rect 16660 10362 16684 10364
rect 16740 10362 16764 10364
rect 16820 10362 16826 10364
rect 16580 10310 16582 10362
rect 16762 10310 16764 10362
rect 16518 10308 16524 10310
rect 16580 10308 16604 10310
rect 16660 10308 16684 10310
rect 16740 10308 16764 10310
rect 16820 10308 16826 10310
rect 16518 10299 16826 10308
rect 16488 9920 16540 9926
rect 16488 9862 16540 9868
rect 16500 9722 16528 9862
rect 16488 9716 16540 9722
rect 16488 9658 16540 9664
rect 16302 9616 16358 9625
rect 16302 9551 16358 9560
rect 16518 9276 16826 9285
rect 16518 9274 16524 9276
rect 16580 9274 16604 9276
rect 16660 9274 16684 9276
rect 16740 9274 16764 9276
rect 16820 9274 16826 9276
rect 16580 9222 16582 9274
rect 16762 9222 16764 9274
rect 16518 9220 16524 9222
rect 16580 9220 16604 9222
rect 16660 9220 16684 9222
rect 16740 9220 16764 9222
rect 16820 9220 16826 9222
rect 16518 9211 16826 9220
rect 16868 9178 16896 13194
rect 17144 12918 17172 13330
rect 17132 12912 17184 12918
rect 17132 12854 17184 12860
rect 17040 12640 17092 12646
rect 17040 12582 17092 12588
rect 16948 11756 17000 11762
rect 16948 11698 17000 11704
rect 16960 11082 16988 11698
rect 16948 11076 17000 11082
rect 16948 11018 17000 11024
rect 16948 10532 17000 10538
rect 16948 10474 17000 10480
rect 16960 10033 16988 10474
rect 16946 10024 17002 10033
rect 16946 9959 17002 9968
rect 16948 9376 17000 9382
rect 16948 9318 17000 9324
rect 16304 9172 16356 9178
rect 16304 9114 16356 9120
rect 16856 9172 16908 9178
rect 16856 9114 16908 9120
rect 16316 8838 16344 9114
rect 16396 8968 16448 8974
rect 16396 8910 16448 8916
rect 16304 8832 16356 8838
rect 16304 8774 16356 8780
rect 16304 8492 16356 8498
rect 16304 8434 16356 8440
rect 16212 7404 16264 7410
rect 16212 7346 16264 7352
rect 16120 6860 16172 6866
rect 16120 6802 16172 6808
rect 16212 6792 16264 6798
rect 16212 6734 16264 6740
rect 16120 6724 16172 6730
rect 16120 6666 16172 6672
rect 16132 5370 16160 6666
rect 16224 5817 16252 6734
rect 16210 5808 16266 5817
rect 16210 5743 16266 5752
rect 16212 5704 16264 5710
rect 16212 5646 16264 5652
rect 16224 5370 16252 5646
rect 16120 5364 16172 5370
rect 16120 5306 16172 5312
rect 16212 5364 16264 5370
rect 16212 5306 16264 5312
rect 16212 5160 16264 5166
rect 16212 5102 16264 5108
rect 16120 5024 16172 5030
rect 16120 4966 16172 4972
rect 16028 4684 16080 4690
rect 16028 4626 16080 4632
rect 16040 4434 16068 4626
rect 16132 4622 16160 4966
rect 16120 4616 16172 4622
rect 16120 4558 16172 4564
rect 16224 4457 16252 5102
rect 16210 4448 16266 4457
rect 16040 4406 16160 4434
rect 16132 4078 16160 4406
rect 16210 4383 16266 4392
rect 16120 4072 16172 4078
rect 16120 4014 16172 4020
rect 16212 4072 16264 4078
rect 16212 4014 16264 4020
rect 15936 3936 15988 3942
rect 15936 3878 15988 3884
rect 16224 3738 16252 4014
rect 16316 3738 16344 8434
rect 16408 7954 16436 8910
rect 16518 8188 16826 8197
rect 16518 8186 16524 8188
rect 16580 8186 16604 8188
rect 16660 8186 16684 8188
rect 16740 8186 16764 8188
rect 16820 8186 16826 8188
rect 16580 8134 16582 8186
rect 16762 8134 16764 8186
rect 16518 8132 16524 8134
rect 16580 8132 16604 8134
rect 16660 8132 16684 8134
rect 16740 8132 16764 8134
rect 16820 8132 16826 8134
rect 16518 8123 16826 8132
rect 16868 7970 16896 9114
rect 16960 9081 16988 9318
rect 16946 9072 17002 9081
rect 16946 9007 17002 9016
rect 16948 8356 17000 8362
rect 16948 8298 17000 8304
rect 16960 8265 16988 8298
rect 16946 8256 17002 8265
rect 16946 8191 17002 8200
rect 16396 7948 16448 7954
rect 16868 7942 16988 7970
rect 16396 7890 16448 7896
rect 16856 7880 16908 7886
rect 16856 7822 16908 7828
rect 16488 7812 16540 7818
rect 16488 7754 16540 7760
rect 16394 7712 16450 7721
rect 16394 7647 16450 7656
rect 16408 7546 16436 7647
rect 16396 7540 16448 7546
rect 16396 7482 16448 7488
rect 16500 7188 16528 7754
rect 16408 7160 16528 7188
rect 16408 5778 16436 7160
rect 16518 7100 16826 7109
rect 16518 7098 16524 7100
rect 16580 7098 16604 7100
rect 16660 7098 16684 7100
rect 16740 7098 16764 7100
rect 16820 7098 16826 7100
rect 16580 7046 16582 7098
rect 16762 7046 16764 7098
rect 16518 7044 16524 7046
rect 16580 7044 16604 7046
rect 16660 7044 16684 7046
rect 16740 7044 16764 7046
rect 16820 7044 16826 7046
rect 16518 7035 16826 7044
rect 16868 7002 16896 7822
rect 16856 6996 16908 7002
rect 16856 6938 16908 6944
rect 16856 6860 16908 6866
rect 16856 6802 16908 6808
rect 16672 6792 16724 6798
rect 16672 6734 16724 6740
rect 16684 6186 16712 6734
rect 16672 6180 16724 6186
rect 16672 6122 16724 6128
rect 16518 6012 16826 6021
rect 16518 6010 16524 6012
rect 16580 6010 16604 6012
rect 16660 6010 16684 6012
rect 16740 6010 16764 6012
rect 16820 6010 16826 6012
rect 16580 5958 16582 6010
rect 16762 5958 16764 6010
rect 16518 5956 16524 5958
rect 16580 5956 16604 5958
rect 16660 5956 16684 5958
rect 16740 5956 16764 5958
rect 16820 5956 16826 5958
rect 16518 5947 16826 5956
rect 16868 5914 16896 6802
rect 16960 6798 16988 7942
rect 17052 6866 17080 12582
rect 17144 12306 17172 12854
rect 17132 12300 17184 12306
rect 17132 12242 17184 12248
rect 17132 12096 17184 12102
rect 17132 12038 17184 12044
rect 17144 11257 17172 12038
rect 17130 11248 17186 11257
rect 17130 11183 17186 11192
rect 17132 11076 17184 11082
rect 17132 11018 17184 11024
rect 17144 10554 17172 11018
rect 17236 10674 17264 13631
rect 17408 13388 17460 13394
rect 17408 13330 17460 13336
rect 17420 12918 17448 13330
rect 17498 13152 17554 13161
rect 17498 13087 17554 13096
rect 17408 12912 17460 12918
rect 17408 12854 17460 12860
rect 17316 12844 17368 12850
rect 17316 12786 17368 12792
rect 17328 12434 17356 12786
rect 17328 12406 17448 12434
rect 17316 12368 17368 12374
rect 17316 12310 17368 12316
rect 17328 11762 17356 12310
rect 17316 11756 17368 11762
rect 17316 11698 17368 11704
rect 17224 10668 17276 10674
rect 17224 10610 17276 10616
rect 17144 10526 17264 10554
rect 17132 10464 17184 10470
rect 17132 10406 17184 10412
rect 17144 7818 17172 10406
rect 17236 10033 17264 10526
rect 17316 10056 17368 10062
rect 17222 10024 17278 10033
rect 17316 9998 17368 10004
rect 17222 9959 17278 9968
rect 17328 9518 17356 9998
rect 17316 9512 17368 9518
rect 17222 9480 17278 9489
rect 17316 9454 17368 9460
rect 17222 9415 17278 9424
rect 17236 8430 17264 9415
rect 17328 9178 17356 9454
rect 17316 9172 17368 9178
rect 17316 9114 17368 9120
rect 17224 8424 17276 8430
rect 17224 8366 17276 8372
rect 17316 8424 17368 8430
rect 17316 8366 17368 8372
rect 17328 8129 17356 8366
rect 17420 8294 17448 12406
rect 17512 10742 17540 13087
rect 17604 12374 17632 14282
rect 17776 14272 17828 14278
rect 17776 14214 17828 14220
rect 17788 13326 17816 14214
rect 17880 13530 17908 16400
rect 18328 14952 18380 14958
rect 18328 14894 18380 14900
rect 18340 14618 18368 14894
rect 18328 14612 18380 14618
rect 18328 14554 18380 14560
rect 18696 14408 18748 14414
rect 18142 14376 18198 14385
rect 18696 14350 18748 14356
rect 18142 14311 18144 14320
rect 18196 14311 18198 14320
rect 18604 14340 18656 14346
rect 18144 14282 18196 14288
rect 18604 14282 18656 14288
rect 18420 13932 18472 13938
rect 18420 13874 18472 13880
rect 18328 13864 18380 13870
rect 18328 13806 18380 13812
rect 18052 13728 18104 13734
rect 18052 13670 18104 13676
rect 17868 13524 17920 13530
rect 17868 13466 17920 13472
rect 17776 13320 17828 13326
rect 17776 13262 17828 13268
rect 17776 13184 17828 13190
rect 17776 13126 17828 13132
rect 17592 12368 17644 12374
rect 17592 12310 17644 12316
rect 17684 12232 17736 12238
rect 17684 12174 17736 12180
rect 17592 12164 17644 12170
rect 17592 12106 17644 12112
rect 17604 11801 17632 12106
rect 17590 11792 17646 11801
rect 17590 11727 17646 11736
rect 17696 11558 17724 12174
rect 17788 11762 17816 13126
rect 17866 12608 17922 12617
rect 17866 12543 17922 12552
rect 17776 11756 17828 11762
rect 17776 11698 17828 11704
rect 17684 11552 17736 11558
rect 17684 11494 17736 11500
rect 17696 11257 17724 11494
rect 17682 11248 17738 11257
rect 17682 11183 17738 11192
rect 17684 11144 17736 11150
rect 17788 11121 17816 11698
rect 17684 11086 17736 11092
rect 17774 11112 17830 11121
rect 17696 10985 17724 11086
rect 17774 11047 17830 11056
rect 17682 10976 17738 10985
rect 17682 10911 17738 10920
rect 17776 10804 17828 10810
rect 17776 10746 17828 10752
rect 17500 10736 17552 10742
rect 17500 10678 17552 10684
rect 17512 9722 17540 10678
rect 17592 10600 17644 10606
rect 17592 10542 17644 10548
rect 17684 10600 17736 10606
rect 17684 10542 17736 10548
rect 17604 10198 17632 10542
rect 17696 10441 17724 10542
rect 17682 10432 17738 10441
rect 17682 10367 17738 10376
rect 17696 10266 17724 10367
rect 17684 10260 17736 10266
rect 17684 10202 17736 10208
rect 17592 10192 17644 10198
rect 17590 10160 17592 10169
rect 17644 10160 17646 10169
rect 17590 10095 17646 10104
rect 17682 10024 17738 10033
rect 17682 9959 17738 9968
rect 17500 9716 17552 9722
rect 17500 9658 17552 9664
rect 17592 9580 17644 9586
rect 17592 9522 17644 9528
rect 17500 9376 17552 9382
rect 17500 9318 17552 9324
rect 17512 8838 17540 9318
rect 17604 8945 17632 9522
rect 17590 8936 17646 8945
rect 17590 8871 17646 8880
rect 17500 8832 17552 8838
rect 17500 8774 17552 8780
rect 17512 8498 17540 8774
rect 17500 8492 17552 8498
rect 17500 8434 17552 8440
rect 17408 8288 17460 8294
rect 17408 8230 17460 8236
rect 17314 8120 17370 8129
rect 17314 8055 17370 8064
rect 17420 7954 17448 8230
rect 17408 7948 17460 7954
rect 17408 7890 17460 7896
rect 17500 7948 17552 7954
rect 17500 7890 17552 7896
rect 17132 7812 17184 7818
rect 17132 7754 17184 7760
rect 17224 7744 17276 7750
rect 17224 7686 17276 7692
rect 17316 7744 17368 7750
rect 17316 7686 17368 7692
rect 17132 7336 17184 7342
rect 17132 7278 17184 7284
rect 17144 7002 17172 7278
rect 17132 6996 17184 7002
rect 17132 6938 17184 6944
rect 17040 6860 17092 6866
rect 17040 6802 17092 6808
rect 16948 6792 17000 6798
rect 16948 6734 17000 6740
rect 17040 6724 17092 6730
rect 17040 6666 17092 6672
rect 16946 6216 17002 6225
rect 16946 6151 17002 6160
rect 16856 5908 16908 5914
rect 16856 5850 16908 5856
rect 16868 5778 16896 5850
rect 16396 5772 16448 5778
rect 16396 5714 16448 5720
rect 16856 5772 16908 5778
rect 16856 5714 16908 5720
rect 16764 5636 16816 5642
rect 16764 5578 16816 5584
rect 16580 5568 16632 5574
rect 16580 5510 16632 5516
rect 16592 5012 16620 5510
rect 16776 5166 16804 5578
rect 16960 5166 16988 6151
rect 17052 5710 17080 6666
rect 17236 6254 17264 7686
rect 17328 7546 17356 7686
rect 17512 7585 17540 7890
rect 17498 7576 17554 7585
rect 17316 7540 17368 7546
rect 17498 7511 17554 7520
rect 17316 7482 17368 7488
rect 17604 7478 17632 8871
rect 17592 7472 17644 7478
rect 17592 7414 17644 7420
rect 17408 7404 17460 7410
rect 17408 7346 17460 7352
rect 17316 6860 17368 6866
rect 17316 6802 17368 6808
rect 17132 6248 17184 6254
rect 17132 6190 17184 6196
rect 17224 6248 17276 6254
rect 17224 6190 17276 6196
rect 17040 5704 17092 5710
rect 17144 5681 17172 6190
rect 17040 5646 17092 5652
rect 17130 5672 17186 5681
rect 17130 5607 17186 5616
rect 17224 5636 17276 5642
rect 17224 5578 17276 5584
rect 17040 5568 17092 5574
rect 17038 5536 17040 5545
rect 17092 5536 17094 5545
rect 17038 5471 17094 5480
rect 16764 5160 16816 5166
rect 16948 5160 17000 5166
rect 16764 5102 16816 5108
rect 16854 5128 16910 5137
rect 16948 5102 17000 5108
rect 16854 5063 16910 5072
rect 16408 4984 16620 5012
rect 16408 4146 16436 4984
rect 16518 4924 16826 4933
rect 16518 4922 16524 4924
rect 16580 4922 16604 4924
rect 16660 4922 16684 4924
rect 16740 4922 16764 4924
rect 16820 4922 16826 4924
rect 16580 4870 16582 4922
rect 16762 4870 16764 4922
rect 16518 4868 16524 4870
rect 16580 4868 16604 4870
rect 16660 4868 16684 4870
rect 16740 4868 16764 4870
rect 16820 4868 16826 4870
rect 16518 4859 16826 4868
rect 16762 4720 16818 4729
rect 16762 4655 16818 4664
rect 16580 4548 16632 4554
rect 16580 4490 16632 4496
rect 16396 4140 16448 4146
rect 16396 4082 16448 4088
rect 16592 3992 16620 4490
rect 16776 4486 16804 4655
rect 16868 4622 16896 5063
rect 17052 4826 17080 5471
rect 17132 5364 17184 5370
rect 17132 5306 17184 5312
rect 17040 4820 17092 4826
rect 17040 4762 17092 4768
rect 16946 4720 17002 4729
rect 16946 4655 17002 4664
rect 16856 4616 16908 4622
rect 16856 4558 16908 4564
rect 16764 4480 16816 4486
rect 16764 4422 16816 4428
rect 16764 4140 16816 4146
rect 16764 4082 16816 4088
rect 16776 4010 16804 4082
rect 16960 4010 16988 4655
rect 17040 4616 17092 4622
rect 17040 4558 17092 4564
rect 16408 3964 16620 3992
rect 16764 4004 16816 4010
rect 16212 3732 16264 3738
rect 16212 3674 16264 3680
rect 16304 3732 16356 3738
rect 16304 3674 16356 3680
rect 15934 3496 15990 3505
rect 15934 3431 15990 3440
rect 16118 3496 16174 3505
rect 16118 3431 16174 3440
rect 15948 3176 15976 3431
rect 16132 3398 16160 3431
rect 16408 3398 16436 3964
rect 16764 3946 16816 3952
rect 16948 4004 17000 4010
rect 16948 3946 17000 3952
rect 16856 3936 16908 3942
rect 16856 3878 16908 3884
rect 16518 3836 16826 3845
rect 16518 3834 16524 3836
rect 16580 3834 16604 3836
rect 16660 3834 16684 3836
rect 16740 3834 16764 3836
rect 16820 3834 16826 3836
rect 16580 3782 16582 3834
rect 16762 3782 16764 3834
rect 16518 3780 16524 3782
rect 16580 3780 16604 3782
rect 16660 3780 16684 3782
rect 16740 3780 16764 3782
rect 16820 3780 16826 3782
rect 16518 3771 16826 3780
rect 16670 3632 16726 3641
rect 16670 3567 16726 3576
rect 16684 3534 16712 3567
rect 16672 3528 16724 3534
rect 16672 3470 16724 3476
rect 16764 3528 16816 3534
rect 16764 3470 16816 3476
rect 16120 3392 16172 3398
rect 16120 3334 16172 3340
rect 16396 3392 16448 3398
rect 16776 3369 16804 3470
rect 16396 3334 16448 3340
rect 16762 3360 16818 3369
rect 16762 3295 16818 3304
rect 16210 3224 16266 3233
rect 16868 3194 16896 3878
rect 16948 3392 17000 3398
rect 16946 3360 16948 3369
rect 17000 3360 17002 3369
rect 16946 3295 17002 3304
rect 17052 3194 17080 4558
rect 17144 4321 17172 5306
rect 17130 4312 17186 4321
rect 17130 4247 17186 4256
rect 17132 4140 17184 4146
rect 17132 4082 17184 4088
rect 17144 3670 17172 4082
rect 17132 3664 17184 3670
rect 17132 3606 17184 3612
rect 15948 3148 16160 3176
rect 16210 3159 16212 3168
rect 16028 3052 16080 3058
rect 16132 3040 16160 3148
rect 16264 3159 16266 3168
rect 16856 3188 16908 3194
rect 16212 3130 16264 3136
rect 16856 3130 16908 3136
rect 17040 3188 17092 3194
rect 17040 3130 17092 3136
rect 17236 3126 17264 5578
rect 17328 5234 17356 6802
rect 17420 6458 17448 7346
rect 17696 6882 17724 9959
rect 17512 6854 17724 6882
rect 17408 6452 17460 6458
rect 17408 6394 17460 6400
rect 17408 6316 17460 6322
rect 17408 6258 17460 6264
rect 17316 5228 17368 5234
rect 17316 5170 17368 5176
rect 17314 4992 17370 5001
rect 17314 4927 17370 4936
rect 17328 4010 17356 4927
rect 17420 4214 17448 6258
rect 17512 5710 17540 6854
rect 17592 6792 17644 6798
rect 17592 6734 17644 6740
rect 17604 6186 17632 6734
rect 17684 6656 17736 6662
rect 17682 6624 17684 6633
rect 17736 6624 17738 6633
rect 17682 6559 17738 6568
rect 17788 6474 17816 10746
rect 17880 10062 17908 12543
rect 18064 12442 18092 13670
rect 18234 13288 18290 13297
rect 18234 13223 18290 13232
rect 18248 12918 18276 13223
rect 18236 12912 18288 12918
rect 18236 12854 18288 12860
rect 18052 12436 18104 12442
rect 18052 12378 18104 12384
rect 18064 11082 18092 12378
rect 18142 12336 18198 12345
rect 18142 12271 18144 12280
rect 18196 12271 18198 12280
rect 18144 12242 18196 12248
rect 18236 12232 18288 12238
rect 18236 12174 18288 12180
rect 18248 11830 18276 12174
rect 18236 11824 18288 11830
rect 18236 11766 18288 11772
rect 18236 11280 18288 11286
rect 18236 11222 18288 11228
rect 18052 11076 18104 11082
rect 18052 11018 18104 11024
rect 17958 10704 18014 10713
rect 17958 10639 18014 10648
rect 18052 10668 18104 10674
rect 17972 10130 18000 10639
rect 18052 10610 18104 10616
rect 17960 10124 18012 10130
rect 17960 10066 18012 10072
rect 17868 10056 17920 10062
rect 17868 9998 17920 10004
rect 17972 9738 18000 10066
rect 17880 9722 18000 9738
rect 18064 9722 18092 10610
rect 18144 10600 18196 10606
rect 18144 10542 18196 10548
rect 18156 9761 18184 10542
rect 18142 9752 18198 9761
rect 17868 9716 18000 9722
rect 17920 9710 18000 9716
rect 18052 9716 18104 9722
rect 17868 9658 17920 9664
rect 18142 9687 18198 9696
rect 18052 9658 18104 9664
rect 17868 9512 17920 9518
rect 17866 9480 17868 9489
rect 17920 9480 17922 9489
rect 17866 9415 17922 9424
rect 17960 9444 18012 9450
rect 17880 8401 17908 9415
rect 17960 9386 18012 9392
rect 17866 8392 17922 8401
rect 17866 8327 17922 8336
rect 17868 8288 17920 8294
rect 17868 8230 17920 8236
rect 17880 7546 17908 8230
rect 17868 7540 17920 7546
rect 17868 7482 17920 7488
rect 17868 7404 17920 7410
rect 17868 7346 17920 7352
rect 17880 6934 17908 7346
rect 17868 6928 17920 6934
rect 17868 6870 17920 6876
rect 17972 6644 18000 9386
rect 18052 8628 18104 8634
rect 18052 8570 18104 8576
rect 18064 7002 18092 8570
rect 18248 8498 18276 11222
rect 18340 10577 18368 13806
rect 18432 12073 18460 13874
rect 18512 12912 18564 12918
rect 18512 12854 18564 12860
rect 18418 12064 18474 12073
rect 18418 11999 18474 12008
rect 18420 11824 18472 11830
rect 18420 11766 18472 11772
rect 18432 10713 18460 11766
rect 18524 11529 18552 12854
rect 18616 12345 18644 14282
rect 18708 12434 18736 14350
rect 18708 12406 18828 12434
rect 18602 12336 18658 12345
rect 18602 12271 18658 12280
rect 18510 11520 18566 11529
rect 18510 11455 18566 11464
rect 18604 11144 18656 11150
rect 18604 11086 18656 11092
rect 18512 11076 18564 11082
rect 18512 11018 18564 11024
rect 18418 10704 18474 10713
rect 18418 10639 18474 10648
rect 18326 10568 18382 10577
rect 18326 10503 18382 10512
rect 18236 8492 18288 8498
rect 18236 8434 18288 8440
rect 18340 8378 18368 10503
rect 18420 9648 18472 9654
rect 18420 9590 18472 9596
rect 18432 9353 18460 9590
rect 18418 9344 18474 9353
rect 18418 9279 18474 9288
rect 18418 8800 18474 8809
rect 18418 8735 18474 8744
rect 18432 8634 18460 8735
rect 18420 8628 18472 8634
rect 18420 8570 18472 8576
rect 18418 8528 18474 8537
rect 18418 8463 18474 8472
rect 18248 8350 18368 8378
rect 18248 8022 18276 8350
rect 18328 8288 18380 8294
rect 18328 8230 18380 8236
rect 18236 8016 18288 8022
rect 18236 7958 18288 7964
rect 18144 7948 18196 7954
rect 18144 7890 18196 7896
rect 18156 7342 18184 7890
rect 18236 7880 18288 7886
rect 18236 7822 18288 7828
rect 18144 7336 18196 7342
rect 18144 7278 18196 7284
rect 18156 7002 18184 7278
rect 18052 6996 18104 7002
rect 18052 6938 18104 6944
rect 18144 6996 18196 7002
rect 18144 6938 18196 6944
rect 18142 6896 18198 6905
rect 18142 6831 18198 6840
rect 18052 6656 18104 6662
rect 17972 6616 18052 6644
rect 18052 6598 18104 6604
rect 17696 6446 17816 6474
rect 17592 6180 17644 6186
rect 17592 6122 17644 6128
rect 17592 5840 17644 5846
rect 17590 5808 17592 5817
rect 17644 5808 17646 5817
rect 17590 5743 17646 5752
rect 17500 5704 17552 5710
rect 17696 5658 17724 6446
rect 17774 6352 17830 6361
rect 17774 6287 17830 6296
rect 17500 5646 17552 5652
rect 17512 5166 17540 5646
rect 17604 5642 17724 5658
rect 17604 5636 17736 5642
rect 17604 5630 17684 5636
rect 17604 5409 17632 5630
rect 17684 5578 17736 5584
rect 17682 5536 17738 5545
rect 17682 5471 17738 5480
rect 17590 5400 17646 5409
rect 17590 5335 17646 5344
rect 17500 5160 17552 5166
rect 17500 5102 17552 5108
rect 17592 5024 17644 5030
rect 17592 4966 17644 4972
rect 17498 4856 17554 4865
rect 17498 4791 17554 4800
rect 17512 4486 17540 4791
rect 17500 4480 17552 4486
rect 17500 4422 17552 4428
rect 17408 4208 17460 4214
rect 17408 4150 17460 4156
rect 17316 4004 17368 4010
rect 17316 3946 17368 3952
rect 17316 3664 17368 3670
rect 17314 3632 17316 3641
rect 17368 3632 17370 3641
rect 17512 3618 17540 4422
rect 17604 4282 17632 4966
rect 17696 4282 17724 5471
rect 17788 4826 17816 6287
rect 17868 6180 17920 6186
rect 17868 6122 17920 6128
rect 17880 5914 17908 6122
rect 18050 6080 18106 6089
rect 18050 6015 18106 6024
rect 17868 5908 17920 5914
rect 17868 5850 17920 5856
rect 17880 5778 17908 5850
rect 17868 5772 17920 5778
rect 17868 5714 17920 5720
rect 17866 5264 17922 5273
rect 17866 5199 17922 5208
rect 17960 5228 18012 5234
rect 17776 4820 17828 4826
rect 17776 4762 17828 4768
rect 17592 4276 17644 4282
rect 17592 4218 17644 4224
rect 17684 4276 17736 4282
rect 17684 4218 17736 4224
rect 17682 4176 17738 4185
rect 17682 4111 17738 4120
rect 17696 3738 17724 4111
rect 17774 4040 17830 4049
rect 17774 3975 17830 3984
rect 17684 3732 17736 3738
rect 17684 3674 17736 3680
rect 17314 3567 17370 3576
rect 17420 3590 17540 3618
rect 17224 3120 17276 3126
rect 17130 3088 17186 3097
rect 16396 3052 16448 3058
rect 16132 3012 16396 3040
rect 16028 2994 16080 3000
rect 17224 3062 17276 3068
rect 17130 3023 17132 3032
rect 16396 2994 16448 3000
rect 17184 3023 17186 3032
rect 17132 2994 17184 3000
rect 15764 2746 15884 2774
rect 15764 2650 15792 2746
rect 15752 2644 15804 2650
rect 15752 2586 15804 2592
rect 15660 2100 15712 2106
rect 15660 2042 15712 2048
rect 16040 1902 16068 2994
rect 16578 2952 16634 2961
rect 16578 2887 16580 2896
rect 16632 2887 16634 2896
rect 16580 2858 16632 2864
rect 17316 2848 17368 2854
rect 17316 2790 17368 2796
rect 16518 2748 16826 2757
rect 16518 2746 16524 2748
rect 16580 2746 16604 2748
rect 16660 2746 16684 2748
rect 16740 2746 16764 2748
rect 16820 2746 16826 2748
rect 16580 2694 16582 2746
rect 16762 2694 16764 2746
rect 16518 2692 16524 2694
rect 16580 2692 16604 2694
rect 16660 2692 16684 2694
rect 16740 2692 16764 2694
rect 16820 2692 16826 2694
rect 16302 2680 16358 2689
rect 16518 2683 16826 2692
rect 16302 2615 16358 2624
rect 16120 2508 16172 2514
rect 16120 2450 16172 2456
rect 16132 1970 16160 2450
rect 16316 2428 16344 2615
rect 17328 2553 17356 2790
rect 17038 2544 17094 2553
rect 17038 2479 17094 2488
rect 17314 2544 17370 2553
rect 17420 2514 17448 3590
rect 17788 3534 17816 3975
rect 17880 3738 17908 5199
rect 17960 5170 18012 5176
rect 17868 3732 17920 3738
rect 17868 3674 17920 3680
rect 17500 3528 17552 3534
rect 17500 3470 17552 3476
rect 17776 3528 17828 3534
rect 17972 3505 18000 5170
rect 18064 4010 18092 6015
rect 18156 4826 18184 6831
rect 18248 5914 18276 7822
rect 18340 7546 18368 8230
rect 18432 8090 18460 8463
rect 18420 8084 18472 8090
rect 18420 8026 18472 8032
rect 18524 7954 18552 11018
rect 18512 7948 18564 7954
rect 18512 7890 18564 7896
rect 18510 7848 18566 7857
rect 18510 7783 18566 7792
rect 18328 7540 18380 7546
rect 18328 7482 18380 7488
rect 18418 7168 18474 7177
rect 18418 7103 18474 7112
rect 18236 5908 18288 5914
rect 18236 5850 18288 5856
rect 18432 4826 18460 7103
rect 18524 6798 18552 7783
rect 18512 6792 18564 6798
rect 18512 6734 18564 6740
rect 18616 6730 18644 11086
rect 18696 10464 18748 10470
rect 18696 10406 18748 10412
rect 18604 6724 18656 6730
rect 18604 6666 18656 6672
rect 18602 6624 18658 6633
rect 18602 6559 18658 6568
rect 18510 5808 18566 5817
rect 18510 5743 18566 5752
rect 18144 4820 18196 4826
rect 18144 4762 18196 4768
rect 18420 4820 18472 4826
rect 18420 4762 18472 4768
rect 18236 4616 18288 4622
rect 18234 4584 18236 4593
rect 18288 4584 18290 4593
rect 18234 4519 18290 4528
rect 18418 4448 18474 4457
rect 18418 4383 18474 4392
rect 18234 4312 18290 4321
rect 18234 4247 18290 4256
rect 18248 4146 18276 4247
rect 18236 4140 18288 4146
rect 18236 4082 18288 4088
rect 18052 4004 18104 4010
rect 18052 3946 18104 3952
rect 18050 3904 18106 3913
rect 18050 3839 18106 3848
rect 17776 3470 17828 3476
rect 17958 3496 18014 3505
rect 17314 2479 17370 2488
rect 17408 2508 17460 2514
rect 17052 2446 17080 2479
rect 17408 2450 17460 2456
rect 16396 2440 16448 2446
rect 16316 2400 16396 2428
rect 16396 2382 16448 2388
rect 17040 2440 17092 2446
rect 17040 2382 17092 2388
rect 16856 2304 16908 2310
rect 17040 2304 17092 2310
rect 16856 2246 16908 2252
rect 16960 2264 17040 2292
rect 16868 1970 16896 2246
rect 16120 1964 16172 1970
rect 16120 1906 16172 1912
rect 16856 1964 16908 1970
rect 16856 1906 16908 1912
rect 16028 1896 16080 1902
rect 16028 1838 16080 1844
rect 16132 800 16160 1906
rect 16960 800 16988 2264
rect 17040 2246 17092 2252
rect 17512 1970 17540 3470
rect 17958 3431 18014 3440
rect 18064 3194 18092 3839
rect 18236 3528 18288 3534
rect 18236 3470 18288 3476
rect 18248 3233 18276 3470
rect 18234 3224 18290 3233
rect 18052 3188 18104 3194
rect 18432 3194 18460 4383
rect 18524 3738 18552 5743
rect 18616 4010 18644 6559
rect 18708 5370 18736 10406
rect 18800 8838 18828 12406
rect 18972 11008 19024 11014
rect 18972 10950 19024 10956
rect 18788 8832 18840 8838
rect 18788 8774 18840 8780
rect 18696 5364 18748 5370
rect 18696 5306 18748 5312
rect 18800 4690 18828 8774
rect 18984 7750 19012 10950
rect 18972 7744 19024 7750
rect 18972 7686 19024 7692
rect 18984 5302 19012 7686
rect 18972 5296 19024 5302
rect 18972 5238 19024 5244
rect 18788 4684 18840 4690
rect 18788 4626 18840 4632
rect 18604 4004 18656 4010
rect 18604 3946 18656 3952
rect 18512 3732 18564 3738
rect 18512 3674 18564 3680
rect 18234 3159 18290 3168
rect 18420 3188 18472 3194
rect 18052 3130 18104 3136
rect 18420 3130 18472 3136
rect 18418 3088 18474 3097
rect 17592 3052 17644 3058
rect 17592 2994 17644 3000
rect 17960 3052 18012 3058
rect 18418 3023 18474 3032
rect 17960 2994 18012 3000
rect 17604 2582 17632 2994
rect 17684 2848 17736 2854
rect 17682 2816 17684 2825
rect 17736 2816 17738 2825
rect 17682 2751 17738 2760
rect 17592 2576 17644 2582
rect 17592 2518 17644 2524
rect 17972 2417 18000 2994
rect 18432 2650 18460 3023
rect 18420 2644 18472 2650
rect 18420 2586 18472 2592
rect 18236 2440 18288 2446
rect 17958 2408 18014 2417
rect 18236 2382 18288 2388
rect 17958 2343 18014 2352
rect 17776 2304 17828 2310
rect 17776 2246 17828 2252
rect 17500 1964 17552 1970
rect 17500 1906 17552 1912
rect 17788 800 17816 2246
rect 18248 2106 18276 2382
rect 18604 2372 18656 2378
rect 18604 2314 18656 2320
rect 18236 2100 18288 2106
rect 18236 2042 18288 2048
rect 18616 800 18644 2314
rect 1214 0 1270 800
rect 2042 0 2098 800
rect 2870 0 2926 800
rect 3698 0 3754 800
rect 4526 0 4582 800
rect 5354 0 5410 800
rect 6182 0 6238 800
rect 7010 0 7066 800
rect 7838 0 7894 800
rect 8666 0 8722 800
rect 9494 0 9550 800
rect 10322 0 10378 800
rect 11150 0 11206 800
rect 11978 0 12034 800
rect 12806 0 12862 800
rect 13634 0 13690 800
rect 14462 0 14518 800
rect 15290 0 15346 800
rect 16118 0 16174 800
rect 16946 0 17002 800
rect 17774 0 17830 800
rect 18602 0 18658 800
<< via2 >>
rect 1858 14864 1914 14920
rect 2134 15408 2190 15464
rect 1950 14184 2006 14240
rect 1950 13932 2006 13968
rect 3054 15136 3110 15192
rect 2778 14864 2834 14920
rect 2226 14048 2282 14104
rect 2962 14592 3018 14648
rect 1950 13912 1952 13932
rect 1952 13912 2004 13932
rect 2004 13912 2006 13932
rect 2778 13912 2834 13968
rect 3974 15000 4030 15056
rect 3180 14714 3236 14716
rect 3260 14714 3316 14716
rect 3340 14714 3396 14716
rect 3420 14714 3476 14716
rect 3180 14662 3226 14714
rect 3226 14662 3236 14714
rect 3260 14662 3290 14714
rect 3290 14662 3302 14714
rect 3302 14662 3316 14714
rect 3340 14662 3354 14714
rect 3354 14662 3366 14714
rect 3366 14662 3396 14714
rect 3420 14662 3430 14714
rect 3430 14662 3476 14714
rect 3180 14660 3236 14662
rect 3260 14660 3316 14662
rect 3340 14660 3396 14662
rect 3420 14660 3476 14662
rect 3514 14456 3570 14512
rect 3514 14048 3570 14104
rect 3054 13912 3110 13968
rect 3422 13776 3478 13832
rect 3180 13626 3236 13628
rect 3260 13626 3316 13628
rect 3340 13626 3396 13628
rect 3420 13626 3476 13628
rect 3180 13574 3226 13626
rect 3226 13574 3236 13626
rect 3260 13574 3290 13626
rect 3290 13574 3302 13626
rect 3302 13574 3316 13626
rect 3340 13574 3354 13626
rect 3354 13574 3366 13626
rect 3366 13574 3396 13626
rect 3420 13574 3430 13626
rect 3430 13574 3476 13626
rect 3180 13572 3236 13574
rect 3260 13572 3316 13574
rect 3340 13572 3396 13574
rect 3420 13572 3476 13574
rect 2870 13504 2926 13560
rect 1950 13388 2006 13424
rect 1950 13368 1952 13388
rect 1952 13368 2004 13388
rect 2004 13368 2006 13388
rect 2686 13132 2688 13152
rect 2688 13132 2740 13152
rect 2740 13132 2742 13152
rect 2686 13096 2742 13132
rect 1674 12280 1730 12336
rect 1398 10004 1400 10024
rect 1400 10004 1452 10024
rect 1452 10004 1454 10024
rect 1398 9968 1454 10004
rect 1490 7792 1546 7848
rect 2042 11192 2098 11248
rect 1950 10920 2006 10976
rect 1950 10104 2006 10160
rect 1950 9560 2006 9616
rect 1950 9288 2006 9344
rect 1950 8472 2006 8528
rect 2226 11636 2228 11656
rect 2228 11636 2280 11656
rect 2280 11636 2282 11656
rect 2226 11600 2282 11636
rect 2226 11092 2228 11112
rect 2228 11092 2280 11112
rect 2280 11092 2282 11112
rect 2226 11056 2282 11092
rect 2134 9832 2190 9888
rect 2226 9696 2282 9752
rect 2226 8336 2282 8392
rect 2410 10512 2466 10568
rect 2502 8744 2558 8800
rect 2778 12416 2834 12472
rect 2778 12008 2834 12064
rect 2778 11736 2834 11792
rect 3238 12824 3294 12880
rect 3180 12538 3236 12540
rect 3260 12538 3316 12540
rect 3340 12538 3396 12540
rect 3420 12538 3476 12540
rect 3180 12486 3226 12538
rect 3226 12486 3236 12538
rect 3260 12486 3290 12538
rect 3290 12486 3302 12538
rect 3302 12486 3316 12538
rect 3340 12486 3354 12538
rect 3354 12486 3366 12538
rect 3366 12486 3396 12538
rect 3420 12486 3430 12538
rect 3430 12486 3476 12538
rect 3180 12484 3236 12486
rect 3260 12484 3316 12486
rect 3340 12484 3396 12486
rect 3420 12484 3476 12486
rect 3146 12180 3148 12200
rect 3148 12180 3200 12200
rect 3200 12180 3202 12200
rect 3146 12144 3202 12180
rect 3054 11872 3110 11928
rect 3180 11450 3236 11452
rect 3260 11450 3316 11452
rect 3340 11450 3396 11452
rect 3420 11450 3476 11452
rect 3180 11398 3226 11450
rect 3226 11398 3236 11450
rect 3260 11398 3290 11450
rect 3290 11398 3302 11450
rect 3302 11398 3316 11450
rect 3340 11398 3354 11450
rect 3354 11398 3366 11450
rect 3366 11398 3396 11450
rect 3420 11398 3430 11450
rect 3430 11398 3476 11450
rect 3180 11396 3236 11398
rect 3260 11396 3316 11398
rect 3340 11396 3396 11398
rect 3420 11396 3476 11398
rect 2778 11228 2780 11248
rect 2780 11228 2832 11248
rect 2832 11228 2834 11248
rect 2778 11192 2834 11228
rect 2870 10784 2926 10840
rect 2594 8472 2650 8528
rect 2778 10240 2834 10296
rect 2778 9424 2834 9480
rect 2962 9152 3018 9208
rect 2870 9016 2926 9072
rect 2778 8880 2834 8936
rect 1674 7656 1730 7712
rect 1490 6704 1546 6760
rect 1490 6160 1546 6216
rect 1398 5888 1454 5944
rect 1490 5072 1546 5128
rect 1306 4120 1362 4176
rect 1490 3984 1546 4040
rect 1950 6160 2006 6216
rect 2318 6704 2374 6760
rect 2410 6452 2466 6488
rect 2410 6432 2412 6452
rect 2412 6432 2464 6452
rect 2464 6432 2466 6452
rect 2686 7520 2742 7576
rect 2962 8880 3018 8936
rect 2962 8064 3018 8120
rect 2962 7540 3018 7576
rect 2962 7520 2964 7540
rect 2964 7520 3016 7540
rect 3016 7520 3018 7540
rect 3146 10512 3202 10568
rect 4066 14320 4122 14376
rect 3974 13232 4030 13288
rect 3882 12960 3938 13016
rect 5078 14864 5134 14920
rect 5078 14320 5134 14376
rect 4342 13912 4398 13968
rect 5170 14184 5226 14240
rect 4618 13776 4674 13832
rect 4158 12144 4214 12200
rect 4250 12008 4306 12064
rect 4158 11772 4160 11792
rect 4160 11772 4212 11792
rect 4212 11772 4214 11792
rect 4158 11736 4214 11772
rect 3974 11464 4030 11520
rect 3606 10784 3662 10840
rect 3180 10362 3236 10364
rect 3260 10362 3316 10364
rect 3340 10362 3396 10364
rect 3420 10362 3476 10364
rect 3180 10310 3226 10362
rect 3226 10310 3236 10362
rect 3260 10310 3290 10362
rect 3290 10310 3302 10362
rect 3302 10310 3316 10362
rect 3340 10310 3354 10362
rect 3354 10310 3366 10362
rect 3366 10310 3396 10362
rect 3420 10310 3430 10362
rect 3430 10310 3476 10362
rect 3180 10308 3236 10310
rect 3260 10308 3316 10310
rect 3340 10308 3396 10310
rect 3420 10308 3476 10310
rect 3330 9968 3386 10024
rect 3974 11192 4030 11248
rect 3882 10684 3884 10704
rect 3884 10684 3936 10704
rect 3936 10684 3938 10704
rect 3882 10648 3938 10684
rect 3180 9274 3236 9276
rect 3260 9274 3316 9276
rect 3340 9274 3396 9276
rect 3420 9274 3476 9276
rect 3180 9222 3226 9274
rect 3226 9222 3236 9274
rect 3260 9222 3290 9274
rect 3290 9222 3302 9274
rect 3302 9222 3316 9274
rect 3340 9222 3354 9274
rect 3354 9222 3366 9274
rect 3366 9222 3396 9274
rect 3420 9222 3430 9274
rect 3430 9222 3476 9274
rect 3180 9220 3236 9222
rect 3260 9220 3316 9222
rect 3340 9220 3396 9222
rect 3420 9220 3476 9222
rect 3238 8608 3294 8664
rect 3180 8186 3236 8188
rect 3260 8186 3316 8188
rect 3340 8186 3396 8188
rect 3420 8186 3476 8188
rect 3180 8134 3226 8186
rect 3226 8134 3236 8186
rect 3260 8134 3290 8186
rect 3290 8134 3302 8186
rect 3302 8134 3316 8186
rect 3340 8134 3354 8186
rect 3354 8134 3366 8186
rect 3366 8134 3396 8186
rect 3420 8134 3430 8186
rect 3430 8134 3476 8186
rect 3180 8132 3236 8134
rect 3260 8132 3316 8134
rect 3340 8132 3396 8134
rect 3420 8132 3476 8134
rect 3698 8472 3754 8528
rect 2870 7112 2926 7168
rect 3054 7248 3110 7304
rect 2962 6976 3018 7032
rect 1858 5616 1914 5672
rect 2134 5616 2190 5672
rect 2318 5480 2374 5536
rect 2226 4820 2282 4856
rect 2226 4800 2228 4820
rect 2228 4800 2280 4820
rect 2280 4800 2282 4820
rect 1858 4528 1914 4584
rect 3180 7098 3236 7100
rect 3260 7098 3316 7100
rect 3340 7098 3396 7100
rect 3420 7098 3476 7100
rect 3180 7046 3226 7098
rect 3226 7046 3236 7098
rect 3260 7046 3290 7098
rect 3290 7046 3302 7098
rect 3302 7046 3316 7098
rect 3340 7046 3354 7098
rect 3354 7046 3366 7098
rect 3366 7046 3396 7098
rect 3420 7046 3430 7098
rect 3430 7046 3476 7098
rect 3180 7044 3236 7046
rect 3260 7044 3316 7046
rect 3340 7044 3396 7046
rect 3420 7044 3476 7046
rect 3330 6432 3386 6488
rect 2870 6160 2926 6216
rect 3422 6296 3478 6352
rect 3180 6010 3236 6012
rect 3260 6010 3316 6012
rect 3340 6010 3396 6012
rect 3420 6010 3476 6012
rect 3180 5958 3226 6010
rect 3226 5958 3236 6010
rect 3260 5958 3290 6010
rect 3290 5958 3302 6010
rect 3302 5958 3316 6010
rect 3340 5958 3354 6010
rect 3354 5958 3366 6010
rect 3366 5958 3396 6010
rect 3420 5958 3430 6010
rect 3430 5958 3476 6010
rect 3180 5956 3236 5958
rect 3260 5956 3316 5958
rect 3340 5956 3396 5958
rect 3420 5956 3476 5958
rect 2778 5364 2834 5400
rect 2778 5344 2780 5364
rect 2780 5344 2832 5364
rect 2832 5344 2834 5364
rect 2502 4528 2558 4584
rect 2226 3712 2282 3768
rect 2778 4256 2834 4312
rect 2686 3984 2742 4040
rect 1950 3440 2006 3496
rect 1490 3188 1546 3224
rect 1490 3168 1492 3188
rect 1492 3168 1544 3188
rect 1544 3168 1546 3188
rect 2318 3168 2374 3224
rect 1858 2916 1914 2952
rect 1858 2896 1860 2916
rect 1860 2896 1912 2916
rect 1912 2896 1914 2916
rect 3238 5616 3294 5672
rect 3422 5480 3478 5536
rect 3514 5228 3570 5264
rect 3514 5208 3516 5228
rect 3516 5208 3568 5228
rect 3568 5208 3570 5228
rect 3422 5092 3478 5128
rect 3422 5072 3424 5092
rect 3424 5072 3476 5092
rect 3476 5072 3478 5092
rect 3180 4922 3236 4924
rect 3260 4922 3316 4924
rect 3340 4922 3396 4924
rect 3420 4922 3476 4924
rect 3180 4870 3226 4922
rect 3226 4870 3236 4922
rect 3260 4870 3290 4922
rect 3290 4870 3302 4922
rect 3302 4870 3316 4922
rect 3340 4870 3354 4922
rect 3354 4870 3366 4922
rect 3366 4870 3396 4922
rect 3420 4870 3430 4922
rect 3430 4870 3476 4922
rect 3180 4868 3236 4870
rect 3260 4868 3316 4870
rect 3340 4868 3396 4870
rect 3420 4868 3476 4870
rect 3330 4664 3386 4720
rect 2778 3476 2780 3496
rect 2780 3476 2832 3496
rect 2832 3476 2834 3496
rect 2778 3440 2834 3476
rect 1490 2644 1546 2680
rect 1490 2624 1492 2644
rect 1492 2624 1544 2644
rect 1544 2624 1546 2644
rect 1858 2352 1914 2408
rect 4158 10784 4214 10840
rect 3974 8880 4030 8936
rect 3790 7248 3846 7304
rect 3422 3984 3478 4040
rect 3180 3834 3236 3836
rect 3260 3834 3316 3836
rect 3340 3834 3396 3836
rect 3420 3834 3476 3836
rect 3180 3782 3226 3834
rect 3226 3782 3236 3834
rect 3260 3782 3290 3834
rect 3290 3782 3302 3834
rect 3302 3782 3316 3834
rect 3340 3782 3354 3834
rect 3354 3782 3366 3834
rect 3366 3782 3396 3834
rect 3420 3782 3430 3834
rect 3430 3782 3476 3834
rect 3180 3780 3236 3782
rect 3260 3780 3316 3782
rect 3340 3780 3396 3782
rect 3420 3780 3476 3782
rect 3180 2746 3236 2748
rect 3260 2746 3316 2748
rect 3340 2746 3396 2748
rect 3420 2746 3476 2748
rect 3180 2694 3226 2746
rect 3226 2694 3236 2746
rect 3260 2694 3290 2746
rect 3290 2694 3302 2746
rect 3302 2694 3316 2746
rect 3340 2694 3354 2746
rect 3354 2694 3366 2746
rect 3366 2694 3396 2746
rect 3420 2694 3430 2746
rect 3430 2694 3476 2746
rect 3180 2692 3236 2694
rect 3260 2692 3316 2694
rect 3340 2692 3396 2694
rect 3420 2692 3476 2694
rect 3974 6976 4030 7032
rect 3974 6840 4030 6896
rect 5078 13368 5134 13424
rect 5404 14170 5460 14172
rect 5484 14170 5540 14172
rect 5564 14170 5620 14172
rect 5644 14170 5700 14172
rect 5404 14118 5450 14170
rect 5450 14118 5460 14170
rect 5484 14118 5514 14170
rect 5514 14118 5526 14170
rect 5526 14118 5540 14170
rect 5564 14118 5578 14170
rect 5578 14118 5590 14170
rect 5590 14118 5620 14170
rect 5644 14118 5654 14170
rect 5654 14118 5700 14170
rect 5404 14116 5460 14118
rect 5484 14116 5540 14118
rect 5564 14116 5620 14118
rect 5644 14116 5700 14118
rect 5262 13776 5318 13832
rect 5262 13132 5264 13152
rect 5264 13132 5316 13152
rect 5316 13132 5318 13152
rect 5262 13096 5318 13132
rect 5404 13082 5460 13084
rect 5484 13082 5540 13084
rect 5564 13082 5620 13084
rect 5644 13082 5700 13084
rect 5404 13030 5450 13082
rect 5450 13030 5460 13082
rect 5484 13030 5514 13082
rect 5514 13030 5526 13082
rect 5526 13030 5540 13082
rect 5564 13030 5578 13082
rect 5578 13030 5590 13082
rect 5590 13030 5620 13082
rect 5644 13030 5654 13082
rect 5654 13030 5700 13082
rect 5404 13028 5460 13030
rect 5484 13028 5540 13030
rect 5564 13028 5620 13030
rect 5644 13028 5700 13030
rect 5170 12724 5172 12744
rect 5172 12724 5224 12744
rect 5224 12724 5226 12744
rect 5170 12688 5226 12724
rect 5538 12552 5594 12608
rect 5998 12144 6054 12200
rect 5404 11994 5460 11996
rect 5484 11994 5540 11996
rect 5564 11994 5620 11996
rect 5644 11994 5700 11996
rect 5404 11942 5450 11994
rect 5450 11942 5460 11994
rect 5484 11942 5514 11994
rect 5514 11942 5526 11994
rect 5526 11942 5540 11994
rect 5564 11942 5578 11994
rect 5578 11942 5590 11994
rect 5590 11942 5620 11994
rect 5644 11942 5654 11994
rect 5654 11942 5700 11994
rect 5404 11940 5460 11942
rect 5484 11940 5540 11942
rect 5564 11940 5620 11942
rect 5644 11940 5700 11942
rect 5630 11736 5686 11792
rect 4710 11464 4766 11520
rect 4894 11056 4950 11112
rect 4342 8472 4398 8528
rect 3974 6296 4030 6352
rect 4066 5344 4122 5400
rect 3790 4664 3846 4720
rect 3790 4276 3846 4312
rect 3790 4256 3792 4276
rect 3792 4256 3844 4276
rect 3844 4256 3846 4276
rect 3974 5208 4030 5264
rect 3882 3188 3938 3224
rect 3882 3168 3884 3188
rect 3884 3168 3936 3188
rect 3936 3168 3938 3188
rect 4802 9832 4858 9888
rect 4986 10956 4988 10976
rect 4988 10956 5040 10976
rect 5040 10956 5042 10976
rect 4986 10920 5042 10956
rect 4986 10412 4988 10432
rect 4988 10412 5040 10432
rect 5040 10412 5042 10432
rect 4986 10376 5042 10412
rect 5814 11756 5870 11792
rect 5814 11736 5816 11756
rect 5816 11736 5868 11756
rect 5868 11736 5870 11756
rect 5722 11192 5778 11248
rect 5906 11620 5962 11656
rect 5906 11600 5908 11620
rect 5908 11600 5960 11620
rect 5960 11600 5962 11620
rect 5814 11056 5870 11112
rect 5404 10906 5460 10908
rect 5484 10906 5540 10908
rect 5564 10906 5620 10908
rect 5644 10906 5700 10908
rect 5404 10854 5450 10906
rect 5450 10854 5460 10906
rect 5484 10854 5514 10906
rect 5514 10854 5526 10906
rect 5526 10854 5540 10906
rect 5564 10854 5578 10906
rect 5578 10854 5590 10906
rect 5590 10854 5620 10906
rect 5644 10854 5654 10906
rect 5654 10854 5700 10906
rect 5404 10852 5460 10854
rect 5484 10852 5540 10854
rect 5564 10852 5620 10854
rect 5644 10852 5700 10854
rect 5262 10784 5318 10840
rect 5722 10668 5778 10704
rect 5722 10648 5724 10668
rect 5724 10648 5776 10668
rect 5776 10648 5778 10668
rect 5262 10104 5318 10160
rect 7628 14714 7684 14716
rect 7708 14714 7764 14716
rect 7788 14714 7844 14716
rect 7868 14714 7924 14716
rect 7628 14662 7674 14714
rect 7674 14662 7684 14714
rect 7708 14662 7738 14714
rect 7738 14662 7750 14714
rect 7750 14662 7764 14714
rect 7788 14662 7802 14714
rect 7802 14662 7814 14714
rect 7814 14662 7844 14714
rect 7868 14662 7878 14714
rect 7878 14662 7924 14714
rect 7628 14660 7684 14662
rect 7708 14660 7764 14662
rect 7788 14660 7844 14662
rect 7868 14660 7924 14662
rect 6458 12008 6514 12064
rect 6274 11464 6330 11520
rect 6458 11328 6514 11384
rect 5906 10512 5962 10568
rect 5404 9818 5460 9820
rect 5484 9818 5540 9820
rect 5564 9818 5620 9820
rect 5644 9818 5700 9820
rect 5404 9766 5450 9818
rect 5450 9766 5460 9818
rect 5484 9766 5514 9818
rect 5514 9766 5526 9818
rect 5526 9766 5540 9818
rect 5564 9766 5578 9818
rect 5578 9766 5590 9818
rect 5590 9766 5620 9818
rect 5644 9766 5654 9818
rect 5654 9766 5700 9818
rect 5404 9764 5460 9766
rect 5484 9764 5540 9766
rect 5564 9764 5620 9766
rect 5644 9764 5700 9766
rect 5354 9152 5410 9208
rect 4434 6740 4436 6760
rect 4436 6740 4488 6760
rect 4488 6740 4490 6760
rect 4434 6704 4490 6740
rect 4250 5480 4306 5536
rect 4250 4820 4306 4856
rect 4250 4800 4252 4820
rect 4252 4800 4304 4820
rect 4304 4800 4306 4820
rect 4158 4392 4214 4448
rect 4802 7792 4858 7848
rect 4894 7384 4950 7440
rect 5404 8730 5460 8732
rect 5484 8730 5540 8732
rect 5564 8730 5620 8732
rect 5644 8730 5700 8732
rect 5404 8678 5450 8730
rect 5450 8678 5460 8730
rect 5484 8678 5514 8730
rect 5514 8678 5526 8730
rect 5526 8678 5540 8730
rect 5564 8678 5578 8730
rect 5578 8678 5590 8730
rect 5590 8678 5620 8730
rect 5644 8678 5654 8730
rect 5654 8678 5700 8730
rect 5404 8676 5460 8678
rect 5484 8676 5540 8678
rect 5564 8676 5620 8678
rect 5644 8676 5700 8678
rect 4894 6432 4950 6488
rect 4986 6296 5042 6352
rect 5404 7642 5460 7644
rect 5484 7642 5540 7644
rect 5564 7642 5620 7644
rect 5644 7642 5700 7644
rect 5404 7590 5450 7642
rect 5450 7590 5460 7642
rect 5484 7590 5514 7642
rect 5514 7590 5526 7642
rect 5526 7590 5540 7642
rect 5564 7590 5578 7642
rect 5578 7590 5590 7642
rect 5590 7590 5620 7642
rect 5644 7590 5654 7642
rect 5654 7590 5700 7642
rect 5404 7588 5460 7590
rect 5484 7588 5540 7590
rect 5564 7588 5620 7590
rect 5644 7588 5700 7590
rect 5906 9832 5962 9888
rect 5906 9016 5962 9072
rect 5906 6976 5962 7032
rect 5262 6604 5264 6624
rect 5264 6604 5316 6624
rect 5316 6604 5318 6624
rect 5262 6568 5318 6604
rect 5404 6554 5460 6556
rect 5484 6554 5540 6556
rect 5564 6554 5620 6556
rect 5644 6554 5700 6556
rect 5404 6502 5450 6554
rect 5450 6502 5460 6554
rect 5484 6502 5514 6554
rect 5514 6502 5526 6554
rect 5526 6502 5540 6554
rect 5564 6502 5578 6554
rect 5578 6502 5590 6554
rect 5590 6502 5620 6554
rect 5644 6502 5654 6554
rect 5654 6502 5700 6554
rect 5404 6500 5460 6502
rect 5484 6500 5540 6502
rect 5564 6500 5620 6502
rect 5644 6500 5700 6502
rect 5354 6296 5410 6352
rect 4802 5616 4858 5672
rect 4894 5344 4950 5400
rect 5262 6160 5318 6216
rect 5446 5888 5502 5944
rect 5404 5466 5460 5468
rect 5484 5466 5540 5468
rect 5564 5466 5620 5468
rect 5644 5466 5700 5468
rect 5404 5414 5450 5466
rect 5450 5414 5460 5466
rect 5484 5414 5514 5466
rect 5514 5414 5526 5466
rect 5526 5414 5540 5466
rect 5564 5414 5578 5466
rect 5578 5414 5590 5466
rect 5590 5414 5620 5466
rect 5644 5414 5654 5466
rect 5654 5414 5700 5466
rect 5404 5412 5460 5414
rect 5484 5412 5540 5414
rect 5564 5412 5620 5414
rect 5644 5412 5700 5414
rect 5078 4564 5080 4584
rect 5080 4564 5132 4584
rect 5132 4564 5134 4584
rect 5078 4528 5134 4564
rect 4986 4120 5042 4176
rect 4710 3476 4712 3496
rect 4712 3476 4764 3496
rect 4764 3476 4766 3496
rect 4710 3440 4766 3476
rect 5404 4378 5460 4380
rect 5484 4378 5540 4380
rect 5564 4378 5620 4380
rect 5644 4378 5700 4380
rect 5404 4326 5450 4378
rect 5450 4326 5460 4378
rect 5484 4326 5514 4378
rect 5514 4326 5526 4378
rect 5526 4326 5540 4378
rect 5564 4326 5578 4378
rect 5578 4326 5590 4378
rect 5590 4326 5620 4378
rect 5644 4326 5654 4378
rect 5654 4326 5700 4378
rect 5404 4324 5460 4326
rect 5484 4324 5540 4326
rect 5564 4324 5620 4326
rect 5644 4324 5700 4326
rect 5404 3290 5460 3292
rect 5484 3290 5540 3292
rect 5564 3290 5620 3292
rect 5644 3290 5700 3292
rect 5404 3238 5450 3290
rect 5450 3238 5460 3290
rect 5484 3238 5514 3290
rect 5514 3238 5526 3290
rect 5526 3238 5540 3290
rect 5564 3238 5578 3290
rect 5578 3238 5590 3290
rect 5590 3238 5620 3290
rect 5644 3238 5654 3290
rect 5654 3238 5700 3290
rect 5404 3236 5460 3238
rect 5484 3236 5540 3238
rect 5564 3236 5620 3238
rect 5644 3236 5700 3238
rect 5906 6024 5962 6080
rect 5906 5228 5962 5264
rect 5906 5208 5908 5228
rect 5908 5208 5960 5228
rect 5960 5208 5962 5228
rect 5814 5072 5870 5128
rect 6182 10512 6238 10568
rect 6182 5516 6184 5536
rect 6184 5516 6236 5536
rect 6236 5516 6238 5536
rect 6182 5480 6238 5516
rect 6550 9424 6606 9480
rect 6458 9016 6514 9072
rect 6734 10240 6790 10296
rect 6918 9696 6974 9752
rect 6734 9016 6790 9072
rect 6642 8780 6644 8800
rect 6644 8780 6696 8800
rect 6696 8780 6698 8800
rect 6642 8744 6698 8780
rect 6458 7384 6514 7440
rect 6458 6840 6514 6896
rect 6458 5208 6514 5264
rect 6826 8608 6882 8664
rect 7194 10784 7250 10840
rect 6734 6840 6790 6896
rect 6642 6296 6698 6352
rect 6826 5480 6882 5536
rect 7628 13626 7684 13628
rect 7708 13626 7764 13628
rect 7788 13626 7844 13628
rect 7868 13626 7924 13628
rect 7628 13574 7674 13626
rect 7674 13574 7684 13626
rect 7708 13574 7738 13626
rect 7738 13574 7750 13626
rect 7750 13574 7764 13626
rect 7788 13574 7802 13626
rect 7802 13574 7814 13626
rect 7814 13574 7844 13626
rect 7868 13574 7878 13626
rect 7878 13574 7924 13626
rect 7628 13572 7684 13574
rect 7708 13572 7764 13574
rect 7788 13572 7844 13574
rect 7868 13572 7924 13574
rect 8758 14320 8814 14376
rect 7628 12538 7684 12540
rect 7708 12538 7764 12540
rect 7788 12538 7844 12540
rect 7868 12538 7924 12540
rect 7628 12486 7674 12538
rect 7674 12486 7684 12538
rect 7708 12486 7738 12538
rect 7738 12486 7750 12538
rect 7750 12486 7764 12538
rect 7788 12486 7802 12538
rect 7802 12486 7814 12538
rect 7814 12486 7844 12538
rect 7868 12486 7878 12538
rect 7878 12486 7924 12538
rect 7628 12484 7684 12486
rect 7708 12484 7764 12486
rect 7788 12484 7844 12486
rect 7868 12484 7924 12486
rect 8482 13368 8538 13424
rect 8482 12552 8538 12608
rect 8574 12280 8630 12336
rect 7628 11450 7684 11452
rect 7708 11450 7764 11452
rect 7788 11450 7844 11452
rect 7868 11450 7924 11452
rect 7628 11398 7674 11450
rect 7674 11398 7684 11450
rect 7708 11398 7738 11450
rect 7738 11398 7750 11450
rect 7750 11398 7764 11450
rect 7788 11398 7802 11450
rect 7802 11398 7814 11450
rect 7814 11398 7844 11450
rect 7868 11398 7878 11450
rect 7878 11398 7924 11450
rect 7628 11396 7684 11398
rect 7708 11396 7764 11398
rect 7788 11396 7844 11398
rect 7868 11396 7924 11398
rect 7628 10362 7684 10364
rect 7708 10362 7764 10364
rect 7788 10362 7844 10364
rect 7868 10362 7924 10364
rect 7628 10310 7674 10362
rect 7674 10310 7684 10362
rect 7708 10310 7738 10362
rect 7738 10310 7750 10362
rect 7750 10310 7764 10362
rect 7788 10310 7802 10362
rect 7802 10310 7814 10362
rect 7814 10310 7844 10362
rect 7868 10310 7878 10362
rect 7878 10310 7924 10362
rect 7628 10308 7684 10310
rect 7708 10308 7764 10310
rect 7788 10308 7844 10310
rect 7868 10308 7924 10310
rect 7194 8064 7250 8120
rect 7102 5344 7158 5400
rect 7102 4800 7158 4856
rect 6918 4256 6974 4312
rect 7628 9274 7684 9276
rect 7708 9274 7764 9276
rect 7788 9274 7844 9276
rect 7868 9274 7924 9276
rect 7628 9222 7674 9274
rect 7674 9222 7684 9274
rect 7708 9222 7738 9274
rect 7738 9222 7750 9274
rect 7750 9222 7764 9274
rect 7788 9222 7802 9274
rect 7802 9222 7814 9274
rect 7814 9222 7844 9274
rect 7868 9222 7878 9274
rect 7878 9222 7924 9274
rect 7628 9220 7684 9222
rect 7708 9220 7764 9222
rect 7788 9220 7844 9222
rect 7868 9220 7924 9222
rect 8022 8628 8078 8664
rect 8022 8608 8024 8628
rect 8024 8608 8076 8628
rect 8076 8608 8078 8628
rect 8114 8372 8116 8392
rect 8116 8372 8168 8392
rect 8168 8372 8170 8392
rect 7628 8186 7684 8188
rect 7708 8186 7764 8188
rect 7788 8186 7844 8188
rect 7868 8186 7924 8188
rect 7628 8134 7674 8186
rect 7674 8134 7684 8186
rect 7708 8134 7738 8186
rect 7738 8134 7750 8186
rect 7750 8134 7764 8186
rect 7788 8134 7802 8186
rect 7802 8134 7814 8186
rect 7814 8134 7844 8186
rect 7868 8134 7878 8186
rect 7878 8134 7924 8186
rect 7628 8132 7684 8134
rect 7708 8132 7764 8134
rect 7788 8132 7844 8134
rect 7868 8132 7924 8134
rect 8114 8336 8170 8372
rect 8114 8200 8170 8256
rect 7628 7098 7684 7100
rect 7708 7098 7764 7100
rect 7788 7098 7844 7100
rect 7868 7098 7924 7100
rect 7628 7046 7674 7098
rect 7674 7046 7684 7098
rect 7708 7046 7738 7098
rect 7738 7046 7750 7098
rect 7750 7046 7764 7098
rect 7788 7046 7802 7098
rect 7802 7046 7814 7098
rect 7814 7046 7844 7098
rect 7868 7046 7878 7098
rect 7878 7046 7924 7098
rect 7628 7044 7684 7046
rect 7708 7044 7764 7046
rect 7788 7044 7844 7046
rect 7868 7044 7924 7046
rect 7746 6860 7802 6896
rect 7746 6840 7748 6860
rect 7748 6840 7800 6860
rect 7800 6840 7802 6860
rect 7470 6432 7526 6488
rect 8022 6296 8078 6352
rect 7628 6010 7684 6012
rect 7708 6010 7764 6012
rect 7788 6010 7844 6012
rect 7868 6010 7924 6012
rect 7628 5958 7674 6010
rect 7674 5958 7684 6010
rect 7708 5958 7738 6010
rect 7738 5958 7750 6010
rect 7750 5958 7764 6010
rect 7788 5958 7802 6010
rect 7802 5958 7814 6010
rect 7814 5958 7844 6010
rect 7868 5958 7878 6010
rect 7878 5958 7924 6010
rect 7628 5956 7684 5958
rect 7708 5956 7764 5958
rect 7788 5956 7844 5958
rect 7868 5956 7924 5958
rect 7286 5616 7342 5672
rect 8758 13232 8814 13288
rect 9852 14170 9908 14172
rect 9932 14170 9988 14172
rect 10012 14170 10068 14172
rect 10092 14170 10148 14172
rect 9852 14118 9898 14170
rect 9898 14118 9908 14170
rect 9932 14118 9962 14170
rect 9962 14118 9974 14170
rect 9974 14118 9988 14170
rect 10012 14118 10026 14170
rect 10026 14118 10038 14170
rect 10038 14118 10068 14170
rect 10092 14118 10102 14170
rect 10102 14118 10148 14170
rect 9852 14116 9908 14118
rect 9932 14116 9988 14118
rect 10012 14116 10068 14118
rect 10092 14116 10148 14118
rect 8942 12280 8998 12336
rect 8942 12008 8998 12064
rect 8850 11192 8906 11248
rect 8942 11056 8998 11112
rect 8850 10512 8906 10568
rect 8758 8472 8814 8528
rect 8666 8200 8722 8256
rect 8942 8880 8998 8936
rect 9402 12688 9458 12744
rect 9218 9832 9274 9888
rect 9126 8880 9182 8936
rect 8574 6976 8630 7032
rect 8298 5636 8354 5672
rect 8298 5616 8300 5636
rect 8300 5616 8352 5636
rect 8352 5616 8354 5636
rect 7628 4922 7684 4924
rect 7708 4922 7764 4924
rect 7788 4922 7844 4924
rect 7868 4922 7924 4924
rect 7628 4870 7674 4922
rect 7674 4870 7684 4922
rect 7708 4870 7738 4922
rect 7738 4870 7750 4922
rect 7750 4870 7764 4922
rect 7788 4870 7802 4922
rect 7802 4870 7814 4922
rect 7814 4870 7844 4922
rect 7868 4870 7878 4922
rect 7878 4870 7924 4922
rect 7628 4868 7684 4870
rect 7708 4868 7764 4870
rect 7788 4868 7844 4870
rect 7868 4868 7924 4870
rect 7470 4800 7526 4856
rect 8850 7404 8906 7440
rect 8850 7384 8852 7404
rect 8852 7384 8904 7404
rect 8904 7384 8906 7404
rect 8482 5480 8538 5536
rect 7470 4392 7526 4448
rect 7470 4120 7526 4176
rect 9310 9288 9366 9344
rect 9678 12860 9680 12880
rect 9680 12860 9732 12880
rect 9732 12860 9734 12880
rect 9678 12824 9734 12860
rect 9586 10804 9642 10840
rect 9586 10784 9588 10804
rect 9588 10784 9640 10804
rect 9640 10784 9642 10804
rect 9852 13082 9908 13084
rect 9932 13082 9988 13084
rect 10012 13082 10068 13084
rect 10092 13082 10148 13084
rect 9852 13030 9898 13082
rect 9898 13030 9908 13082
rect 9932 13030 9962 13082
rect 9962 13030 9974 13082
rect 9974 13030 9988 13082
rect 10012 13030 10026 13082
rect 10026 13030 10038 13082
rect 10038 13030 10068 13082
rect 10092 13030 10102 13082
rect 10102 13030 10148 13082
rect 9852 13028 9908 13030
rect 9932 13028 9988 13030
rect 10012 13028 10068 13030
rect 10092 13028 10148 13030
rect 10230 12824 10286 12880
rect 9852 11994 9908 11996
rect 9932 11994 9988 11996
rect 10012 11994 10068 11996
rect 10092 11994 10148 11996
rect 9852 11942 9898 11994
rect 9898 11942 9908 11994
rect 9932 11942 9962 11994
rect 9962 11942 9974 11994
rect 9974 11942 9988 11994
rect 10012 11942 10026 11994
rect 10026 11942 10038 11994
rect 10038 11942 10068 11994
rect 10092 11942 10102 11994
rect 10102 11942 10148 11994
rect 9852 11940 9908 11942
rect 9932 11940 9988 11942
rect 10012 11940 10068 11942
rect 10092 11940 10148 11942
rect 9852 10906 9908 10908
rect 9932 10906 9988 10908
rect 10012 10906 10068 10908
rect 10092 10906 10148 10908
rect 9852 10854 9898 10906
rect 9898 10854 9908 10906
rect 9932 10854 9962 10906
rect 9962 10854 9974 10906
rect 9974 10854 9988 10906
rect 10012 10854 10026 10906
rect 10026 10854 10038 10906
rect 10038 10854 10068 10906
rect 10092 10854 10102 10906
rect 10102 10854 10148 10906
rect 9852 10852 9908 10854
rect 9932 10852 9988 10854
rect 10012 10852 10068 10854
rect 10092 10852 10148 10854
rect 10230 10784 10286 10840
rect 10046 10376 10102 10432
rect 10230 9832 10286 9888
rect 9852 9818 9908 9820
rect 9932 9818 9988 9820
rect 10012 9818 10068 9820
rect 10092 9818 10148 9820
rect 9852 9766 9898 9818
rect 9898 9766 9908 9818
rect 9932 9766 9962 9818
rect 9962 9766 9974 9818
rect 9974 9766 9988 9818
rect 10012 9766 10026 9818
rect 10026 9766 10038 9818
rect 10038 9766 10068 9818
rect 10092 9766 10102 9818
rect 10102 9766 10148 9818
rect 9852 9764 9908 9766
rect 9932 9764 9988 9766
rect 10012 9764 10068 9766
rect 10092 9764 10148 9766
rect 9678 9560 9734 9616
rect 9310 7520 9366 7576
rect 9218 6840 9274 6896
rect 8942 5652 8944 5672
rect 8944 5652 8996 5672
rect 8996 5652 8998 5672
rect 8942 5616 8998 5652
rect 9954 9324 9956 9344
rect 9956 9324 10008 9344
rect 10008 9324 10010 9344
rect 9954 9288 10010 9324
rect 10046 9152 10102 9208
rect 10322 9696 10378 9752
rect 9852 8730 9908 8732
rect 9932 8730 9988 8732
rect 10012 8730 10068 8732
rect 10092 8730 10148 8732
rect 9852 8678 9898 8730
rect 9898 8678 9908 8730
rect 9932 8678 9962 8730
rect 9962 8678 9974 8730
rect 9974 8678 9988 8730
rect 10012 8678 10026 8730
rect 10026 8678 10038 8730
rect 10038 8678 10068 8730
rect 10092 8678 10102 8730
rect 10102 8678 10148 8730
rect 9852 8676 9908 8678
rect 9932 8676 9988 8678
rect 10012 8676 10068 8678
rect 10092 8676 10148 8678
rect 9862 8356 9918 8392
rect 9862 8336 9864 8356
rect 9864 8336 9916 8356
rect 9916 8336 9918 8356
rect 10046 7792 10102 7848
rect 9852 7642 9908 7644
rect 9932 7642 9988 7644
rect 10012 7642 10068 7644
rect 10092 7642 10148 7644
rect 9852 7590 9898 7642
rect 9898 7590 9908 7642
rect 9932 7590 9962 7642
rect 9962 7590 9974 7642
rect 9974 7590 9988 7642
rect 10012 7590 10026 7642
rect 10026 7590 10038 7642
rect 10038 7590 10068 7642
rect 10092 7590 10102 7642
rect 10102 7590 10148 7642
rect 9852 7588 9908 7590
rect 9932 7588 9988 7590
rect 10012 7588 10068 7590
rect 10092 7588 10148 7590
rect 9310 5772 9366 5808
rect 9310 5752 9312 5772
rect 9312 5752 9364 5772
rect 9364 5752 9366 5772
rect 9126 4936 9182 4992
rect 8298 4392 8354 4448
rect 7628 3834 7684 3836
rect 7708 3834 7764 3836
rect 7788 3834 7844 3836
rect 7868 3834 7924 3836
rect 7628 3782 7674 3834
rect 7674 3782 7684 3834
rect 7708 3782 7738 3834
rect 7738 3782 7750 3834
rect 7750 3782 7764 3834
rect 7788 3782 7802 3834
rect 7802 3782 7814 3834
rect 7814 3782 7844 3834
rect 7868 3782 7878 3834
rect 7878 3782 7924 3834
rect 7628 3780 7684 3782
rect 7708 3780 7764 3782
rect 7788 3780 7844 3782
rect 7868 3780 7924 3782
rect 7628 2746 7684 2748
rect 7708 2746 7764 2748
rect 7788 2746 7844 2748
rect 7868 2746 7924 2748
rect 7628 2694 7674 2746
rect 7674 2694 7684 2746
rect 7708 2694 7738 2746
rect 7738 2694 7750 2746
rect 7750 2694 7764 2746
rect 7788 2694 7802 2746
rect 7802 2694 7814 2746
rect 7814 2694 7844 2746
rect 7868 2694 7878 2746
rect 7878 2694 7924 2746
rect 7628 2692 7684 2694
rect 7708 2692 7764 2694
rect 7788 2692 7844 2694
rect 7868 2692 7924 2694
rect 3606 2352 3662 2408
rect 2594 2080 2650 2136
rect 2226 1808 2282 1864
rect 2778 1536 2834 1592
rect 5404 2202 5460 2204
rect 5484 2202 5540 2204
rect 5564 2202 5620 2204
rect 5644 2202 5700 2204
rect 5404 2150 5450 2202
rect 5450 2150 5460 2202
rect 5484 2150 5514 2202
rect 5514 2150 5526 2202
rect 5526 2150 5540 2202
rect 5564 2150 5578 2202
rect 5578 2150 5590 2202
rect 5590 2150 5620 2202
rect 5644 2150 5654 2202
rect 5654 2150 5700 2202
rect 5404 2148 5460 2150
rect 5484 2148 5540 2150
rect 5564 2148 5620 2150
rect 5644 2148 5700 2150
rect 9218 4528 9274 4584
rect 8206 3576 8262 3632
rect 9770 6840 9826 6896
rect 10598 10376 10654 10432
rect 10874 11600 10930 11656
rect 10690 9560 10746 9616
rect 10598 8880 10654 8936
rect 12076 14714 12132 14716
rect 12156 14714 12212 14716
rect 12236 14714 12292 14716
rect 12316 14714 12372 14716
rect 12076 14662 12122 14714
rect 12122 14662 12132 14714
rect 12156 14662 12186 14714
rect 12186 14662 12198 14714
rect 12198 14662 12212 14714
rect 12236 14662 12250 14714
rect 12250 14662 12262 14714
rect 12262 14662 12292 14714
rect 12316 14662 12326 14714
rect 12326 14662 12372 14714
rect 12076 14660 12132 14662
rect 12156 14660 12212 14662
rect 12236 14660 12292 14662
rect 12316 14660 12372 14662
rect 11978 14456 12034 14512
rect 12076 13626 12132 13628
rect 12156 13626 12212 13628
rect 12236 13626 12292 13628
rect 12316 13626 12372 13628
rect 12076 13574 12122 13626
rect 12122 13574 12132 13626
rect 12156 13574 12186 13626
rect 12186 13574 12198 13626
rect 12198 13574 12212 13626
rect 12236 13574 12250 13626
rect 12250 13574 12262 13626
rect 12262 13574 12292 13626
rect 12316 13574 12326 13626
rect 12326 13574 12372 13626
rect 12076 13572 12132 13574
rect 12156 13572 12212 13574
rect 12236 13572 12292 13574
rect 12316 13572 12372 13574
rect 11242 11872 11298 11928
rect 11610 11500 11612 11520
rect 11612 11500 11664 11520
rect 11664 11500 11666 11520
rect 11610 11464 11666 11500
rect 11794 11464 11850 11520
rect 10874 9288 10930 9344
rect 10690 8744 10746 8800
rect 10138 7112 10194 7168
rect 9852 6554 9908 6556
rect 9932 6554 9988 6556
rect 10012 6554 10068 6556
rect 10092 6554 10148 6556
rect 9852 6502 9898 6554
rect 9898 6502 9908 6554
rect 9932 6502 9962 6554
rect 9962 6502 9974 6554
rect 9974 6502 9988 6554
rect 10012 6502 10026 6554
rect 10026 6502 10038 6554
rect 10038 6502 10068 6554
rect 10092 6502 10102 6554
rect 10102 6502 10148 6554
rect 9852 6500 9908 6502
rect 9932 6500 9988 6502
rect 10012 6500 10068 6502
rect 10092 6500 10148 6502
rect 10046 6296 10102 6352
rect 10230 6296 10286 6352
rect 10046 6024 10102 6080
rect 9852 5466 9908 5468
rect 9932 5466 9988 5468
rect 10012 5466 10068 5468
rect 10092 5466 10148 5468
rect 9852 5414 9898 5466
rect 9898 5414 9908 5466
rect 9932 5414 9962 5466
rect 9962 5414 9974 5466
rect 9974 5414 9988 5466
rect 10012 5414 10026 5466
rect 10026 5414 10038 5466
rect 10038 5414 10068 5466
rect 10092 5414 10102 5466
rect 10102 5414 10148 5466
rect 9852 5412 9908 5414
rect 9932 5412 9988 5414
rect 10012 5412 10068 5414
rect 10092 5412 10148 5414
rect 11150 9560 11206 9616
rect 11334 9152 11390 9208
rect 11334 8880 11390 8936
rect 11518 9560 11574 9616
rect 10966 8200 11022 8256
rect 10874 5616 10930 5672
rect 10782 4684 10838 4720
rect 10782 4664 10784 4684
rect 10784 4664 10836 4684
rect 10836 4664 10838 4684
rect 9852 4378 9908 4380
rect 9932 4378 9988 4380
rect 10012 4378 10068 4380
rect 10092 4378 10148 4380
rect 9852 4326 9898 4378
rect 9898 4326 9908 4378
rect 9932 4326 9962 4378
rect 9962 4326 9974 4378
rect 9974 4326 9988 4378
rect 10012 4326 10026 4378
rect 10026 4326 10038 4378
rect 10038 4326 10068 4378
rect 10092 4326 10102 4378
rect 10102 4326 10148 4378
rect 9852 4324 9908 4326
rect 9932 4324 9988 4326
rect 10012 4324 10068 4326
rect 10092 4324 10148 4326
rect 10782 3984 10838 4040
rect 9852 3290 9908 3292
rect 9932 3290 9988 3292
rect 10012 3290 10068 3292
rect 10092 3290 10148 3292
rect 9852 3238 9898 3290
rect 9898 3238 9908 3290
rect 9932 3238 9962 3290
rect 9962 3238 9974 3290
rect 9974 3238 9988 3290
rect 10012 3238 10026 3290
rect 10026 3238 10038 3290
rect 10038 3238 10068 3290
rect 10092 3238 10102 3290
rect 10102 3238 10148 3290
rect 9852 3236 9908 3238
rect 9932 3236 9988 3238
rect 10012 3236 10068 3238
rect 10092 3236 10148 3238
rect 10966 5208 11022 5264
rect 11150 6976 11206 7032
rect 11426 6432 11482 6488
rect 11242 4664 11298 4720
rect 11426 5208 11482 5264
rect 11426 4936 11482 4992
rect 11150 4528 11206 4584
rect 11150 3032 11206 3088
rect 12076 12538 12132 12540
rect 12156 12538 12212 12540
rect 12236 12538 12292 12540
rect 12316 12538 12372 12540
rect 12076 12486 12122 12538
rect 12122 12486 12132 12538
rect 12156 12486 12186 12538
rect 12186 12486 12198 12538
rect 12198 12486 12212 12538
rect 12236 12486 12250 12538
rect 12250 12486 12262 12538
rect 12262 12486 12292 12538
rect 12316 12486 12326 12538
rect 12326 12486 12372 12538
rect 12076 12484 12132 12486
rect 12156 12484 12212 12486
rect 12236 12484 12292 12486
rect 12316 12484 12372 12486
rect 12076 11450 12132 11452
rect 12156 11450 12212 11452
rect 12236 11450 12292 11452
rect 12316 11450 12372 11452
rect 12076 11398 12122 11450
rect 12122 11398 12132 11450
rect 12156 11398 12186 11450
rect 12186 11398 12198 11450
rect 12198 11398 12212 11450
rect 12236 11398 12250 11450
rect 12250 11398 12262 11450
rect 12262 11398 12292 11450
rect 12316 11398 12326 11450
rect 12326 11398 12372 11450
rect 12076 11396 12132 11398
rect 12156 11396 12212 11398
rect 12236 11396 12292 11398
rect 12316 11396 12372 11398
rect 12076 10362 12132 10364
rect 12156 10362 12212 10364
rect 12236 10362 12292 10364
rect 12316 10362 12372 10364
rect 12076 10310 12122 10362
rect 12122 10310 12132 10362
rect 12156 10310 12186 10362
rect 12186 10310 12198 10362
rect 12198 10310 12212 10362
rect 12236 10310 12250 10362
rect 12250 10310 12262 10362
rect 12262 10310 12292 10362
rect 12316 10310 12326 10362
rect 12326 10310 12372 10362
rect 12076 10308 12132 10310
rect 12156 10308 12212 10310
rect 12236 10308 12292 10310
rect 12316 10308 12372 10310
rect 12076 9274 12132 9276
rect 12156 9274 12212 9276
rect 12236 9274 12292 9276
rect 12316 9274 12372 9276
rect 12076 9222 12122 9274
rect 12122 9222 12132 9274
rect 12156 9222 12186 9274
rect 12186 9222 12198 9274
rect 12198 9222 12212 9274
rect 12236 9222 12250 9274
rect 12250 9222 12262 9274
rect 12262 9222 12292 9274
rect 12316 9222 12326 9274
rect 12326 9222 12372 9274
rect 12076 9220 12132 9222
rect 12156 9220 12212 9222
rect 12236 9220 12292 9222
rect 12316 9220 12372 9222
rect 12622 10240 12678 10296
rect 12622 9968 12678 10024
rect 13082 11736 13138 11792
rect 12070 8336 12126 8392
rect 12076 8186 12132 8188
rect 12156 8186 12212 8188
rect 12236 8186 12292 8188
rect 12316 8186 12372 8188
rect 12076 8134 12122 8186
rect 12122 8134 12132 8186
rect 12156 8134 12186 8186
rect 12186 8134 12198 8186
rect 12198 8134 12212 8186
rect 12236 8134 12250 8186
rect 12250 8134 12262 8186
rect 12262 8134 12292 8186
rect 12316 8134 12326 8186
rect 12326 8134 12372 8186
rect 12076 8132 12132 8134
rect 12156 8132 12212 8134
rect 12236 8132 12292 8134
rect 12316 8132 12372 8134
rect 12070 7792 12126 7848
rect 12076 7098 12132 7100
rect 12156 7098 12212 7100
rect 12236 7098 12292 7100
rect 12316 7098 12372 7100
rect 12076 7046 12122 7098
rect 12122 7046 12132 7098
rect 12156 7046 12186 7098
rect 12186 7046 12198 7098
rect 12198 7046 12212 7098
rect 12236 7046 12250 7098
rect 12250 7046 12262 7098
rect 12262 7046 12292 7098
rect 12316 7046 12326 7098
rect 12326 7046 12372 7098
rect 12076 7044 12132 7046
rect 12156 7044 12212 7046
rect 12236 7044 12292 7046
rect 12316 7044 12372 7046
rect 11978 6840 12034 6896
rect 12438 6704 12494 6760
rect 12254 6160 12310 6216
rect 12076 6010 12132 6012
rect 12156 6010 12212 6012
rect 12236 6010 12292 6012
rect 12316 6010 12372 6012
rect 12076 5958 12122 6010
rect 12122 5958 12132 6010
rect 12156 5958 12186 6010
rect 12186 5958 12198 6010
rect 12198 5958 12212 6010
rect 12236 5958 12250 6010
rect 12250 5958 12262 6010
rect 12262 5958 12292 6010
rect 12316 5958 12326 6010
rect 12326 5958 12372 6010
rect 12076 5956 12132 5958
rect 12156 5956 12212 5958
rect 12236 5956 12292 5958
rect 12316 5956 12372 5958
rect 12622 7656 12678 7712
rect 12070 5616 12126 5672
rect 12254 5344 12310 5400
rect 11794 4820 11850 4856
rect 11794 4800 11796 4820
rect 11796 4800 11848 4820
rect 11848 4800 11850 4820
rect 12076 4922 12132 4924
rect 12156 4922 12212 4924
rect 12236 4922 12292 4924
rect 12316 4922 12372 4924
rect 12076 4870 12122 4922
rect 12122 4870 12132 4922
rect 12156 4870 12186 4922
rect 12186 4870 12198 4922
rect 12198 4870 12212 4922
rect 12236 4870 12250 4922
rect 12250 4870 12262 4922
rect 12262 4870 12292 4922
rect 12316 4870 12326 4922
rect 12326 4870 12372 4922
rect 12076 4868 12132 4870
rect 12156 4868 12212 4870
rect 12236 4868 12292 4870
rect 12316 4868 12372 4870
rect 11978 4020 11980 4040
rect 11980 4020 12032 4040
rect 12032 4020 12034 4040
rect 11978 3984 12034 4020
rect 12076 3834 12132 3836
rect 12156 3834 12212 3836
rect 12236 3834 12292 3836
rect 12316 3834 12372 3836
rect 12076 3782 12122 3834
rect 12122 3782 12132 3834
rect 12156 3782 12186 3834
rect 12186 3782 12198 3834
rect 12198 3782 12212 3834
rect 12236 3782 12250 3834
rect 12250 3782 12262 3834
rect 12262 3782 12292 3834
rect 12316 3782 12326 3834
rect 12326 3782 12372 3834
rect 12076 3780 12132 3782
rect 12156 3780 12212 3782
rect 12236 3780 12292 3782
rect 12316 3780 12372 3782
rect 12076 2746 12132 2748
rect 12156 2746 12212 2748
rect 12236 2746 12292 2748
rect 12316 2746 12372 2748
rect 12076 2694 12122 2746
rect 12122 2694 12132 2746
rect 12156 2694 12186 2746
rect 12186 2694 12198 2746
rect 12198 2694 12212 2746
rect 12236 2694 12250 2746
rect 12250 2694 12262 2746
rect 12262 2694 12292 2746
rect 12316 2694 12326 2746
rect 12326 2694 12372 2746
rect 12076 2692 12132 2694
rect 12156 2692 12212 2694
rect 12236 2692 12292 2694
rect 12316 2692 12372 2694
rect 12990 9968 13046 10024
rect 12714 6876 12716 6896
rect 12716 6876 12768 6896
rect 12768 6876 12770 6896
rect 12714 6840 12770 6876
rect 13450 14456 13506 14512
rect 16524 14714 16580 14716
rect 16604 14714 16660 14716
rect 16684 14714 16740 14716
rect 16764 14714 16820 14716
rect 16524 14662 16570 14714
rect 16570 14662 16580 14714
rect 16604 14662 16634 14714
rect 16634 14662 16646 14714
rect 16646 14662 16660 14714
rect 16684 14662 16698 14714
rect 16698 14662 16710 14714
rect 16710 14662 16740 14714
rect 16764 14662 16774 14714
rect 16774 14662 16820 14714
rect 16524 14660 16580 14662
rect 16604 14660 16660 14662
rect 16684 14660 16740 14662
rect 16764 14660 16820 14662
rect 13450 10512 13506 10568
rect 13450 9424 13506 9480
rect 13726 10104 13782 10160
rect 14300 14170 14356 14172
rect 14380 14170 14436 14172
rect 14460 14170 14516 14172
rect 14540 14170 14596 14172
rect 14300 14118 14346 14170
rect 14346 14118 14356 14170
rect 14380 14118 14410 14170
rect 14410 14118 14422 14170
rect 14422 14118 14436 14170
rect 14460 14118 14474 14170
rect 14474 14118 14486 14170
rect 14486 14118 14516 14170
rect 14540 14118 14550 14170
rect 14550 14118 14596 14170
rect 14300 14116 14356 14118
rect 14380 14116 14436 14118
rect 14460 14116 14516 14118
rect 14540 14116 14596 14118
rect 14094 12688 14150 12744
rect 14300 13082 14356 13084
rect 14380 13082 14436 13084
rect 14460 13082 14516 13084
rect 14540 13082 14596 13084
rect 14300 13030 14346 13082
rect 14346 13030 14356 13082
rect 14380 13030 14410 13082
rect 14410 13030 14422 13082
rect 14422 13030 14436 13082
rect 14460 13030 14474 13082
rect 14474 13030 14486 13082
rect 14486 13030 14516 13082
rect 14540 13030 14550 13082
rect 14550 13030 14596 13082
rect 14300 13028 14356 13030
rect 14380 13028 14436 13030
rect 14460 13028 14516 13030
rect 14540 13028 14596 13030
rect 15382 13912 15438 13968
rect 15290 13368 15346 13424
rect 14738 12824 14794 12880
rect 14094 12008 14150 12064
rect 14300 11994 14356 11996
rect 14380 11994 14436 11996
rect 14460 11994 14516 11996
rect 14540 11994 14596 11996
rect 14300 11942 14346 11994
rect 14346 11942 14356 11994
rect 14380 11942 14410 11994
rect 14410 11942 14422 11994
rect 14422 11942 14436 11994
rect 14460 11942 14474 11994
rect 14474 11942 14486 11994
rect 14486 11942 14516 11994
rect 14540 11942 14550 11994
rect 14550 11942 14596 11994
rect 14300 11940 14356 11942
rect 14380 11940 14436 11942
rect 14460 11940 14516 11942
rect 14540 11940 14596 11942
rect 14094 11600 14150 11656
rect 13634 9424 13690 9480
rect 13542 8780 13544 8800
rect 13544 8780 13596 8800
rect 13596 8780 13598 8800
rect 13358 8472 13414 8528
rect 12990 7248 13046 7304
rect 12806 6024 12862 6080
rect 13266 5652 13268 5672
rect 13268 5652 13320 5672
rect 13320 5652 13322 5672
rect 12806 4392 12862 4448
rect 12990 4392 13046 4448
rect 13266 5616 13322 5652
rect 13174 4392 13230 4448
rect 13542 8744 13598 8780
rect 13634 7928 13690 7984
rect 13818 7248 13874 7304
rect 12990 3576 13046 3632
rect 13082 3440 13138 3496
rect 13910 6432 13966 6488
rect 13910 5516 13912 5536
rect 13912 5516 13964 5536
rect 13964 5516 13966 5536
rect 13910 5480 13966 5516
rect 13910 5364 13966 5400
rect 13910 5344 13912 5364
rect 13912 5344 13964 5364
rect 13964 5344 13966 5364
rect 14300 10906 14356 10908
rect 14380 10906 14436 10908
rect 14460 10906 14516 10908
rect 14540 10906 14596 10908
rect 14300 10854 14346 10906
rect 14346 10854 14356 10906
rect 14380 10854 14410 10906
rect 14410 10854 14422 10906
rect 14422 10854 14436 10906
rect 14460 10854 14474 10906
rect 14474 10854 14486 10906
rect 14486 10854 14516 10906
rect 14540 10854 14550 10906
rect 14550 10854 14596 10906
rect 14300 10852 14356 10854
rect 14380 10852 14436 10854
rect 14460 10852 14516 10854
rect 14540 10852 14596 10854
rect 14094 9832 14150 9888
rect 14300 9818 14356 9820
rect 14380 9818 14436 9820
rect 14460 9818 14516 9820
rect 14540 9818 14596 9820
rect 14300 9766 14346 9818
rect 14346 9766 14356 9818
rect 14380 9766 14410 9818
rect 14410 9766 14422 9818
rect 14422 9766 14436 9818
rect 14460 9766 14474 9818
rect 14474 9766 14486 9818
rect 14486 9766 14516 9818
rect 14540 9766 14550 9818
rect 14550 9766 14596 9818
rect 14300 9764 14356 9766
rect 14380 9764 14436 9766
rect 14460 9764 14516 9766
rect 14540 9764 14596 9766
rect 14300 8730 14356 8732
rect 14380 8730 14436 8732
rect 14460 8730 14516 8732
rect 14540 8730 14596 8732
rect 14300 8678 14346 8730
rect 14346 8678 14356 8730
rect 14380 8678 14410 8730
rect 14410 8678 14422 8730
rect 14422 8678 14436 8730
rect 14460 8678 14474 8730
rect 14474 8678 14486 8730
rect 14486 8678 14516 8730
rect 14540 8678 14550 8730
rect 14550 8678 14596 8730
rect 14300 8676 14356 8678
rect 14380 8676 14436 8678
rect 14460 8676 14516 8678
rect 14540 8676 14596 8678
rect 14300 7642 14356 7644
rect 14380 7642 14436 7644
rect 14460 7642 14516 7644
rect 14540 7642 14596 7644
rect 14300 7590 14346 7642
rect 14346 7590 14356 7642
rect 14380 7590 14410 7642
rect 14410 7590 14422 7642
rect 14422 7590 14436 7642
rect 14460 7590 14474 7642
rect 14474 7590 14486 7642
rect 14486 7590 14516 7642
rect 14540 7590 14550 7642
rect 14550 7590 14596 7642
rect 14300 7588 14356 7590
rect 14380 7588 14436 7590
rect 14460 7588 14516 7590
rect 14540 7588 14596 7590
rect 14300 6554 14356 6556
rect 14380 6554 14436 6556
rect 14460 6554 14516 6556
rect 14540 6554 14596 6556
rect 14300 6502 14346 6554
rect 14346 6502 14356 6554
rect 14380 6502 14410 6554
rect 14410 6502 14422 6554
rect 14422 6502 14436 6554
rect 14460 6502 14474 6554
rect 14474 6502 14486 6554
rect 14486 6502 14516 6554
rect 14540 6502 14550 6554
rect 14550 6502 14596 6554
rect 14300 6500 14356 6502
rect 14380 6500 14436 6502
rect 14460 6500 14516 6502
rect 14540 6500 14596 6502
rect 14370 6160 14426 6216
rect 14300 5466 14356 5468
rect 14380 5466 14436 5468
rect 14460 5466 14516 5468
rect 14540 5466 14596 5468
rect 14300 5414 14346 5466
rect 14346 5414 14356 5466
rect 14380 5414 14410 5466
rect 14410 5414 14422 5466
rect 14422 5414 14436 5466
rect 14460 5414 14474 5466
rect 14474 5414 14486 5466
rect 14486 5414 14516 5466
rect 14540 5414 14550 5466
rect 14550 5414 14596 5466
rect 14300 5412 14356 5414
rect 14380 5412 14436 5414
rect 14460 5412 14516 5414
rect 14540 5412 14596 5414
rect 14002 4392 14058 4448
rect 14300 4378 14356 4380
rect 14380 4378 14436 4380
rect 14460 4378 14516 4380
rect 14540 4378 14596 4380
rect 14300 4326 14346 4378
rect 14346 4326 14356 4378
rect 14380 4326 14410 4378
rect 14410 4326 14422 4378
rect 14422 4326 14436 4378
rect 14460 4326 14474 4378
rect 14474 4326 14486 4378
rect 14486 4326 14516 4378
rect 14540 4326 14550 4378
rect 14550 4326 14596 4378
rect 14300 4324 14356 4326
rect 14380 4324 14436 4326
rect 14460 4324 14516 4326
rect 14540 4324 14596 4326
rect 15198 12824 15254 12880
rect 15934 14184 15990 14240
rect 17222 13640 17278 13696
rect 16524 13626 16580 13628
rect 16604 13626 16660 13628
rect 16684 13626 16740 13628
rect 16764 13626 16820 13628
rect 16524 13574 16570 13626
rect 16570 13574 16580 13626
rect 16604 13574 16634 13626
rect 16634 13574 16646 13626
rect 16646 13574 16660 13626
rect 16684 13574 16698 13626
rect 16698 13574 16710 13626
rect 16710 13574 16740 13626
rect 16764 13574 16774 13626
rect 16774 13574 16820 13626
rect 16524 13572 16580 13574
rect 16604 13572 16660 13574
rect 16684 13572 16740 13574
rect 16764 13572 16820 13574
rect 16486 12860 16488 12880
rect 16488 12860 16540 12880
rect 16540 12860 16542 12880
rect 16486 12824 16542 12860
rect 16524 12538 16580 12540
rect 16604 12538 16660 12540
rect 16684 12538 16740 12540
rect 16764 12538 16820 12540
rect 16524 12486 16570 12538
rect 16570 12486 16580 12538
rect 16604 12486 16634 12538
rect 16634 12486 16646 12538
rect 16646 12486 16660 12538
rect 16684 12486 16698 12538
rect 16698 12486 16710 12538
rect 16710 12486 16740 12538
rect 16764 12486 16774 12538
rect 16774 12486 16820 12538
rect 16524 12484 16580 12486
rect 16604 12484 16660 12486
rect 16684 12484 16740 12486
rect 16764 12484 16820 12486
rect 15658 11736 15714 11792
rect 15198 9832 15254 9888
rect 15106 9696 15162 9752
rect 15106 9016 15162 9072
rect 15658 10376 15714 10432
rect 15106 8336 15162 8392
rect 15198 7384 15254 7440
rect 14830 5616 14886 5672
rect 14830 5208 14886 5264
rect 14738 4664 14794 4720
rect 14094 3712 14150 3768
rect 13634 3460 13690 3496
rect 13634 3440 13636 3460
rect 13636 3440 13688 3460
rect 13688 3440 13690 3460
rect 13174 3188 13230 3224
rect 13174 3168 13176 3188
rect 13176 3168 13228 3188
rect 13228 3168 13230 3188
rect 13082 2916 13138 2952
rect 13082 2896 13084 2916
rect 13084 2896 13136 2916
rect 13136 2896 13138 2916
rect 13818 3168 13874 3224
rect 14002 3168 14058 3224
rect 14300 3290 14356 3292
rect 14380 3290 14436 3292
rect 14460 3290 14516 3292
rect 14540 3290 14596 3292
rect 14300 3238 14346 3290
rect 14346 3238 14356 3290
rect 14380 3238 14410 3290
rect 14410 3238 14422 3290
rect 14422 3238 14436 3290
rect 14460 3238 14474 3290
rect 14474 3238 14486 3290
rect 14486 3238 14516 3290
rect 14540 3238 14550 3290
rect 14550 3238 14596 3290
rect 14300 3236 14356 3238
rect 14380 3236 14436 3238
rect 14460 3236 14516 3238
rect 14540 3236 14596 3238
rect 13542 2760 13598 2816
rect 13542 2624 13598 2680
rect 8114 1944 8170 2000
rect 9852 2202 9908 2204
rect 9932 2202 9988 2204
rect 10012 2202 10068 2204
rect 10092 2202 10148 2204
rect 9852 2150 9898 2202
rect 9898 2150 9908 2202
rect 9932 2150 9962 2202
rect 9962 2150 9974 2202
rect 9974 2150 9988 2202
rect 10012 2150 10026 2202
rect 10026 2150 10038 2202
rect 10038 2150 10068 2202
rect 10092 2150 10102 2202
rect 10102 2150 10148 2202
rect 9852 2148 9908 2150
rect 9932 2148 9988 2150
rect 10012 2148 10068 2150
rect 10092 2148 10148 2150
rect 13726 2488 13782 2544
rect 13910 2488 13966 2544
rect 14922 3340 14924 3360
rect 14924 3340 14976 3360
rect 14976 3340 14978 3360
rect 14922 3304 14978 3340
rect 15106 5480 15162 5536
rect 15198 5344 15254 5400
rect 15658 8472 15714 8528
rect 15566 7928 15622 7984
rect 15934 10104 15990 10160
rect 16026 8880 16082 8936
rect 16762 11600 16818 11656
rect 16524 11450 16580 11452
rect 16604 11450 16660 11452
rect 16684 11450 16740 11452
rect 16764 11450 16820 11452
rect 16524 11398 16570 11450
rect 16570 11398 16580 11450
rect 16604 11398 16634 11450
rect 16634 11398 16646 11450
rect 16646 11398 16660 11450
rect 16684 11398 16698 11450
rect 16698 11398 16710 11450
rect 16710 11398 16740 11450
rect 16764 11398 16774 11450
rect 16774 11398 16820 11450
rect 16524 11396 16580 11398
rect 16604 11396 16660 11398
rect 16684 11396 16740 11398
rect 16764 11396 16820 11398
rect 15934 7692 15936 7712
rect 15936 7692 15988 7712
rect 15988 7692 15990 7712
rect 15566 6568 15622 6624
rect 15474 6024 15530 6080
rect 15934 7656 15990 7692
rect 15566 5072 15622 5128
rect 15382 4392 15438 4448
rect 15290 3984 15346 4040
rect 15474 3712 15530 3768
rect 14646 2352 14702 2408
rect 15842 5072 15898 5128
rect 15750 2896 15806 2952
rect 14300 2202 14356 2204
rect 14380 2202 14436 2204
rect 14460 2202 14516 2204
rect 14540 2202 14596 2204
rect 14300 2150 14346 2202
rect 14346 2150 14356 2202
rect 14380 2150 14410 2202
rect 14410 2150 14422 2202
rect 14422 2150 14436 2202
rect 14460 2150 14474 2202
rect 14474 2150 14486 2202
rect 14486 2150 14516 2202
rect 14540 2150 14550 2202
rect 14550 2150 14596 2202
rect 14300 2148 14356 2150
rect 14380 2148 14436 2150
rect 14460 2148 14516 2150
rect 14540 2148 14596 2150
rect 14002 1944 14058 2000
rect 16118 7928 16174 7984
rect 16118 7656 16174 7712
rect 16524 10362 16580 10364
rect 16604 10362 16660 10364
rect 16684 10362 16740 10364
rect 16764 10362 16820 10364
rect 16524 10310 16570 10362
rect 16570 10310 16580 10362
rect 16604 10310 16634 10362
rect 16634 10310 16646 10362
rect 16646 10310 16660 10362
rect 16684 10310 16698 10362
rect 16698 10310 16710 10362
rect 16710 10310 16740 10362
rect 16764 10310 16774 10362
rect 16774 10310 16820 10362
rect 16524 10308 16580 10310
rect 16604 10308 16660 10310
rect 16684 10308 16740 10310
rect 16764 10308 16820 10310
rect 16302 9560 16358 9616
rect 16524 9274 16580 9276
rect 16604 9274 16660 9276
rect 16684 9274 16740 9276
rect 16764 9274 16820 9276
rect 16524 9222 16570 9274
rect 16570 9222 16580 9274
rect 16604 9222 16634 9274
rect 16634 9222 16646 9274
rect 16646 9222 16660 9274
rect 16684 9222 16698 9274
rect 16698 9222 16710 9274
rect 16710 9222 16740 9274
rect 16764 9222 16774 9274
rect 16774 9222 16820 9274
rect 16524 9220 16580 9222
rect 16604 9220 16660 9222
rect 16684 9220 16740 9222
rect 16764 9220 16820 9222
rect 16946 9968 17002 10024
rect 16210 5752 16266 5808
rect 16210 4392 16266 4448
rect 16524 8186 16580 8188
rect 16604 8186 16660 8188
rect 16684 8186 16740 8188
rect 16764 8186 16820 8188
rect 16524 8134 16570 8186
rect 16570 8134 16580 8186
rect 16604 8134 16634 8186
rect 16634 8134 16646 8186
rect 16646 8134 16660 8186
rect 16684 8134 16698 8186
rect 16698 8134 16710 8186
rect 16710 8134 16740 8186
rect 16764 8134 16774 8186
rect 16774 8134 16820 8186
rect 16524 8132 16580 8134
rect 16604 8132 16660 8134
rect 16684 8132 16740 8134
rect 16764 8132 16820 8134
rect 16946 9016 17002 9072
rect 16946 8200 17002 8256
rect 16394 7656 16450 7712
rect 16524 7098 16580 7100
rect 16604 7098 16660 7100
rect 16684 7098 16740 7100
rect 16764 7098 16820 7100
rect 16524 7046 16570 7098
rect 16570 7046 16580 7098
rect 16604 7046 16634 7098
rect 16634 7046 16646 7098
rect 16646 7046 16660 7098
rect 16684 7046 16698 7098
rect 16698 7046 16710 7098
rect 16710 7046 16740 7098
rect 16764 7046 16774 7098
rect 16774 7046 16820 7098
rect 16524 7044 16580 7046
rect 16604 7044 16660 7046
rect 16684 7044 16740 7046
rect 16764 7044 16820 7046
rect 16524 6010 16580 6012
rect 16604 6010 16660 6012
rect 16684 6010 16740 6012
rect 16764 6010 16820 6012
rect 16524 5958 16570 6010
rect 16570 5958 16580 6010
rect 16604 5958 16634 6010
rect 16634 5958 16646 6010
rect 16646 5958 16660 6010
rect 16684 5958 16698 6010
rect 16698 5958 16710 6010
rect 16710 5958 16740 6010
rect 16764 5958 16774 6010
rect 16774 5958 16820 6010
rect 16524 5956 16580 5958
rect 16604 5956 16660 5958
rect 16684 5956 16740 5958
rect 16764 5956 16820 5958
rect 17130 11192 17186 11248
rect 17498 13096 17554 13152
rect 17222 9968 17278 10024
rect 17222 9424 17278 9480
rect 18142 14340 18198 14376
rect 18142 14320 18144 14340
rect 18144 14320 18196 14340
rect 18196 14320 18198 14340
rect 17590 11736 17646 11792
rect 17866 12552 17922 12608
rect 17682 11192 17738 11248
rect 17774 11056 17830 11112
rect 17682 10920 17738 10976
rect 17682 10376 17738 10432
rect 17590 10140 17592 10160
rect 17592 10140 17644 10160
rect 17644 10140 17646 10160
rect 17590 10104 17646 10140
rect 17682 9968 17738 10024
rect 17590 8880 17646 8936
rect 17314 8064 17370 8120
rect 16946 6160 17002 6216
rect 17498 7520 17554 7576
rect 17130 5616 17186 5672
rect 17038 5516 17040 5536
rect 17040 5516 17092 5536
rect 17092 5516 17094 5536
rect 17038 5480 17094 5516
rect 16854 5072 16910 5128
rect 16524 4922 16580 4924
rect 16604 4922 16660 4924
rect 16684 4922 16740 4924
rect 16764 4922 16820 4924
rect 16524 4870 16570 4922
rect 16570 4870 16580 4922
rect 16604 4870 16634 4922
rect 16634 4870 16646 4922
rect 16646 4870 16660 4922
rect 16684 4870 16698 4922
rect 16698 4870 16710 4922
rect 16710 4870 16740 4922
rect 16764 4870 16774 4922
rect 16774 4870 16820 4922
rect 16524 4868 16580 4870
rect 16604 4868 16660 4870
rect 16684 4868 16740 4870
rect 16764 4868 16820 4870
rect 16762 4664 16818 4720
rect 16946 4664 17002 4720
rect 15934 3440 15990 3496
rect 16118 3440 16174 3496
rect 16524 3834 16580 3836
rect 16604 3834 16660 3836
rect 16684 3834 16740 3836
rect 16764 3834 16820 3836
rect 16524 3782 16570 3834
rect 16570 3782 16580 3834
rect 16604 3782 16634 3834
rect 16634 3782 16646 3834
rect 16646 3782 16660 3834
rect 16684 3782 16698 3834
rect 16698 3782 16710 3834
rect 16710 3782 16740 3834
rect 16764 3782 16774 3834
rect 16774 3782 16820 3834
rect 16524 3780 16580 3782
rect 16604 3780 16660 3782
rect 16684 3780 16740 3782
rect 16764 3780 16820 3782
rect 16670 3576 16726 3632
rect 16762 3304 16818 3360
rect 16210 3188 16266 3224
rect 16946 3340 16948 3360
rect 16948 3340 17000 3360
rect 17000 3340 17002 3360
rect 16946 3304 17002 3340
rect 17130 4256 17186 4312
rect 16210 3168 16212 3188
rect 16212 3168 16264 3188
rect 16264 3168 16266 3188
rect 17314 4936 17370 4992
rect 17682 6604 17684 6624
rect 17684 6604 17736 6624
rect 17736 6604 17738 6624
rect 17682 6568 17738 6604
rect 18234 13232 18290 13288
rect 18142 12300 18198 12336
rect 18142 12280 18144 12300
rect 18144 12280 18196 12300
rect 18196 12280 18198 12300
rect 17958 10648 18014 10704
rect 18142 9696 18198 9752
rect 17866 9460 17868 9480
rect 17868 9460 17920 9480
rect 17920 9460 17922 9480
rect 17866 9424 17922 9460
rect 17866 8336 17922 8392
rect 18418 12008 18474 12064
rect 18602 12280 18658 12336
rect 18510 11464 18566 11520
rect 18418 10648 18474 10704
rect 18326 10512 18382 10568
rect 18418 9288 18474 9344
rect 18418 8744 18474 8800
rect 18418 8472 18474 8528
rect 18142 6840 18198 6896
rect 17590 5788 17592 5808
rect 17592 5788 17644 5808
rect 17644 5788 17646 5808
rect 17590 5752 17646 5788
rect 17774 6296 17830 6352
rect 17682 5480 17738 5536
rect 17590 5344 17646 5400
rect 17498 4800 17554 4856
rect 17314 3612 17316 3632
rect 17316 3612 17368 3632
rect 17368 3612 17370 3632
rect 18050 6024 18106 6080
rect 17866 5208 17922 5264
rect 17682 4120 17738 4176
rect 17774 3984 17830 4040
rect 17314 3576 17370 3612
rect 17130 3052 17186 3088
rect 17130 3032 17132 3052
rect 17132 3032 17184 3052
rect 17184 3032 17186 3052
rect 16578 2916 16634 2952
rect 16578 2896 16580 2916
rect 16580 2896 16632 2916
rect 16632 2896 16634 2916
rect 16524 2746 16580 2748
rect 16604 2746 16660 2748
rect 16684 2746 16740 2748
rect 16764 2746 16820 2748
rect 16524 2694 16570 2746
rect 16570 2694 16580 2746
rect 16604 2694 16634 2746
rect 16634 2694 16646 2746
rect 16646 2694 16660 2746
rect 16684 2694 16698 2746
rect 16698 2694 16710 2746
rect 16710 2694 16740 2746
rect 16764 2694 16774 2746
rect 16774 2694 16820 2746
rect 16524 2692 16580 2694
rect 16604 2692 16660 2694
rect 16684 2692 16740 2694
rect 16764 2692 16820 2694
rect 16302 2624 16358 2680
rect 17038 2488 17094 2544
rect 17314 2488 17370 2544
rect 18510 7792 18566 7848
rect 18418 7112 18474 7168
rect 18602 6568 18658 6624
rect 18510 5752 18566 5808
rect 18234 4564 18236 4584
rect 18236 4564 18288 4584
rect 18288 4564 18290 4584
rect 18234 4528 18290 4564
rect 18418 4392 18474 4448
rect 18234 4256 18290 4312
rect 18050 3848 18106 3904
rect 17958 3440 18014 3496
rect 18234 3168 18290 3224
rect 18418 3032 18474 3088
rect 17682 2796 17684 2816
rect 17684 2796 17736 2816
rect 17736 2796 17738 2816
rect 17682 2760 17738 2796
rect 17958 2352 18014 2408
<< metal3 >>
rect 0 15466 800 15496
rect 2129 15466 2195 15469
rect 0 15464 2195 15466
rect 0 15408 2134 15464
rect 2190 15408 2195 15464
rect 0 15406 2195 15408
rect 0 15376 800 15406
rect 2129 15403 2195 15406
rect 0 15194 800 15224
rect 3049 15194 3115 15197
rect 0 15192 3115 15194
rect 0 15136 3054 15192
rect 3110 15136 3115 15192
rect 0 15134 3115 15136
rect 0 15104 800 15134
rect 3049 15131 3115 15134
rect 3969 15058 4035 15061
rect 13670 15058 13676 15060
rect 3969 15056 13676 15058
rect 3969 15000 3974 15056
rect 4030 15000 13676 15056
rect 3969 14998 13676 15000
rect 3969 14995 4035 14998
rect 13670 14996 13676 14998
rect 13740 14996 13746 15060
rect 0 14922 800 14952
rect 1853 14922 1919 14925
rect 0 14920 1919 14922
rect 0 14864 1858 14920
rect 1914 14864 1919 14920
rect 0 14862 1919 14864
rect 0 14832 800 14862
rect 1853 14859 1919 14862
rect 2773 14922 2839 14925
rect 5073 14922 5139 14925
rect 2773 14920 5139 14922
rect 2773 14864 2778 14920
rect 2834 14864 5078 14920
rect 5134 14864 5139 14920
rect 2773 14862 5139 14864
rect 2773 14859 2839 14862
rect 5073 14859 5139 14862
rect 3170 14720 3486 14721
rect 0 14650 800 14680
rect 3170 14656 3176 14720
rect 3240 14656 3256 14720
rect 3320 14656 3336 14720
rect 3400 14656 3416 14720
rect 3480 14656 3486 14720
rect 3170 14655 3486 14656
rect 7618 14720 7934 14721
rect 7618 14656 7624 14720
rect 7688 14656 7704 14720
rect 7768 14656 7784 14720
rect 7848 14656 7864 14720
rect 7928 14656 7934 14720
rect 7618 14655 7934 14656
rect 12066 14720 12382 14721
rect 12066 14656 12072 14720
rect 12136 14656 12152 14720
rect 12216 14656 12232 14720
rect 12296 14656 12312 14720
rect 12376 14656 12382 14720
rect 12066 14655 12382 14656
rect 16514 14720 16830 14721
rect 16514 14656 16520 14720
rect 16584 14656 16600 14720
rect 16664 14656 16680 14720
rect 16744 14656 16760 14720
rect 16824 14656 16830 14720
rect 16514 14655 16830 14656
rect 2957 14650 3023 14653
rect 0 14648 3023 14650
rect 0 14592 2962 14648
rect 3018 14592 3023 14648
rect 0 14590 3023 14592
rect 0 14560 800 14590
rect 2957 14587 3023 14590
rect 3509 14514 3575 14517
rect 11973 14514 12039 14517
rect 3509 14512 12039 14514
rect 3509 14456 3514 14512
rect 3570 14456 11978 14512
rect 12034 14456 12039 14512
rect 3509 14454 12039 14456
rect 3509 14451 3575 14454
rect 11973 14451 12039 14454
rect 13445 14514 13511 14517
rect 19200 14514 20000 14544
rect 13445 14512 20000 14514
rect 13445 14456 13450 14512
rect 13506 14456 20000 14512
rect 13445 14454 20000 14456
rect 13445 14451 13511 14454
rect 19200 14424 20000 14454
rect 0 14378 800 14408
rect 4061 14378 4127 14381
rect 0 14376 4127 14378
rect 0 14320 4066 14376
rect 4122 14320 4127 14376
rect 0 14318 4127 14320
rect 0 14288 800 14318
rect 4061 14315 4127 14318
rect 5073 14378 5139 14381
rect 8753 14378 8819 14381
rect 18137 14378 18203 14381
rect 5073 14376 6010 14378
rect 5073 14320 5078 14376
rect 5134 14320 6010 14376
rect 5073 14318 6010 14320
rect 5073 14315 5139 14318
rect 1945 14242 2011 14245
rect 5165 14242 5231 14245
rect 1945 14240 5231 14242
rect 1945 14184 1950 14240
rect 2006 14184 5170 14240
rect 5226 14184 5231 14240
rect 1945 14182 5231 14184
rect 5950 14242 6010 14318
rect 8753 14376 18203 14378
rect 8753 14320 8758 14376
rect 8814 14320 18142 14376
rect 18198 14320 18203 14376
rect 8753 14318 18203 14320
rect 8753 14315 8819 14318
rect 18137 14315 18203 14318
rect 15929 14242 15995 14245
rect 19200 14242 20000 14272
rect 5950 14182 9322 14242
rect 1945 14179 2011 14182
rect 5165 14179 5231 14182
rect 5394 14176 5710 14177
rect 0 14106 800 14136
rect 5394 14112 5400 14176
rect 5464 14112 5480 14176
rect 5544 14112 5560 14176
rect 5624 14112 5640 14176
rect 5704 14112 5710 14176
rect 5394 14111 5710 14112
rect 2221 14106 2287 14109
rect 0 14104 2287 14106
rect 0 14048 2226 14104
rect 2282 14048 2287 14104
rect 0 14046 2287 14048
rect 0 14016 800 14046
rect 2221 14043 2287 14046
rect 2998 14044 3004 14108
rect 3068 14106 3074 14108
rect 3509 14106 3575 14109
rect 3068 14104 3575 14106
rect 3068 14048 3514 14104
rect 3570 14048 3575 14104
rect 3068 14046 3575 14048
rect 3068 14044 3074 14046
rect 3509 14043 3575 14046
rect 1945 13970 2011 13973
rect 2773 13970 2839 13973
rect 1945 13968 2839 13970
rect 1945 13912 1950 13968
rect 2006 13912 2778 13968
rect 2834 13912 2839 13968
rect 1945 13910 2839 13912
rect 1945 13907 2011 13910
rect 2773 13907 2839 13910
rect 3049 13970 3115 13973
rect 4337 13970 4403 13973
rect 9070 13970 9076 13972
rect 3049 13968 3618 13970
rect 3049 13912 3054 13968
rect 3110 13912 3618 13968
rect 3049 13910 3618 13912
rect 3049 13907 3115 13910
rect 0 13834 800 13864
rect 3417 13834 3483 13837
rect 0 13832 3483 13834
rect 0 13776 3422 13832
rect 3478 13776 3483 13832
rect 0 13774 3483 13776
rect 3558 13834 3618 13910
rect 4337 13968 9076 13970
rect 4337 13912 4342 13968
rect 4398 13912 9076 13968
rect 4337 13910 9076 13912
rect 4337 13907 4403 13910
rect 9070 13908 9076 13910
rect 9140 13908 9146 13972
rect 9262 13970 9322 14182
rect 15929 14240 20000 14242
rect 15929 14184 15934 14240
rect 15990 14184 20000 14240
rect 15929 14182 20000 14184
rect 15929 14179 15995 14182
rect 9842 14176 10158 14177
rect 9842 14112 9848 14176
rect 9912 14112 9928 14176
rect 9992 14112 10008 14176
rect 10072 14112 10088 14176
rect 10152 14112 10158 14176
rect 9842 14111 10158 14112
rect 14290 14176 14606 14177
rect 14290 14112 14296 14176
rect 14360 14112 14376 14176
rect 14440 14112 14456 14176
rect 14520 14112 14536 14176
rect 14600 14112 14606 14176
rect 19200 14152 20000 14182
rect 14290 14111 14606 14112
rect 10358 13970 10364 13972
rect 9262 13910 10364 13970
rect 10358 13908 10364 13910
rect 10428 13908 10434 13972
rect 15377 13970 15443 13973
rect 19200 13970 20000 14000
rect 15377 13968 20000 13970
rect 15377 13912 15382 13968
rect 15438 13912 20000 13968
rect 15377 13910 20000 13912
rect 15377 13907 15443 13910
rect 19200 13880 20000 13910
rect 4613 13834 4679 13837
rect 5257 13834 5323 13837
rect 13854 13834 13860 13836
rect 3558 13832 13860 13834
rect 3558 13776 4618 13832
rect 4674 13776 5262 13832
rect 5318 13776 13860 13832
rect 3558 13774 13860 13776
rect 0 13744 800 13774
rect 3417 13771 3483 13774
rect 4613 13771 4679 13774
rect 5257 13771 5323 13774
rect 13854 13772 13860 13774
rect 13924 13772 13930 13836
rect 17217 13698 17283 13701
rect 19200 13698 20000 13728
rect 17217 13696 20000 13698
rect 17217 13640 17222 13696
rect 17278 13640 20000 13696
rect 17217 13638 20000 13640
rect 17217 13635 17283 13638
rect 3170 13632 3486 13633
rect 0 13562 800 13592
rect 3170 13568 3176 13632
rect 3240 13568 3256 13632
rect 3320 13568 3336 13632
rect 3400 13568 3416 13632
rect 3480 13568 3486 13632
rect 3170 13567 3486 13568
rect 7618 13632 7934 13633
rect 7618 13568 7624 13632
rect 7688 13568 7704 13632
rect 7768 13568 7784 13632
rect 7848 13568 7864 13632
rect 7928 13568 7934 13632
rect 7618 13567 7934 13568
rect 12066 13632 12382 13633
rect 12066 13568 12072 13632
rect 12136 13568 12152 13632
rect 12216 13568 12232 13632
rect 12296 13568 12312 13632
rect 12376 13568 12382 13632
rect 12066 13567 12382 13568
rect 16514 13632 16830 13633
rect 16514 13568 16520 13632
rect 16584 13568 16600 13632
rect 16664 13568 16680 13632
rect 16744 13568 16760 13632
rect 16824 13568 16830 13632
rect 19200 13608 20000 13638
rect 16514 13567 16830 13568
rect 2865 13562 2931 13565
rect 0 13560 2931 13562
rect 0 13504 2870 13560
rect 2926 13504 2931 13560
rect 0 13502 2931 13504
rect 0 13472 800 13502
rect 2865 13499 2931 13502
rect 1945 13426 2011 13429
rect 5073 13426 5139 13429
rect 1945 13424 5139 13426
rect 1945 13368 1950 13424
rect 2006 13368 5078 13424
rect 5134 13368 5139 13424
rect 1945 13366 5139 13368
rect 1945 13363 2011 13366
rect 5073 13363 5139 13366
rect 8477 13426 8543 13429
rect 11830 13426 11836 13428
rect 8477 13424 11836 13426
rect 8477 13368 8482 13424
rect 8538 13368 11836 13424
rect 8477 13366 11836 13368
rect 8477 13363 8543 13366
rect 11830 13364 11836 13366
rect 11900 13364 11906 13428
rect 15285 13426 15351 13429
rect 19200 13426 20000 13456
rect 15285 13424 20000 13426
rect 15285 13368 15290 13424
rect 15346 13368 20000 13424
rect 15285 13366 20000 13368
rect 15285 13363 15351 13366
rect 19200 13336 20000 13366
rect 0 13290 800 13320
rect 3969 13290 4035 13293
rect 0 13288 4035 13290
rect 0 13232 3974 13288
rect 4030 13232 4035 13288
rect 0 13230 4035 13232
rect 0 13200 800 13230
rect 3969 13227 4035 13230
rect 8753 13290 8819 13293
rect 18229 13290 18295 13293
rect 8753 13288 18295 13290
rect 8753 13232 8758 13288
rect 8814 13232 18234 13288
rect 18290 13232 18295 13288
rect 8753 13230 18295 13232
rect 8753 13227 8819 13230
rect 18229 13227 18295 13230
rect 2681 13154 2747 13157
rect 5257 13154 5323 13157
rect 2681 13152 5323 13154
rect 2681 13096 2686 13152
rect 2742 13096 5262 13152
rect 5318 13096 5323 13152
rect 2681 13094 5323 13096
rect 2681 13091 2747 13094
rect 5257 13091 5323 13094
rect 17493 13154 17559 13157
rect 19200 13154 20000 13184
rect 17493 13152 20000 13154
rect 17493 13096 17498 13152
rect 17554 13096 20000 13152
rect 17493 13094 20000 13096
rect 17493 13091 17559 13094
rect 5394 13088 5710 13089
rect 0 13018 800 13048
rect 5394 13024 5400 13088
rect 5464 13024 5480 13088
rect 5544 13024 5560 13088
rect 5624 13024 5640 13088
rect 5704 13024 5710 13088
rect 5394 13023 5710 13024
rect 9842 13088 10158 13089
rect 9842 13024 9848 13088
rect 9912 13024 9928 13088
rect 9992 13024 10008 13088
rect 10072 13024 10088 13088
rect 10152 13024 10158 13088
rect 9842 13023 10158 13024
rect 14290 13088 14606 13089
rect 14290 13024 14296 13088
rect 14360 13024 14376 13088
rect 14440 13024 14456 13088
rect 14520 13024 14536 13088
rect 14600 13024 14606 13088
rect 19200 13064 20000 13094
rect 14290 13023 14606 13024
rect 3877 13018 3943 13021
rect 0 13016 3943 13018
rect 0 12960 3882 13016
rect 3938 12960 3943 13016
rect 0 12958 3943 12960
rect 0 12928 800 12958
rect 3877 12955 3943 12958
rect 3233 12882 3299 12885
rect 9673 12882 9739 12885
rect 3233 12880 9739 12882
rect 3233 12824 3238 12880
rect 3294 12824 9678 12880
rect 9734 12824 9739 12880
rect 3233 12822 9739 12824
rect 3233 12819 3299 12822
rect 9673 12819 9739 12822
rect 10225 12882 10291 12885
rect 14733 12882 14799 12885
rect 10225 12880 14799 12882
rect 10225 12824 10230 12880
rect 10286 12824 14738 12880
rect 14794 12824 14799 12880
rect 10225 12822 14799 12824
rect 10225 12819 10291 12822
rect 14733 12819 14799 12822
rect 15193 12882 15259 12885
rect 16481 12882 16547 12885
rect 19200 12882 20000 12912
rect 15193 12880 20000 12882
rect 15193 12824 15198 12880
rect 15254 12824 16486 12880
rect 16542 12824 20000 12880
rect 15193 12822 20000 12824
rect 15193 12819 15259 12822
rect 16481 12819 16547 12822
rect 19200 12792 20000 12822
rect 0 12746 800 12776
rect 5165 12746 5231 12749
rect 7414 12746 7420 12748
rect 0 12686 4216 12746
rect 0 12656 800 12686
rect 4156 12610 4216 12686
rect 5165 12744 7420 12746
rect 5165 12688 5170 12744
rect 5226 12688 7420 12744
rect 5165 12686 7420 12688
rect 5165 12683 5231 12686
rect 7414 12684 7420 12686
rect 7484 12684 7490 12748
rect 9254 12684 9260 12748
rect 9324 12746 9330 12748
rect 9397 12746 9463 12749
rect 14089 12746 14155 12749
rect 9324 12744 9463 12746
rect 9324 12688 9402 12744
rect 9458 12688 9463 12744
rect 9324 12686 9463 12688
rect 9324 12684 9330 12686
rect 9397 12683 9463 12686
rect 9630 12744 14155 12746
rect 9630 12688 14094 12744
rect 14150 12688 14155 12744
rect 9630 12686 14155 12688
rect 5533 12610 5599 12613
rect 4156 12608 5599 12610
rect 4156 12552 5538 12608
rect 5594 12552 5599 12608
rect 4156 12550 5599 12552
rect 5533 12547 5599 12550
rect 8477 12610 8543 12613
rect 9630 12610 9690 12686
rect 14089 12683 14155 12686
rect 8477 12608 9690 12610
rect 8477 12552 8482 12608
rect 8538 12552 9690 12608
rect 8477 12550 9690 12552
rect 17861 12610 17927 12613
rect 19200 12610 20000 12640
rect 17861 12608 20000 12610
rect 17861 12552 17866 12608
rect 17922 12552 20000 12608
rect 17861 12550 20000 12552
rect 8477 12547 8543 12550
rect 17861 12547 17927 12550
rect 3170 12544 3486 12545
rect 0 12474 800 12504
rect 3170 12480 3176 12544
rect 3240 12480 3256 12544
rect 3320 12480 3336 12544
rect 3400 12480 3416 12544
rect 3480 12480 3486 12544
rect 3170 12479 3486 12480
rect 7618 12544 7934 12545
rect 7618 12480 7624 12544
rect 7688 12480 7704 12544
rect 7768 12480 7784 12544
rect 7848 12480 7864 12544
rect 7928 12480 7934 12544
rect 7618 12479 7934 12480
rect 12066 12544 12382 12545
rect 12066 12480 12072 12544
rect 12136 12480 12152 12544
rect 12216 12480 12232 12544
rect 12296 12480 12312 12544
rect 12376 12480 12382 12544
rect 12066 12479 12382 12480
rect 16514 12544 16830 12545
rect 16514 12480 16520 12544
rect 16584 12480 16600 12544
rect 16664 12480 16680 12544
rect 16744 12480 16760 12544
rect 16824 12480 16830 12544
rect 19200 12520 20000 12550
rect 16514 12479 16830 12480
rect 2773 12474 2839 12477
rect 0 12472 2839 12474
rect 0 12416 2778 12472
rect 2834 12416 2839 12472
rect 0 12414 2839 12416
rect 0 12384 800 12414
rect 2773 12411 2839 12414
rect 1669 12338 1735 12341
rect 8569 12338 8635 12341
rect 1669 12336 8635 12338
rect 1669 12280 1674 12336
rect 1730 12280 8574 12336
rect 8630 12280 8635 12336
rect 1669 12278 8635 12280
rect 1669 12275 1735 12278
rect 8569 12275 8635 12278
rect 8937 12338 9003 12341
rect 18137 12338 18203 12341
rect 8937 12336 18203 12338
rect 8937 12280 8942 12336
rect 8998 12280 18142 12336
rect 18198 12280 18203 12336
rect 8937 12278 18203 12280
rect 8937 12275 9003 12278
rect 18137 12275 18203 12278
rect 18597 12338 18663 12341
rect 19200 12338 20000 12368
rect 18597 12336 20000 12338
rect 18597 12280 18602 12336
rect 18658 12280 20000 12336
rect 18597 12278 20000 12280
rect 18597 12275 18663 12278
rect 19200 12248 20000 12278
rect 0 12202 800 12232
rect 3141 12202 3207 12205
rect 0 12200 3207 12202
rect 0 12144 3146 12200
rect 3202 12144 3207 12200
rect 0 12142 3207 12144
rect 0 12112 800 12142
rect 3141 12139 3207 12142
rect 4153 12202 4219 12205
rect 4286 12202 4292 12204
rect 4153 12200 4292 12202
rect 4153 12144 4158 12200
rect 4214 12144 4292 12200
rect 4153 12142 4292 12144
rect 4153 12139 4219 12142
rect 4286 12140 4292 12142
rect 4356 12202 4362 12204
rect 5993 12202 6059 12205
rect 4356 12200 10058 12202
rect 4356 12144 5998 12200
rect 6054 12168 10058 12200
rect 6054 12144 10426 12168
rect 4356 12142 10426 12144
rect 4356 12140 4362 12142
rect 5993 12139 6059 12142
rect 9998 12108 10426 12142
rect 2773 12066 2839 12069
rect 4245 12066 4311 12069
rect 2773 12064 4311 12066
rect 2773 12008 2778 12064
rect 2834 12008 4250 12064
rect 4306 12008 4311 12064
rect 2773 12006 4311 12008
rect 2773 12003 2839 12006
rect 4245 12003 4311 12006
rect 6453 12066 6519 12069
rect 8937 12066 9003 12069
rect 6453 12064 9003 12066
rect 6453 12008 6458 12064
rect 6514 12008 8942 12064
rect 8998 12008 9003 12064
rect 6453 12006 9003 12008
rect 10366 12066 10426 12108
rect 12934 12066 12940 12068
rect 10366 12006 12940 12066
rect 6453 12003 6519 12006
rect 8937 12003 9003 12006
rect 12934 12004 12940 12006
rect 13004 12066 13010 12068
rect 14089 12066 14155 12069
rect 13004 12064 14155 12066
rect 13004 12008 14094 12064
rect 14150 12008 14155 12064
rect 13004 12006 14155 12008
rect 13004 12004 13010 12006
rect 14089 12003 14155 12006
rect 18413 12066 18479 12069
rect 19200 12066 20000 12096
rect 18413 12064 20000 12066
rect 18413 12008 18418 12064
rect 18474 12008 20000 12064
rect 18413 12006 20000 12008
rect 18413 12003 18479 12006
rect 5394 12000 5710 12001
rect 0 11930 800 11960
rect 5394 11936 5400 12000
rect 5464 11936 5480 12000
rect 5544 11936 5560 12000
rect 5624 11936 5640 12000
rect 5704 11936 5710 12000
rect 5394 11935 5710 11936
rect 9842 12000 10158 12001
rect 9842 11936 9848 12000
rect 9912 11936 9928 12000
rect 9992 11936 10008 12000
rect 10072 11936 10088 12000
rect 10152 11936 10158 12000
rect 9842 11935 10158 11936
rect 14290 12000 14606 12001
rect 14290 11936 14296 12000
rect 14360 11936 14376 12000
rect 14440 11936 14456 12000
rect 14520 11936 14536 12000
rect 14600 11936 14606 12000
rect 19200 11976 20000 12006
rect 14290 11935 14606 11936
rect 3049 11930 3115 11933
rect 0 11928 3115 11930
rect 0 11872 3054 11928
rect 3110 11872 3115 11928
rect 0 11870 3115 11872
rect 0 11840 800 11870
rect 3049 11867 3115 11870
rect 11237 11932 11303 11933
rect 11237 11928 11284 11932
rect 11348 11930 11354 11932
rect 13486 11930 13492 11932
rect 11237 11872 11242 11928
rect 11237 11868 11284 11872
rect 11348 11870 11394 11930
rect 12758 11870 13492 11930
rect 11348 11868 11354 11870
rect 11237 11867 11303 11868
rect 2773 11794 2839 11797
rect 1350 11792 2839 11794
rect 1350 11736 2778 11792
rect 2834 11736 2839 11792
rect 1350 11734 2839 11736
rect 0 11658 800 11688
rect 1350 11658 1410 11734
rect 2773 11731 2839 11734
rect 4153 11794 4219 11797
rect 5206 11794 5212 11796
rect 4153 11792 5212 11794
rect 4153 11736 4158 11792
rect 4214 11736 5212 11792
rect 4153 11734 5212 11736
rect 4153 11731 4219 11734
rect 5206 11732 5212 11734
rect 5276 11794 5282 11796
rect 5625 11794 5691 11797
rect 5276 11792 5691 11794
rect 5276 11736 5630 11792
rect 5686 11736 5691 11792
rect 5276 11734 5691 11736
rect 5276 11732 5282 11734
rect 5625 11731 5691 11734
rect 5809 11794 5875 11797
rect 12758 11794 12818 11870
rect 13486 11868 13492 11870
rect 13556 11868 13562 11932
rect 13077 11794 13143 11797
rect 15653 11794 15719 11797
rect 5809 11792 12818 11794
rect 5809 11736 5814 11792
rect 5870 11736 12818 11792
rect 5809 11734 12818 11736
rect 12942 11792 15719 11794
rect 12942 11736 13082 11792
rect 13138 11736 15658 11792
rect 15714 11736 15719 11792
rect 12942 11734 15719 11736
rect 5809 11731 5875 11734
rect 0 11598 1410 11658
rect 2221 11658 2287 11661
rect 5901 11658 5967 11661
rect 2221 11656 5967 11658
rect 2221 11600 2226 11656
rect 2282 11600 5906 11656
rect 5962 11600 5967 11656
rect 2221 11598 5967 11600
rect 0 11568 800 11598
rect 2221 11595 2287 11598
rect 5901 11595 5967 11598
rect 10869 11658 10935 11661
rect 12942 11658 13002 11734
rect 13077 11731 13143 11734
rect 15653 11731 15719 11734
rect 17585 11794 17651 11797
rect 19200 11794 20000 11824
rect 17585 11792 20000 11794
rect 17585 11736 17590 11792
rect 17646 11736 20000 11792
rect 17585 11734 20000 11736
rect 17585 11731 17651 11734
rect 19200 11704 20000 11734
rect 10869 11656 13002 11658
rect 10869 11600 10874 11656
rect 10930 11600 13002 11656
rect 10869 11598 13002 11600
rect 14089 11658 14155 11661
rect 16757 11658 16823 11661
rect 14089 11656 16823 11658
rect 14089 11600 14094 11656
rect 14150 11600 16762 11656
rect 16818 11600 16823 11656
rect 14089 11598 16823 11600
rect 10869 11595 10935 11598
rect 14089 11595 14155 11598
rect 16757 11595 16823 11598
rect 0 11386 800 11416
rect 2224 11386 2284 11595
rect 3969 11522 4035 11525
rect 4705 11522 4771 11525
rect 6269 11522 6335 11525
rect 11605 11524 11671 11525
rect 11605 11522 11652 11524
rect 3969 11520 6335 11522
rect 3969 11464 3974 11520
rect 4030 11464 4710 11520
rect 4766 11464 6274 11520
rect 6330 11464 6335 11520
rect 3969 11462 6335 11464
rect 11560 11520 11652 11522
rect 11716 11522 11722 11524
rect 11789 11522 11855 11525
rect 11716 11520 11855 11522
rect 11560 11464 11610 11520
rect 11716 11464 11794 11520
rect 11850 11464 11855 11520
rect 11560 11462 11652 11464
rect 3969 11459 4035 11462
rect 4705 11459 4771 11462
rect 6269 11459 6335 11462
rect 11605 11460 11652 11462
rect 11716 11462 11855 11464
rect 11716 11460 11722 11462
rect 11605 11459 11671 11460
rect 11789 11459 11855 11462
rect 18505 11522 18571 11525
rect 19200 11522 20000 11552
rect 18505 11520 20000 11522
rect 18505 11464 18510 11520
rect 18566 11464 20000 11520
rect 18505 11462 20000 11464
rect 18505 11459 18571 11462
rect 3170 11456 3486 11457
rect 3170 11392 3176 11456
rect 3240 11392 3256 11456
rect 3320 11392 3336 11456
rect 3400 11392 3416 11456
rect 3480 11392 3486 11456
rect 3170 11391 3486 11392
rect 7618 11456 7934 11457
rect 7618 11392 7624 11456
rect 7688 11392 7704 11456
rect 7768 11392 7784 11456
rect 7848 11392 7864 11456
rect 7928 11392 7934 11456
rect 7618 11391 7934 11392
rect 12066 11456 12382 11457
rect 12066 11392 12072 11456
rect 12136 11392 12152 11456
rect 12216 11392 12232 11456
rect 12296 11392 12312 11456
rect 12376 11392 12382 11456
rect 12066 11391 12382 11392
rect 16514 11456 16830 11457
rect 16514 11392 16520 11456
rect 16584 11392 16600 11456
rect 16664 11392 16680 11456
rect 16744 11392 16760 11456
rect 16824 11392 16830 11456
rect 19200 11432 20000 11462
rect 16514 11391 16830 11392
rect 6453 11386 6519 11389
rect 0 11326 2284 11386
rect 3742 11384 6519 11386
rect 3742 11328 6458 11384
rect 6514 11328 6519 11384
rect 3742 11326 6519 11328
rect 0 11296 800 11326
rect 2037 11250 2103 11253
rect 2773 11250 2839 11253
rect 3742 11250 3802 11326
rect 6453 11323 6519 11326
rect 2037 11248 2514 11250
rect 2037 11192 2042 11248
rect 2098 11192 2514 11248
rect 2037 11190 2514 11192
rect 2037 11187 2103 11190
rect 0 11114 800 11144
rect 2221 11114 2287 11117
rect 0 11112 2287 11114
rect 0 11056 2226 11112
rect 2282 11056 2287 11112
rect 0 11054 2287 11056
rect 2454 11114 2514 11190
rect 2773 11248 3802 11250
rect 2773 11192 2778 11248
rect 2834 11192 3802 11248
rect 2773 11190 3802 11192
rect 3969 11250 4035 11253
rect 5717 11250 5783 11253
rect 3969 11248 5783 11250
rect 3969 11192 3974 11248
rect 4030 11192 5722 11248
rect 5778 11192 5783 11248
rect 3969 11190 5783 11192
rect 2773 11187 2839 11190
rect 3969 11187 4035 11190
rect 5717 11187 5783 11190
rect 8845 11250 8911 11253
rect 14038 11250 14044 11252
rect 8845 11248 14044 11250
rect 8845 11192 8850 11248
rect 8906 11192 14044 11248
rect 8845 11190 14044 11192
rect 8845 11187 8911 11190
rect 14038 11188 14044 11190
rect 14108 11188 14114 11252
rect 16246 11188 16252 11252
rect 16316 11250 16322 11252
rect 17125 11250 17191 11253
rect 16316 11248 17191 11250
rect 16316 11192 17130 11248
rect 17186 11192 17191 11248
rect 16316 11190 17191 11192
rect 16316 11188 16322 11190
rect 17125 11187 17191 11190
rect 17677 11250 17743 11253
rect 19200 11250 20000 11280
rect 17677 11248 20000 11250
rect 17677 11192 17682 11248
rect 17738 11192 20000 11248
rect 17677 11190 20000 11192
rect 17677 11187 17743 11190
rect 19200 11160 20000 11190
rect 4889 11114 4955 11117
rect 5809 11114 5875 11117
rect 2454 11112 5875 11114
rect 2454 11056 4894 11112
rect 4950 11056 5814 11112
rect 5870 11056 5875 11112
rect 2454 11054 5875 11056
rect 0 11024 800 11054
rect 2221 11051 2287 11054
rect 4889 11051 4955 11054
rect 5809 11051 5875 11054
rect 8937 11114 9003 11117
rect 10726 11114 10732 11116
rect 8937 11112 10732 11114
rect 8937 11056 8942 11112
rect 8998 11056 10732 11112
rect 8937 11054 10732 11056
rect 8937 11051 9003 11054
rect 10726 11052 10732 11054
rect 10796 11052 10802 11116
rect 17769 11114 17835 11117
rect 17902 11114 17908 11116
rect 17769 11112 17908 11114
rect 17769 11056 17774 11112
rect 17830 11056 17908 11112
rect 17769 11054 17908 11056
rect 17769 11051 17835 11054
rect 17902 11052 17908 11054
rect 17972 11052 17978 11116
rect 1945 10978 2011 10981
rect 4981 10978 5047 10981
rect 1945 10976 5047 10978
rect 1945 10920 1950 10976
rect 2006 10920 4986 10976
rect 5042 10920 5047 10976
rect 1945 10918 5047 10920
rect 1945 10915 2011 10918
rect 4981 10915 5047 10918
rect 17677 10978 17743 10981
rect 19200 10978 20000 11008
rect 17677 10976 20000 10978
rect 17677 10920 17682 10976
rect 17738 10920 20000 10976
rect 17677 10918 20000 10920
rect 17677 10915 17743 10918
rect 5394 10912 5710 10913
rect 0 10842 800 10872
rect 5394 10848 5400 10912
rect 5464 10848 5480 10912
rect 5544 10848 5560 10912
rect 5624 10848 5640 10912
rect 5704 10848 5710 10912
rect 5394 10847 5710 10848
rect 9842 10912 10158 10913
rect 9842 10848 9848 10912
rect 9912 10848 9928 10912
rect 9992 10848 10008 10912
rect 10072 10848 10088 10912
rect 10152 10848 10158 10912
rect 9842 10847 10158 10848
rect 14290 10912 14606 10913
rect 14290 10848 14296 10912
rect 14360 10848 14376 10912
rect 14440 10848 14456 10912
rect 14520 10848 14536 10912
rect 14600 10848 14606 10912
rect 19200 10888 20000 10918
rect 14290 10847 14606 10848
rect 2865 10842 2931 10845
rect 0 10840 2931 10842
rect 0 10784 2870 10840
rect 2926 10784 2931 10840
rect 0 10782 2931 10784
rect 0 10752 800 10782
rect 2865 10779 2931 10782
rect 3601 10842 3667 10845
rect 4153 10842 4219 10845
rect 5257 10842 5323 10845
rect 3601 10840 5323 10842
rect 3601 10784 3606 10840
rect 3662 10784 4158 10840
rect 4214 10784 5262 10840
rect 5318 10784 5323 10840
rect 3601 10782 5323 10784
rect 3601 10779 3667 10782
rect 4153 10779 4219 10782
rect 5257 10779 5323 10782
rect 7189 10842 7255 10845
rect 9581 10842 9647 10845
rect 7189 10840 9647 10842
rect 7189 10784 7194 10840
rect 7250 10784 9586 10840
rect 9642 10784 9647 10840
rect 7189 10782 9647 10784
rect 7189 10779 7255 10782
rect 9581 10779 9647 10782
rect 10225 10842 10291 10845
rect 10542 10842 10548 10844
rect 10225 10840 10548 10842
rect 10225 10784 10230 10840
rect 10286 10784 10548 10840
rect 10225 10782 10548 10784
rect 10225 10779 10291 10782
rect 10542 10780 10548 10782
rect 10612 10780 10618 10844
rect 3734 10644 3740 10708
rect 3804 10706 3810 10708
rect 3877 10706 3943 10709
rect 3804 10704 3943 10706
rect 3804 10648 3882 10704
rect 3938 10648 3943 10704
rect 3804 10646 3943 10648
rect 3804 10644 3810 10646
rect 3877 10643 3943 10646
rect 5717 10706 5783 10709
rect 17953 10706 18019 10709
rect 5717 10704 18019 10706
rect 5717 10648 5722 10704
rect 5778 10648 17958 10704
rect 18014 10648 18019 10704
rect 5717 10646 18019 10648
rect 5717 10643 5783 10646
rect 17953 10643 18019 10646
rect 18413 10706 18479 10709
rect 19200 10706 20000 10736
rect 18413 10704 20000 10706
rect 18413 10648 18418 10704
rect 18474 10648 20000 10704
rect 18413 10646 20000 10648
rect 18413 10643 18479 10646
rect 19200 10616 20000 10646
rect 0 10570 800 10600
rect 2405 10570 2471 10573
rect 0 10568 2471 10570
rect 0 10512 2410 10568
rect 2466 10512 2471 10568
rect 0 10510 2471 10512
rect 0 10480 800 10510
rect 2405 10507 2471 10510
rect 3141 10570 3207 10573
rect 5901 10570 5967 10573
rect 3141 10568 5967 10570
rect 3141 10512 3146 10568
rect 3202 10512 5906 10568
rect 5962 10512 5967 10568
rect 3141 10510 5967 10512
rect 3141 10507 3207 10510
rect 5901 10507 5967 10510
rect 6177 10570 6243 10573
rect 8845 10570 8911 10573
rect 13445 10570 13511 10573
rect 18321 10570 18387 10573
rect 6177 10568 13370 10570
rect 6177 10512 6182 10568
rect 6238 10512 8850 10568
rect 8906 10512 13370 10568
rect 6177 10510 13370 10512
rect 6177 10507 6243 10510
rect 8845 10507 8911 10510
rect 4981 10436 5047 10437
rect 4981 10434 5028 10436
rect 4936 10432 5028 10434
rect 4936 10376 4986 10432
rect 4936 10374 5028 10376
rect 4981 10372 5028 10374
rect 5092 10372 5098 10436
rect 10041 10434 10107 10437
rect 10593 10434 10659 10437
rect 10041 10432 10659 10434
rect 10041 10376 10046 10432
rect 10102 10376 10598 10432
rect 10654 10376 10659 10432
rect 10041 10374 10659 10376
rect 13310 10434 13370 10510
rect 13445 10568 18387 10570
rect 13445 10512 13450 10568
rect 13506 10512 18326 10568
rect 18382 10512 18387 10568
rect 13445 10510 18387 10512
rect 13445 10507 13511 10510
rect 18321 10507 18387 10510
rect 15653 10434 15719 10437
rect 13310 10432 15719 10434
rect 13310 10376 15658 10432
rect 15714 10376 15719 10432
rect 13310 10374 15719 10376
rect 4981 10371 5047 10372
rect 10041 10371 10107 10374
rect 10593 10371 10659 10374
rect 15653 10371 15719 10374
rect 17677 10434 17743 10437
rect 19200 10434 20000 10464
rect 17677 10432 20000 10434
rect 17677 10376 17682 10432
rect 17738 10376 20000 10432
rect 17677 10374 20000 10376
rect 17677 10371 17743 10374
rect 3170 10368 3486 10369
rect 0 10298 800 10328
rect 3170 10304 3176 10368
rect 3240 10304 3256 10368
rect 3320 10304 3336 10368
rect 3400 10304 3416 10368
rect 3480 10304 3486 10368
rect 3170 10303 3486 10304
rect 7618 10368 7934 10369
rect 7618 10304 7624 10368
rect 7688 10304 7704 10368
rect 7768 10304 7784 10368
rect 7848 10304 7864 10368
rect 7928 10304 7934 10368
rect 7618 10303 7934 10304
rect 12066 10368 12382 10369
rect 12066 10304 12072 10368
rect 12136 10304 12152 10368
rect 12216 10304 12232 10368
rect 12296 10304 12312 10368
rect 12376 10304 12382 10368
rect 12066 10303 12382 10304
rect 16514 10368 16830 10369
rect 16514 10304 16520 10368
rect 16584 10304 16600 10368
rect 16664 10304 16680 10368
rect 16744 10304 16760 10368
rect 16824 10304 16830 10368
rect 19200 10344 20000 10374
rect 16514 10303 16830 10304
rect 2773 10298 2839 10301
rect 6729 10298 6795 10301
rect 0 10296 2839 10298
rect 0 10240 2778 10296
rect 2834 10240 2839 10296
rect 0 10238 2839 10240
rect 0 10208 800 10238
rect 2773 10235 2839 10238
rect 5030 10296 6795 10298
rect 5030 10240 6734 10296
rect 6790 10240 6795 10296
rect 5030 10238 6795 10240
rect 1945 10162 2011 10165
rect 5030 10162 5090 10238
rect 6729 10235 6795 10238
rect 12617 10298 12683 10301
rect 14958 10298 14964 10300
rect 12617 10296 14964 10298
rect 12617 10240 12622 10296
rect 12678 10240 14964 10296
rect 12617 10238 14964 10240
rect 12617 10235 12683 10238
rect 14958 10236 14964 10238
rect 15028 10236 15034 10300
rect 1945 10160 5090 10162
rect 1945 10104 1950 10160
rect 2006 10104 5090 10160
rect 1945 10102 5090 10104
rect 5257 10162 5323 10165
rect 13721 10162 13787 10165
rect 5257 10160 13787 10162
rect 5257 10104 5262 10160
rect 5318 10104 13726 10160
rect 13782 10104 13787 10160
rect 5257 10102 13787 10104
rect 1945 10099 2011 10102
rect 5257 10099 5323 10102
rect 13721 10099 13787 10102
rect 15929 10162 15995 10165
rect 16982 10162 16988 10164
rect 15929 10160 16988 10162
rect 15929 10104 15934 10160
rect 15990 10104 16988 10160
rect 15929 10102 16988 10104
rect 15929 10099 15995 10102
rect 16982 10100 16988 10102
rect 17052 10100 17058 10164
rect 17585 10162 17651 10165
rect 19200 10162 20000 10192
rect 17585 10160 20000 10162
rect 17585 10104 17590 10160
rect 17646 10104 20000 10160
rect 17585 10102 20000 10104
rect 17585 10099 17651 10102
rect 19200 10072 20000 10102
rect 0 10026 800 10056
rect 1393 10026 1459 10029
rect 0 10024 1459 10026
rect 0 9968 1398 10024
rect 1454 9968 1459 10024
rect 0 9966 1459 9968
rect 0 9936 800 9966
rect 1393 9963 1459 9966
rect 3325 10026 3391 10029
rect 12617 10026 12683 10029
rect 3325 10024 12683 10026
rect 3325 9968 3330 10024
rect 3386 9968 12622 10024
rect 12678 9968 12683 10024
rect 3325 9966 12683 9968
rect 3325 9963 3391 9966
rect 12617 9963 12683 9966
rect 12985 10026 13051 10029
rect 16941 10026 17007 10029
rect 12985 10024 17007 10026
rect 12985 9968 12990 10024
rect 13046 9968 16946 10024
rect 17002 9968 17007 10024
rect 12985 9966 17007 9968
rect 12985 9963 13051 9966
rect 16941 9963 17007 9966
rect 17217 10026 17283 10029
rect 17677 10026 17743 10029
rect 17217 10024 17743 10026
rect 17217 9968 17222 10024
rect 17278 9968 17682 10024
rect 17738 9968 17743 10024
rect 17217 9966 17743 9968
rect 17217 9963 17283 9966
rect 17677 9963 17743 9966
rect 2129 9890 2195 9893
rect 4797 9890 4863 9893
rect 2129 9888 4863 9890
rect 2129 9832 2134 9888
rect 2190 9832 4802 9888
rect 4858 9832 4863 9888
rect 2129 9830 4863 9832
rect 2129 9827 2195 9830
rect 4797 9827 4863 9830
rect 5901 9890 5967 9893
rect 9213 9890 9279 9893
rect 5901 9888 9279 9890
rect 5901 9832 5906 9888
rect 5962 9832 9218 9888
rect 9274 9832 9279 9888
rect 5901 9830 9279 9832
rect 5901 9827 5967 9830
rect 9213 9827 9279 9830
rect 10225 9890 10291 9893
rect 14089 9890 14155 9893
rect 10225 9888 14155 9890
rect 10225 9832 10230 9888
rect 10286 9832 14094 9888
rect 14150 9832 14155 9888
rect 10225 9830 14155 9832
rect 10225 9827 10291 9830
rect 14089 9827 14155 9830
rect 15193 9890 15259 9893
rect 19200 9890 20000 9920
rect 15193 9888 20000 9890
rect 15193 9832 15198 9888
rect 15254 9832 20000 9888
rect 15193 9830 20000 9832
rect 15193 9827 15259 9830
rect 5394 9824 5710 9825
rect 0 9754 800 9784
rect 5394 9760 5400 9824
rect 5464 9760 5480 9824
rect 5544 9760 5560 9824
rect 5624 9760 5640 9824
rect 5704 9760 5710 9824
rect 5394 9759 5710 9760
rect 9842 9824 10158 9825
rect 9842 9760 9848 9824
rect 9912 9760 9928 9824
rect 9992 9760 10008 9824
rect 10072 9760 10088 9824
rect 10152 9760 10158 9824
rect 9842 9759 10158 9760
rect 14290 9824 14606 9825
rect 14290 9760 14296 9824
rect 14360 9760 14376 9824
rect 14440 9760 14456 9824
rect 14520 9760 14536 9824
rect 14600 9760 14606 9824
rect 19200 9800 20000 9830
rect 14290 9759 14606 9760
rect 2221 9754 2287 9757
rect 0 9752 2287 9754
rect 0 9696 2226 9752
rect 2282 9696 2287 9752
rect 0 9694 2287 9696
rect 0 9664 800 9694
rect 2221 9691 2287 9694
rect 6913 9754 6979 9757
rect 7414 9754 7420 9756
rect 6913 9752 7420 9754
rect 6913 9696 6918 9752
rect 6974 9696 7420 9752
rect 6913 9694 7420 9696
rect 6913 9691 6979 9694
rect 7414 9692 7420 9694
rect 7484 9692 7490 9756
rect 10317 9754 10383 9757
rect 10542 9754 10548 9756
rect 10317 9752 10548 9754
rect 10317 9696 10322 9752
rect 10378 9696 10548 9752
rect 10317 9694 10548 9696
rect 10317 9691 10383 9694
rect 10542 9692 10548 9694
rect 10612 9692 10618 9756
rect 15101 9754 15167 9757
rect 18137 9754 18203 9757
rect 15101 9752 18203 9754
rect 15101 9696 15106 9752
rect 15162 9696 18142 9752
rect 18198 9696 18203 9752
rect 15101 9694 18203 9696
rect 15101 9691 15167 9694
rect 18137 9691 18203 9694
rect 1945 9618 2011 9621
rect 9673 9618 9739 9621
rect 10685 9618 10751 9621
rect 1945 9616 10751 9618
rect 1945 9560 1950 9616
rect 2006 9560 9678 9616
rect 9734 9560 10690 9616
rect 10746 9560 10751 9616
rect 1945 9558 10751 9560
rect 1945 9555 2011 9558
rect 9673 9555 9739 9558
rect 10685 9555 10751 9558
rect 11145 9618 11211 9621
rect 11513 9618 11579 9621
rect 11145 9616 11579 9618
rect 11145 9560 11150 9616
rect 11206 9560 11518 9616
rect 11574 9560 11579 9616
rect 11145 9558 11579 9560
rect 11145 9555 11211 9558
rect 11513 9555 11579 9558
rect 16297 9618 16363 9621
rect 19200 9618 20000 9648
rect 16297 9616 20000 9618
rect 16297 9560 16302 9616
rect 16358 9560 20000 9616
rect 16297 9558 20000 9560
rect 16297 9555 16363 9558
rect 19200 9528 20000 9558
rect 0 9482 800 9512
rect 2773 9482 2839 9485
rect 0 9480 2839 9482
rect 0 9424 2778 9480
rect 2834 9424 2839 9480
rect 0 9422 2839 9424
rect 0 9392 800 9422
rect 2773 9419 2839 9422
rect 6545 9482 6611 9485
rect 13445 9482 13511 9485
rect 6545 9480 13511 9482
rect 6545 9424 6550 9480
rect 6606 9424 13450 9480
rect 13506 9424 13511 9480
rect 6545 9422 13511 9424
rect 6545 9419 6611 9422
rect 13445 9419 13511 9422
rect 13629 9482 13695 9485
rect 17217 9482 17283 9485
rect 17861 9484 17927 9485
rect 17861 9482 17908 9484
rect 13629 9480 17283 9482
rect 13629 9424 13634 9480
rect 13690 9424 17222 9480
rect 17278 9424 17283 9480
rect 13629 9422 17283 9424
rect 17816 9480 17908 9482
rect 17816 9424 17866 9480
rect 17816 9422 17908 9424
rect 13629 9419 13695 9422
rect 17217 9419 17283 9422
rect 17861 9420 17908 9422
rect 17972 9420 17978 9484
rect 17861 9419 17927 9420
rect 1945 9346 2011 9349
rect 2078 9346 2084 9348
rect 1945 9344 2084 9346
rect 1945 9288 1950 9344
rect 2006 9288 2084 9344
rect 1945 9286 2084 9288
rect 1945 9283 2011 9286
rect 2078 9284 2084 9286
rect 2148 9284 2154 9348
rect 9305 9346 9371 9349
rect 9949 9346 10015 9349
rect 10869 9346 10935 9349
rect 9305 9344 10935 9346
rect 9305 9288 9310 9344
rect 9366 9288 9954 9344
rect 10010 9288 10874 9344
rect 10930 9288 10935 9344
rect 9305 9286 10935 9288
rect 9305 9283 9371 9286
rect 9949 9283 10015 9286
rect 10869 9283 10935 9286
rect 18413 9346 18479 9349
rect 19200 9346 20000 9376
rect 18413 9344 20000 9346
rect 18413 9288 18418 9344
rect 18474 9288 20000 9344
rect 18413 9286 20000 9288
rect 18413 9283 18479 9286
rect 3170 9280 3486 9281
rect 0 9210 800 9240
rect 3170 9216 3176 9280
rect 3240 9216 3256 9280
rect 3320 9216 3336 9280
rect 3400 9216 3416 9280
rect 3480 9216 3486 9280
rect 3170 9215 3486 9216
rect 7618 9280 7934 9281
rect 7618 9216 7624 9280
rect 7688 9216 7704 9280
rect 7768 9216 7784 9280
rect 7848 9216 7864 9280
rect 7928 9216 7934 9280
rect 7618 9215 7934 9216
rect 12066 9280 12382 9281
rect 12066 9216 12072 9280
rect 12136 9216 12152 9280
rect 12216 9216 12232 9280
rect 12296 9216 12312 9280
rect 12376 9216 12382 9280
rect 12066 9215 12382 9216
rect 16514 9280 16830 9281
rect 16514 9216 16520 9280
rect 16584 9216 16600 9280
rect 16664 9216 16680 9280
rect 16744 9216 16760 9280
rect 16824 9216 16830 9280
rect 19200 9256 20000 9286
rect 16514 9215 16830 9216
rect 2957 9210 3023 9213
rect 0 9208 3023 9210
rect 0 9152 2962 9208
rect 3018 9152 3023 9208
rect 0 9150 3023 9152
rect 0 9120 800 9150
rect 2957 9147 3023 9150
rect 4838 9148 4844 9212
rect 4908 9210 4914 9212
rect 5349 9210 5415 9213
rect 4908 9208 5415 9210
rect 4908 9152 5354 9208
rect 5410 9152 5415 9208
rect 4908 9150 5415 9152
rect 4908 9148 4914 9150
rect 5349 9147 5415 9150
rect 10041 9210 10107 9213
rect 11329 9210 11395 9213
rect 10041 9208 11395 9210
rect 10041 9152 10046 9208
rect 10102 9152 11334 9208
rect 11390 9152 11395 9208
rect 10041 9150 11395 9152
rect 10041 9147 10107 9150
rect 11329 9147 11395 9150
rect 2865 9074 2931 9077
rect 5901 9074 5967 9077
rect 2865 9072 5967 9074
rect 2865 9016 2870 9072
rect 2926 9016 5906 9072
rect 5962 9016 5967 9072
rect 2865 9014 5967 9016
rect 2865 9011 2931 9014
rect 5901 9011 5967 9014
rect 6453 9076 6519 9077
rect 6453 9072 6500 9076
rect 6564 9074 6570 9076
rect 6729 9074 6795 9077
rect 15101 9074 15167 9077
rect 6453 9016 6458 9072
rect 6453 9012 6500 9016
rect 6564 9014 6610 9074
rect 6729 9072 15167 9074
rect 6729 9016 6734 9072
rect 6790 9016 15106 9072
rect 15162 9016 15167 9072
rect 6729 9014 15167 9016
rect 6564 9012 6570 9014
rect 6453 9011 6519 9012
rect 6729 9011 6795 9014
rect 15101 9011 15167 9014
rect 16941 9074 17007 9077
rect 19200 9074 20000 9104
rect 16941 9072 20000 9074
rect 16941 9016 16946 9072
rect 17002 9016 20000 9072
rect 16941 9014 20000 9016
rect 16941 9011 17007 9014
rect 19200 8984 20000 9014
rect 0 8938 800 8968
rect 2773 8938 2839 8941
rect 0 8936 2839 8938
rect 0 8880 2778 8936
rect 2834 8880 2839 8936
rect 0 8878 2839 8880
rect 0 8848 800 8878
rect 2773 8875 2839 8878
rect 2957 8938 3023 8941
rect 3969 8938 4035 8941
rect 8937 8938 9003 8941
rect 2957 8936 4035 8938
rect 2957 8880 2962 8936
rect 3018 8880 3974 8936
rect 4030 8880 4035 8936
rect 2957 8878 4035 8880
rect 2957 8875 3023 8878
rect 3969 8875 4035 8878
rect 5214 8936 9003 8938
rect 5214 8880 8942 8936
rect 8998 8880 9003 8936
rect 5214 8878 9003 8880
rect 2497 8802 2563 8805
rect 5214 8802 5274 8878
rect 8937 8875 9003 8878
rect 9121 8938 9187 8941
rect 10593 8938 10659 8941
rect 9121 8936 10659 8938
rect 9121 8880 9126 8936
rect 9182 8880 10598 8936
rect 10654 8880 10659 8936
rect 9121 8878 10659 8880
rect 9121 8875 9187 8878
rect 10593 8875 10659 8878
rect 11329 8938 11395 8941
rect 16021 8938 16087 8941
rect 17585 8938 17651 8941
rect 11329 8936 17651 8938
rect 11329 8880 11334 8936
rect 11390 8880 16026 8936
rect 16082 8880 17590 8936
rect 17646 8880 17651 8936
rect 11329 8878 17651 8880
rect 11329 8875 11395 8878
rect 16021 8875 16087 8878
rect 17585 8875 17651 8878
rect 2497 8800 5274 8802
rect 2497 8744 2502 8800
rect 2558 8744 5274 8800
rect 2497 8742 5274 8744
rect 6637 8802 6703 8805
rect 7046 8802 7052 8804
rect 6637 8800 7052 8802
rect 6637 8744 6642 8800
rect 6698 8744 7052 8800
rect 6637 8742 7052 8744
rect 2497 8739 2563 8742
rect 6637 8739 6703 8742
rect 7046 8740 7052 8742
rect 7116 8740 7122 8804
rect 10685 8802 10751 8805
rect 13537 8802 13603 8805
rect 10685 8800 13603 8802
rect 10685 8744 10690 8800
rect 10746 8744 13542 8800
rect 13598 8744 13603 8800
rect 10685 8742 13603 8744
rect 10685 8739 10751 8742
rect 13537 8739 13603 8742
rect 18413 8802 18479 8805
rect 19200 8802 20000 8832
rect 18413 8800 20000 8802
rect 18413 8744 18418 8800
rect 18474 8744 20000 8800
rect 18413 8742 20000 8744
rect 18413 8739 18479 8742
rect 5394 8736 5710 8737
rect 0 8666 800 8696
rect 5394 8672 5400 8736
rect 5464 8672 5480 8736
rect 5544 8672 5560 8736
rect 5624 8672 5640 8736
rect 5704 8672 5710 8736
rect 5394 8671 5710 8672
rect 9842 8736 10158 8737
rect 9842 8672 9848 8736
rect 9912 8672 9928 8736
rect 9992 8672 10008 8736
rect 10072 8672 10088 8736
rect 10152 8672 10158 8736
rect 9842 8671 10158 8672
rect 14290 8736 14606 8737
rect 14290 8672 14296 8736
rect 14360 8672 14376 8736
rect 14440 8672 14456 8736
rect 14520 8672 14536 8736
rect 14600 8672 14606 8736
rect 19200 8712 20000 8742
rect 14290 8671 14606 8672
rect 3233 8666 3299 8669
rect 0 8664 3299 8666
rect 0 8608 3238 8664
rect 3294 8608 3299 8664
rect 0 8606 3299 8608
rect 0 8576 800 8606
rect 3233 8603 3299 8606
rect 6821 8666 6887 8669
rect 8017 8666 8083 8669
rect 6821 8664 8083 8666
rect 6821 8608 6826 8664
rect 6882 8608 8022 8664
rect 8078 8608 8083 8664
rect 6821 8606 8083 8608
rect 6821 8603 6887 8606
rect 8017 8603 8083 8606
rect 1945 8530 2011 8533
rect 2262 8530 2268 8532
rect 1945 8528 2268 8530
rect 1945 8472 1950 8528
rect 2006 8472 2268 8528
rect 1945 8470 2268 8472
rect 1945 8467 2011 8470
rect 2262 8468 2268 8470
rect 2332 8468 2338 8532
rect 2589 8528 2655 8533
rect 2589 8472 2594 8528
rect 2650 8472 2655 8528
rect 2589 8467 2655 8472
rect 3693 8530 3759 8533
rect 4337 8530 4403 8533
rect 3693 8528 4403 8530
rect 3693 8472 3698 8528
rect 3754 8472 4342 8528
rect 4398 8472 4403 8528
rect 3693 8470 4403 8472
rect 3693 8467 3759 8470
rect 4337 8467 4403 8470
rect 8753 8530 8819 8533
rect 13353 8530 13419 8533
rect 15653 8530 15719 8533
rect 8753 8528 15719 8530
rect 8753 8472 8758 8528
rect 8814 8472 13358 8528
rect 13414 8472 15658 8528
rect 15714 8472 15719 8528
rect 8753 8470 15719 8472
rect 8753 8467 8819 8470
rect 13353 8467 13419 8470
rect 15653 8467 15719 8470
rect 18413 8530 18479 8533
rect 19200 8530 20000 8560
rect 18413 8528 20000 8530
rect 18413 8472 18418 8528
rect 18474 8472 20000 8528
rect 18413 8470 20000 8472
rect 18413 8467 18479 8470
rect 0 8394 800 8424
rect 2221 8394 2287 8397
rect 0 8392 2287 8394
rect 0 8336 2226 8392
rect 2282 8336 2287 8392
rect 0 8334 2287 8336
rect 2592 8394 2652 8467
rect 19200 8440 20000 8470
rect 8109 8396 8175 8397
rect 6862 8394 6868 8396
rect 2592 8334 6868 8394
rect 0 8304 800 8334
rect 2221 8331 2287 8334
rect 6862 8332 6868 8334
rect 6932 8332 6938 8396
rect 8109 8394 8156 8396
rect 8064 8392 8156 8394
rect 8064 8336 8114 8392
rect 8064 8334 8156 8336
rect 8109 8332 8156 8334
rect 8220 8332 8226 8396
rect 9857 8394 9923 8397
rect 12065 8394 12131 8397
rect 9857 8392 12131 8394
rect 9857 8336 9862 8392
rect 9918 8336 12070 8392
rect 12126 8336 12131 8392
rect 9857 8334 12131 8336
rect 8109 8331 8175 8332
rect 9857 8331 9923 8334
rect 12065 8331 12131 8334
rect 15101 8394 15167 8397
rect 17861 8394 17927 8397
rect 15101 8392 17927 8394
rect 15101 8336 15106 8392
rect 15162 8336 17866 8392
rect 17922 8336 17927 8392
rect 15101 8334 17927 8336
rect 15101 8331 15167 8334
rect 17861 8331 17927 8334
rect 8109 8258 8175 8261
rect 8661 8258 8727 8261
rect 10542 8258 10548 8260
rect 8109 8256 10548 8258
rect 8109 8200 8114 8256
rect 8170 8200 8666 8256
rect 8722 8200 10548 8256
rect 8109 8198 10548 8200
rect 8109 8195 8175 8198
rect 8661 8195 8727 8198
rect 10542 8196 10548 8198
rect 10612 8258 10618 8260
rect 10961 8258 11027 8261
rect 10612 8256 11027 8258
rect 10612 8200 10966 8256
rect 11022 8200 11027 8256
rect 10612 8198 11027 8200
rect 10612 8196 10618 8198
rect 10961 8195 11027 8198
rect 16941 8258 17007 8261
rect 19200 8258 20000 8288
rect 16941 8256 20000 8258
rect 16941 8200 16946 8256
rect 17002 8200 20000 8256
rect 16941 8198 20000 8200
rect 16941 8195 17007 8198
rect 3170 8192 3486 8193
rect 0 8122 800 8152
rect 3170 8128 3176 8192
rect 3240 8128 3256 8192
rect 3320 8128 3336 8192
rect 3400 8128 3416 8192
rect 3480 8128 3486 8192
rect 3170 8127 3486 8128
rect 7618 8192 7934 8193
rect 7618 8128 7624 8192
rect 7688 8128 7704 8192
rect 7768 8128 7784 8192
rect 7848 8128 7864 8192
rect 7928 8128 7934 8192
rect 7618 8127 7934 8128
rect 12066 8192 12382 8193
rect 12066 8128 12072 8192
rect 12136 8128 12152 8192
rect 12216 8128 12232 8192
rect 12296 8128 12312 8192
rect 12376 8128 12382 8192
rect 12066 8127 12382 8128
rect 16514 8192 16830 8193
rect 16514 8128 16520 8192
rect 16584 8128 16600 8192
rect 16664 8128 16680 8192
rect 16744 8128 16760 8192
rect 16824 8128 16830 8192
rect 19200 8168 20000 8198
rect 16514 8127 16830 8128
rect 2957 8122 3023 8125
rect 0 8120 3023 8122
rect 0 8064 2962 8120
rect 3018 8064 3023 8120
rect 0 8062 3023 8064
rect 0 8032 800 8062
rect 2957 8059 3023 8062
rect 6126 8060 6132 8124
rect 6196 8122 6202 8124
rect 7189 8122 7255 8125
rect 17309 8124 17375 8125
rect 17309 8122 17356 8124
rect 6196 8120 7255 8122
rect 6196 8064 7194 8120
rect 7250 8064 7255 8120
rect 6196 8062 7255 8064
rect 17264 8120 17356 8122
rect 17264 8064 17314 8120
rect 17264 8062 17356 8064
rect 6196 8060 6202 8062
rect 7189 8059 7255 8062
rect 17309 8060 17356 8062
rect 17420 8060 17426 8124
rect 17309 8059 17375 8060
rect 13629 7986 13695 7989
rect 15561 7986 15627 7989
rect 13629 7984 15627 7986
rect 13629 7928 13634 7984
rect 13690 7928 15566 7984
rect 15622 7928 15627 7984
rect 13629 7926 15627 7928
rect 13629 7923 13695 7926
rect 15561 7923 15627 7926
rect 16113 7986 16179 7989
rect 19200 7986 20000 8016
rect 16113 7984 20000 7986
rect 16113 7928 16118 7984
rect 16174 7928 20000 7984
rect 16113 7926 20000 7928
rect 16113 7923 16179 7926
rect 19200 7896 20000 7926
rect 0 7850 800 7880
rect 1485 7850 1551 7853
rect 0 7848 1551 7850
rect 0 7792 1490 7848
rect 1546 7792 1551 7848
rect 0 7790 1551 7792
rect 0 7760 800 7790
rect 1485 7787 1551 7790
rect 4797 7850 4863 7853
rect 10041 7850 10107 7853
rect 4797 7848 10107 7850
rect 4797 7792 4802 7848
rect 4858 7792 10046 7848
rect 10102 7792 10107 7848
rect 4797 7790 10107 7792
rect 4797 7787 4863 7790
rect 10041 7787 10107 7790
rect 12065 7850 12131 7853
rect 18505 7850 18571 7853
rect 12065 7848 18571 7850
rect 12065 7792 12070 7848
rect 12126 7792 18510 7848
rect 18566 7792 18571 7848
rect 12065 7790 18571 7792
rect 12065 7787 12131 7790
rect 12620 7717 12680 7790
rect 18505 7787 18571 7790
rect 1669 7714 1735 7717
rect 3550 7714 3556 7716
rect 1669 7712 3556 7714
rect 1669 7656 1674 7712
rect 1730 7656 3556 7712
rect 1669 7654 3556 7656
rect 1669 7651 1735 7654
rect 3550 7652 3556 7654
rect 3620 7652 3626 7716
rect 12617 7712 12683 7717
rect 15929 7716 15995 7717
rect 12617 7656 12622 7712
rect 12678 7656 12683 7712
rect 12617 7651 12683 7656
rect 15878 7652 15884 7716
rect 15948 7714 15995 7716
rect 16113 7714 16179 7717
rect 16246 7714 16252 7716
rect 15948 7712 16040 7714
rect 15990 7656 16040 7712
rect 15948 7654 16040 7656
rect 16113 7712 16252 7714
rect 16113 7656 16118 7712
rect 16174 7656 16252 7712
rect 16113 7654 16252 7656
rect 15948 7652 15995 7654
rect 15929 7651 15995 7652
rect 16113 7651 16179 7654
rect 16246 7652 16252 7654
rect 16316 7652 16322 7716
rect 16389 7714 16455 7717
rect 19200 7714 20000 7744
rect 16389 7712 20000 7714
rect 16389 7656 16394 7712
rect 16450 7656 20000 7712
rect 16389 7654 20000 7656
rect 16389 7651 16455 7654
rect 5394 7648 5710 7649
rect 0 7578 800 7608
rect 5394 7584 5400 7648
rect 5464 7584 5480 7648
rect 5544 7584 5560 7648
rect 5624 7584 5640 7648
rect 5704 7584 5710 7648
rect 5394 7583 5710 7584
rect 9842 7648 10158 7649
rect 9842 7584 9848 7648
rect 9912 7584 9928 7648
rect 9992 7584 10008 7648
rect 10072 7584 10088 7648
rect 10152 7584 10158 7648
rect 9842 7583 10158 7584
rect 14290 7648 14606 7649
rect 14290 7584 14296 7648
rect 14360 7584 14376 7648
rect 14440 7584 14456 7648
rect 14520 7584 14536 7648
rect 14600 7584 14606 7648
rect 19200 7624 20000 7654
rect 14290 7583 14606 7584
rect 2681 7578 2747 7581
rect 0 7576 2747 7578
rect 0 7520 2686 7576
rect 2742 7520 2747 7576
rect 0 7518 2747 7520
rect 0 7488 800 7518
rect 2681 7515 2747 7518
rect 2814 7516 2820 7580
rect 2884 7578 2890 7580
rect 2957 7578 3023 7581
rect 9305 7578 9371 7581
rect 17493 7578 17559 7581
rect 2884 7576 3023 7578
rect 2884 7520 2962 7576
rect 3018 7520 3023 7576
rect 2884 7518 3023 7520
rect 2884 7516 2890 7518
rect 2957 7515 3023 7518
rect 5812 7576 9371 7578
rect 5812 7520 9310 7576
rect 9366 7520 9371 7576
rect 5812 7518 9371 7520
rect 4889 7442 4955 7445
rect 5812 7442 5872 7518
rect 9305 7515 9371 7518
rect 14966 7576 17559 7578
rect 14966 7520 17498 7576
rect 17554 7520 17559 7576
rect 14966 7518 17559 7520
rect 4889 7440 5872 7442
rect 4889 7384 4894 7440
rect 4950 7384 5872 7440
rect 4889 7382 5872 7384
rect 6453 7442 6519 7445
rect 8845 7442 8911 7445
rect 14966 7442 15026 7518
rect 17493 7515 17559 7518
rect 6453 7440 15026 7442
rect 6453 7384 6458 7440
rect 6514 7384 8850 7440
rect 8906 7384 15026 7440
rect 6453 7382 15026 7384
rect 15193 7442 15259 7445
rect 19200 7442 20000 7472
rect 15193 7440 20000 7442
rect 15193 7384 15198 7440
rect 15254 7384 20000 7440
rect 15193 7382 20000 7384
rect 4889 7379 4955 7382
rect 6453 7379 6519 7382
rect 8845 7379 8911 7382
rect 15193 7379 15259 7382
rect 19200 7352 20000 7382
rect 0 7306 800 7336
rect 3049 7306 3115 7309
rect 3785 7306 3851 7309
rect 12985 7306 13051 7309
rect 0 7246 1410 7306
rect 0 7216 800 7246
rect 1350 7170 1410 7246
rect 3049 7304 13051 7306
rect 3049 7248 3054 7304
rect 3110 7248 3790 7304
rect 3846 7248 12990 7304
rect 13046 7248 13051 7304
rect 3049 7246 13051 7248
rect 3049 7243 3115 7246
rect 3785 7243 3851 7246
rect 12985 7243 13051 7246
rect 13813 7306 13879 7309
rect 17902 7306 17908 7308
rect 13813 7304 17908 7306
rect 13813 7248 13818 7304
rect 13874 7248 17908 7304
rect 13813 7246 17908 7248
rect 13813 7243 13879 7246
rect 17902 7244 17908 7246
rect 17972 7244 17978 7308
rect 2865 7170 2931 7173
rect 1350 7168 2931 7170
rect 1350 7112 2870 7168
rect 2926 7112 2931 7168
rect 1350 7110 2931 7112
rect 2865 7107 2931 7110
rect 10133 7170 10199 7173
rect 10542 7170 10548 7172
rect 10133 7168 10548 7170
rect 10133 7112 10138 7168
rect 10194 7112 10548 7168
rect 10133 7110 10548 7112
rect 10133 7107 10199 7110
rect 10542 7108 10548 7110
rect 10612 7108 10618 7172
rect 18413 7170 18479 7173
rect 19200 7170 20000 7200
rect 18413 7168 20000 7170
rect 18413 7112 18418 7168
rect 18474 7112 20000 7168
rect 18413 7110 20000 7112
rect 18413 7107 18479 7110
rect 3170 7104 3486 7105
rect 0 7034 800 7064
rect 3170 7040 3176 7104
rect 3240 7040 3256 7104
rect 3320 7040 3336 7104
rect 3400 7040 3416 7104
rect 3480 7040 3486 7104
rect 3170 7039 3486 7040
rect 7618 7104 7934 7105
rect 7618 7040 7624 7104
rect 7688 7040 7704 7104
rect 7768 7040 7784 7104
rect 7848 7040 7864 7104
rect 7928 7040 7934 7104
rect 7618 7039 7934 7040
rect 12066 7104 12382 7105
rect 12066 7040 12072 7104
rect 12136 7040 12152 7104
rect 12216 7040 12232 7104
rect 12296 7040 12312 7104
rect 12376 7040 12382 7104
rect 12066 7039 12382 7040
rect 16514 7104 16830 7105
rect 16514 7040 16520 7104
rect 16584 7040 16600 7104
rect 16664 7040 16680 7104
rect 16744 7040 16760 7104
rect 16824 7040 16830 7104
rect 19200 7080 20000 7110
rect 16514 7039 16830 7040
rect 2957 7034 3023 7037
rect 0 7032 3023 7034
rect 0 6976 2962 7032
rect 3018 6976 3023 7032
rect 0 6974 3023 6976
rect 0 6944 800 6974
rect 2957 6971 3023 6974
rect 3969 7034 4035 7037
rect 5901 7034 5967 7037
rect 3969 7032 5967 7034
rect 3969 6976 3974 7032
rect 4030 6976 5906 7032
rect 5962 6976 5967 7032
rect 3969 6974 5967 6976
rect 3969 6971 4035 6974
rect 5901 6971 5967 6974
rect 8569 7034 8635 7037
rect 11145 7034 11211 7037
rect 8569 7032 11211 7034
rect 8569 6976 8574 7032
rect 8630 6976 11150 7032
rect 11206 6976 11211 7032
rect 8569 6974 11211 6976
rect 8569 6971 8635 6974
rect 11145 6971 11211 6974
rect 2998 6836 3004 6900
rect 3068 6898 3074 6900
rect 3969 6898 4035 6901
rect 3068 6896 4035 6898
rect 3068 6840 3974 6896
rect 4030 6840 4035 6896
rect 3068 6838 4035 6840
rect 3068 6836 3074 6838
rect 3969 6835 4035 6838
rect 5022 6836 5028 6900
rect 5092 6898 5098 6900
rect 6453 6898 6519 6901
rect 6729 6900 6795 6901
rect 6678 6898 6684 6900
rect 5092 6896 6519 6898
rect 5092 6840 6458 6896
rect 6514 6840 6519 6896
rect 5092 6838 6519 6840
rect 6638 6838 6684 6898
rect 6748 6896 6795 6900
rect 6790 6840 6795 6896
rect 5092 6836 5098 6838
rect 6453 6835 6519 6838
rect 6678 6836 6684 6838
rect 6748 6836 6795 6840
rect 6729 6835 6795 6836
rect 7741 6898 7807 6901
rect 9213 6900 9279 6901
rect 8150 6898 8156 6900
rect 7741 6896 8156 6898
rect 7741 6840 7746 6896
rect 7802 6840 8156 6896
rect 7741 6838 8156 6840
rect 7741 6835 7807 6838
rect 8150 6836 8156 6838
rect 8220 6836 8226 6900
rect 9213 6896 9260 6900
rect 9324 6898 9330 6900
rect 9765 6898 9831 6901
rect 11973 6898 12039 6901
rect 12709 6900 12775 6901
rect 12709 6898 12756 6900
rect 9213 6840 9218 6896
rect 9213 6836 9260 6840
rect 9324 6838 9370 6898
rect 9765 6896 12039 6898
rect 9765 6840 9770 6896
rect 9826 6840 11978 6896
rect 12034 6840 12039 6896
rect 9765 6838 12039 6840
rect 12664 6896 12756 6898
rect 12664 6840 12714 6896
rect 12664 6838 12756 6840
rect 9324 6836 9330 6838
rect 9213 6835 9279 6836
rect 9765 6835 9831 6838
rect 11973 6835 12039 6838
rect 12709 6836 12756 6838
rect 12820 6836 12826 6900
rect 18137 6898 18203 6901
rect 19200 6898 20000 6928
rect 18137 6896 20000 6898
rect 18137 6840 18142 6896
rect 18198 6840 20000 6896
rect 18137 6838 20000 6840
rect 12709 6835 12775 6836
rect 18137 6835 18203 6838
rect 19200 6808 20000 6838
rect 0 6762 800 6792
rect 1485 6762 1551 6765
rect 0 6760 1551 6762
rect 0 6704 1490 6760
rect 1546 6704 1551 6760
rect 0 6702 1551 6704
rect 0 6672 800 6702
rect 1485 6699 1551 6702
rect 2313 6762 2379 6765
rect 2630 6762 2636 6764
rect 2313 6760 2636 6762
rect 2313 6704 2318 6760
rect 2374 6704 2636 6760
rect 2313 6702 2636 6704
rect 2313 6699 2379 6702
rect 2630 6700 2636 6702
rect 2700 6762 2706 6764
rect 4286 6762 4292 6764
rect 2700 6702 4292 6762
rect 2700 6700 2706 6702
rect 4286 6700 4292 6702
rect 4356 6700 4362 6764
rect 4429 6762 4495 6765
rect 12433 6762 12499 6765
rect 4429 6760 12499 6762
rect 4429 6704 4434 6760
rect 4490 6704 12438 6760
rect 12494 6704 12499 6760
rect 4429 6702 12499 6704
rect 4429 6699 4495 6702
rect 12433 6699 12499 6702
rect 2262 6564 2268 6628
rect 2332 6626 2338 6628
rect 5257 6626 5323 6629
rect 2332 6624 5323 6626
rect 2332 6568 5262 6624
rect 5318 6568 5323 6624
rect 2332 6566 5323 6568
rect 2332 6564 2338 6566
rect 5257 6563 5323 6566
rect 15561 6626 15627 6629
rect 17677 6626 17743 6629
rect 15561 6624 17743 6626
rect 15561 6568 15566 6624
rect 15622 6568 17682 6624
rect 17738 6568 17743 6624
rect 15561 6566 17743 6568
rect 15561 6563 15627 6566
rect 17677 6563 17743 6566
rect 18597 6626 18663 6629
rect 19200 6626 20000 6656
rect 18597 6624 20000 6626
rect 18597 6568 18602 6624
rect 18658 6568 20000 6624
rect 18597 6566 20000 6568
rect 18597 6563 18663 6566
rect 5394 6560 5710 6561
rect 0 6490 800 6520
rect 5394 6496 5400 6560
rect 5464 6496 5480 6560
rect 5544 6496 5560 6560
rect 5624 6496 5640 6560
rect 5704 6496 5710 6560
rect 5394 6495 5710 6496
rect 9842 6560 10158 6561
rect 9842 6496 9848 6560
rect 9912 6496 9928 6560
rect 9992 6496 10008 6560
rect 10072 6496 10088 6560
rect 10152 6496 10158 6560
rect 9842 6495 10158 6496
rect 14290 6560 14606 6561
rect 14290 6496 14296 6560
rect 14360 6496 14376 6560
rect 14440 6496 14456 6560
rect 14520 6496 14536 6560
rect 14600 6496 14606 6560
rect 19200 6536 20000 6566
rect 14290 6495 14606 6496
rect 2405 6490 2471 6493
rect 0 6488 2471 6490
rect 0 6432 2410 6488
rect 2466 6432 2471 6488
rect 0 6430 2471 6432
rect 0 6400 800 6430
rect 2405 6427 2471 6430
rect 3325 6490 3391 6493
rect 3918 6490 3924 6492
rect 3325 6488 3924 6490
rect 3325 6432 3330 6488
rect 3386 6432 3924 6488
rect 3325 6430 3924 6432
rect 3325 6427 3391 6430
rect 3918 6428 3924 6430
rect 3988 6490 3994 6492
rect 4889 6490 4955 6493
rect 3988 6488 4955 6490
rect 3988 6432 4894 6488
rect 4950 6432 4955 6488
rect 3988 6430 4955 6432
rect 3988 6428 3994 6430
rect 4889 6427 4955 6430
rect 7465 6490 7531 6493
rect 11421 6490 11487 6493
rect 13905 6490 13971 6493
rect 7465 6488 9690 6490
rect 7465 6432 7470 6488
rect 7526 6432 9690 6488
rect 7465 6430 9690 6432
rect 7465 6427 7531 6430
rect 3417 6354 3483 6357
rect 3969 6354 4035 6357
rect 3417 6352 4035 6354
rect 3417 6296 3422 6352
rect 3478 6296 3974 6352
rect 4030 6296 4035 6352
rect 3417 6294 4035 6296
rect 3417 6291 3483 6294
rect 3969 6291 4035 6294
rect 4981 6354 5047 6357
rect 5349 6354 5415 6357
rect 4981 6352 5415 6354
rect 4981 6296 4986 6352
rect 5042 6296 5354 6352
rect 5410 6296 5415 6352
rect 4981 6294 5415 6296
rect 4981 6291 5047 6294
rect 5349 6291 5415 6294
rect 6637 6354 6703 6357
rect 8017 6354 8083 6357
rect 6637 6352 8083 6354
rect 6637 6296 6642 6352
rect 6698 6296 8022 6352
rect 8078 6296 8083 6352
rect 6637 6294 8083 6296
rect 9630 6354 9690 6430
rect 11421 6488 13971 6490
rect 11421 6432 11426 6488
rect 11482 6432 13910 6488
rect 13966 6432 13971 6488
rect 11421 6430 13971 6432
rect 11421 6427 11487 6430
rect 13905 6427 13971 6430
rect 10041 6354 10107 6357
rect 9630 6352 10107 6354
rect 9630 6296 10046 6352
rect 10102 6296 10107 6352
rect 9630 6294 10107 6296
rect 6637 6291 6703 6294
rect 8017 6291 8083 6294
rect 10041 6291 10107 6294
rect 10225 6354 10291 6357
rect 17769 6354 17835 6357
rect 19200 6354 20000 6384
rect 10225 6352 12450 6354
rect 10225 6296 10230 6352
rect 10286 6296 12450 6352
rect 10225 6294 12450 6296
rect 10225 6291 10291 6294
rect 0 6218 800 6248
rect 1485 6218 1551 6221
rect 0 6216 1551 6218
rect 0 6160 1490 6216
rect 1546 6160 1551 6216
rect 0 6158 1551 6160
rect 0 6128 800 6158
rect 1485 6155 1551 6158
rect 1945 6218 2011 6221
rect 2078 6218 2084 6220
rect 1945 6216 2084 6218
rect 1945 6160 1950 6216
rect 2006 6160 2084 6216
rect 1945 6158 2084 6160
rect 1945 6155 2011 6158
rect 2078 6156 2084 6158
rect 2148 6156 2154 6220
rect 2865 6218 2931 6221
rect 5257 6218 5323 6221
rect 12249 6218 12315 6221
rect 2865 6216 5090 6218
rect 2865 6160 2870 6216
rect 2926 6160 5090 6216
rect 2865 6158 5090 6160
rect 2865 6155 2931 6158
rect 5030 6082 5090 6158
rect 5257 6216 12315 6218
rect 5257 6160 5262 6216
rect 5318 6160 12254 6216
rect 12310 6160 12315 6216
rect 5257 6158 12315 6160
rect 12390 6218 12450 6294
rect 17769 6352 20000 6354
rect 17769 6296 17774 6352
rect 17830 6296 20000 6352
rect 17769 6294 20000 6296
rect 17769 6291 17835 6294
rect 19200 6264 20000 6294
rect 14365 6218 14431 6221
rect 16941 6218 17007 6221
rect 12390 6216 17007 6218
rect 12390 6160 14370 6216
rect 14426 6160 16946 6216
rect 17002 6160 17007 6216
rect 12390 6158 17007 6160
rect 5257 6155 5323 6158
rect 12249 6155 12315 6158
rect 14365 6155 14431 6158
rect 16941 6155 17007 6158
rect 5901 6082 5967 6085
rect 5030 6080 5967 6082
rect 5030 6024 5906 6080
rect 5962 6024 5967 6080
rect 5030 6022 5967 6024
rect 5901 6019 5967 6022
rect 10041 6082 10107 6085
rect 11278 6082 11284 6084
rect 10041 6080 11284 6082
rect 10041 6024 10046 6080
rect 10102 6024 11284 6080
rect 10041 6022 11284 6024
rect 10041 6019 10107 6022
rect 11278 6020 11284 6022
rect 11348 6020 11354 6084
rect 12801 6082 12867 6085
rect 15469 6082 15535 6085
rect 12801 6080 15535 6082
rect 12801 6024 12806 6080
rect 12862 6024 15474 6080
rect 15530 6024 15535 6080
rect 12801 6022 15535 6024
rect 12801 6019 12867 6022
rect 15469 6019 15535 6022
rect 18045 6082 18111 6085
rect 19200 6082 20000 6112
rect 18045 6080 20000 6082
rect 18045 6024 18050 6080
rect 18106 6024 20000 6080
rect 18045 6022 20000 6024
rect 18045 6019 18111 6022
rect 3170 6016 3486 6017
rect 0 5946 800 5976
rect 3170 5952 3176 6016
rect 3240 5952 3256 6016
rect 3320 5952 3336 6016
rect 3400 5952 3416 6016
rect 3480 5952 3486 6016
rect 3170 5951 3486 5952
rect 7618 6016 7934 6017
rect 7618 5952 7624 6016
rect 7688 5952 7704 6016
rect 7768 5952 7784 6016
rect 7848 5952 7864 6016
rect 7928 5952 7934 6016
rect 7618 5951 7934 5952
rect 12066 6016 12382 6017
rect 12066 5952 12072 6016
rect 12136 5952 12152 6016
rect 12216 5952 12232 6016
rect 12296 5952 12312 6016
rect 12376 5952 12382 6016
rect 12066 5951 12382 5952
rect 16514 6016 16830 6017
rect 16514 5952 16520 6016
rect 16584 5952 16600 6016
rect 16664 5952 16680 6016
rect 16744 5952 16760 6016
rect 16824 5952 16830 6016
rect 19200 5992 20000 6022
rect 16514 5951 16830 5952
rect 1393 5946 1459 5949
rect 0 5944 1459 5946
rect 0 5888 1398 5944
rect 1454 5888 1459 5944
rect 0 5886 1459 5888
rect 0 5856 800 5886
rect 1393 5883 1459 5886
rect 5441 5946 5507 5949
rect 5942 5946 5948 5948
rect 5441 5944 5948 5946
rect 5441 5888 5446 5944
rect 5502 5888 5948 5944
rect 5441 5886 5948 5888
rect 5441 5883 5507 5886
rect 5942 5884 5948 5886
rect 6012 5884 6018 5948
rect 4838 5810 4844 5812
rect 2730 5750 4844 5810
rect 0 5674 800 5704
rect 1853 5674 1919 5677
rect 0 5672 1919 5674
rect 0 5616 1858 5672
rect 1914 5616 1919 5672
rect 0 5614 1919 5616
rect 0 5584 800 5614
rect 1853 5611 1919 5614
rect 2129 5674 2195 5677
rect 2730 5674 2790 5750
rect 4838 5748 4844 5750
rect 4908 5748 4914 5812
rect 9305 5810 9371 5813
rect 4984 5808 9371 5810
rect 4984 5752 9310 5808
rect 9366 5752 9371 5808
rect 4984 5750 9371 5752
rect 2129 5672 2790 5674
rect 2129 5616 2134 5672
rect 2190 5616 2790 5672
rect 2129 5614 2790 5616
rect 3233 5674 3299 5677
rect 4797 5674 4863 5677
rect 3233 5672 4863 5674
rect 3233 5616 3238 5672
rect 3294 5616 4802 5672
rect 4858 5616 4863 5672
rect 3233 5614 4863 5616
rect 2129 5611 2195 5614
rect 3233 5611 3299 5614
rect 4797 5611 4863 5614
rect 2313 5538 2379 5541
rect 3417 5538 3483 5541
rect 2313 5536 3483 5538
rect 2313 5480 2318 5536
rect 2374 5480 3422 5536
rect 3478 5480 3483 5536
rect 2313 5478 3483 5480
rect 2313 5475 2379 5478
rect 3417 5475 3483 5478
rect 3550 5476 3556 5540
rect 3620 5538 3626 5540
rect 4245 5538 4311 5541
rect 4984 5538 5044 5750
rect 9305 5747 9371 5750
rect 16205 5810 16271 5813
rect 17585 5810 17651 5813
rect 16205 5808 17651 5810
rect 16205 5752 16210 5808
rect 16266 5752 17590 5808
rect 17646 5752 17651 5808
rect 16205 5750 17651 5752
rect 16205 5747 16271 5750
rect 17585 5747 17651 5750
rect 18505 5810 18571 5813
rect 19200 5810 20000 5840
rect 18505 5808 20000 5810
rect 18505 5752 18510 5808
rect 18566 5752 20000 5808
rect 18505 5750 20000 5752
rect 18505 5747 18571 5750
rect 19200 5720 20000 5750
rect 6862 5612 6868 5676
rect 6932 5674 6938 5676
rect 7281 5674 7347 5677
rect 8293 5674 8359 5677
rect 6932 5672 8359 5674
rect 6932 5616 7286 5672
rect 7342 5616 8298 5672
rect 8354 5616 8359 5672
rect 6932 5614 8359 5616
rect 6932 5612 6938 5614
rect 7281 5611 7347 5614
rect 8293 5611 8359 5614
rect 8937 5674 9003 5677
rect 10869 5674 10935 5677
rect 8937 5672 10935 5674
rect 8937 5616 8942 5672
rect 8998 5616 10874 5672
rect 10930 5616 10935 5672
rect 8937 5614 10935 5616
rect 8937 5611 9003 5614
rect 10869 5611 10935 5614
rect 12065 5674 12131 5677
rect 13261 5674 13327 5677
rect 12065 5672 13327 5674
rect 12065 5616 12070 5672
rect 12126 5616 13266 5672
rect 13322 5616 13327 5672
rect 12065 5614 13327 5616
rect 12065 5611 12131 5614
rect 13261 5611 13327 5614
rect 14825 5674 14891 5677
rect 17125 5674 17191 5677
rect 14825 5672 17191 5674
rect 14825 5616 14830 5672
rect 14886 5616 17130 5672
rect 17186 5616 17191 5672
rect 14825 5614 17191 5616
rect 14825 5611 14891 5614
rect 17125 5611 17191 5614
rect 3620 5478 3986 5538
rect 3620 5476 3626 5478
rect 0 5402 800 5432
rect 2773 5402 2839 5405
rect 0 5400 2839 5402
rect 0 5344 2778 5400
rect 2834 5344 2839 5400
rect 0 5342 2839 5344
rect 0 5312 800 5342
rect 2773 5339 2839 5342
rect 3926 5269 3986 5478
rect 4245 5536 5044 5538
rect 4245 5480 4250 5536
rect 4306 5480 5044 5536
rect 4245 5478 5044 5480
rect 6177 5538 6243 5541
rect 6678 5538 6684 5540
rect 6177 5536 6684 5538
rect 6177 5480 6182 5536
rect 6238 5480 6684 5536
rect 6177 5478 6684 5480
rect 4245 5475 4311 5478
rect 6177 5475 6243 5478
rect 6678 5476 6684 5478
rect 6748 5476 6754 5540
rect 6821 5538 6887 5541
rect 7046 5538 7052 5540
rect 6821 5536 7052 5538
rect 6821 5480 6826 5536
rect 6882 5480 7052 5536
rect 6821 5478 7052 5480
rect 6821 5475 6887 5478
rect 7046 5476 7052 5478
rect 7116 5538 7122 5540
rect 8477 5538 8543 5541
rect 7116 5536 8543 5538
rect 7116 5480 8482 5536
rect 8538 5480 8543 5536
rect 7116 5478 8543 5480
rect 7116 5476 7122 5478
rect 8477 5475 8543 5478
rect 11278 5476 11284 5540
rect 11348 5538 11354 5540
rect 13905 5538 13971 5541
rect 11348 5536 13971 5538
rect 11348 5480 13910 5536
rect 13966 5480 13971 5536
rect 11348 5478 13971 5480
rect 11348 5476 11354 5478
rect 13905 5475 13971 5478
rect 15101 5538 15167 5541
rect 17033 5540 17099 5541
rect 15878 5538 15884 5540
rect 15101 5536 15884 5538
rect 15101 5480 15106 5536
rect 15162 5480 15884 5536
rect 15101 5478 15884 5480
rect 15101 5475 15167 5478
rect 15878 5476 15884 5478
rect 15948 5476 15954 5540
rect 16982 5538 16988 5540
rect 16942 5478 16988 5538
rect 17052 5536 17099 5540
rect 17094 5480 17099 5536
rect 16982 5476 16988 5478
rect 17052 5476 17099 5480
rect 17033 5475 17099 5476
rect 17677 5538 17743 5541
rect 19200 5538 20000 5568
rect 17677 5536 20000 5538
rect 17677 5480 17682 5536
rect 17738 5480 20000 5536
rect 17677 5478 20000 5480
rect 17677 5475 17743 5478
rect 5394 5472 5710 5473
rect 5394 5408 5400 5472
rect 5464 5408 5480 5472
rect 5544 5408 5560 5472
rect 5624 5408 5640 5472
rect 5704 5408 5710 5472
rect 5394 5407 5710 5408
rect 9842 5472 10158 5473
rect 9842 5408 9848 5472
rect 9912 5408 9928 5472
rect 9992 5408 10008 5472
rect 10072 5408 10088 5472
rect 10152 5408 10158 5472
rect 9842 5407 10158 5408
rect 14290 5472 14606 5473
rect 14290 5408 14296 5472
rect 14360 5408 14376 5472
rect 14440 5408 14456 5472
rect 14520 5408 14536 5472
rect 14600 5408 14606 5472
rect 19200 5448 20000 5478
rect 14290 5407 14606 5408
rect 4061 5402 4127 5405
rect 4889 5402 4955 5405
rect 5022 5402 5028 5404
rect 4061 5400 4170 5402
rect 4061 5344 4066 5400
rect 4122 5344 4170 5400
rect 4061 5339 4170 5344
rect 4889 5400 5028 5402
rect 4889 5344 4894 5400
rect 4950 5344 5028 5400
rect 4889 5342 5028 5344
rect 4889 5339 4955 5342
rect 5022 5340 5028 5342
rect 5092 5340 5098 5404
rect 6494 5340 6500 5404
rect 6564 5402 6570 5404
rect 7097 5402 7163 5405
rect 6564 5400 7163 5402
rect 6564 5344 7102 5400
rect 7158 5344 7163 5400
rect 6564 5342 7163 5344
rect 6564 5340 6570 5342
rect 7097 5339 7163 5342
rect 12249 5402 12315 5405
rect 13905 5402 13971 5405
rect 12249 5400 13971 5402
rect 12249 5344 12254 5400
rect 12310 5344 13910 5400
rect 13966 5344 13971 5400
rect 12249 5342 13971 5344
rect 12249 5339 12315 5342
rect 13905 5339 13971 5342
rect 15193 5402 15259 5405
rect 17585 5402 17651 5405
rect 15193 5400 17651 5402
rect 15193 5344 15198 5400
rect 15254 5344 17590 5400
rect 17646 5344 17651 5400
rect 15193 5342 17651 5344
rect 15193 5339 15259 5342
rect 17585 5339 17651 5342
rect 3509 5268 3575 5269
rect 3509 5266 3556 5268
rect 3464 5264 3556 5266
rect 3464 5208 3514 5264
rect 3464 5206 3556 5208
rect 3509 5204 3556 5206
rect 3620 5204 3626 5268
rect 3926 5264 4035 5269
rect 3926 5208 3974 5264
rect 4030 5208 4035 5264
rect 3926 5206 4035 5208
rect 4110 5266 4170 5339
rect 5901 5266 5967 5269
rect 6126 5266 6132 5268
rect 4110 5264 6132 5266
rect 4110 5208 5906 5264
rect 5962 5208 6132 5264
rect 4110 5206 6132 5208
rect 3509 5203 3575 5204
rect 3969 5203 4035 5206
rect 5901 5203 5967 5206
rect 6126 5204 6132 5206
rect 6196 5204 6202 5268
rect 6453 5266 6519 5269
rect 10961 5266 11027 5269
rect 6453 5264 11027 5266
rect 6453 5208 6458 5264
rect 6514 5208 10966 5264
rect 11022 5208 11027 5264
rect 6453 5206 11027 5208
rect 6453 5203 6519 5206
rect 10961 5203 11027 5206
rect 11421 5266 11487 5269
rect 14825 5266 14891 5269
rect 11421 5264 14891 5266
rect 11421 5208 11426 5264
rect 11482 5208 14830 5264
rect 14886 5208 14891 5264
rect 11421 5206 14891 5208
rect 11421 5203 11487 5206
rect 14825 5203 14891 5206
rect 17861 5266 17927 5269
rect 19200 5266 20000 5296
rect 17861 5264 20000 5266
rect 17861 5208 17866 5264
rect 17922 5208 20000 5264
rect 17861 5206 20000 5208
rect 17861 5203 17927 5206
rect 19200 5176 20000 5206
rect 0 5130 800 5160
rect 1485 5130 1551 5133
rect 0 5128 1551 5130
rect 0 5072 1490 5128
rect 1546 5072 1551 5128
rect 0 5070 1551 5072
rect 0 5040 800 5070
rect 1485 5067 1551 5070
rect 2814 5068 2820 5132
rect 2884 5130 2890 5132
rect 3417 5130 3483 5133
rect 5809 5130 5875 5133
rect 15561 5130 15627 5133
rect 2884 5128 3618 5130
rect 2884 5072 3422 5128
rect 3478 5072 3618 5128
rect 2884 5070 3618 5072
rect 2884 5068 2890 5070
rect 3417 5067 3483 5070
rect 3170 4928 3486 4929
rect 0 4858 800 4888
rect 3170 4864 3176 4928
rect 3240 4864 3256 4928
rect 3320 4864 3336 4928
rect 3400 4864 3416 4928
rect 3480 4864 3486 4928
rect 3170 4863 3486 4864
rect 2221 4858 2287 4861
rect 0 4856 2287 4858
rect 0 4800 2226 4856
rect 2282 4800 2287 4856
rect 0 4798 2287 4800
rect 0 4768 800 4798
rect 2221 4795 2287 4798
rect 3325 4722 3391 4725
rect 3558 4722 3618 5070
rect 5809 5128 15627 5130
rect 5809 5072 5814 5128
rect 5870 5072 15566 5128
rect 15622 5072 15627 5128
rect 5809 5070 15627 5072
rect 5809 5067 5875 5070
rect 15561 5067 15627 5070
rect 15837 5130 15903 5133
rect 16849 5130 16915 5133
rect 15837 5128 16915 5130
rect 15837 5072 15842 5128
rect 15898 5072 16854 5128
rect 16910 5072 16915 5128
rect 15837 5070 16915 5072
rect 15837 5067 15903 5070
rect 16849 5067 16915 5070
rect 9121 4994 9187 4997
rect 11421 4994 11487 4997
rect 9121 4992 11487 4994
rect 9121 4936 9126 4992
rect 9182 4936 11426 4992
rect 11482 4936 11487 4992
rect 9121 4934 11487 4936
rect 9121 4931 9187 4934
rect 11421 4931 11487 4934
rect 17309 4994 17375 4997
rect 19200 4994 20000 5024
rect 17309 4992 20000 4994
rect 17309 4936 17314 4992
rect 17370 4936 20000 4992
rect 17309 4934 20000 4936
rect 17309 4931 17375 4934
rect 7618 4928 7934 4929
rect 7618 4864 7624 4928
rect 7688 4864 7704 4928
rect 7768 4864 7784 4928
rect 7848 4864 7864 4928
rect 7928 4864 7934 4928
rect 7618 4863 7934 4864
rect 12066 4928 12382 4929
rect 12066 4864 12072 4928
rect 12136 4864 12152 4928
rect 12216 4864 12232 4928
rect 12296 4864 12312 4928
rect 12376 4864 12382 4928
rect 12066 4863 12382 4864
rect 16514 4928 16830 4929
rect 16514 4864 16520 4928
rect 16584 4864 16600 4928
rect 16664 4864 16680 4928
rect 16744 4864 16760 4928
rect 16824 4864 16830 4928
rect 19200 4904 20000 4934
rect 16514 4863 16830 4864
rect 4245 4858 4311 4861
rect 4838 4858 4844 4860
rect 4245 4856 4844 4858
rect 4245 4800 4250 4856
rect 4306 4800 4844 4856
rect 4245 4798 4844 4800
rect 4245 4795 4311 4798
rect 4838 4796 4844 4798
rect 4908 4796 4914 4860
rect 7097 4858 7163 4861
rect 7465 4858 7531 4861
rect 11789 4860 11855 4861
rect 11789 4858 11836 4860
rect 7097 4856 7531 4858
rect 7097 4800 7102 4856
rect 7158 4800 7470 4856
rect 7526 4800 7531 4856
rect 7097 4798 7531 4800
rect 11744 4856 11836 4858
rect 11744 4800 11794 4856
rect 11744 4798 11836 4800
rect 7097 4795 7163 4798
rect 7465 4795 7531 4798
rect 11789 4796 11836 4798
rect 11900 4796 11906 4860
rect 17350 4796 17356 4860
rect 17420 4858 17426 4860
rect 17493 4858 17559 4861
rect 17420 4856 17559 4858
rect 17420 4800 17498 4856
rect 17554 4800 17559 4856
rect 17420 4798 17559 4800
rect 17420 4796 17426 4798
rect 11789 4795 11855 4796
rect 17493 4795 17559 4798
rect 3325 4720 3618 4722
rect 3325 4664 3330 4720
rect 3386 4664 3618 4720
rect 3325 4662 3618 4664
rect 3785 4722 3851 4725
rect 10777 4724 10843 4725
rect 3918 4722 3924 4724
rect 3785 4720 3924 4722
rect 3785 4664 3790 4720
rect 3846 4664 3924 4720
rect 3785 4662 3924 4664
rect 3325 4659 3391 4662
rect 3785 4659 3851 4662
rect 3918 4660 3924 4662
rect 3988 4660 3994 4724
rect 10726 4660 10732 4724
rect 10796 4722 10843 4724
rect 11237 4722 11303 4725
rect 10796 4720 11303 4722
rect 10838 4664 11242 4720
rect 11298 4664 11303 4720
rect 10796 4662 11303 4664
rect 10796 4660 10843 4662
rect 10777 4659 10843 4660
rect 11237 4659 11303 4662
rect 14733 4722 14799 4725
rect 16757 4722 16823 4725
rect 14733 4720 16823 4722
rect 14733 4664 14738 4720
rect 14794 4664 16762 4720
rect 16818 4664 16823 4720
rect 14733 4662 16823 4664
rect 14733 4659 14799 4662
rect 16757 4659 16823 4662
rect 16941 4722 17007 4725
rect 19200 4722 20000 4752
rect 16941 4720 20000 4722
rect 16941 4664 16946 4720
rect 17002 4664 20000 4720
rect 16941 4662 20000 4664
rect 16941 4659 17007 4662
rect 19200 4632 20000 4662
rect 0 4586 800 4616
rect 1853 4586 1919 4589
rect 0 4584 1919 4586
rect 0 4528 1858 4584
rect 1914 4528 1919 4584
rect 0 4526 1919 4528
rect 0 4496 800 4526
rect 1853 4523 1919 4526
rect 2497 4586 2563 4589
rect 5073 4586 5139 4589
rect 2497 4584 5139 4586
rect 2497 4528 2502 4584
rect 2558 4528 5078 4584
rect 5134 4528 5139 4584
rect 2497 4526 5139 4528
rect 2497 4523 2563 4526
rect 5073 4523 5139 4526
rect 5942 4524 5948 4588
rect 6012 4586 6018 4588
rect 9213 4586 9279 4589
rect 6012 4584 9279 4586
rect 6012 4528 9218 4584
rect 9274 4528 9279 4584
rect 6012 4526 9279 4528
rect 6012 4524 6018 4526
rect 9213 4523 9279 4526
rect 11145 4586 11211 4589
rect 18229 4586 18295 4589
rect 11145 4584 18295 4586
rect 11145 4528 11150 4584
rect 11206 4528 18234 4584
rect 18290 4528 18295 4584
rect 11145 4526 18295 4528
rect 11145 4523 11211 4526
rect 18229 4523 18295 4526
rect 2078 4388 2084 4452
rect 2148 4450 2154 4452
rect 4153 4450 4219 4453
rect 2148 4448 4219 4450
rect 2148 4392 4158 4448
rect 4214 4392 4219 4448
rect 2148 4390 4219 4392
rect 2148 4388 2154 4390
rect 4153 4387 4219 4390
rect 7465 4450 7531 4453
rect 8293 4450 8359 4453
rect 12801 4452 12867 4453
rect 12985 4452 13051 4453
rect 12750 4450 12756 4452
rect 7465 4448 8359 4450
rect 7465 4392 7470 4448
rect 7526 4392 8298 4448
rect 8354 4392 8359 4448
rect 7465 4390 8359 4392
rect 12710 4390 12756 4450
rect 12820 4448 12867 4452
rect 12862 4392 12867 4448
rect 7465 4387 7531 4390
rect 8293 4387 8359 4390
rect 12750 4388 12756 4390
rect 12820 4388 12867 4392
rect 12934 4388 12940 4452
rect 13004 4450 13051 4452
rect 13169 4450 13235 4453
rect 13997 4450 14063 4453
rect 13004 4448 13096 4450
rect 13046 4392 13096 4448
rect 13004 4390 13096 4392
rect 13169 4448 14063 4450
rect 13169 4392 13174 4448
rect 13230 4392 14002 4448
rect 14058 4392 14063 4448
rect 13169 4390 14063 4392
rect 13004 4388 13051 4390
rect 12801 4387 12867 4388
rect 12985 4387 13051 4388
rect 13169 4387 13235 4390
rect 13997 4387 14063 4390
rect 15377 4450 15443 4453
rect 16205 4450 16271 4453
rect 15377 4448 16271 4450
rect 15377 4392 15382 4448
rect 15438 4392 16210 4448
rect 16266 4392 16271 4448
rect 15377 4390 16271 4392
rect 15377 4387 15443 4390
rect 16205 4387 16271 4390
rect 18413 4450 18479 4453
rect 19200 4450 20000 4480
rect 18413 4448 20000 4450
rect 18413 4392 18418 4448
rect 18474 4392 20000 4448
rect 18413 4390 20000 4392
rect 18413 4387 18479 4390
rect 5394 4384 5710 4385
rect 0 4314 800 4344
rect 5394 4320 5400 4384
rect 5464 4320 5480 4384
rect 5544 4320 5560 4384
rect 5624 4320 5640 4384
rect 5704 4320 5710 4384
rect 5394 4319 5710 4320
rect 9842 4384 10158 4385
rect 9842 4320 9848 4384
rect 9912 4320 9928 4384
rect 9992 4320 10008 4384
rect 10072 4320 10088 4384
rect 10152 4320 10158 4384
rect 9842 4319 10158 4320
rect 14290 4384 14606 4385
rect 14290 4320 14296 4384
rect 14360 4320 14376 4384
rect 14440 4320 14456 4384
rect 14520 4320 14536 4384
rect 14600 4320 14606 4384
rect 19200 4360 20000 4390
rect 14290 4319 14606 4320
rect 2773 4314 2839 4317
rect 3785 4316 3851 4317
rect 6913 4316 6979 4317
rect 0 4312 2839 4314
rect 0 4256 2778 4312
rect 2834 4256 2839 4312
rect 0 4254 2839 4256
rect 0 4224 800 4254
rect 2773 4251 2839 4254
rect 3734 4252 3740 4316
rect 3804 4314 3851 4316
rect 3804 4312 3896 4314
rect 3846 4256 3896 4312
rect 3804 4254 3896 4256
rect 3804 4252 3851 4254
rect 6862 4252 6868 4316
rect 6932 4314 6979 4316
rect 6932 4312 7024 4314
rect 6974 4256 7024 4312
rect 6932 4254 7024 4256
rect 17125 4312 17191 4317
rect 17125 4256 17130 4312
rect 17186 4256 17191 4312
rect 6932 4252 6979 4254
rect 3785 4251 3851 4252
rect 6913 4251 6979 4252
rect 17125 4251 17191 4256
rect 17902 4252 17908 4316
rect 17972 4314 17978 4316
rect 18229 4314 18295 4317
rect 17972 4312 18295 4314
rect 17972 4256 18234 4312
rect 18290 4256 18295 4312
rect 17972 4254 18295 4256
rect 17972 4252 17978 4254
rect 18229 4251 18295 4254
rect 1301 4178 1367 4181
rect 4981 4178 5047 4181
rect 7465 4180 7531 4181
rect 1301 4176 5047 4178
rect 1301 4120 1306 4176
rect 1362 4120 4986 4176
rect 5042 4120 5047 4176
rect 1301 4118 5047 4120
rect 1301 4115 1367 4118
rect 4981 4115 5047 4118
rect 7414 4116 7420 4180
rect 7484 4178 7531 4180
rect 17128 4178 17188 4251
rect 7484 4176 7576 4178
rect 7526 4120 7576 4176
rect 7484 4118 7576 4120
rect 14598 4118 17188 4178
rect 17677 4178 17743 4181
rect 19200 4178 20000 4208
rect 17677 4176 20000 4178
rect 17677 4120 17682 4176
rect 17738 4120 20000 4176
rect 17677 4118 20000 4120
rect 7484 4116 7531 4118
rect 7465 4115 7531 4116
rect 0 4042 800 4072
rect 1485 4042 1551 4045
rect 2681 4044 2747 4045
rect 2630 4042 2636 4044
rect 0 4040 1551 4042
rect 0 3984 1490 4040
rect 1546 3984 1551 4040
rect 0 3982 1551 3984
rect 2590 3982 2636 4042
rect 2700 4042 2747 4044
rect 3417 4042 3483 4045
rect 2700 4040 3483 4042
rect 2742 3984 3422 4040
rect 3478 3984 3483 4040
rect 0 3952 800 3982
rect 1485 3979 1551 3982
rect 2630 3980 2636 3982
rect 2700 3982 3483 3984
rect 2700 3980 2747 3982
rect 2681 3979 2747 3980
rect 3417 3979 3483 3982
rect 7230 3980 7236 4044
rect 7300 4042 7306 4044
rect 10777 4042 10843 4045
rect 7300 4040 10843 4042
rect 7300 3984 10782 4040
rect 10838 3984 10843 4040
rect 7300 3982 10843 3984
rect 7300 3980 7306 3982
rect 10777 3979 10843 3982
rect 11973 4042 12039 4045
rect 14598 4042 14658 4118
rect 17677 4115 17743 4118
rect 19200 4088 20000 4118
rect 11973 4040 14658 4042
rect 11973 3984 11978 4040
rect 12034 3984 14658 4040
rect 11973 3982 14658 3984
rect 15285 4042 15351 4045
rect 17769 4042 17835 4045
rect 15285 4040 17835 4042
rect 15285 3984 15290 4040
rect 15346 3984 17774 4040
rect 17830 3984 17835 4040
rect 15285 3982 17835 3984
rect 11973 3979 12039 3982
rect 15285 3979 15351 3982
rect 17769 3979 17835 3982
rect 18045 3906 18111 3909
rect 19200 3906 20000 3936
rect 18045 3904 20000 3906
rect 18045 3848 18050 3904
rect 18106 3848 20000 3904
rect 18045 3846 20000 3848
rect 18045 3843 18111 3846
rect 3170 3840 3486 3841
rect 0 3770 800 3800
rect 3170 3776 3176 3840
rect 3240 3776 3256 3840
rect 3320 3776 3336 3840
rect 3400 3776 3416 3840
rect 3480 3776 3486 3840
rect 3170 3775 3486 3776
rect 7618 3840 7934 3841
rect 7618 3776 7624 3840
rect 7688 3776 7704 3840
rect 7768 3776 7784 3840
rect 7848 3776 7864 3840
rect 7928 3776 7934 3840
rect 7618 3775 7934 3776
rect 12066 3840 12382 3841
rect 12066 3776 12072 3840
rect 12136 3776 12152 3840
rect 12216 3776 12232 3840
rect 12296 3776 12312 3840
rect 12376 3776 12382 3840
rect 12066 3775 12382 3776
rect 16514 3840 16830 3841
rect 16514 3776 16520 3840
rect 16584 3776 16600 3840
rect 16664 3776 16680 3840
rect 16744 3776 16760 3840
rect 16824 3776 16830 3840
rect 19200 3816 20000 3846
rect 16514 3775 16830 3776
rect 2221 3770 2287 3773
rect 14089 3770 14155 3773
rect 15469 3770 15535 3773
rect 0 3768 2287 3770
rect 0 3712 2226 3768
rect 2282 3712 2287 3768
rect 0 3710 2287 3712
rect 0 3680 800 3710
rect 2221 3707 2287 3710
rect 12758 3768 15535 3770
rect 12758 3712 14094 3768
rect 14150 3712 15474 3768
rect 15530 3712 15535 3768
rect 12758 3710 15535 3712
rect 8201 3634 8267 3637
rect 12758 3634 12818 3710
rect 14089 3707 14155 3710
rect 15469 3707 15535 3710
rect 8201 3632 12818 3634
rect 8201 3576 8206 3632
rect 8262 3576 12818 3632
rect 8201 3574 12818 3576
rect 12985 3634 13051 3637
rect 16665 3634 16731 3637
rect 12985 3632 16731 3634
rect 12985 3576 12990 3632
rect 13046 3576 16670 3632
rect 16726 3576 16731 3632
rect 12985 3574 16731 3576
rect 8201 3571 8267 3574
rect 12985 3571 13051 3574
rect 16665 3571 16731 3574
rect 17309 3634 17375 3637
rect 19200 3634 20000 3664
rect 17309 3632 20000 3634
rect 17309 3576 17314 3632
rect 17370 3576 20000 3632
rect 17309 3574 20000 3576
rect 17309 3571 17375 3574
rect 19200 3544 20000 3574
rect 0 3498 800 3528
rect 1945 3498 2011 3501
rect 0 3496 2011 3498
rect 0 3440 1950 3496
rect 2006 3440 2011 3496
rect 0 3438 2011 3440
rect 0 3408 800 3438
rect 1945 3435 2011 3438
rect 2773 3498 2839 3501
rect 4705 3498 4771 3501
rect 2773 3496 4771 3498
rect 2773 3440 2778 3496
rect 2834 3440 4710 3496
rect 4766 3440 4771 3496
rect 2773 3438 4771 3440
rect 2773 3435 2839 3438
rect 4705 3435 4771 3438
rect 9070 3436 9076 3500
rect 9140 3498 9146 3500
rect 13077 3498 13143 3501
rect 9140 3496 13143 3498
rect 9140 3440 13082 3496
rect 13138 3440 13143 3496
rect 9140 3438 13143 3440
rect 9140 3436 9146 3438
rect 13077 3435 13143 3438
rect 13629 3498 13695 3501
rect 15929 3498 15995 3501
rect 13629 3496 15995 3498
rect 13629 3440 13634 3496
rect 13690 3440 15934 3496
rect 15990 3440 15995 3496
rect 13629 3438 15995 3440
rect 13629 3435 13695 3438
rect 15929 3435 15995 3438
rect 16113 3498 16179 3501
rect 17953 3498 18019 3501
rect 16113 3496 18019 3498
rect 16113 3440 16118 3496
rect 16174 3440 17958 3496
rect 18014 3440 18019 3496
rect 16113 3438 18019 3440
rect 16113 3435 16179 3438
rect 17953 3435 18019 3438
rect 14917 3362 14983 3365
rect 16757 3362 16823 3365
rect 14917 3360 16823 3362
rect 14917 3304 14922 3360
rect 14978 3304 16762 3360
rect 16818 3304 16823 3360
rect 14917 3302 16823 3304
rect 14917 3299 14983 3302
rect 16757 3299 16823 3302
rect 16941 3362 17007 3365
rect 19200 3362 20000 3392
rect 16941 3360 20000 3362
rect 16941 3304 16946 3360
rect 17002 3304 20000 3360
rect 16941 3302 20000 3304
rect 16941 3299 17007 3302
rect 5394 3296 5710 3297
rect 0 3226 800 3256
rect 5394 3232 5400 3296
rect 5464 3232 5480 3296
rect 5544 3232 5560 3296
rect 5624 3232 5640 3296
rect 5704 3232 5710 3296
rect 5394 3231 5710 3232
rect 9842 3296 10158 3297
rect 9842 3232 9848 3296
rect 9912 3232 9928 3296
rect 9992 3232 10008 3296
rect 10072 3232 10088 3296
rect 10152 3232 10158 3296
rect 9842 3231 10158 3232
rect 14290 3296 14606 3297
rect 14290 3232 14296 3296
rect 14360 3232 14376 3296
rect 14440 3232 14456 3296
rect 14520 3232 14536 3296
rect 14600 3232 14606 3296
rect 19200 3272 20000 3302
rect 14290 3231 14606 3232
rect 1485 3226 1551 3229
rect 0 3224 1551 3226
rect 0 3168 1490 3224
rect 1546 3168 1551 3224
rect 0 3166 1551 3168
rect 0 3136 800 3166
rect 1485 3163 1551 3166
rect 2313 3226 2379 3229
rect 3877 3226 3943 3229
rect 5206 3226 5212 3228
rect 2313 3224 5212 3226
rect 2313 3168 2318 3224
rect 2374 3168 3882 3224
rect 3938 3168 5212 3224
rect 2313 3166 5212 3168
rect 2313 3163 2379 3166
rect 3877 3163 3943 3166
rect 5206 3164 5212 3166
rect 5276 3164 5282 3228
rect 10358 3164 10364 3228
rect 10428 3226 10434 3228
rect 13169 3226 13235 3229
rect 13813 3228 13879 3229
rect 13997 3228 14063 3229
rect 13813 3226 13860 3228
rect 10428 3224 13235 3226
rect 10428 3168 13174 3224
rect 13230 3168 13235 3224
rect 10428 3166 13235 3168
rect 13768 3224 13860 3226
rect 13768 3168 13818 3224
rect 13768 3166 13860 3168
rect 10428 3164 10434 3166
rect 13169 3163 13235 3166
rect 13813 3164 13860 3166
rect 13924 3164 13930 3228
rect 13997 3224 14044 3228
rect 14108 3226 14114 3228
rect 16205 3226 16271 3229
rect 18229 3226 18295 3229
rect 13997 3168 14002 3224
rect 13997 3164 14044 3168
rect 14108 3166 14154 3226
rect 16205 3224 18295 3226
rect 16205 3168 16210 3224
rect 16266 3168 18234 3224
rect 18290 3168 18295 3224
rect 16205 3166 18295 3168
rect 14108 3164 14114 3166
rect 13813 3163 13879 3164
rect 13997 3163 14063 3164
rect 16205 3163 16271 3166
rect 18229 3163 18295 3166
rect 11145 3090 11211 3093
rect 17125 3090 17191 3093
rect 11145 3088 17191 3090
rect 11145 3032 11150 3088
rect 11206 3032 17130 3088
rect 17186 3032 17191 3088
rect 11145 3030 17191 3032
rect 11145 3027 11211 3030
rect 17125 3027 17191 3030
rect 18413 3090 18479 3093
rect 19200 3090 20000 3120
rect 18413 3088 20000 3090
rect 18413 3032 18418 3088
rect 18474 3032 20000 3088
rect 18413 3030 20000 3032
rect 18413 3027 18479 3030
rect 19200 3000 20000 3030
rect 0 2954 800 2984
rect 1853 2954 1919 2957
rect 0 2952 1919 2954
rect 0 2896 1858 2952
rect 1914 2896 1919 2952
rect 0 2894 1919 2896
rect 0 2864 800 2894
rect 1853 2891 1919 2894
rect 13077 2954 13143 2957
rect 15745 2954 15811 2957
rect 13077 2952 15811 2954
rect 13077 2896 13082 2952
rect 13138 2896 15750 2952
rect 15806 2896 15811 2952
rect 13077 2894 15811 2896
rect 13077 2891 13143 2894
rect 15745 2891 15811 2894
rect 16246 2892 16252 2956
rect 16316 2954 16322 2956
rect 16573 2954 16639 2957
rect 16316 2952 16639 2954
rect 16316 2896 16578 2952
rect 16634 2896 16639 2952
rect 16316 2894 16639 2896
rect 16316 2892 16322 2894
rect 13537 2818 13603 2821
rect 16254 2818 16314 2892
rect 16573 2891 16639 2894
rect 13537 2816 16314 2818
rect 13537 2760 13542 2816
rect 13598 2760 16314 2816
rect 13537 2758 16314 2760
rect 17677 2818 17743 2821
rect 19200 2818 20000 2848
rect 17677 2816 20000 2818
rect 17677 2760 17682 2816
rect 17738 2760 20000 2816
rect 17677 2758 20000 2760
rect 13537 2755 13603 2758
rect 17677 2755 17743 2758
rect 3170 2752 3486 2753
rect 0 2682 800 2712
rect 3170 2688 3176 2752
rect 3240 2688 3256 2752
rect 3320 2688 3336 2752
rect 3400 2688 3416 2752
rect 3480 2688 3486 2752
rect 3170 2687 3486 2688
rect 7618 2752 7934 2753
rect 7618 2688 7624 2752
rect 7688 2688 7704 2752
rect 7768 2688 7784 2752
rect 7848 2688 7864 2752
rect 7928 2688 7934 2752
rect 7618 2687 7934 2688
rect 12066 2752 12382 2753
rect 12066 2688 12072 2752
rect 12136 2688 12152 2752
rect 12216 2688 12232 2752
rect 12296 2688 12312 2752
rect 12376 2688 12382 2752
rect 12066 2687 12382 2688
rect 16514 2752 16830 2753
rect 16514 2688 16520 2752
rect 16584 2688 16600 2752
rect 16664 2688 16680 2752
rect 16744 2688 16760 2752
rect 16824 2688 16830 2752
rect 19200 2728 20000 2758
rect 16514 2687 16830 2688
rect 1485 2682 1551 2685
rect 13537 2684 13603 2685
rect 13486 2682 13492 2684
rect 0 2680 1551 2682
rect 0 2624 1490 2680
rect 1546 2624 1551 2680
rect 0 2622 1551 2624
rect 13446 2622 13492 2682
rect 13556 2680 13603 2684
rect 13598 2624 13603 2680
rect 0 2592 800 2622
rect 1485 2619 1551 2622
rect 13486 2620 13492 2622
rect 13556 2620 13603 2624
rect 15878 2620 15884 2684
rect 15948 2682 15954 2684
rect 16297 2682 16363 2685
rect 15948 2680 16363 2682
rect 15948 2624 16302 2680
rect 16358 2624 16363 2680
rect 15948 2622 16363 2624
rect 15948 2620 15954 2622
rect 13537 2619 13603 2620
rect 16297 2619 16363 2622
rect 13721 2548 13787 2549
rect 13670 2484 13676 2548
rect 13740 2546 13787 2548
rect 13905 2546 13971 2549
rect 14958 2546 14964 2548
rect 13740 2544 13832 2546
rect 13782 2488 13832 2544
rect 13740 2486 13832 2488
rect 13905 2544 14964 2546
rect 13905 2488 13910 2544
rect 13966 2488 14964 2544
rect 13905 2486 14964 2488
rect 13740 2484 13787 2486
rect 13721 2483 13787 2484
rect 13905 2483 13971 2486
rect 14958 2484 14964 2486
rect 15028 2546 15034 2548
rect 17033 2546 17099 2549
rect 15028 2544 17099 2546
rect 15028 2488 17038 2544
rect 17094 2488 17099 2544
rect 15028 2486 17099 2488
rect 15028 2484 15034 2486
rect 17033 2483 17099 2486
rect 17309 2546 17375 2549
rect 19200 2546 20000 2576
rect 17309 2544 20000 2546
rect 17309 2488 17314 2544
rect 17370 2488 20000 2544
rect 17309 2486 20000 2488
rect 17309 2483 17375 2486
rect 19200 2456 20000 2486
rect 0 2410 800 2440
rect 1853 2410 1919 2413
rect 0 2408 1919 2410
rect 0 2352 1858 2408
rect 1914 2352 1919 2408
rect 0 2350 1919 2352
rect 0 2320 800 2350
rect 1853 2347 1919 2350
rect 3601 2410 3667 2413
rect 11646 2410 11652 2412
rect 3601 2408 11652 2410
rect 3601 2352 3606 2408
rect 3662 2352 11652 2408
rect 3601 2350 11652 2352
rect 3601 2347 3667 2350
rect 11646 2348 11652 2350
rect 11716 2348 11722 2412
rect 14641 2410 14707 2413
rect 17953 2410 18019 2413
rect 14641 2408 18019 2410
rect 14641 2352 14646 2408
rect 14702 2352 17958 2408
rect 18014 2352 18019 2408
rect 14641 2350 18019 2352
rect 14641 2347 14707 2350
rect 17953 2347 18019 2350
rect 5394 2208 5710 2209
rect 0 2138 800 2168
rect 5394 2144 5400 2208
rect 5464 2144 5480 2208
rect 5544 2144 5560 2208
rect 5624 2144 5640 2208
rect 5704 2144 5710 2208
rect 5394 2143 5710 2144
rect 9842 2208 10158 2209
rect 9842 2144 9848 2208
rect 9912 2144 9928 2208
rect 9992 2144 10008 2208
rect 10072 2144 10088 2208
rect 10152 2144 10158 2208
rect 9842 2143 10158 2144
rect 14290 2208 14606 2209
rect 14290 2144 14296 2208
rect 14360 2144 14376 2208
rect 14440 2144 14456 2208
rect 14520 2144 14536 2208
rect 14600 2144 14606 2208
rect 14290 2143 14606 2144
rect 2589 2138 2655 2141
rect 0 2136 2655 2138
rect 0 2080 2594 2136
rect 2650 2080 2655 2136
rect 0 2078 2655 2080
rect 0 2048 800 2078
rect 2589 2075 2655 2078
rect 8109 2002 8175 2005
rect 13997 2002 14063 2005
rect 8109 2000 14063 2002
rect 8109 1944 8114 2000
rect 8170 1944 14002 2000
rect 14058 1944 14063 2000
rect 8109 1942 14063 1944
rect 8109 1939 8175 1942
rect 13997 1939 14063 1942
rect 0 1866 800 1896
rect 2221 1866 2287 1869
rect 0 1864 2287 1866
rect 0 1808 2226 1864
rect 2282 1808 2287 1864
rect 0 1806 2287 1808
rect 0 1776 800 1806
rect 2221 1803 2287 1806
rect 0 1594 800 1624
rect 2773 1594 2839 1597
rect 0 1592 2839 1594
rect 0 1536 2778 1592
rect 2834 1536 2839 1592
rect 0 1534 2839 1536
rect 0 1504 800 1534
rect 2773 1531 2839 1534
<< via3 >>
rect 13676 14996 13740 15060
rect 3176 14716 3240 14720
rect 3176 14660 3180 14716
rect 3180 14660 3236 14716
rect 3236 14660 3240 14716
rect 3176 14656 3240 14660
rect 3256 14716 3320 14720
rect 3256 14660 3260 14716
rect 3260 14660 3316 14716
rect 3316 14660 3320 14716
rect 3256 14656 3320 14660
rect 3336 14716 3400 14720
rect 3336 14660 3340 14716
rect 3340 14660 3396 14716
rect 3396 14660 3400 14716
rect 3336 14656 3400 14660
rect 3416 14716 3480 14720
rect 3416 14660 3420 14716
rect 3420 14660 3476 14716
rect 3476 14660 3480 14716
rect 3416 14656 3480 14660
rect 7624 14716 7688 14720
rect 7624 14660 7628 14716
rect 7628 14660 7684 14716
rect 7684 14660 7688 14716
rect 7624 14656 7688 14660
rect 7704 14716 7768 14720
rect 7704 14660 7708 14716
rect 7708 14660 7764 14716
rect 7764 14660 7768 14716
rect 7704 14656 7768 14660
rect 7784 14716 7848 14720
rect 7784 14660 7788 14716
rect 7788 14660 7844 14716
rect 7844 14660 7848 14716
rect 7784 14656 7848 14660
rect 7864 14716 7928 14720
rect 7864 14660 7868 14716
rect 7868 14660 7924 14716
rect 7924 14660 7928 14716
rect 7864 14656 7928 14660
rect 12072 14716 12136 14720
rect 12072 14660 12076 14716
rect 12076 14660 12132 14716
rect 12132 14660 12136 14716
rect 12072 14656 12136 14660
rect 12152 14716 12216 14720
rect 12152 14660 12156 14716
rect 12156 14660 12212 14716
rect 12212 14660 12216 14716
rect 12152 14656 12216 14660
rect 12232 14716 12296 14720
rect 12232 14660 12236 14716
rect 12236 14660 12292 14716
rect 12292 14660 12296 14716
rect 12232 14656 12296 14660
rect 12312 14716 12376 14720
rect 12312 14660 12316 14716
rect 12316 14660 12372 14716
rect 12372 14660 12376 14716
rect 12312 14656 12376 14660
rect 16520 14716 16584 14720
rect 16520 14660 16524 14716
rect 16524 14660 16580 14716
rect 16580 14660 16584 14716
rect 16520 14656 16584 14660
rect 16600 14716 16664 14720
rect 16600 14660 16604 14716
rect 16604 14660 16660 14716
rect 16660 14660 16664 14716
rect 16600 14656 16664 14660
rect 16680 14716 16744 14720
rect 16680 14660 16684 14716
rect 16684 14660 16740 14716
rect 16740 14660 16744 14716
rect 16680 14656 16744 14660
rect 16760 14716 16824 14720
rect 16760 14660 16764 14716
rect 16764 14660 16820 14716
rect 16820 14660 16824 14716
rect 16760 14656 16824 14660
rect 5400 14172 5464 14176
rect 5400 14116 5404 14172
rect 5404 14116 5460 14172
rect 5460 14116 5464 14172
rect 5400 14112 5464 14116
rect 5480 14172 5544 14176
rect 5480 14116 5484 14172
rect 5484 14116 5540 14172
rect 5540 14116 5544 14172
rect 5480 14112 5544 14116
rect 5560 14172 5624 14176
rect 5560 14116 5564 14172
rect 5564 14116 5620 14172
rect 5620 14116 5624 14172
rect 5560 14112 5624 14116
rect 5640 14172 5704 14176
rect 5640 14116 5644 14172
rect 5644 14116 5700 14172
rect 5700 14116 5704 14172
rect 5640 14112 5704 14116
rect 3004 14044 3068 14108
rect 9076 13908 9140 13972
rect 9848 14172 9912 14176
rect 9848 14116 9852 14172
rect 9852 14116 9908 14172
rect 9908 14116 9912 14172
rect 9848 14112 9912 14116
rect 9928 14172 9992 14176
rect 9928 14116 9932 14172
rect 9932 14116 9988 14172
rect 9988 14116 9992 14172
rect 9928 14112 9992 14116
rect 10008 14172 10072 14176
rect 10008 14116 10012 14172
rect 10012 14116 10068 14172
rect 10068 14116 10072 14172
rect 10008 14112 10072 14116
rect 10088 14172 10152 14176
rect 10088 14116 10092 14172
rect 10092 14116 10148 14172
rect 10148 14116 10152 14172
rect 10088 14112 10152 14116
rect 14296 14172 14360 14176
rect 14296 14116 14300 14172
rect 14300 14116 14356 14172
rect 14356 14116 14360 14172
rect 14296 14112 14360 14116
rect 14376 14172 14440 14176
rect 14376 14116 14380 14172
rect 14380 14116 14436 14172
rect 14436 14116 14440 14172
rect 14376 14112 14440 14116
rect 14456 14172 14520 14176
rect 14456 14116 14460 14172
rect 14460 14116 14516 14172
rect 14516 14116 14520 14172
rect 14456 14112 14520 14116
rect 14536 14172 14600 14176
rect 14536 14116 14540 14172
rect 14540 14116 14596 14172
rect 14596 14116 14600 14172
rect 14536 14112 14600 14116
rect 10364 13908 10428 13972
rect 13860 13772 13924 13836
rect 3176 13628 3240 13632
rect 3176 13572 3180 13628
rect 3180 13572 3236 13628
rect 3236 13572 3240 13628
rect 3176 13568 3240 13572
rect 3256 13628 3320 13632
rect 3256 13572 3260 13628
rect 3260 13572 3316 13628
rect 3316 13572 3320 13628
rect 3256 13568 3320 13572
rect 3336 13628 3400 13632
rect 3336 13572 3340 13628
rect 3340 13572 3396 13628
rect 3396 13572 3400 13628
rect 3336 13568 3400 13572
rect 3416 13628 3480 13632
rect 3416 13572 3420 13628
rect 3420 13572 3476 13628
rect 3476 13572 3480 13628
rect 3416 13568 3480 13572
rect 7624 13628 7688 13632
rect 7624 13572 7628 13628
rect 7628 13572 7684 13628
rect 7684 13572 7688 13628
rect 7624 13568 7688 13572
rect 7704 13628 7768 13632
rect 7704 13572 7708 13628
rect 7708 13572 7764 13628
rect 7764 13572 7768 13628
rect 7704 13568 7768 13572
rect 7784 13628 7848 13632
rect 7784 13572 7788 13628
rect 7788 13572 7844 13628
rect 7844 13572 7848 13628
rect 7784 13568 7848 13572
rect 7864 13628 7928 13632
rect 7864 13572 7868 13628
rect 7868 13572 7924 13628
rect 7924 13572 7928 13628
rect 7864 13568 7928 13572
rect 12072 13628 12136 13632
rect 12072 13572 12076 13628
rect 12076 13572 12132 13628
rect 12132 13572 12136 13628
rect 12072 13568 12136 13572
rect 12152 13628 12216 13632
rect 12152 13572 12156 13628
rect 12156 13572 12212 13628
rect 12212 13572 12216 13628
rect 12152 13568 12216 13572
rect 12232 13628 12296 13632
rect 12232 13572 12236 13628
rect 12236 13572 12292 13628
rect 12292 13572 12296 13628
rect 12232 13568 12296 13572
rect 12312 13628 12376 13632
rect 12312 13572 12316 13628
rect 12316 13572 12372 13628
rect 12372 13572 12376 13628
rect 12312 13568 12376 13572
rect 16520 13628 16584 13632
rect 16520 13572 16524 13628
rect 16524 13572 16580 13628
rect 16580 13572 16584 13628
rect 16520 13568 16584 13572
rect 16600 13628 16664 13632
rect 16600 13572 16604 13628
rect 16604 13572 16660 13628
rect 16660 13572 16664 13628
rect 16600 13568 16664 13572
rect 16680 13628 16744 13632
rect 16680 13572 16684 13628
rect 16684 13572 16740 13628
rect 16740 13572 16744 13628
rect 16680 13568 16744 13572
rect 16760 13628 16824 13632
rect 16760 13572 16764 13628
rect 16764 13572 16820 13628
rect 16820 13572 16824 13628
rect 16760 13568 16824 13572
rect 11836 13364 11900 13428
rect 5400 13084 5464 13088
rect 5400 13028 5404 13084
rect 5404 13028 5460 13084
rect 5460 13028 5464 13084
rect 5400 13024 5464 13028
rect 5480 13084 5544 13088
rect 5480 13028 5484 13084
rect 5484 13028 5540 13084
rect 5540 13028 5544 13084
rect 5480 13024 5544 13028
rect 5560 13084 5624 13088
rect 5560 13028 5564 13084
rect 5564 13028 5620 13084
rect 5620 13028 5624 13084
rect 5560 13024 5624 13028
rect 5640 13084 5704 13088
rect 5640 13028 5644 13084
rect 5644 13028 5700 13084
rect 5700 13028 5704 13084
rect 5640 13024 5704 13028
rect 9848 13084 9912 13088
rect 9848 13028 9852 13084
rect 9852 13028 9908 13084
rect 9908 13028 9912 13084
rect 9848 13024 9912 13028
rect 9928 13084 9992 13088
rect 9928 13028 9932 13084
rect 9932 13028 9988 13084
rect 9988 13028 9992 13084
rect 9928 13024 9992 13028
rect 10008 13084 10072 13088
rect 10008 13028 10012 13084
rect 10012 13028 10068 13084
rect 10068 13028 10072 13084
rect 10008 13024 10072 13028
rect 10088 13084 10152 13088
rect 10088 13028 10092 13084
rect 10092 13028 10148 13084
rect 10148 13028 10152 13084
rect 10088 13024 10152 13028
rect 14296 13084 14360 13088
rect 14296 13028 14300 13084
rect 14300 13028 14356 13084
rect 14356 13028 14360 13084
rect 14296 13024 14360 13028
rect 14376 13084 14440 13088
rect 14376 13028 14380 13084
rect 14380 13028 14436 13084
rect 14436 13028 14440 13084
rect 14376 13024 14440 13028
rect 14456 13084 14520 13088
rect 14456 13028 14460 13084
rect 14460 13028 14516 13084
rect 14516 13028 14520 13084
rect 14456 13024 14520 13028
rect 14536 13084 14600 13088
rect 14536 13028 14540 13084
rect 14540 13028 14596 13084
rect 14596 13028 14600 13084
rect 14536 13024 14600 13028
rect 7420 12684 7484 12748
rect 9260 12684 9324 12748
rect 3176 12540 3240 12544
rect 3176 12484 3180 12540
rect 3180 12484 3236 12540
rect 3236 12484 3240 12540
rect 3176 12480 3240 12484
rect 3256 12540 3320 12544
rect 3256 12484 3260 12540
rect 3260 12484 3316 12540
rect 3316 12484 3320 12540
rect 3256 12480 3320 12484
rect 3336 12540 3400 12544
rect 3336 12484 3340 12540
rect 3340 12484 3396 12540
rect 3396 12484 3400 12540
rect 3336 12480 3400 12484
rect 3416 12540 3480 12544
rect 3416 12484 3420 12540
rect 3420 12484 3476 12540
rect 3476 12484 3480 12540
rect 3416 12480 3480 12484
rect 7624 12540 7688 12544
rect 7624 12484 7628 12540
rect 7628 12484 7684 12540
rect 7684 12484 7688 12540
rect 7624 12480 7688 12484
rect 7704 12540 7768 12544
rect 7704 12484 7708 12540
rect 7708 12484 7764 12540
rect 7764 12484 7768 12540
rect 7704 12480 7768 12484
rect 7784 12540 7848 12544
rect 7784 12484 7788 12540
rect 7788 12484 7844 12540
rect 7844 12484 7848 12540
rect 7784 12480 7848 12484
rect 7864 12540 7928 12544
rect 7864 12484 7868 12540
rect 7868 12484 7924 12540
rect 7924 12484 7928 12540
rect 7864 12480 7928 12484
rect 12072 12540 12136 12544
rect 12072 12484 12076 12540
rect 12076 12484 12132 12540
rect 12132 12484 12136 12540
rect 12072 12480 12136 12484
rect 12152 12540 12216 12544
rect 12152 12484 12156 12540
rect 12156 12484 12212 12540
rect 12212 12484 12216 12540
rect 12152 12480 12216 12484
rect 12232 12540 12296 12544
rect 12232 12484 12236 12540
rect 12236 12484 12292 12540
rect 12292 12484 12296 12540
rect 12232 12480 12296 12484
rect 12312 12540 12376 12544
rect 12312 12484 12316 12540
rect 12316 12484 12372 12540
rect 12372 12484 12376 12540
rect 12312 12480 12376 12484
rect 16520 12540 16584 12544
rect 16520 12484 16524 12540
rect 16524 12484 16580 12540
rect 16580 12484 16584 12540
rect 16520 12480 16584 12484
rect 16600 12540 16664 12544
rect 16600 12484 16604 12540
rect 16604 12484 16660 12540
rect 16660 12484 16664 12540
rect 16600 12480 16664 12484
rect 16680 12540 16744 12544
rect 16680 12484 16684 12540
rect 16684 12484 16740 12540
rect 16740 12484 16744 12540
rect 16680 12480 16744 12484
rect 16760 12540 16824 12544
rect 16760 12484 16764 12540
rect 16764 12484 16820 12540
rect 16820 12484 16824 12540
rect 16760 12480 16824 12484
rect 4292 12140 4356 12204
rect 12940 12004 13004 12068
rect 5400 11996 5464 12000
rect 5400 11940 5404 11996
rect 5404 11940 5460 11996
rect 5460 11940 5464 11996
rect 5400 11936 5464 11940
rect 5480 11996 5544 12000
rect 5480 11940 5484 11996
rect 5484 11940 5540 11996
rect 5540 11940 5544 11996
rect 5480 11936 5544 11940
rect 5560 11996 5624 12000
rect 5560 11940 5564 11996
rect 5564 11940 5620 11996
rect 5620 11940 5624 11996
rect 5560 11936 5624 11940
rect 5640 11996 5704 12000
rect 5640 11940 5644 11996
rect 5644 11940 5700 11996
rect 5700 11940 5704 11996
rect 5640 11936 5704 11940
rect 9848 11996 9912 12000
rect 9848 11940 9852 11996
rect 9852 11940 9908 11996
rect 9908 11940 9912 11996
rect 9848 11936 9912 11940
rect 9928 11996 9992 12000
rect 9928 11940 9932 11996
rect 9932 11940 9988 11996
rect 9988 11940 9992 11996
rect 9928 11936 9992 11940
rect 10008 11996 10072 12000
rect 10008 11940 10012 11996
rect 10012 11940 10068 11996
rect 10068 11940 10072 11996
rect 10008 11936 10072 11940
rect 10088 11996 10152 12000
rect 10088 11940 10092 11996
rect 10092 11940 10148 11996
rect 10148 11940 10152 11996
rect 10088 11936 10152 11940
rect 14296 11996 14360 12000
rect 14296 11940 14300 11996
rect 14300 11940 14356 11996
rect 14356 11940 14360 11996
rect 14296 11936 14360 11940
rect 14376 11996 14440 12000
rect 14376 11940 14380 11996
rect 14380 11940 14436 11996
rect 14436 11940 14440 11996
rect 14376 11936 14440 11940
rect 14456 11996 14520 12000
rect 14456 11940 14460 11996
rect 14460 11940 14516 11996
rect 14516 11940 14520 11996
rect 14456 11936 14520 11940
rect 14536 11996 14600 12000
rect 14536 11940 14540 11996
rect 14540 11940 14596 11996
rect 14596 11940 14600 11996
rect 14536 11936 14600 11940
rect 11284 11928 11348 11932
rect 11284 11872 11298 11928
rect 11298 11872 11348 11928
rect 11284 11868 11348 11872
rect 5212 11732 5276 11796
rect 13492 11868 13556 11932
rect 11652 11520 11716 11524
rect 11652 11464 11666 11520
rect 11666 11464 11716 11520
rect 11652 11460 11716 11464
rect 3176 11452 3240 11456
rect 3176 11396 3180 11452
rect 3180 11396 3236 11452
rect 3236 11396 3240 11452
rect 3176 11392 3240 11396
rect 3256 11452 3320 11456
rect 3256 11396 3260 11452
rect 3260 11396 3316 11452
rect 3316 11396 3320 11452
rect 3256 11392 3320 11396
rect 3336 11452 3400 11456
rect 3336 11396 3340 11452
rect 3340 11396 3396 11452
rect 3396 11396 3400 11452
rect 3336 11392 3400 11396
rect 3416 11452 3480 11456
rect 3416 11396 3420 11452
rect 3420 11396 3476 11452
rect 3476 11396 3480 11452
rect 3416 11392 3480 11396
rect 7624 11452 7688 11456
rect 7624 11396 7628 11452
rect 7628 11396 7684 11452
rect 7684 11396 7688 11452
rect 7624 11392 7688 11396
rect 7704 11452 7768 11456
rect 7704 11396 7708 11452
rect 7708 11396 7764 11452
rect 7764 11396 7768 11452
rect 7704 11392 7768 11396
rect 7784 11452 7848 11456
rect 7784 11396 7788 11452
rect 7788 11396 7844 11452
rect 7844 11396 7848 11452
rect 7784 11392 7848 11396
rect 7864 11452 7928 11456
rect 7864 11396 7868 11452
rect 7868 11396 7924 11452
rect 7924 11396 7928 11452
rect 7864 11392 7928 11396
rect 12072 11452 12136 11456
rect 12072 11396 12076 11452
rect 12076 11396 12132 11452
rect 12132 11396 12136 11452
rect 12072 11392 12136 11396
rect 12152 11452 12216 11456
rect 12152 11396 12156 11452
rect 12156 11396 12212 11452
rect 12212 11396 12216 11452
rect 12152 11392 12216 11396
rect 12232 11452 12296 11456
rect 12232 11396 12236 11452
rect 12236 11396 12292 11452
rect 12292 11396 12296 11452
rect 12232 11392 12296 11396
rect 12312 11452 12376 11456
rect 12312 11396 12316 11452
rect 12316 11396 12372 11452
rect 12372 11396 12376 11452
rect 12312 11392 12376 11396
rect 16520 11452 16584 11456
rect 16520 11396 16524 11452
rect 16524 11396 16580 11452
rect 16580 11396 16584 11452
rect 16520 11392 16584 11396
rect 16600 11452 16664 11456
rect 16600 11396 16604 11452
rect 16604 11396 16660 11452
rect 16660 11396 16664 11452
rect 16600 11392 16664 11396
rect 16680 11452 16744 11456
rect 16680 11396 16684 11452
rect 16684 11396 16740 11452
rect 16740 11396 16744 11452
rect 16680 11392 16744 11396
rect 16760 11452 16824 11456
rect 16760 11396 16764 11452
rect 16764 11396 16820 11452
rect 16820 11396 16824 11452
rect 16760 11392 16824 11396
rect 14044 11188 14108 11252
rect 16252 11188 16316 11252
rect 10732 11052 10796 11116
rect 17908 11052 17972 11116
rect 5400 10908 5464 10912
rect 5400 10852 5404 10908
rect 5404 10852 5460 10908
rect 5460 10852 5464 10908
rect 5400 10848 5464 10852
rect 5480 10908 5544 10912
rect 5480 10852 5484 10908
rect 5484 10852 5540 10908
rect 5540 10852 5544 10908
rect 5480 10848 5544 10852
rect 5560 10908 5624 10912
rect 5560 10852 5564 10908
rect 5564 10852 5620 10908
rect 5620 10852 5624 10908
rect 5560 10848 5624 10852
rect 5640 10908 5704 10912
rect 5640 10852 5644 10908
rect 5644 10852 5700 10908
rect 5700 10852 5704 10908
rect 5640 10848 5704 10852
rect 9848 10908 9912 10912
rect 9848 10852 9852 10908
rect 9852 10852 9908 10908
rect 9908 10852 9912 10908
rect 9848 10848 9912 10852
rect 9928 10908 9992 10912
rect 9928 10852 9932 10908
rect 9932 10852 9988 10908
rect 9988 10852 9992 10908
rect 9928 10848 9992 10852
rect 10008 10908 10072 10912
rect 10008 10852 10012 10908
rect 10012 10852 10068 10908
rect 10068 10852 10072 10908
rect 10008 10848 10072 10852
rect 10088 10908 10152 10912
rect 10088 10852 10092 10908
rect 10092 10852 10148 10908
rect 10148 10852 10152 10908
rect 10088 10848 10152 10852
rect 14296 10908 14360 10912
rect 14296 10852 14300 10908
rect 14300 10852 14356 10908
rect 14356 10852 14360 10908
rect 14296 10848 14360 10852
rect 14376 10908 14440 10912
rect 14376 10852 14380 10908
rect 14380 10852 14436 10908
rect 14436 10852 14440 10908
rect 14376 10848 14440 10852
rect 14456 10908 14520 10912
rect 14456 10852 14460 10908
rect 14460 10852 14516 10908
rect 14516 10852 14520 10908
rect 14456 10848 14520 10852
rect 14536 10908 14600 10912
rect 14536 10852 14540 10908
rect 14540 10852 14596 10908
rect 14596 10852 14600 10908
rect 14536 10848 14600 10852
rect 10548 10780 10612 10844
rect 3740 10644 3804 10708
rect 5028 10432 5092 10436
rect 5028 10376 5042 10432
rect 5042 10376 5092 10432
rect 5028 10372 5092 10376
rect 3176 10364 3240 10368
rect 3176 10308 3180 10364
rect 3180 10308 3236 10364
rect 3236 10308 3240 10364
rect 3176 10304 3240 10308
rect 3256 10364 3320 10368
rect 3256 10308 3260 10364
rect 3260 10308 3316 10364
rect 3316 10308 3320 10364
rect 3256 10304 3320 10308
rect 3336 10364 3400 10368
rect 3336 10308 3340 10364
rect 3340 10308 3396 10364
rect 3396 10308 3400 10364
rect 3336 10304 3400 10308
rect 3416 10364 3480 10368
rect 3416 10308 3420 10364
rect 3420 10308 3476 10364
rect 3476 10308 3480 10364
rect 3416 10304 3480 10308
rect 7624 10364 7688 10368
rect 7624 10308 7628 10364
rect 7628 10308 7684 10364
rect 7684 10308 7688 10364
rect 7624 10304 7688 10308
rect 7704 10364 7768 10368
rect 7704 10308 7708 10364
rect 7708 10308 7764 10364
rect 7764 10308 7768 10364
rect 7704 10304 7768 10308
rect 7784 10364 7848 10368
rect 7784 10308 7788 10364
rect 7788 10308 7844 10364
rect 7844 10308 7848 10364
rect 7784 10304 7848 10308
rect 7864 10364 7928 10368
rect 7864 10308 7868 10364
rect 7868 10308 7924 10364
rect 7924 10308 7928 10364
rect 7864 10304 7928 10308
rect 12072 10364 12136 10368
rect 12072 10308 12076 10364
rect 12076 10308 12132 10364
rect 12132 10308 12136 10364
rect 12072 10304 12136 10308
rect 12152 10364 12216 10368
rect 12152 10308 12156 10364
rect 12156 10308 12212 10364
rect 12212 10308 12216 10364
rect 12152 10304 12216 10308
rect 12232 10364 12296 10368
rect 12232 10308 12236 10364
rect 12236 10308 12292 10364
rect 12292 10308 12296 10364
rect 12232 10304 12296 10308
rect 12312 10364 12376 10368
rect 12312 10308 12316 10364
rect 12316 10308 12372 10364
rect 12372 10308 12376 10364
rect 12312 10304 12376 10308
rect 16520 10364 16584 10368
rect 16520 10308 16524 10364
rect 16524 10308 16580 10364
rect 16580 10308 16584 10364
rect 16520 10304 16584 10308
rect 16600 10364 16664 10368
rect 16600 10308 16604 10364
rect 16604 10308 16660 10364
rect 16660 10308 16664 10364
rect 16600 10304 16664 10308
rect 16680 10364 16744 10368
rect 16680 10308 16684 10364
rect 16684 10308 16740 10364
rect 16740 10308 16744 10364
rect 16680 10304 16744 10308
rect 16760 10364 16824 10368
rect 16760 10308 16764 10364
rect 16764 10308 16820 10364
rect 16820 10308 16824 10364
rect 16760 10304 16824 10308
rect 14964 10236 15028 10300
rect 16988 10100 17052 10164
rect 5400 9820 5464 9824
rect 5400 9764 5404 9820
rect 5404 9764 5460 9820
rect 5460 9764 5464 9820
rect 5400 9760 5464 9764
rect 5480 9820 5544 9824
rect 5480 9764 5484 9820
rect 5484 9764 5540 9820
rect 5540 9764 5544 9820
rect 5480 9760 5544 9764
rect 5560 9820 5624 9824
rect 5560 9764 5564 9820
rect 5564 9764 5620 9820
rect 5620 9764 5624 9820
rect 5560 9760 5624 9764
rect 5640 9820 5704 9824
rect 5640 9764 5644 9820
rect 5644 9764 5700 9820
rect 5700 9764 5704 9820
rect 5640 9760 5704 9764
rect 9848 9820 9912 9824
rect 9848 9764 9852 9820
rect 9852 9764 9908 9820
rect 9908 9764 9912 9820
rect 9848 9760 9912 9764
rect 9928 9820 9992 9824
rect 9928 9764 9932 9820
rect 9932 9764 9988 9820
rect 9988 9764 9992 9820
rect 9928 9760 9992 9764
rect 10008 9820 10072 9824
rect 10008 9764 10012 9820
rect 10012 9764 10068 9820
rect 10068 9764 10072 9820
rect 10008 9760 10072 9764
rect 10088 9820 10152 9824
rect 10088 9764 10092 9820
rect 10092 9764 10148 9820
rect 10148 9764 10152 9820
rect 10088 9760 10152 9764
rect 14296 9820 14360 9824
rect 14296 9764 14300 9820
rect 14300 9764 14356 9820
rect 14356 9764 14360 9820
rect 14296 9760 14360 9764
rect 14376 9820 14440 9824
rect 14376 9764 14380 9820
rect 14380 9764 14436 9820
rect 14436 9764 14440 9820
rect 14376 9760 14440 9764
rect 14456 9820 14520 9824
rect 14456 9764 14460 9820
rect 14460 9764 14516 9820
rect 14516 9764 14520 9820
rect 14456 9760 14520 9764
rect 14536 9820 14600 9824
rect 14536 9764 14540 9820
rect 14540 9764 14596 9820
rect 14596 9764 14600 9820
rect 14536 9760 14600 9764
rect 7420 9692 7484 9756
rect 10548 9692 10612 9756
rect 17908 9480 17972 9484
rect 17908 9424 17922 9480
rect 17922 9424 17972 9480
rect 17908 9420 17972 9424
rect 2084 9284 2148 9348
rect 3176 9276 3240 9280
rect 3176 9220 3180 9276
rect 3180 9220 3236 9276
rect 3236 9220 3240 9276
rect 3176 9216 3240 9220
rect 3256 9276 3320 9280
rect 3256 9220 3260 9276
rect 3260 9220 3316 9276
rect 3316 9220 3320 9276
rect 3256 9216 3320 9220
rect 3336 9276 3400 9280
rect 3336 9220 3340 9276
rect 3340 9220 3396 9276
rect 3396 9220 3400 9276
rect 3336 9216 3400 9220
rect 3416 9276 3480 9280
rect 3416 9220 3420 9276
rect 3420 9220 3476 9276
rect 3476 9220 3480 9276
rect 3416 9216 3480 9220
rect 7624 9276 7688 9280
rect 7624 9220 7628 9276
rect 7628 9220 7684 9276
rect 7684 9220 7688 9276
rect 7624 9216 7688 9220
rect 7704 9276 7768 9280
rect 7704 9220 7708 9276
rect 7708 9220 7764 9276
rect 7764 9220 7768 9276
rect 7704 9216 7768 9220
rect 7784 9276 7848 9280
rect 7784 9220 7788 9276
rect 7788 9220 7844 9276
rect 7844 9220 7848 9276
rect 7784 9216 7848 9220
rect 7864 9276 7928 9280
rect 7864 9220 7868 9276
rect 7868 9220 7924 9276
rect 7924 9220 7928 9276
rect 7864 9216 7928 9220
rect 12072 9276 12136 9280
rect 12072 9220 12076 9276
rect 12076 9220 12132 9276
rect 12132 9220 12136 9276
rect 12072 9216 12136 9220
rect 12152 9276 12216 9280
rect 12152 9220 12156 9276
rect 12156 9220 12212 9276
rect 12212 9220 12216 9276
rect 12152 9216 12216 9220
rect 12232 9276 12296 9280
rect 12232 9220 12236 9276
rect 12236 9220 12292 9276
rect 12292 9220 12296 9276
rect 12232 9216 12296 9220
rect 12312 9276 12376 9280
rect 12312 9220 12316 9276
rect 12316 9220 12372 9276
rect 12372 9220 12376 9276
rect 12312 9216 12376 9220
rect 16520 9276 16584 9280
rect 16520 9220 16524 9276
rect 16524 9220 16580 9276
rect 16580 9220 16584 9276
rect 16520 9216 16584 9220
rect 16600 9276 16664 9280
rect 16600 9220 16604 9276
rect 16604 9220 16660 9276
rect 16660 9220 16664 9276
rect 16600 9216 16664 9220
rect 16680 9276 16744 9280
rect 16680 9220 16684 9276
rect 16684 9220 16740 9276
rect 16740 9220 16744 9276
rect 16680 9216 16744 9220
rect 16760 9276 16824 9280
rect 16760 9220 16764 9276
rect 16764 9220 16820 9276
rect 16820 9220 16824 9276
rect 16760 9216 16824 9220
rect 4844 9148 4908 9212
rect 6500 9072 6564 9076
rect 6500 9016 6514 9072
rect 6514 9016 6564 9072
rect 6500 9012 6564 9016
rect 7052 8740 7116 8804
rect 5400 8732 5464 8736
rect 5400 8676 5404 8732
rect 5404 8676 5460 8732
rect 5460 8676 5464 8732
rect 5400 8672 5464 8676
rect 5480 8732 5544 8736
rect 5480 8676 5484 8732
rect 5484 8676 5540 8732
rect 5540 8676 5544 8732
rect 5480 8672 5544 8676
rect 5560 8732 5624 8736
rect 5560 8676 5564 8732
rect 5564 8676 5620 8732
rect 5620 8676 5624 8732
rect 5560 8672 5624 8676
rect 5640 8732 5704 8736
rect 5640 8676 5644 8732
rect 5644 8676 5700 8732
rect 5700 8676 5704 8732
rect 5640 8672 5704 8676
rect 9848 8732 9912 8736
rect 9848 8676 9852 8732
rect 9852 8676 9908 8732
rect 9908 8676 9912 8732
rect 9848 8672 9912 8676
rect 9928 8732 9992 8736
rect 9928 8676 9932 8732
rect 9932 8676 9988 8732
rect 9988 8676 9992 8732
rect 9928 8672 9992 8676
rect 10008 8732 10072 8736
rect 10008 8676 10012 8732
rect 10012 8676 10068 8732
rect 10068 8676 10072 8732
rect 10008 8672 10072 8676
rect 10088 8732 10152 8736
rect 10088 8676 10092 8732
rect 10092 8676 10148 8732
rect 10148 8676 10152 8732
rect 10088 8672 10152 8676
rect 14296 8732 14360 8736
rect 14296 8676 14300 8732
rect 14300 8676 14356 8732
rect 14356 8676 14360 8732
rect 14296 8672 14360 8676
rect 14376 8732 14440 8736
rect 14376 8676 14380 8732
rect 14380 8676 14436 8732
rect 14436 8676 14440 8732
rect 14376 8672 14440 8676
rect 14456 8732 14520 8736
rect 14456 8676 14460 8732
rect 14460 8676 14516 8732
rect 14516 8676 14520 8732
rect 14456 8672 14520 8676
rect 14536 8732 14600 8736
rect 14536 8676 14540 8732
rect 14540 8676 14596 8732
rect 14596 8676 14600 8732
rect 14536 8672 14600 8676
rect 2268 8468 2332 8532
rect 6868 8332 6932 8396
rect 8156 8392 8220 8396
rect 8156 8336 8170 8392
rect 8170 8336 8220 8392
rect 8156 8332 8220 8336
rect 10548 8196 10612 8260
rect 3176 8188 3240 8192
rect 3176 8132 3180 8188
rect 3180 8132 3236 8188
rect 3236 8132 3240 8188
rect 3176 8128 3240 8132
rect 3256 8188 3320 8192
rect 3256 8132 3260 8188
rect 3260 8132 3316 8188
rect 3316 8132 3320 8188
rect 3256 8128 3320 8132
rect 3336 8188 3400 8192
rect 3336 8132 3340 8188
rect 3340 8132 3396 8188
rect 3396 8132 3400 8188
rect 3336 8128 3400 8132
rect 3416 8188 3480 8192
rect 3416 8132 3420 8188
rect 3420 8132 3476 8188
rect 3476 8132 3480 8188
rect 3416 8128 3480 8132
rect 7624 8188 7688 8192
rect 7624 8132 7628 8188
rect 7628 8132 7684 8188
rect 7684 8132 7688 8188
rect 7624 8128 7688 8132
rect 7704 8188 7768 8192
rect 7704 8132 7708 8188
rect 7708 8132 7764 8188
rect 7764 8132 7768 8188
rect 7704 8128 7768 8132
rect 7784 8188 7848 8192
rect 7784 8132 7788 8188
rect 7788 8132 7844 8188
rect 7844 8132 7848 8188
rect 7784 8128 7848 8132
rect 7864 8188 7928 8192
rect 7864 8132 7868 8188
rect 7868 8132 7924 8188
rect 7924 8132 7928 8188
rect 7864 8128 7928 8132
rect 12072 8188 12136 8192
rect 12072 8132 12076 8188
rect 12076 8132 12132 8188
rect 12132 8132 12136 8188
rect 12072 8128 12136 8132
rect 12152 8188 12216 8192
rect 12152 8132 12156 8188
rect 12156 8132 12212 8188
rect 12212 8132 12216 8188
rect 12152 8128 12216 8132
rect 12232 8188 12296 8192
rect 12232 8132 12236 8188
rect 12236 8132 12292 8188
rect 12292 8132 12296 8188
rect 12232 8128 12296 8132
rect 12312 8188 12376 8192
rect 12312 8132 12316 8188
rect 12316 8132 12372 8188
rect 12372 8132 12376 8188
rect 12312 8128 12376 8132
rect 16520 8188 16584 8192
rect 16520 8132 16524 8188
rect 16524 8132 16580 8188
rect 16580 8132 16584 8188
rect 16520 8128 16584 8132
rect 16600 8188 16664 8192
rect 16600 8132 16604 8188
rect 16604 8132 16660 8188
rect 16660 8132 16664 8188
rect 16600 8128 16664 8132
rect 16680 8188 16744 8192
rect 16680 8132 16684 8188
rect 16684 8132 16740 8188
rect 16740 8132 16744 8188
rect 16680 8128 16744 8132
rect 16760 8188 16824 8192
rect 16760 8132 16764 8188
rect 16764 8132 16820 8188
rect 16820 8132 16824 8188
rect 16760 8128 16824 8132
rect 6132 8060 6196 8124
rect 17356 8120 17420 8124
rect 17356 8064 17370 8120
rect 17370 8064 17420 8120
rect 17356 8060 17420 8064
rect 3556 7652 3620 7716
rect 15884 7712 15948 7716
rect 15884 7656 15934 7712
rect 15934 7656 15948 7712
rect 15884 7652 15948 7656
rect 16252 7652 16316 7716
rect 5400 7644 5464 7648
rect 5400 7588 5404 7644
rect 5404 7588 5460 7644
rect 5460 7588 5464 7644
rect 5400 7584 5464 7588
rect 5480 7644 5544 7648
rect 5480 7588 5484 7644
rect 5484 7588 5540 7644
rect 5540 7588 5544 7644
rect 5480 7584 5544 7588
rect 5560 7644 5624 7648
rect 5560 7588 5564 7644
rect 5564 7588 5620 7644
rect 5620 7588 5624 7644
rect 5560 7584 5624 7588
rect 5640 7644 5704 7648
rect 5640 7588 5644 7644
rect 5644 7588 5700 7644
rect 5700 7588 5704 7644
rect 5640 7584 5704 7588
rect 9848 7644 9912 7648
rect 9848 7588 9852 7644
rect 9852 7588 9908 7644
rect 9908 7588 9912 7644
rect 9848 7584 9912 7588
rect 9928 7644 9992 7648
rect 9928 7588 9932 7644
rect 9932 7588 9988 7644
rect 9988 7588 9992 7644
rect 9928 7584 9992 7588
rect 10008 7644 10072 7648
rect 10008 7588 10012 7644
rect 10012 7588 10068 7644
rect 10068 7588 10072 7644
rect 10008 7584 10072 7588
rect 10088 7644 10152 7648
rect 10088 7588 10092 7644
rect 10092 7588 10148 7644
rect 10148 7588 10152 7644
rect 10088 7584 10152 7588
rect 14296 7644 14360 7648
rect 14296 7588 14300 7644
rect 14300 7588 14356 7644
rect 14356 7588 14360 7644
rect 14296 7584 14360 7588
rect 14376 7644 14440 7648
rect 14376 7588 14380 7644
rect 14380 7588 14436 7644
rect 14436 7588 14440 7644
rect 14376 7584 14440 7588
rect 14456 7644 14520 7648
rect 14456 7588 14460 7644
rect 14460 7588 14516 7644
rect 14516 7588 14520 7644
rect 14456 7584 14520 7588
rect 14536 7644 14600 7648
rect 14536 7588 14540 7644
rect 14540 7588 14596 7644
rect 14596 7588 14600 7644
rect 14536 7584 14600 7588
rect 2820 7516 2884 7580
rect 17908 7244 17972 7308
rect 10548 7108 10612 7172
rect 3176 7100 3240 7104
rect 3176 7044 3180 7100
rect 3180 7044 3236 7100
rect 3236 7044 3240 7100
rect 3176 7040 3240 7044
rect 3256 7100 3320 7104
rect 3256 7044 3260 7100
rect 3260 7044 3316 7100
rect 3316 7044 3320 7100
rect 3256 7040 3320 7044
rect 3336 7100 3400 7104
rect 3336 7044 3340 7100
rect 3340 7044 3396 7100
rect 3396 7044 3400 7100
rect 3336 7040 3400 7044
rect 3416 7100 3480 7104
rect 3416 7044 3420 7100
rect 3420 7044 3476 7100
rect 3476 7044 3480 7100
rect 3416 7040 3480 7044
rect 7624 7100 7688 7104
rect 7624 7044 7628 7100
rect 7628 7044 7684 7100
rect 7684 7044 7688 7100
rect 7624 7040 7688 7044
rect 7704 7100 7768 7104
rect 7704 7044 7708 7100
rect 7708 7044 7764 7100
rect 7764 7044 7768 7100
rect 7704 7040 7768 7044
rect 7784 7100 7848 7104
rect 7784 7044 7788 7100
rect 7788 7044 7844 7100
rect 7844 7044 7848 7100
rect 7784 7040 7848 7044
rect 7864 7100 7928 7104
rect 7864 7044 7868 7100
rect 7868 7044 7924 7100
rect 7924 7044 7928 7100
rect 7864 7040 7928 7044
rect 12072 7100 12136 7104
rect 12072 7044 12076 7100
rect 12076 7044 12132 7100
rect 12132 7044 12136 7100
rect 12072 7040 12136 7044
rect 12152 7100 12216 7104
rect 12152 7044 12156 7100
rect 12156 7044 12212 7100
rect 12212 7044 12216 7100
rect 12152 7040 12216 7044
rect 12232 7100 12296 7104
rect 12232 7044 12236 7100
rect 12236 7044 12292 7100
rect 12292 7044 12296 7100
rect 12232 7040 12296 7044
rect 12312 7100 12376 7104
rect 12312 7044 12316 7100
rect 12316 7044 12372 7100
rect 12372 7044 12376 7100
rect 12312 7040 12376 7044
rect 16520 7100 16584 7104
rect 16520 7044 16524 7100
rect 16524 7044 16580 7100
rect 16580 7044 16584 7100
rect 16520 7040 16584 7044
rect 16600 7100 16664 7104
rect 16600 7044 16604 7100
rect 16604 7044 16660 7100
rect 16660 7044 16664 7100
rect 16600 7040 16664 7044
rect 16680 7100 16744 7104
rect 16680 7044 16684 7100
rect 16684 7044 16740 7100
rect 16740 7044 16744 7100
rect 16680 7040 16744 7044
rect 16760 7100 16824 7104
rect 16760 7044 16764 7100
rect 16764 7044 16820 7100
rect 16820 7044 16824 7100
rect 16760 7040 16824 7044
rect 3004 6836 3068 6900
rect 5028 6836 5092 6900
rect 6684 6896 6748 6900
rect 6684 6840 6734 6896
rect 6734 6840 6748 6896
rect 6684 6836 6748 6840
rect 8156 6836 8220 6900
rect 9260 6896 9324 6900
rect 9260 6840 9274 6896
rect 9274 6840 9324 6896
rect 9260 6836 9324 6840
rect 12756 6896 12820 6900
rect 12756 6840 12770 6896
rect 12770 6840 12820 6896
rect 12756 6836 12820 6840
rect 2636 6700 2700 6764
rect 4292 6700 4356 6764
rect 2268 6564 2332 6628
rect 5400 6556 5464 6560
rect 5400 6500 5404 6556
rect 5404 6500 5460 6556
rect 5460 6500 5464 6556
rect 5400 6496 5464 6500
rect 5480 6556 5544 6560
rect 5480 6500 5484 6556
rect 5484 6500 5540 6556
rect 5540 6500 5544 6556
rect 5480 6496 5544 6500
rect 5560 6556 5624 6560
rect 5560 6500 5564 6556
rect 5564 6500 5620 6556
rect 5620 6500 5624 6556
rect 5560 6496 5624 6500
rect 5640 6556 5704 6560
rect 5640 6500 5644 6556
rect 5644 6500 5700 6556
rect 5700 6500 5704 6556
rect 5640 6496 5704 6500
rect 9848 6556 9912 6560
rect 9848 6500 9852 6556
rect 9852 6500 9908 6556
rect 9908 6500 9912 6556
rect 9848 6496 9912 6500
rect 9928 6556 9992 6560
rect 9928 6500 9932 6556
rect 9932 6500 9988 6556
rect 9988 6500 9992 6556
rect 9928 6496 9992 6500
rect 10008 6556 10072 6560
rect 10008 6500 10012 6556
rect 10012 6500 10068 6556
rect 10068 6500 10072 6556
rect 10008 6496 10072 6500
rect 10088 6556 10152 6560
rect 10088 6500 10092 6556
rect 10092 6500 10148 6556
rect 10148 6500 10152 6556
rect 10088 6496 10152 6500
rect 14296 6556 14360 6560
rect 14296 6500 14300 6556
rect 14300 6500 14356 6556
rect 14356 6500 14360 6556
rect 14296 6496 14360 6500
rect 14376 6556 14440 6560
rect 14376 6500 14380 6556
rect 14380 6500 14436 6556
rect 14436 6500 14440 6556
rect 14376 6496 14440 6500
rect 14456 6556 14520 6560
rect 14456 6500 14460 6556
rect 14460 6500 14516 6556
rect 14516 6500 14520 6556
rect 14456 6496 14520 6500
rect 14536 6556 14600 6560
rect 14536 6500 14540 6556
rect 14540 6500 14596 6556
rect 14596 6500 14600 6556
rect 14536 6496 14600 6500
rect 3924 6428 3988 6492
rect 2084 6156 2148 6220
rect 11284 6020 11348 6084
rect 3176 6012 3240 6016
rect 3176 5956 3180 6012
rect 3180 5956 3236 6012
rect 3236 5956 3240 6012
rect 3176 5952 3240 5956
rect 3256 6012 3320 6016
rect 3256 5956 3260 6012
rect 3260 5956 3316 6012
rect 3316 5956 3320 6012
rect 3256 5952 3320 5956
rect 3336 6012 3400 6016
rect 3336 5956 3340 6012
rect 3340 5956 3396 6012
rect 3396 5956 3400 6012
rect 3336 5952 3400 5956
rect 3416 6012 3480 6016
rect 3416 5956 3420 6012
rect 3420 5956 3476 6012
rect 3476 5956 3480 6012
rect 3416 5952 3480 5956
rect 7624 6012 7688 6016
rect 7624 5956 7628 6012
rect 7628 5956 7684 6012
rect 7684 5956 7688 6012
rect 7624 5952 7688 5956
rect 7704 6012 7768 6016
rect 7704 5956 7708 6012
rect 7708 5956 7764 6012
rect 7764 5956 7768 6012
rect 7704 5952 7768 5956
rect 7784 6012 7848 6016
rect 7784 5956 7788 6012
rect 7788 5956 7844 6012
rect 7844 5956 7848 6012
rect 7784 5952 7848 5956
rect 7864 6012 7928 6016
rect 7864 5956 7868 6012
rect 7868 5956 7924 6012
rect 7924 5956 7928 6012
rect 7864 5952 7928 5956
rect 12072 6012 12136 6016
rect 12072 5956 12076 6012
rect 12076 5956 12132 6012
rect 12132 5956 12136 6012
rect 12072 5952 12136 5956
rect 12152 6012 12216 6016
rect 12152 5956 12156 6012
rect 12156 5956 12212 6012
rect 12212 5956 12216 6012
rect 12152 5952 12216 5956
rect 12232 6012 12296 6016
rect 12232 5956 12236 6012
rect 12236 5956 12292 6012
rect 12292 5956 12296 6012
rect 12232 5952 12296 5956
rect 12312 6012 12376 6016
rect 12312 5956 12316 6012
rect 12316 5956 12372 6012
rect 12372 5956 12376 6012
rect 12312 5952 12376 5956
rect 16520 6012 16584 6016
rect 16520 5956 16524 6012
rect 16524 5956 16580 6012
rect 16580 5956 16584 6012
rect 16520 5952 16584 5956
rect 16600 6012 16664 6016
rect 16600 5956 16604 6012
rect 16604 5956 16660 6012
rect 16660 5956 16664 6012
rect 16600 5952 16664 5956
rect 16680 6012 16744 6016
rect 16680 5956 16684 6012
rect 16684 5956 16740 6012
rect 16740 5956 16744 6012
rect 16680 5952 16744 5956
rect 16760 6012 16824 6016
rect 16760 5956 16764 6012
rect 16764 5956 16820 6012
rect 16820 5956 16824 6012
rect 16760 5952 16824 5956
rect 5948 5884 6012 5948
rect 4844 5748 4908 5812
rect 3556 5476 3620 5540
rect 6868 5612 6932 5676
rect 6684 5476 6748 5540
rect 7052 5476 7116 5540
rect 11284 5476 11348 5540
rect 15884 5476 15948 5540
rect 16988 5536 17052 5540
rect 16988 5480 17038 5536
rect 17038 5480 17052 5536
rect 16988 5476 17052 5480
rect 5400 5468 5464 5472
rect 5400 5412 5404 5468
rect 5404 5412 5460 5468
rect 5460 5412 5464 5468
rect 5400 5408 5464 5412
rect 5480 5468 5544 5472
rect 5480 5412 5484 5468
rect 5484 5412 5540 5468
rect 5540 5412 5544 5468
rect 5480 5408 5544 5412
rect 5560 5468 5624 5472
rect 5560 5412 5564 5468
rect 5564 5412 5620 5468
rect 5620 5412 5624 5468
rect 5560 5408 5624 5412
rect 5640 5468 5704 5472
rect 5640 5412 5644 5468
rect 5644 5412 5700 5468
rect 5700 5412 5704 5468
rect 5640 5408 5704 5412
rect 9848 5468 9912 5472
rect 9848 5412 9852 5468
rect 9852 5412 9908 5468
rect 9908 5412 9912 5468
rect 9848 5408 9912 5412
rect 9928 5468 9992 5472
rect 9928 5412 9932 5468
rect 9932 5412 9988 5468
rect 9988 5412 9992 5468
rect 9928 5408 9992 5412
rect 10008 5468 10072 5472
rect 10008 5412 10012 5468
rect 10012 5412 10068 5468
rect 10068 5412 10072 5468
rect 10008 5408 10072 5412
rect 10088 5468 10152 5472
rect 10088 5412 10092 5468
rect 10092 5412 10148 5468
rect 10148 5412 10152 5468
rect 10088 5408 10152 5412
rect 14296 5468 14360 5472
rect 14296 5412 14300 5468
rect 14300 5412 14356 5468
rect 14356 5412 14360 5468
rect 14296 5408 14360 5412
rect 14376 5468 14440 5472
rect 14376 5412 14380 5468
rect 14380 5412 14436 5468
rect 14436 5412 14440 5468
rect 14376 5408 14440 5412
rect 14456 5468 14520 5472
rect 14456 5412 14460 5468
rect 14460 5412 14516 5468
rect 14516 5412 14520 5468
rect 14456 5408 14520 5412
rect 14536 5468 14600 5472
rect 14536 5412 14540 5468
rect 14540 5412 14596 5468
rect 14596 5412 14600 5468
rect 14536 5408 14600 5412
rect 5028 5340 5092 5404
rect 6500 5340 6564 5404
rect 3556 5264 3620 5268
rect 3556 5208 3570 5264
rect 3570 5208 3620 5264
rect 3556 5204 3620 5208
rect 6132 5204 6196 5268
rect 2820 5068 2884 5132
rect 3176 4924 3240 4928
rect 3176 4868 3180 4924
rect 3180 4868 3236 4924
rect 3236 4868 3240 4924
rect 3176 4864 3240 4868
rect 3256 4924 3320 4928
rect 3256 4868 3260 4924
rect 3260 4868 3316 4924
rect 3316 4868 3320 4924
rect 3256 4864 3320 4868
rect 3336 4924 3400 4928
rect 3336 4868 3340 4924
rect 3340 4868 3396 4924
rect 3396 4868 3400 4924
rect 3336 4864 3400 4868
rect 3416 4924 3480 4928
rect 3416 4868 3420 4924
rect 3420 4868 3476 4924
rect 3476 4868 3480 4924
rect 3416 4864 3480 4868
rect 7624 4924 7688 4928
rect 7624 4868 7628 4924
rect 7628 4868 7684 4924
rect 7684 4868 7688 4924
rect 7624 4864 7688 4868
rect 7704 4924 7768 4928
rect 7704 4868 7708 4924
rect 7708 4868 7764 4924
rect 7764 4868 7768 4924
rect 7704 4864 7768 4868
rect 7784 4924 7848 4928
rect 7784 4868 7788 4924
rect 7788 4868 7844 4924
rect 7844 4868 7848 4924
rect 7784 4864 7848 4868
rect 7864 4924 7928 4928
rect 7864 4868 7868 4924
rect 7868 4868 7924 4924
rect 7924 4868 7928 4924
rect 7864 4864 7928 4868
rect 12072 4924 12136 4928
rect 12072 4868 12076 4924
rect 12076 4868 12132 4924
rect 12132 4868 12136 4924
rect 12072 4864 12136 4868
rect 12152 4924 12216 4928
rect 12152 4868 12156 4924
rect 12156 4868 12212 4924
rect 12212 4868 12216 4924
rect 12152 4864 12216 4868
rect 12232 4924 12296 4928
rect 12232 4868 12236 4924
rect 12236 4868 12292 4924
rect 12292 4868 12296 4924
rect 12232 4864 12296 4868
rect 12312 4924 12376 4928
rect 12312 4868 12316 4924
rect 12316 4868 12372 4924
rect 12372 4868 12376 4924
rect 12312 4864 12376 4868
rect 16520 4924 16584 4928
rect 16520 4868 16524 4924
rect 16524 4868 16580 4924
rect 16580 4868 16584 4924
rect 16520 4864 16584 4868
rect 16600 4924 16664 4928
rect 16600 4868 16604 4924
rect 16604 4868 16660 4924
rect 16660 4868 16664 4924
rect 16600 4864 16664 4868
rect 16680 4924 16744 4928
rect 16680 4868 16684 4924
rect 16684 4868 16740 4924
rect 16740 4868 16744 4924
rect 16680 4864 16744 4868
rect 16760 4924 16824 4928
rect 16760 4868 16764 4924
rect 16764 4868 16820 4924
rect 16820 4868 16824 4924
rect 16760 4864 16824 4868
rect 4844 4796 4908 4860
rect 11836 4856 11900 4860
rect 11836 4800 11850 4856
rect 11850 4800 11900 4856
rect 11836 4796 11900 4800
rect 17356 4796 17420 4860
rect 3924 4660 3988 4724
rect 10732 4720 10796 4724
rect 10732 4664 10782 4720
rect 10782 4664 10796 4720
rect 10732 4660 10796 4664
rect 5948 4524 6012 4588
rect 2084 4388 2148 4452
rect 12756 4448 12820 4452
rect 12756 4392 12806 4448
rect 12806 4392 12820 4448
rect 12756 4388 12820 4392
rect 12940 4448 13004 4452
rect 12940 4392 12990 4448
rect 12990 4392 13004 4448
rect 12940 4388 13004 4392
rect 5400 4380 5464 4384
rect 5400 4324 5404 4380
rect 5404 4324 5460 4380
rect 5460 4324 5464 4380
rect 5400 4320 5464 4324
rect 5480 4380 5544 4384
rect 5480 4324 5484 4380
rect 5484 4324 5540 4380
rect 5540 4324 5544 4380
rect 5480 4320 5544 4324
rect 5560 4380 5624 4384
rect 5560 4324 5564 4380
rect 5564 4324 5620 4380
rect 5620 4324 5624 4380
rect 5560 4320 5624 4324
rect 5640 4380 5704 4384
rect 5640 4324 5644 4380
rect 5644 4324 5700 4380
rect 5700 4324 5704 4380
rect 5640 4320 5704 4324
rect 9848 4380 9912 4384
rect 9848 4324 9852 4380
rect 9852 4324 9908 4380
rect 9908 4324 9912 4380
rect 9848 4320 9912 4324
rect 9928 4380 9992 4384
rect 9928 4324 9932 4380
rect 9932 4324 9988 4380
rect 9988 4324 9992 4380
rect 9928 4320 9992 4324
rect 10008 4380 10072 4384
rect 10008 4324 10012 4380
rect 10012 4324 10068 4380
rect 10068 4324 10072 4380
rect 10008 4320 10072 4324
rect 10088 4380 10152 4384
rect 10088 4324 10092 4380
rect 10092 4324 10148 4380
rect 10148 4324 10152 4380
rect 10088 4320 10152 4324
rect 14296 4380 14360 4384
rect 14296 4324 14300 4380
rect 14300 4324 14356 4380
rect 14356 4324 14360 4380
rect 14296 4320 14360 4324
rect 14376 4380 14440 4384
rect 14376 4324 14380 4380
rect 14380 4324 14436 4380
rect 14436 4324 14440 4380
rect 14376 4320 14440 4324
rect 14456 4380 14520 4384
rect 14456 4324 14460 4380
rect 14460 4324 14516 4380
rect 14516 4324 14520 4380
rect 14456 4320 14520 4324
rect 14536 4380 14600 4384
rect 14536 4324 14540 4380
rect 14540 4324 14596 4380
rect 14596 4324 14600 4380
rect 14536 4320 14600 4324
rect 3740 4312 3804 4316
rect 3740 4256 3790 4312
rect 3790 4256 3804 4312
rect 3740 4252 3804 4256
rect 6868 4312 6932 4316
rect 6868 4256 6918 4312
rect 6918 4256 6932 4312
rect 6868 4252 6932 4256
rect 17908 4252 17972 4316
rect 7420 4176 7484 4180
rect 7420 4120 7470 4176
rect 7470 4120 7484 4176
rect 7420 4116 7484 4120
rect 2636 4040 2700 4044
rect 2636 3984 2686 4040
rect 2686 3984 2700 4040
rect 2636 3980 2700 3984
rect 7236 3980 7300 4044
rect 3176 3836 3240 3840
rect 3176 3780 3180 3836
rect 3180 3780 3236 3836
rect 3236 3780 3240 3836
rect 3176 3776 3240 3780
rect 3256 3836 3320 3840
rect 3256 3780 3260 3836
rect 3260 3780 3316 3836
rect 3316 3780 3320 3836
rect 3256 3776 3320 3780
rect 3336 3836 3400 3840
rect 3336 3780 3340 3836
rect 3340 3780 3396 3836
rect 3396 3780 3400 3836
rect 3336 3776 3400 3780
rect 3416 3836 3480 3840
rect 3416 3780 3420 3836
rect 3420 3780 3476 3836
rect 3476 3780 3480 3836
rect 3416 3776 3480 3780
rect 7624 3836 7688 3840
rect 7624 3780 7628 3836
rect 7628 3780 7684 3836
rect 7684 3780 7688 3836
rect 7624 3776 7688 3780
rect 7704 3836 7768 3840
rect 7704 3780 7708 3836
rect 7708 3780 7764 3836
rect 7764 3780 7768 3836
rect 7704 3776 7768 3780
rect 7784 3836 7848 3840
rect 7784 3780 7788 3836
rect 7788 3780 7844 3836
rect 7844 3780 7848 3836
rect 7784 3776 7848 3780
rect 7864 3836 7928 3840
rect 7864 3780 7868 3836
rect 7868 3780 7924 3836
rect 7924 3780 7928 3836
rect 7864 3776 7928 3780
rect 12072 3836 12136 3840
rect 12072 3780 12076 3836
rect 12076 3780 12132 3836
rect 12132 3780 12136 3836
rect 12072 3776 12136 3780
rect 12152 3836 12216 3840
rect 12152 3780 12156 3836
rect 12156 3780 12212 3836
rect 12212 3780 12216 3836
rect 12152 3776 12216 3780
rect 12232 3836 12296 3840
rect 12232 3780 12236 3836
rect 12236 3780 12292 3836
rect 12292 3780 12296 3836
rect 12232 3776 12296 3780
rect 12312 3836 12376 3840
rect 12312 3780 12316 3836
rect 12316 3780 12372 3836
rect 12372 3780 12376 3836
rect 12312 3776 12376 3780
rect 16520 3836 16584 3840
rect 16520 3780 16524 3836
rect 16524 3780 16580 3836
rect 16580 3780 16584 3836
rect 16520 3776 16584 3780
rect 16600 3836 16664 3840
rect 16600 3780 16604 3836
rect 16604 3780 16660 3836
rect 16660 3780 16664 3836
rect 16600 3776 16664 3780
rect 16680 3836 16744 3840
rect 16680 3780 16684 3836
rect 16684 3780 16740 3836
rect 16740 3780 16744 3836
rect 16680 3776 16744 3780
rect 16760 3836 16824 3840
rect 16760 3780 16764 3836
rect 16764 3780 16820 3836
rect 16820 3780 16824 3836
rect 16760 3776 16824 3780
rect 9076 3436 9140 3500
rect 5400 3292 5464 3296
rect 5400 3236 5404 3292
rect 5404 3236 5460 3292
rect 5460 3236 5464 3292
rect 5400 3232 5464 3236
rect 5480 3292 5544 3296
rect 5480 3236 5484 3292
rect 5484 3236 5540 3292
rect 5540 3236 5544 3292
rect 5480 3232 5544 3236
rect 5560 3292 5624 3296
rect 5560 3236 5564 3292
rect 5564 3236 5620 3292
rect 5620 3236 5624 3292
rect 5560 3232 5624 3236
rect 5640 3292 5704 3296
rect 5640 3236 5644 3292
rect 5644 3236 5700 3292
rect 5700 3236 5704 3292
rect 5640 3232 5704 3236
rect 9848 3292 9912 3296
rect 9848 3236 9852 3292
rect 9852 3236 9908 3292
rect 9908 3236 9912 3292
rect 9848 3232 9912 3236
rect 9928 3292 9992 3296
rect 9928 3236 9932 3292
rect 9932 3236 9988 3292
rect 9988 3236 9992 3292
rect 9928 3232 9992 3236
rect 10008 3292 10072 3296
rect 10008 3236 10012 3292
rect 10012 3236 10068 3292
rect 10068 3236 10072 3292
rect 10008 3232 10072 3236
rect 10088 3292 10152 3296
rect 10088 3236 10092 3292
rect 10092 3236 10148 3292
rect 10148 3236 10152 3292
rect 10088 3232 10152 3236
rect 14296 3292 14360 3296
rect 14296 3236 14300 3292
rect 14300 3236 14356 3292
rect 14356 3236 14360 3292
rect 14296 3232 14360 3236
rect 14376 3292 14440 3296
rect 14376 3236 14380 3292
rect 14380 3236 14436 3292
rect 14436 3236 14440 3292
rect 14376 3232 14440 3236
rect 14456 3292 14520 3296
rect 14456 3236 14460 3292
rect 14460 3236 14516 3292
rect 14516 3236 14520 3292
rect 14456 3232 14520 3236
rect 14536 3292 14600 3296
rect 14536 3236 14540 3292
rect 14540 3236 14596 3292
rect 14596 3236 14600 3292
rect 14536 3232 14600 3236
rect 5212 3164 5276 3228
rect 10364 3164 10428 3228
rect 13860 3224 13924 3228
rect 13860 3168 13874 3224
rect 13874 3168 13924 3224
rect 13860 3164 13924 3168
rect 14044 3224 14108 3228
rect 14044 3168 14058 3224
rect 14058 3168 14108 3224
rect 14044 3164 14108 3168
rect 16252 2892 16316 2956
rect 3176 2748 3240 2752
rect 3176 2692 3180 2748
rect 3180 2692 3236 2748
rect 3236 2692 3240 2748
rect 3176 2688 3240 2692
rect 3256 2748 3320 2752
rect 3256 2692 3260 2748
rect 3260 2692 3316 2748
rect 3316 2692 3320 2748
rect 3256 2688 3320 2692
rect 3336 2748 3400 2752
rect 3336 2692 3340 2748
rect 3340 2692 3396 2748
rect 3396 2692 3400 2748
rect 3336 2688 3400 2692
rect 3416 2748 3480 2752
rect 3416 2692 3420 2748
rect 3420 2692 3476 2748
rect 3476 2692 3480 2748
rect 3416 2688 3480 2692
rect 7624 2748 7688 2752
rect 7624 2692 7628 2748
rect 7628 2692 7684 2748
rect 7684 2692 7688 2748
rect 7624 2688 7688 2692
rect 7704 2748 7768 2752
rect 7704 2692 7708 2748
rect 7708 2692 7764 2748
rect 7764 2692 7768 2748
rect 7704 2688 7768 2692
rect 7784 2748 7848 2752
rect 7784 2692 7788 2748
rect 7788 2692 7844 2748
rect 7844 2692 7848 2748
rect 7784 2688 7848 2692
rect 7864 2748 7928 2752
rect 7864 2692 7868 2748
rect 7868 2692 7924 2748
rect 7924 2692 7928 2748
rect 7864 2688 7928 2692
rect 12072 2748 12136 2752
rect 12072 2692 12076 2748
rect 12076 2692 12132 2748
rect 12132 2692 12136 2748
rect 12072 2688 12136 2692
rect 12152 2748 12216 2752
rect 12152 2692 12156 2748
rect 12156 2692 12212 2748
rect 12212 2692 12216 2748
rect 12152 2688 12216 2692
rect 12232 2748 12296 2752
rect 12232 2692 12236 2748
rect 12236 2692 12292 2748
rect 12292 2692 12296 2748
rect 12232 2688 12296 2692
rect 12312 2748 12376 2752
rect 12312 2692 12316 2748
rect 12316 2692 12372 2748
rect 12372 2692 12376 2748
rect 12312 2688 12376 2692
rect 16520 2748 16584 2752
rect 16520 2692 16524 2748
rect 16524 2692 16580 2748
rect 16580 2692 16584 2748
rect 16520 2688 16584 2692
rect 16600 2748 16664 2752
rect 16600 2692 16604 2748
rect 16604 2692 16660 2748
rect 16660 2692 16664 2748
rect 16600 2688 16664 2692
rect 16680 2748 16744 2752
rect 16680 2692 16684 2748
rect 16684 2692 16740 2748
rect 16740 2692 16744 2748
rect 16680 2688 16744 2692
rect 16760 2748 16824 2752
rect 16760 2692 16764 2748
rect 16764 2692 16820 2748
rect 16820 2692 16824 2748
rect 16760 2688 16824 2692
rect 13492 2680 13556 2684
rect 13492 2624 13542 2680
rect 13542 2624 13556 2680
rect 13492 2620 13556 2624
rect 15884 2620 15948 2684
rect 13676 2544 13740 2548
rect 13676 2488 13726 2544
rect 13726 2488 13740 2544
rect 13676 2484 13740 2488
rect 14964 2484 15028 2548
rect 11652 2348 11716 2412
rect 5400 2204 5464 2208
rect 5400 2148 5404 2204
rect 5404 2148 5460 2204
rect 5460 2148 5464 2204
rect 5400 2144 5464 2148
rect 5480 2204 5544 2208
rect 5480 2148 5484 2204
rect 5484 2148 5540 2204
rect 5540 2148 5544 2204
rect 5480 2144 5544 2148
rect 5560 2204 5624 2208
rect 5560 2148 5564 2204
rect 5564 2148 5620 2204
rect 5620 2148 5624 2204
rect 5560 2144 5624 2148
rect 5640 2204 5704 2208
rect 5640 2148 5644 2204
rect 5644 2148 5700 2204
rect 5700 2148 5704 2204
rect 5640 2144 5704 2148
rect 9848 2204 9912 2208
rect 9848 2148 9852 2204
rect 9852 2148 9908 2204
rect 9908 2148 9912 2204
rect 9848 2144 9912 2148
rect 9928 2204 9992 2208
rect 9928 2148 9932 2204
rect 9932 2148 9988 2204
rect 9988 2148 9992 2204
rect 9928 2144 9992 2148
rect 10008 2204 10072 2208
rect 10008 2148 10012 2204
rect 10012 2148 10068 2204
rect 10068 2148 10072 2204
rect 10008 2144 10072 2148
rect 10088 2204 10152 2208
rect 10088 2148 10092 2204
rect 10092 2148 10148 2204
rect 10148 2148 10152 2204
rect 10088 2144 10152 2148
rect 14296 2204 14360 2208
rect 14296 2148 14300 2204
rect 14300 2148 14356 2204
rect 14356 2148 14360 2204
rect 14296 2144 14360 2148
rect 14376 2204 14440 2208
rect 14376 2148 14380 2204
rect 14380 2148 14436 2204
rect 14436 2148 14440 2204
rect 14376 2144 14440 2148
rect 14456 2204 14520 2208
rect 14456 2148 14460 2204
rect 14460 2148 14516 2204
rect 14516 2148 14520 2204
rect 14456 2144 14520 2148
rect 14536 2204 14600 2208
rect 14536 2148 14540 2204
rect 14540 2148 14596 2204
rect 14596 2148 14600 2204
rect 14536 2144 14600 2148
<< metal4 >>
rect 13675 15060 13741 15061
rect 13675 14996 13676 15060
rect 13740 14996 13741 15060
rect 13675 14995 13741 14996
rect 3168 14720 3488 14736
rect 3168 14656 3176 14720
rect 3240 14656 3256 14720
rect 3320 14656 3336 14720
rect 3400 14656 3416 14720
rect 3480 14656 3488 14720
rect 3003 14108 3069 14109
rect 3003 14044 3004 14108
rect 3068 14044 3069 14108
rect 3003 14043 3069 14044
rect 2083 9348 2149 9349
rect 2083 9284 2084 9348
rect 2148 9284 2149 9348
rect 2083 9283 2149 9284
rect 2086 6221 2146 9283
rect 2267 8532 2333 8533
rect 2267 8468 2268 8532
rect 2332 8468 2333 8532
rect 2267 8467 2333 8468
rect 2270 6629 2330 8467
rect 2819 7580 2885 7581
rect 2819 7516 2820 7580
rect 2884 7516 2885 7580
rect 2819 7515 2885 7516
rect 2635 6764 2701 6765
rect 2635 6700 2636 6764
rect 2700 6700 2701 6764
rect 2635 6699 2701 6700
rect 2267 6628 2333 6629
rect 2267 6564 2268 6628
rect 2332 6564 2333 6628
rect 2267 6563 2333 6564
rect 2083 6220 2149 6221
rect 2083 6156 2084 6220
rect 2148 6156 2149 6220
rect 2083 6155 2149 6156
rect 2086 4453 2146 6155
rect 2083 4452 2149 4453
rect 2083 4388 2084 4452
rect 2148 4388 2149 4452
rect 2083 4387 2149 4388
rect 2638 4045 2698 6699
rect 2822 5133 2882 7515
rect 3006 6901 3066 14043
rect 3168 13632 3488 14656
rect 3168 13568 3176 13632
rect 3240 13568 3256 13632
rect 3320 13568 3336 13632
rect 3400 13568 3416 13632
rect 3480 13568 3488 13632
rect 3168 12544 3488 13568
rect 3168 12480 3176 12544
rect 3240 12480 3256 12544
rect 3320 12480 3336 12544
rect 3400 12480 3416 12544
rect 3480 12480 3488 12544
rect 3168 11456 3488 12480
rect 5392 14176 5712 14736
rect 5392 14112 5400 14176
rect 5464 14112 5480 14176
rect 5544 14112 5560 14176
rect 5624 14112 5640 14176
rect 5704 14112 5712 14176
rect 5392 13088 5712 14112
rect 5392 13024 5400 13088
rect 5464 13024 5480 13088
rect 5544 13024 5560 13088
rect 5624 13024 5640 13088
rect 5704 13024 5712 13088
rect 4291 12204 4357 12205
rect 4291 12140 4292 12204
rect 4356 12140 4357 12204
rect 4291 12139 4357 12140
rect 3168 11392 3176 11456
rect 3240 11392 3256 11456
rect 3320 11392 3336 11456
rect 3400 11392 3416 11456
rect 3480 11392 3488 11456
rect 3168 10368 3488 11392
rect 3739 10708 3805 10709
rect 3739 10644 3740 10708
rect 3804 10644 3805 10708
rect 3739 10643 3805 10644
rect 3168 10304 3176 10368
rect 3240 10304 3256 10368
rect 3320 10304 3336 10368
rect 3400 10304 3416 10368
rect 3480 10304 3488 10368
rect 3168 9280 3488 10304
rect 3168 9216 3176 9280
rect 3240 9216 3256 9280
rect 3320 9216 3336 9280
rect 3400 9216 3416 9280
rect 3480 9216 3488 9280
rect 3168 8192 3488 9216
rect 3168 8128 3176 8192
rect 3240 8128 3256 8192
rect 3320 8128 3336 8192
rect 3400 8128 3416 8192
rect 3480 8128 3488 8192
rect 3168 7104 3488 8128
rect 3555 7716 3621 7717
rect 3555 7652 3556 7716
rect 3620 7652 3621 7716
rect 3555 7651 3621 7652
rect 3168 7040 3176 7104
rect 3240 7040 3256 7104
rect 3320 7040 3336 7104
rect 3400 7040 3416 7104
rect 3480 7040 3488 7104
rect 3003 6900 3069 6901
rect 3003 6836 3004 6900
rect 3068 6836 3069 6900
rect 3003 6835 3069 6836
rect 3168 6016 3488 7040
rect 3168 5952 3176 6016
rect 3240 5952 3256 6016
rect 3320 5952 3336 6016
rect 3400 5952 3416 6016
rect 3480 5952 3488 6016
rect 2819 5132 2885 5133
rect 2819 5068 2820 5132
rect 2884 5068 2885 5132
rect 2819 5067 2885 5068
rect 3168 4928 3488 5952
rect 3558 5541 3618 7651
rect 3555 5540 3621 5541
rect 3555 5476 3556 5540
rect 3620 5476 3621 5540
rect 3555 5475 3621 5476
rect 3555 5268 3621 5269
rect 3555 5204 3556 5268
rect 3620 5266 3621 5268
rect 3742 5266 3802 10643
rect 4294 6765 4354 12139
rect 5392 12000 5712 13024
rect 7616 14720 7936 14736
rect 7616 14656 7624 14720
rect 7688 14656 7704 14720
rect 7768 14656 7784 14720
rect 7848 14656 7864 14720
rect 7928 14656 7936 14720
rect 7616 13632 7936 14656
rect 9840 14176 10160 14736
rect 9840 14112 9848 14176
rect 9912 14112 9928 14176
rect 9992 14112 10008 14176
rect 10072 14112 10088 14176
rect 10152 14112 10160 14176
rect 9075 13972 9141 13973
rect 9075 13908 9076 13972
rect 9140 13908 9141 13972
rect 9075 13907 9141 13908
rect 7616 13568 7624 13632
rect 7688 13568 7704 13632
rect 7768 13568 7784 13632
rect 7848 13568 7864 13632
rect 7928 13568 7936 13632
rect 7419 12748 7485 12749
rect 7419 12684 7420 12748
rect 7484 12684 7485 12748
rect 7419 12683 7485 12684
rect 7422 12450 7482 12683
rect 5392 11936 5400 12000
rect 5464 11936 5480 12000
rect 5544 11936 5560 12000
rect 5624 11936 5640 12000
rect 5704 11936 5712 12000
rect 5211 11796 5277 11797
rect 5211 11732 5212 11796
rect 5276 11732 5277 11796
rect 5211 11731 5277 11732
rect 5027 10436 5093 10437
rect 5027 10372 5028 10436
rect 5092 10372 5093 10436
rect 5027 10371 5093 10372
rect 4843 9212 4909 9213
rect 4843 9148 4844 9212
rect 4908 9148 4909 9212
rect 4843 9147 4909 9148
rect 4291 6764 4357 6765
rect 4291 6700 4292 6764
rect 4356 6700 4357 6764
rect 4291 6699 4357 6700
rect 3923 6492 3989 6493
rect 3923 6428 3924 6492
rect 3988 6428 3989 6492
rect 3923 6427 3989 6428
rect 3620 5206 3802 5266
rect 3620 5204 3621 5206
rect 3555 5203 3621 5204
rect 3168 4864 3176 4928
rect 3240 4864 3256 4928
rect 3320 4864 3336 4928
rect 3400 4864 3416 4928
rect 3480 4864 3488 4928
rect 2635 4044 2701 4045
rect 2635 3980 2636 4044
rect 2700 3980 2701 4044
rect 2635 3979 2701 3980
rect 3168 3840 3488 4864
rect 3742 4317 3802 5206
rect 3926 4725 3986 6427
rect 4846 5813 4906 9147
rect 5030 6901 5090 10371
rect 5027 6900 5093 6901
rect 5027 6836 5028 6900
rect 5092 6836 5093 6900
rect 5027 6835 5093 6836
rect 4843 5812 4909 5813
rect 4843 5748 4844 5812
rect 4908 5748 4909 5812
rect 4843 5747 4909 5748
rect 4846 4861 4906 5747
rect 5030 5405 5090 6835
rect 5027 5404 5093 5405
rect 5027 5340 5028 5404
rect 5092 5340 5093 5404
rect 5027 5339 5093 5340
rect 4843 4860 4909 4861
rect 4843 4796 4844 4860
rect 4908 4796 4909 4860
rect 4843 4795 4909 4796
rect 3923 4724 3989 4725
rect 3923 4660 3924 4724
rect 3988 4660 3989 4724
rect 3923 4659 3989 4660
rect 3739 4316 3805 4317
rect 3739 4252 3740 4316
rect 3804 4252 3805 4316
rect 3739 4251 3805 4252
rect 3168 3776 3176 3840
rect 3240 3776 3256 3840
rect 3320 3776 3336 3840
rect 3400 3776 3416 3840
rect 3480 3776 3488 3840
rect 3168 2752 3488 3776
rect 5214 3229 5274 11731
rect 5392 10912 5712 11936
rect 5392 10848 5400 10912
rect 5464 10848 5480 10912
rect 5544 10848 5560 10912
rect 5624 10848 5640 10912
rect 5704 10848 5712 10912
rect 5392 9824 5712 10848
rect 5392 9760 5400 9824
rect 5464 9760 5480 9824
rect 5544 9760 5560 9824
rect 5624 9760 5640 9824
rect 5704 9760 5712 9824
rect 5392 8736 5712 9760
rect 7238 12390 7482 12450
rect 7616 12544 7936 13568
rect 7616 12480 7624 12544
rect 7688 12480 7704 12544
rect 7768 12480 7784 12544
rect 7848 12480 7864 12544
rect 7928 12480 7936 12544
rect 6499 9076 6565 9077
rect 6499 9012 6500 9076
rect 6564 9012 6565 9076
rect 6499 9011 6565 9012
rect 5392 8672 5400 8736
rect 5464 8672 5480 8736
rect 5544 8672 5560 8736
rect 5624 8672 5640 8736
rect 5704 8672 5712 8736
rect 5392 7648 5712 8672
rect 6131 8124 6197 8125
rect 6131 8060 6132 8124
rect 6196 8060 6197 8124
rect 6131 8059 6197 8060
rect 5392 7584 5400 7648
rect 5464 7584 5480 7648
rect 5544 7584 5560 7648
rect 5624 7584 5640 7648
rect 5704 7584 5712 7648
rect 5392 6560 5712 7584
rect 5392 6496 5400 6560
rect 5464 6496 5480 6560
rect 5544 6496 5560 6560
rect 5624 6496 5640 6560
rect 5704 6496 5712 6560
rect 5392 5472 5712 6496
rect 5947 5948 6013 5949
rect 5947 5884 5948 5948
rect 6012 5884 6013 5948
rect 5947 5883 6013 5884
rect 5392 5408 5400 5472
rect 5464 5408 5480 5472
rect 5544 5408 5560 5472
rect 5624 5408 5640 5472
rect 5704 5408 5712 5472
rect 5392 4384 5712 5408
rect 5950 4589 6010 5883
rect 6134 5269 6194 8059
rect 6502 5405 6562 9011
rect 7051 8804 7117 8805
rect 7051 8740 7052 8804
rect 7116 8740 7117 8804
rect 7051 8739 7117 8740
rect 6867 8396 6933 8397
rect 6867 8332 6868 8396
rect 6932 8332 6933 8396
rect 6867 8331 6933 8332
rect 6683 6900 6749 6901
rect 6683 6836 6684 6900
rect 6748 6836 6749 6900
rect 6683 6835 6749 6836
rect 6686 5541 6746 6835
rect 6870 5677 6930 8331
rect 6867 5676 6933 5677
rect 6867 5612 6868 5676
rect 6932 5612 6933 5676
rect 6867 5611 6933 5612
rect 6683 5540 6749 5541
rect 6683 5476 6684 5540
rect 6748 5476 6749 5540
rect 6683 5475 6749 5476
rect 6499 5404 6565 5405
rect 6499 5340 6500 5404
rect 6564 5340 6565 5404
rect 6499 5339 6565 5340
rect 6131 5268 6197 5269
rect 6131 5204 6132 5268
rect 6196 5204 6197 5268
rect 6131 5203 6197 5204
rect 5947 4588 6013 4589
rect 5947 4524 5948 4588
rect 6012 4524 6013 4588
rect 5947 4523 6013 4524
rect 5392 4320 5400 4384
rect 5464 4320 5480 4384
rect 5544 4320 5560 4384
rect 5624 4320 5640 4384
rect 5704 4320 5712 4384
rect 5392 3296 5712 4320
rect 6870 4317 6930 5611
rect 7054 5541 7114 8739
rect 7051 5540 7117 5541
rect 7051 5476 7052 5540
rect 7116 5476 7117 5540
rect 7051 5475 7117 5476
rect 6867 4316 6933 4317
rect 6867 4252 6868 4316
rect 6932 4252 6933 4316
rect 6867 4251 6933 4252
rect 7238 4045 7298 12390
rect 7616 11456 7936 12480
rect 7616 11392 7624 11456
rect 7688 11392 7704 11456
rect 7768 11392 7784 11456
rect 7848 11392 7864 11456
rect 7928 11392 7936 11456
rect 7616 10368 7936 11392
rect 7616 10304 7624 10368
rect 7688 10304 7704 10368
rect 7768 10304 7784 10368
rect 7848 10304 7864 10368
rect 7928 10304 7936 10368
rect 7419 9756 7485 9757
rect 7419 9692 7420 9756
rect 7484 9692 7485 9756
rect 7419 9691 7485 9692
rect 7422 4181 7482 9691
rect 7616 9280 7936 10304
rect 7616 9216 7624 9280
rect 7688 9216 7704 9280
rect 7768 9216 7784 9280
rect 7848 9216 7864 9280
rect 7928 9216 7936 9280
rect 7616 8192 7936 9216
rect 8155 8396 8221 8397
rect 8155 8332 8156 8396
rect 8220 8332 8221 8396
rect 8155 8331 8221 8332
rect 7616 8128 7624 8192
rect 7688 8128 7704 8192
rect 7768 8128 7784 8192
rect 7848 8128 7864 8192
rect 7928 8128 7936 8192
rect 7616 7104 7936 8128
rect 7616 7040 7624 7104
rect 7688 7040 7704 7104
rect 7768 7040 7784 7104
rect 7848 7040 7864 7104
rect 7928 7040 7936 7104
rect 7616 6016 7936 7040
rect 8158 6901 8218 8331
rect 8155 6900 8221 6901
rect 8155 6836 8156 6900
rect 8220 6836 8221 6900
rect 8155 6835 8221 6836
rect 7616 5952 7624 6016
rect 7688 5952 7704 6016
rect 7768 5952 7784 6016
rect 7848 5952 7864 6016
rect 7928 5952 7936 6016
rect 7616 4928 7936 5952
rect 7616 4864 7624 4928
rect 7688 4864 7704 4928
rect 7768 4864 7784 4928
rect 7848 4864 7864 4928
rect 7928 4864 7936 4928
rect 7419 4180 7485 4181
rect 7419 4116 7420 4180
rect 7484 4116 7485 4180
rect 7419 4115 7485 4116
rect 7235 4044 7301 4045
rect 7235 3980 7236 4044
rect 7300 3980 7301 4044
rect 7235 3979 7301 3980
rect 5392 3232 5400 3296
rect 5464 3232 5480 3296
rect 5544 3232 5560 3296
rect 5624 3232 5640 3296
rect 5704 3232 5712 3296
rect 5211 3228 5277 3229
rect 5211 3164 5212 3228
rect 5276 3164 5277 3228
rect 5211 3163 5277 3164
rect 3168 2688 3176 2752
rect 3240 2688 3256 2752
rect 3320 2688 3336 2752
rect 3400 2688 3416 2752
rect 3480 2688 3488 2752
rect 3168 2128 3488 2688
rect 5392 2208 5712 3232
rect 5392 2144 5400 2208
rect 5464 2144 5480 2208
rect 5544 2144 5560 2208
rect 5624 2144 5640 2208
rect 5704 2144 5712 2208
rect 5392 2128 5712 2144
rect 7616 3840 7936 4864
rect 7616 3776 7624 3840
rect 7688 3776 7704 3840
rect 7768 3776 7784 3840
rect 7848 3776 7864 3840
rect 7928 3776 7936 3840
rect 7616 2752 7936 3776
rect 9078 3501 9138 13907
rect 9840 13088 10160 14112
rect 12064 14720 12384 14736
rect 12064 14656 12072 14720
rect 12136 14656 12152 14720
rect 12216 14656 12232 14720
rect 12296 14656 12312 14720
rect 12376 14656 12384 14720
rect 10363 13972 10429 13973
rect 10363 13908 10364 13972
rect 10428 13908 10429 13972
rect 10363 13907 10429 13908
rect 9840 13024 9848 13088
rect 9912 13024 9928 13088
rect 9992 13024 10008 13088
rect 10072 13024 10088 13088
rect 10152 13024 10160 13088
rect 9259 12748 9325 12749
rect 9259 12684 9260 12748
rect 9324 12684 9325 12748
rect 9259 12683 9325 12684
rect 9262 6901 9322 12683
rect 9840 12000 10160 13024
rect 9840 11936 9848 12000
rect 9912 11936 9928 12000
rect 9992 11936 10008 12000
rect 10072 11936 10088 12000
rect 10152 11936 10160 12000
rect 9840 10912 10160 11936
rect 9840 10848 9848 10912
rect 9912 10848 9928 10912
rect 9992 10848 10008 10912
rect 10072 10848 10088 10912
rect 10152 10848 10160 10912
rect 9840 9824 10160 10848
rect 9840 9760 9848 9824
rect 9912 9760 9928 9824
rect 9992 9760 10008 9824
rect 10072 9760 10088 9824
rect 10152 9760 10160 9824
rect 9840 8736 10160 9760
rect 9840 8672 9848 8736
rect 9912 8672 9928 8736
rect 9992 8672 10008 8736
rect 10072 8672 10088 8736
rect 10152 8672 10160 8736
rect 9840 7648 10160 8672
rect 9840 7584 9848 7648
rect 9912 7584 9928 7648
rect 9992 7584 10008 7648
rect 10072 7584 10088 7648
rect 10152 7584 10160 7648
rect 9259 6900 9325 6901
rect 9259 6836 9260 6900
rect 9324 6836 9325 6900
rect 9259 6835 9325 6836
rect 9840 6560 10160 7584
rect 9840 6496 9848 6560
rect 9912 6496 9928 6560
rect 9992 6496 10008 6560
rect 10072 6496 10088 6560
rect 10152 6496 10160 6560
rect 9840 5472 10160 6496
rect 9840 5408 9848 5472
rect 9912 5408 9928 5472
rect 9992 5408 10008 5472
rect 10072 5408 10088 5472
rect 10152 5408 10160 5472
rect 9840 4384 10160 5408
rect 9840 4320 9848 4384
rect 9912 4320 9928 4384
rect 9992 4320 10008 4384
rect 10072 4320 10088 4384
rect 10152 4320 10160 4384
rect 9075 3500 9141 3501
rect 9075 3436 9076 3500
rect 9140 3436 9141 3500
rect 9075 3435 9141 3436
rect 7616 2688 7624 2752
rect 7688 2688 7704 2752
rect 7768 2688 7784 2752
rect 7848 2688 7864 2752
rect 7928 2688 7936 2752
rect 7616 2128 7936 2688
rect 9840 3296 10160 4320
rect 9840 3232 9848 3296
rect 9912 3232 9928 3296
rect 9992 3232 10008 3296
rect 10072 3232 10088 3296
rect 10152 3232 10160 3296
rect 9840 2208 10160 3232
rect 10366 3229 10426 13907
rect 12064 13632 12384 14656
rect 12064 13568 12072 13632
rect 12136 13568 12152 13632
rect 12216 13568 12232 13632
rect 12296 13568 12312 13632
rect 12376 13568 12384 13632
rect 11835 13428 11901 13429
rect 11835 13364 11836 13428
rect 11900 13364 11901 13428
rect 11835 13363 11901 13364
rect 11283 11932 11349 11933
rect 11283 11868 11284 11932
rect 11348 11868 11349 11932
rect 11283 11867 11349 11868
rect 10731 11116 10797 11117
rect 10731 11052 10732 11116
rect 10796 11052 10797 11116
rect 10731 11051 10797 11052
rect 10547 10844 10613 10845
rect 10547 10780 10548 10844
rect 10612 10780 10613 10844
rect 10547 10779 10613 10780
rect 10550 9757 10610 10779
rect 10547 9756 10613 9757
rect 10547 9692 10548 9756
rect 10612 9692 10613 9756
rect 10547 9691 10613 9692
rect 10547 8260 10613 8261
rect 10547 8196 10548 8260
rect 10612 8196 10613 8260
rect 10547 8195 10613 8196
rect 10550 7173 10610 8195
rect 10547 7172 10613 7173
rect 10547 7108 10548 7172
rect 10612 7108 10613 7172
rect 10547 7107 10613 7108
rect 10734 4725 10794 11051
rect 11286 6085 11346 11867
rect 11651 11524 11717 11525
rect 11651 11460 11652 11524
rect 11716 11460 11717 11524
rect 11651 11459 11717 11460
rect 11283 6084 11349 6085
rect 11283 6020 11284 6084
rect 11348 6020 11349 6084
rect 11283 6019 11349 6020
rect 11286 5541 11346 6019
rect 11283 5540 11349 5541
rect 11283 5476 11284 5540
rect 11348 5476 11349 5540
rect 11283 5475 11349 5476
rect 10731 4724 10797 4725
rect 10731 4660 10732 4724
rect 10796 4660 10797 4724
rect 10731 4659 10797 4660
rect 10363 3228 10429 3229
rect 10363 3164 10364 3228
rect 10428 3164 10429 3228
rect 10363 3163 10429 3164
rect 11654 2413 11714 11459
rect 11838 4861 11898 13363
rect 12064 12544 12384 13568
rect 12064 12480 12072 12544
rect 12136 12480 12152 12544
rect 12216 12480 12232 12544
rect 12296 12480 12312 12544
rect 12376 12480 12384 12544
rect 12064 11456 12384 12480
rect 12939 12068 13005 12069
rect 12939 12004 12940 12068
rect 13004 12004 13005 12068
rect 12939 12003 13005 12004
rect 12064 11392 12072 11456
rect 12136 11392 12152 11456
rect 12216 11392 12232 11456
rect 12296 11392 12312 11456
rect 12376 11392 12384 11456
rect 12064 10368 12384 11392
rect 12064 10304 12072 10368
rect 12136 10304 12152 10368
rect 12216 10304 12232 10368
rect 12296 10304 12312 10368
rect 12376 10304 12384 10368
rect 12064 9280 12384 10304
rect 12064 9216 12072 9280
rect 12136 9216 12152 9280
rect 12216 9216 12232 9280
rect 12296 9216 12312 9280
rect 12376 9216 12384 9280
rect 12064 8192 12384 9216
rect 12064 8128 12072 8192
rect 12136 8128 12152 8192
rect 12216 8128 12232 8192
rect 12296 8128 12312 8192
rect 12376 8128 12384 8192
rect 12064 7104 12384 8128
rect 12064 7040 12072 7104
rect 12136 7040 12152 7104
rect 12216 7040 12232 7104
rect 12296 7040 12312 7104
rect 12376 7040 12384 7104
rect 12064 6016 12384 7040
rect 12755 6900 12821 6901
rect 12755 6836 12756 6900
rect 12820 6836 12821 6900
rect 12755 6835 12821 6836
rect 12064 5952 12072 6016
rect 12136 5952 12152 6016
rect 12216 5952 12232 6016
rect 12296 5952 12312 6016
rect 12376 5952 12384 6016
rect 12064 4928 12384 5952
rect 12064 4864 12072 4928
rect 12136 4864 12152 4928
rect 12216 4864 12232 4928
rect 12296 4864 12312 4928
rect 12376 4864 12384 4928
rect 11835 4860 11901 4861
rect 11835 4796 11836 4860
rect 11900 4796 11901 4860
rect 11835 4795 11901 4796
rect 12064 3840 12384 4864
rect 12758 4453 12818 6835
rect 12942 4453 13002 12003
rect 13491 11932 13557 11933
rect 13491 11868 13492 11932
rect 13556 11868 13557 11932
rect 13491 11867 13557 11868
rect 12755 4452 12821 4453
rect 12755 4388 12756 4452
rect 12820 4388 12821 4452
rect 12755 4387 12821 4388
rect 12939 4452 13005 4453
rect 12939 4388 12940 4452
rect 13004 4388 13005 4452
rect 12939 4387 13005 4388
rect 12064 3776 12072 3840
rect 12136 3776 12152 3840
rect 12216 3776 12232 3840
rect 12296 3776 12312 3840
rect 12376 3776 12384 3840
rect 12064 2752 12384 3776
rect 12064 2688 12072 2752
rect 12136 2688 12152 2752
rect 12216 2688 12232 2752
rect 12296 2688 12312 2752
rect 12376 2688 12384 2752
rect 11651 2412 11717 2413
rect 11651 2348 11652 2412
rect 11716 2348 11717 2412
rect 11651 2347 11717 2348
rect 9840 2144 9848 2208
rect 9912 2144 9928 2208
rect 9992 2144 10008 2208
rect 10072 2144 10088 2208
rect 10152 2144 10160 2208
rect 9840 2128 10160 2144
rect 12064 2128 12384 2688
rect 13494 2685 13554 11867
rect 13491 2684 13557 2685
rect 13491 2620 13492 2684
rect 13556 2620 13557 2684
rect 13491 2619 13557 2620
rect 13678 2549 13738 14995
rect 14288 14176 14608 14736
rect 14288 14112 14296 14176
rect 14360 14112 14376 14176
rect 14440 14112 14456 14176
rect 14520 14112 14536 14176
rect 14600 14112 14608 14176
rect 13859 13836 13925 13837
rect 13859 13772 13860 13836
rect 13924 13772 13925 13836
rect 13859 13771 13925 13772
rect 13862 3229 13922 13771
rect 14288 13088 14608 14112
rect 14288 13024 14296 13088
rect 14360 13024 14376 13088
rect 14440 13024 14456 13088
rect 14520 13024 14536 13088
rect 14600 13024 14608 13088
rect 14288 12000 14608 13024
rect 14288 11936 14296 12000
rect 14360 11936 14376 12000
rect 14440 11936 14456 12000
rect 14520 11936 14536 12000
rect 14600 11936 14608 12000
rect 14043 11252 14109 11253
rect 14043 11188 14044 11252
rect 14108 11188 14109 11252
rect 14043 11187 14109 11188
rect 14046 3229 14106 11187
rect 14288 10912 14608 11936
rect 16512 14720 16832 14736
rect 16512 14656 16520 14720
rect 16584 14656 16600 14720
rect 16664 14656 16680 14720
rect 16744 14656 16760 14720
rect 16824 14656 16832 14720
rect 16512 13632 16832 14656
rect 16512 13568 16520 13632
rect 16584 13568 16600 13632
rect 16664 13568 16680 13632
rect 16744 13568 16760 13632
rect 16824 13568 16832 13632
rect 16512 12544 16832 13568
rect 16512 12480 16520 12544
rect 16584 12480 16600 12544
rect 16664 12480 16680 12544
rect 16744 12480 16760 12544
rect 16824 12480 16832 12544
rect 16512 11456 16832 12480
rect 16512 11392 16520 11456
rect 16584 11392 16600 11456
rect 16664 11392 16680 11456
rect 16744 11392 16760 11456
rect 16824 11392 16832 11456
rect 16251 11252 16317 11253
rect 16251 11188 16252 11252
rect 16316 11188 16317 11252
rect 16251 11187 16317 11188
rect 14288 10848 14296 10912
rect 14360 10848 14376 10912
rect 14440 10848 14456 10912
rect 14520 10848 14536 10912
rect 14600 10848 14608 10912
rect 14288 9824 14608 10848
rect 14963 10300 15029 10301
rect 14963 10236 14964 10300
rect 15028 10236 15029 10300
rect 14963 10235 15029 10236
rect 14288 9760 14296 9824
rect 14360 9760 14376 9824
rect 14440 9760 14456 9824
rect 14520 9760 14536 9824
rect 14600 9760 14608 9824
rect 14288 8736 14608 9760
rect 14288 8672 14296 8736
rect 14360 8672 14376 8736
rect 14440 8672 14456 8736
rect 14520 8672 14536 8736
rect 14600 8672 14608 8736
rect 14288 7648 14608 8672
rect 14288 7584 14296 7648
rect 14360 7584 14376 7648
rect 14440 7584 14456 7648
rect 14520 7584 14536 7648
rect 14600 7584 14608 7648
rect 14288 6560 14608 7584
rect 14288 6496 14296 6560
rect 14360 6496 14376 6560
rect 14440 6496 14456 6560
rect 14520 6496 14536 6560
rect 14600 6496 14608 6560
rect 14288 5472 14608 6496
rect 14288 5408 14296 5472
rect 14360 5408 14376 5472
rect 14440 5408 14456 5472
rect 14520 5408 14536 5472
rect 14600 5408 14608 5472
rect 14288 4384 14608 5408
rect 14288 4320 14296 4384
rect 14360 4320 14376 4384
rect 14440 4320 14456 4384
rect 14520 4320 14536 4384
rect 14600 4320 14608 4384
rect 14288 3296 14608 4320
rect 14288 3232 14296 3296
rect 14360 3232 14376 3296
rect 14440 3232 14456 3296
rect 14520 3232 14536 3296
rect 14600 3232 14608 3296
rect 13859 3228 13925 3229
rect 13859 3164 13860 3228
rect 13924 3164 13925 3228
rect 13859 3163 13925 3164
rect 14043 3228 14109 3229
rect 14043 3164 14044 3228
rect 14108 3164 14109 3228
rect 14043 3163 14109 3164
rect 13675 2548 13741 2549
rect 13675 2484 13676 2548
rect 13740 2484 13741 2548
rect 13675 2483 13741 2484
rect 14288 2208 14608 3232
rect 14966 2549 15026 10235
rect 16254 7717 16314 11187
rect 16512 10368 16832 11392
rect 17907 11116 17973 11117
rect 17907 11052 17908 11116
rect 17972 11052 17973 11116
rect 17907 11051 17973 11052
rect 16512 10304 16520 10368
rect 16584 10304 16600 10368
rect 16664 10304 16680 10368
rect 16744 10304 16760 10368
rect 16824 10304 16832 10368
rect 16512 9280 16832 10304
rect 16987 10164 17053 10165
rect 16987 10100 16988 10164
rect 17052 10100 17053 10164
rect 16987 10099 17053 10100
rect 16512 9216 16520 9280
rect 16584 9216 16600 9280
rect 16664 9216 16680 9280
rect 16744 9216 16760 9280
rect 16824 9216 16832 9280
rect 16512 8192 16832 9216
rect 16512 8128 16520 8192
rect 16584 8128 16600 8192
rect 16664 8128 16680 8192
rect 16744 8128 16760 8192
rect 16824 8128 16832 8192
rect 15883 7716 15949 7717
rect 15883 7652 15884 7716
rect 15948 7652 15949 7716
rect 15883 7651 15949 7652
rect 16251 7716 16317 7717
rect 16251 7652 16252 7716
rect 16316 7652 16317 7716
rect 16251 7651 16317 7652
rect 15886 5541 15946 7651
rect 15883 5540 15949 5541
rect 15883 5476 15884 5540
rect 15948 5476 15949 5540
rect 15883 5475 15949 5476
rect 15886 2685 15946 5475
rect 16254 2957 16314 7651
rect 16512 7104 16832 8128
rect 16512 7040 16520 7104
rect 16584 7040 16600 7104
rect 16664 7040 16680 7104
rect 16744 7040 16760 7104
rect 16824 7040 16832 7104
rect 16512 6016 16832 7040
rect 16512 5952 16520 6016
rect 16584 5952 16600 6016
rect 16664 5952 16680 6016
rect 16744 5952 16760 6016
rect 16824 5952 16832 6016
rect 16512 4928 16832 5952
rect 16990 5541 17050 10099
rect 17910 9485 17970 11051
rect 17907 9484 17973 9485
rect 17907 9420 17908 9484
rect 17972 9420 17973 9484
rect 17907 9419 17973 9420
rect 17355 8124 17421 8125
rect 17355 8060 17356 8124
rect 17420 8060 17421 8124
rect 17355 8059 17421 8060
rect 16987 5540 17053 5541
rect 16987 5476 16988 5540
rect 17052 5476 17053 5540
rect 16987 5475 17053 5476
rect 16512 4864 16520 4928
rect 16584 4864 16600 4928
rect 16664 4864 16680 4928
rect 16744 4864 16760 4928
rect 16824 4864 16832 4928
rect 16512 3840 16832 4864
rect 17358 4861 17418 8059
rect 17907 7308 17973 7309
rect 17907 7244 17908 7308
rect 17972 7244 17973 7308
rect 17907 7243 17973 7244
rect 17355 4860 17421 4861
rect 17355 4796 17356 4860
rect 17420 4796 17421 4860
rect 17355 4795 17421 4796
rect 17910 4317 17970 7243
rect 17907 4316 17973 4317
rect 17907 4252 17908 4316
rect 17972 4252 17973 4316
rect 17907 4251 17973 4252
rect 16512 3776 16520 3840
rect 16584 3776 16600 3840
rect 16664 3776 16680 3840
rect 16744 3776 16760 3840
rect 16824 3776 16832 3840
rect 16251 2956 16317 2957
rect 16251 2892 16252 2956
rect 16316 2892 16317 2956
rect 16251 2891 16317 2892
rect 16512 2752 16832 3776
rect 16512 2688 16520 2752
rect 16584 2688 16600 2752
rect 16664 2688 16680 2752
rect 16744 2688 16760 2752
rect 16824 2688 16832 2752
rect 15883 2684 15949 2685
rect 15883 2620 15884 2684
rect 15948 2620 15949 2684
rect 15883 2619 15949 2620
rect 14963 2548 15029 2549
rect 14963 2484 14964 2548
rect 15028 2484 15029 2548
rect 14963 2483 15029 2484
rect 14288 2144 14296 2208
rect 14360 2144 14376 2208
rect 14440 2144 14456 2208
rect 14520 2144 14536 2208
rect 14600 2144 14608 2208
rect 14288 2128 14608 2144
rect 16512 2128 16832 2688
use sky130_fd_sc_hd__diode_2  ANTENNA__39__A dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 4416 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__40__A
timestamp 1649977179
transform 1 0 4232 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__41__A
timestamp 1649977179
transform 1 0 4048 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__42__A
timestamp 1649977179
transform -1 0 4508 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__43__A
timestamp 1649977179
transform -1 0 3772 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__44__A
timestamp 1649977179
transform 1 0 4416 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__45__A
timestamp 1649977179
transform -1 0 5060 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__46__A
timestamp 1649977179
transform -1 0 3956 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__48__A
timestamp 1649977179
transform -1 0 3312 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__49__A
timestamp 1649977179
transform 1 0 5060 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__50__A
timestamp 1649977179
transform -1 0 4600 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__52__A
timestamp 1649977179
transform 1 0 3864 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__53__A
timestamp 1649977179
transform 1 0 4692 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__61__A
timestamp 1649977179
transform -1 0 13524 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__62__A
timestamp 1649977179
transform -1 0 13616 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__63__A
timestamp 1649977179
transform -1 0 12788 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__64__A
timestamp 1649977179
transform -1 0 12604 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__65__A
timestamp 1649977179
transform 1 0 13616 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__66__A
timestamp 1649977179
transform 1 0 12420 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__68__A
timestamp 1649977179
transform -1 0 13616 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__69__A
timestamp 1649977179
transform 1 0 15824 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__70__A
timestamp 1649977179
transform -1 0 12972 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__71__A
timestamp 1649977179
transform 1 0 11868 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__72__A
timestamp 1649977179
transform -1 0 12788 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__73__A
timestamp 1649977179
transform 1 0 15456 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__74__A
timestamp 1649977179
transform -1 0 13708 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clk_1_N_FTB01_A
timestamp 1649977179
transform 1 0 4968 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clk_1_S_FTB01_A
timestamp 1649977179
transform -1 0 13340 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clk_2_E_FTB01_A
timestamp 1649977179
transform -1 0 13892 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clk_2_W_FTB01_A
timestamp 1649977179
transform 1 0 5152 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clk_3_E_FTB01_A
timestamp 1649977179
transform -1 0 14076 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clk_3_W_FTB01_A
timestamp 1649977179
transform -1 0 5060 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1649977179
transform -1 0 5796 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1649977179
transform -1 0 12880 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1649977179
transform -1 0 5152 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1649977179
transform -1 0 4324 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1649977179
transform -1 0 4324 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1649977179
transform -1 0 5888 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1649977179
transform -1 0 1564 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1649977179
transform -1 0 5152 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1649977179
transform -1 0 3404 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1649977179
transform -1 0 5244 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1649977179
transform -1 0 6348 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1649977179
transform -1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1649977179
transform -1 0 6164 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1649977179
transform -1 0 5980 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1649977179
transform -1 0 5980 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1649977179
transform -1 0 4692 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1649977179
transform -1 0 3404 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1649977179
transform -1 0 1564 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1649977179
transform -1 0 5152 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1649977179
transform -1 0 6532 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1649977179
transform -1 0 3680 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1649977179
transform -1 0 6256 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1649977179
transform -1 0 5704 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1649977179
transform -1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1649977179
transform -1 0 13984 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1649977179
transform -1 0 9936 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1649977179
transform -1 0 8832 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1649977179
transform -1 0 14352 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1649977179
transform -1 0 16560 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1649977179
transform -1 0 16836 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1649977179
transform -1 0 14260 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1649977179
transform -1 0 18216 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1649977179
transform -1 0 13524 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1649977179
transform -1 0 11040 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1649977179
transform -1 0 12052 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1649977179
transform -1 0 15824 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1649977179
transform -1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1649977179
transform -1 0 17664 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1649977179
transform -1 0 14536 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1649977179
transform -1 0 13984 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1649977179
transform -1 0 14444 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1649977179
transform -1 0 11960 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1649977179
transform -1 0 11408 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1649977179
transform -1 0 14260 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1649977179
transform -1 0 5704 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1649977179
transform -1 0 5520 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1649977179
transform -1 0 5612 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1649977179
transform -1 0 5520 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1649977179
transform -1 0 5336 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1649977179
transform -1 0 5704 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform -1 0 13708 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1649977179
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1649977179
transform 1 0 12972 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform -1 0 15732 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1649977179
transform 1 0 13156 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0__S
timestamp 1649977179
transform -1 0 3588 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1__S
timestamp 1649977179
transform 1 0 3680 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 3588 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_2__S
timestamp 1649977179
transform 1 0 3772 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 4048 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 4876 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 5244 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_0__S
timestamp 1649977179
transform -1 0 4140 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_1__S
timestamp 1649977179
transform -1 0 3680 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 3496 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 4232 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 3312 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l4_in_0__S
timestamp 1649977179
transform -1 0 3956 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 8740 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 6808 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 8004 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 8464 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 2668 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 5704 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 5428 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_2__A0
timestamp 1649977179
transform -1 0 5796 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 5428 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0__S
timestamp 1649977179
transform -1 0 6532 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1__S
timestamp 1649977179
transform -1 0 5428 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 6440 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_2__S
timestamp 1649977179
transform -1 0 6716 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 4692 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 7820 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 6808 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 8556 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_0__S
timestamp 1649977179
transform 1 0 5520 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 4692 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_1__S
timestamp 1649977179
transform 1 0 5704 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 4508 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_2__S
timestamp 1649977179
transform 1 0 4784 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 6808 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_3__S
timestamp 1649977179
transform -1 0 6808 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 9568 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 6624 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 6900 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 7820 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 5336 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 4600 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 3680 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 3404 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 5520 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 7084 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 6072 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 5152 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 6440 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_2__A0
timestamp 1649977179
transform -1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 14168 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 14352 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_2__A0
timestamp 1649977179
transform -1 0 14260 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_2__A1
timestamp 1649977179
transform -1 0 13984 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 12052 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 9292 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 11592 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 11684 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 15180 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 16008 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 12788 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 16008 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_2__A1
timestamp 1649977179
transform -1 0 16836 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 14720 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 15364 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_2__A0
timestamp 1649977179
transform -1 0 18584 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 13432 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 14812 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 13248 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 12052 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_2__A1
timestamp 1649977179
transform -1 0 13616 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output52_A
timestamp 1649977179
transform 1 0 12512 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1649977179
transform -1 0 11868 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_W_FTB01_A
timestamp 1649977179
transform 1 0 16376 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_1_N_FTB01_A
timestamp 1649977179
transform 1 0 13616 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_1_S_FTB01_A
timestamp 1649977179
transform 1 0 13248 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_2_E_FTB01_A
timestamp 1649977179
transform -1 0 13156 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_2_W_FTB01_A
timestamp 1649977179
transform 1 0 3496 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_3_E_FTB01_A
timestamp 1649977179
transform 1 0 10764 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_3_W_FTB01_A
timestamp 1649977179
transform 1 0 5060 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2852 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp 1649977179
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 4324 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 4968 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46
timestamp 1649977179
transform 1 0 5336 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51
timestamp 1649977179
transform 1 0 5796 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55
timestamp 1649977179
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61
timestamp 1649977179
transform 1 0 6716 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69
timestamp 1649977179
transform 1 0 7452 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73
timestamp 1649977179
transform 1 0 7820 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 8280 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_89
timestamp 1649977179
transform 1 0 9292 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_96
timestamp 1649977179
transform 1 0 9936 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100
timestamp 1649977179
transform 1 0 10304 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_105
timestamp 1649977179
transform 1 0 10764 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1649977179
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_117 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 11868 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_123
timestamp 1649977179
transform 1 0 12420 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_145
timestamp 1649977179
transform 1 0 14444 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_150
timestamp 1649977179
transform 1 0 14904 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_169
timestamp 1649977179
transform 1 0 16652 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_177
timestamp 1649977179
transform 1 0 17388 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_31 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_43
timestamp 1649977179
transform 1 0 5060 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_1_49
timestamp 1649977179
transform 1 0 5612 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1649977179
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_57
timestamp 1649977179
transform 1 0 6348 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_63
timestamp 1649977179
transform 1 0 6900 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_70
timestamp 1649977179
transform 1 0 7544 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_82
timestamp 1649977179
transform 1 0 8648 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_94
timestamp 1649977179
transform 1 0 9752 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_106
timestamp 1649977179
transform 1 0 10856 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_119
timestamp 1649977179
transform 1 0 12052 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_146
timestamp 1649977179
transform 1 0 14536 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_152
timestamp 1649977179
transform 1 0 15088 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1649977179
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_36
timestamp 1649977179
transform 1 0 4416 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_48
timestamp 1649977179
transform 1 0 5520 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_63
timestamp 1649977179
transform 1 0 6900 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_69
timestamp 1649977179
transform 1 0 7452 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_76 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 8096 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_97
timestamp 1649977179
transform 1 0 10028 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_110
timestamp 1649977179
transform 1 0 11224 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_122
timestamp 1649977179
transform 1 0 12328 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_141
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_160
timestamp 1649977179
transform 1 0 15824 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_38
timestamp 1649977179
transform 1 0 4600 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_50
timestamp 1649977179
transform 1 0 5704 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_61
timestamp 1649977179
transform 1 0 6716 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_77
timestamp 1649977179
transform 1 0 8188 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_80
timestamp 1649977179
transform 1 0 8464 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_94
timestamp 1649977179
transform 1 0 9752 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_98
timestamp 1649977179
transform 1 0 10120 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_106
timestamp 1649977179
transform 1 0 10856 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_116
timestamp 1649977179
transform 1 0 11776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_169
timestamp 1649977179
transform 1 0 16652 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_41
timestamp 1649977179
transform 1 0 4876 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_45
timestamp 1649977179
transform 1 0 5244 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1649977179
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_85
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_113
timestamp 1649977179
transform 1 0 11500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_119
timestamp 1649977179
transform 1 0 12052 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_177
timestamp 1649977179
transform 1 0 17388 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_7
timestamp 1649977179
transform 1 0 1748 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_38
timestamp 1649977179
transform 1 0 4600 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_82
timestamp 1649977179
transform 1 0 8648 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_101
timestamp 1649977179
transform 1 0 10396 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1649977179
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_155
timestamp 1649977179
transform 1 0 15364 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_38
timestamp 1649977179
transform 1 0 4600 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_57
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_98
timestamp 1649977179
transform 1 0 10120 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1649977179
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_62
timestamp 1649977179
transform 1 0 6808 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1649977179
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_88
timestamp 1649977179
transform 1 0 9200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1649977179
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_141
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_57
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_125
timestamp 1649977179
transform 1 0 12604 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_38
timestamp 1649977179
transform 1 0 4600 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_114
timestamp 1649977179
transform 1 0 11592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_136
timestamp 1649977179
transform 1 0 13616 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_150
timestamp 1649977179
transform 1 0 14904 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_185
timestamp 1649977179
transform 1 0 18124 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_27
timestamp 1649977179
transform 1 0 3588 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1649977179
transform 1 0 6532 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_79
timestamp 1649977179
transform 1 0 8372 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_125
timestamp 1649977179
transform 1 0 12604 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_169
timestamp 1649977179
transform 1 0 16652 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_44
timestamp 1649977179
transform 1 0 5152 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_67
timestamp 1649977179
transform 1 0 7268 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_117
timestamp 1649977179
transform 1 0 11868 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_189
timestamp 1649977179
transform 1 0 18492 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_52
timestamp 1649977179
transform 1 0 5888 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_66
timestamp 1649977179
transform 1 0 7176 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_90
timestamp 1649977179
transform 1 0 9384 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_94
timestamp 1649977179
transform 1 0 9752 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1649977179
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_25
timestamp 1649977179
transform 1 0 3404 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_29
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_64
timestamp 1649977179
transform 1 0 6992 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_97
timestamp 1649977179
transform 1 0 10028 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_114
timestamp 1649977179
transform 1 0 11592 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_141
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_17
timestamp 1649977179
transform 1 0 2668 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_66
timestamp 1649977179
transform 1 0 7176 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_74
timestamp 1649977179
transform 1 0 7912 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_91
timestamp 1649977179
transform 1 0 9476 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_95
timestamp 1649977179
transform 1 0 9844 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_113
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_121
timestamp 1649977179
transform 1 0 12236 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_31
timestamp 1649977179
transform 1 0 3956 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_45
timestamp 1649977179
transform 1 0 5244 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_57
timestamp 1649977179
transform 1 0 6348 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_69
timestamp 1649977179
transform 1 0 7452 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_81
timestamp 1649977179
transform 1 0 8556 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_101
timestamp 1649977179
transform 1 0 10396 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_105
timestamp 1649977179
transform 1 0 10764 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1649977179
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_57
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_65
timestamp 1649977179
transform 1 0 7084 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_98
timestamp 1649977179
transform 1 0 10120 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1649977179
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_115
timestamp 1649977179
transform 1 0 11684 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1649977179
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_185
timestamp 1649977179
transform 1 0 18124 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_55
timestamp 1649977179
transform 1 0 6164 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_67
timestamp 1649977179
transform 1 0 7268 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_79
timestamp 1649977179
transform 1 0 8372 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1649977179
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_137
timestamp 1649977179
transform 1 0 13708 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_157
timestamp 1649977179
transform 1 0 15548 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_175
timestamp 1649977179
transform 1 0 17204 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_53
timestamp 1649977179
transform 1 0 5980 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_69
timestamp 1649977179
transform 1 0 7452 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_75
timestamp 1649977179
transform 1 0 8004 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_108
timestamp 1649977179
transform 1 0 11040 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_185
timestamp 1649977179
transform 1 0 18124 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_40
timestamp 1649977179
transform 1 0 4784 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_49
timestamp 1649977179
transform 1 0 5612 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_61
timestamp 1649977179
transform 1 0 6716 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_67
timestamp 1649977179
transform 1 0 7268 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_97
timestamp 1649977179
transform 1 0 10028 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_50
timestamp 1649977179
transform 1 0 5704 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_57
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_61
timestamp 1649977179
transform 1 0 6716 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_129
timestamp 1649977179
transform 1 0 12972 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_185
timestamp 1649977179
transform 1 0 18124 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1649977179
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_50
timestamp 1649977179
transform 1 0 5704 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_61
timestamp 1649977179
transform 1 0 6716 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_73
timestamp 1649977179
transform 1 0 7820 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_81
timestamp 1649977179
transform 1 0 8556 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_105
timestamp 1649977179
transform 1 0 10764 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_129
timestamp 1649977179
transform 1 0 12972 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_143
timestamp 1649977179
transform 1 0 14260 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_185
timestamp 1649977179
transform 1 0 18124 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 18860 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 18860 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 18860 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 18860 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 18860 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 18860 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 18860 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 18860 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 18860 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 18860 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 18860 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 18860 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1649977179
transform 1 0 6256 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1649977179
transform 1 0 11408 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1649977179
transform 1 0 16560 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _32_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 3496 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _33_
timestamp 1649977179
transform -1 0 3404 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _34_
timestamp 1649977179
transform 1 0 11776 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _35_
timestamp 1649977179
transform 1 0 2944 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _36_
timestamp 1649977179
transform 1 0 3036 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _37_
timestamp 1649977179
transform 1 0 2852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _38_
timestamp 1649977179
transform 1 0 2852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _39_
timestamp 1649977179
transform 1 0 3128 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _40_
timestamp 1649977179
transform 1 0 2392 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _41_
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _42_
timestamp 1649977179
transform 1 0 1748 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _43_
timestamp 1649977179
transform 1 0 2668 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _44_
timestamp 1649977179
transform 1 0 2760 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _45_
timestamp 1649977179
transform 1 0 4324 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _46_
timestamp 1649977179
transform 1 0 2116 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _47_
timestamp 1649977179
transform 1 0 3404 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _48_
timestamp 1649977179
transform 1 0 2484 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _49_
timestamp 1649977179
transform 1 0 3956 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _50_
timestamp 1649977179
transform 1 0 4048 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _51_
timestamp 1649977179
transform 1 0 3496 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _52_
timestamp 1649977179
transform 1 0 3312 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _53_
timestamp 1649977179
transform 1 0 3036 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _54_
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _55_
timestamp 1649977179
transform -1 0 16560 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _56_
timestamp 1649977179
transform -1 0 17020 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _57_
timestamp 1649977179
transform -1 0 14444 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _58_
timestamp 1649977179
transform -1 0 14720 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _59_
timestamp 1649977179
transform -1 0 15824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _60_
timestamp 1649977179
transform -1 0 15364 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _61_
timestamp 1649977179
transform -1 0 15548 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _62_
timestamp 1649977179
transform -1 0 16284 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _63_
timestamp 1649977179
transform -1 0 16560 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _64_
timestamp 1649977179
transform -1 0 17112 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _65_
timestamp 1649977179
transform -1 0 13984 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _66_
timestamp 1649977179
transform -1 0 16468 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _67_
timestamp 1649977179
transform -1 0 11408 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _68_
timestamp 1649977179
transform -1 0 13708 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _69_
timestamp 1649977179
transform -1 0 16284 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _70_
timestamp 1649977179
transform 1 0 16468 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _71_
timestamp 1649977179
transform 1 0 18308 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _72_
timestamp 1649977179
transform 1 0 18308 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _73_
timestamp 1649977179
transform -1 0 17664 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _74_
timestamp 1649977179
transform 1 0 18308 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clk_1_N_FTB01
timestamp 1649977179
transform -1 0 4968 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clk_1_S_FTB01
timestamp 1649977179
transform -1 0 15456 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clk_2_E_FTB01
timestamp 1649977179
transform -1 0 15272 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clk_2_W_FTB01
timestamp 1649977179
transform 1 0 4416 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clk_3_E_FTB01
timestamp 1649977179
transform -1 0 14996 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clk_3_W_FTB01
timestamp 1649977179
transform 1 0 5060 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1649977179
transform 1 0 5336 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1649977179
transform 1 0 16008 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1649977179
transform 1 0 4692 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1649977179
transform -1 0 3588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1649977179
transform -1 0 4048 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input6 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 2300 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input7
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input8
timestamp 1649977179
transform -1 0 2300 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input9 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2300 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 1649977179
transform 1 0 2300 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input11
timestamp 1649977179
transform -1 0 2300 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input12
timestamp 1649977179
transform -1 0 2300 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input13
timestamp 1649977179
transform -1 0 2300 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input14
timestamp 1649977179
transform -1 0 2300 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input15
timestamp 1649977179
transform -1 0 3220 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1649977179
transform -1 0 3496 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1649977179
transform -1 0 2944 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1649977179
transform -1 0 3496 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input19
timestamp 1649977179
transform -1 0 3220 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input20
timestamp 1649977179
transform -1 0 2300 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp 1649977179
transform 1 0 3128 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input22
timestamp 1649977179
transform -1 0 2300 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input23
timestamp 1649977179
transform -1 0 3220 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input24
timestamp 1649977179
transform -1 0 2300 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input25
timestamp 1649977179
transform -1 0 18584 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input26
timestamp 1649977179
transform -1 0 18584 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input27
timestamp 1649977179
transform -1 0 18584 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input28
timestamp 1649977179
transform 1 0 17664 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input29
timestamp 1649977179
transform -1 0 14996 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input30
timestamp 1649977179
transform -1 0 17664 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input31
timestamp 1649977179
transform -1 0 13984 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input32
timestamp 1649977179
transform -1 0 17296 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input33
timestamp 1649977179
transform -1 0 13340 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input34
timestamp 1649977179
transform -1 0 11408 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input35
timestamp 1649977179
transform -1 0 12420 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1649977179
transform -1 0 16560 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1649977179
transform 1 0 17940 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1649977179
transform 1 0 16652 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input39
timestamp 1649977179
transform 1 0 17664 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input40
timestamp 1649977179
transform -1 0 18584 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input41
timestamp 1649977179
transform 1 0 17664 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input42
timestamp 1649977179
transform 1 0 17664 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input43
timestamp 1649977179
transform -1 0 18584 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input44
timestamp 1649977179
transform -1 0 17664 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input45
timestamp 1649977179
transform -1 0 2300 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input46
timestamp 1649977179
transform -1 0 3220 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input47
timestamp 1649977179
transform -1 0 2300 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input48
timestamp 1649977179
transform -1 0 3220 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input49
timestamp 1649977179
transform -1 0 4692 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input50
timestamp 1649977179
transform -1 0 2300 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 11500 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 13524 0 -1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 7176 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 15548 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 8832 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 11408 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 9936 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 11408 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 16376 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 9568 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 11684 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 11868 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 10396 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 13984 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 9384 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 8648 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 9568 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 16560 0 -1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 12972 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 7360 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 11960 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 13064 0 -1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 15548 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 9936 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 17204 0 1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 10396 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 12052 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 15916 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 12972 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 12972 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 8004 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 11960 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 13984 0 1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 12328 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 11408 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 7360 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 16008 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 15456 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 17020 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 16652 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 17388 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 16468 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 17480 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 11500 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 6808 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 10120 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 15548 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 17204 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 18124 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 16468 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14536 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 16652 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 16376 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 14168 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 12328 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 14996 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 13524 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 16468 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 14904 0 -1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 8280 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 10396 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1840 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_1_
timestamp 1649977179
transform 1 0 2392 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_2_
timestamp 1649977179
transform 1 0 2392 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 1564 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_1_
timestamp 1649977179
transform -1 0 2300 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_2_
timestamp 1649977179
transform 1 0 4416 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_0.mux_l2_in_3__145 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3588 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_3_
timestamp 1649977179
transform 1 0 2852 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_0_
timestamp 1649977179
transform -1 0 2392 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_1_
timestamp 1649977179
transform 1 0 2300 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l4_in_0_
timestamp 1649977179
transform -1 0 3128 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 3404 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l1_in_0_
timestamp 1649977179
transform 1 0 4692 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_0_
timestamp 1649977179
transform 1 0 4600 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_1_
timestamp 1649977179
transform 1 0 4048 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_2_
timestamp 1649977179
transform -1 0 3680 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_1.mux_l2_in_3__146
timestamp 1649977179
transform 1 0 3128 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_3_
timestamp 1649977179
transform -1 0 2852 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_0_
timestamp 1649977179
transform 1 0 3772 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_1_
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l4_in_0_
timestamp 1649977179
transform -1 0 3772 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 3588 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l1_in_0_
timestamp 1649977179
transform -1 0 9936 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_0_
timestamp 1649977179
transform 1 0 9568 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_1_
timestamp 1649977179
transform 1 0 9016 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_2_
timestamp 1649977179
transform -1 0 7820 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_2.mux_l2_in_3__153
timestamp 1649977179
transform 1 0 8280 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_3_
timestamp 1649977179
transform 1 0 7452 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_0_
timestamp 1649977179
transform 1 0 8924 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_1_
timestamp 1649977179
transform 1 0 6992 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l4_in_0_
timestamp 1649977179
transform 1 0 6624 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 5336 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_0_
timestamp 1649977179
transform -1 0 3128 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_1_
timestamp 1649977179
transform -1 0 3128 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_2_
timestamp 1649977179
transform -1 0 3128 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_0_
timestamp 1649977179
transform 1 0 4692 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_1_
timestamp 1649977179
transform -1 0 3128 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_2_
timestamp 1649977179
transform -1 0 4600 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_3_
timestamp 1649977179
transform -1 0 4048 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_3.mux_l2_in_3__154
timestamp 1649977179
transform 1 0 4508 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_0_
timestamp 1649977179
transform 1 0 4600 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_1_
timestamp 1649977179
transform 1 0 3956 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l4_in_0_
timestamp 1649977179
transform -1 0 3956 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 5244 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_0_
timestamp 1649977179
transform 1 0 5612 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_1_
timestamp 1649977179
transform 1 0 5428 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_2_
timestamp 1649977179
transform -1 0 6532 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_0_
timestamp 1649977179
transform -1 0 5704 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_1_
timestamp 1649977179
transform 1 0 5704 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_2_
timestamp 1649977179
transform 1 0 8004 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_4.mux_l2_in_3__155
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_3_
timestamp 1649977179
transform -1 0 8464 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_0_
timestamp 1649977179
transform -1 0 6256 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_1_
timestamp 1649977179
transform 1 0 7820 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l4_in_0_
timestamp 1649977179
transform -1 0 7820 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 7268 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l1_in_0_
timestamp 1649977179
transform 1 0 5244 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_0_
timestamp 1649977179
transform 1 0 4692 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_1_
timestamp 1649977179
transform 1 0 4876 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_2_
timestamp 1649977179
transform -1 0 4600 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_5.mux_l2_in_3__140
timestamp 1649977179
transform -1 0 6716 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_3_
timestamp 1649977179
transform 1 0 6808 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_0_
timestamp 1649977179
transform -1 0 5428 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_1_
timestamp 1649977179
transform -1 0 6256 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l4_in_0_
timestamp 1649977179
transform -1 0 6348 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 7268 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l1_in_0_
timestamp 1649977179
transform 1 0 8924 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_0_
timestamp 1649977179
transform -1 0 8832 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_1_
timestamp 1649977179
transform 1 0 9752 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_2_
timestamp 1649977179
transform 1 0 8096 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_6.mux_l2_in_3__141
timestamp 1649977179
transform -1 0 8096 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_3_
timestamp 1649977179
transform 1 0 7912 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l3_in_0_
timestamp 1649977179
transform 1 0 9476 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l3_in_1_
timestamp 1649977179
transform 1 0 7176 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l4_in_0_
timestamp 1649977179
transform -1 0 7176 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 7820 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_0_
timestamp 1649977179
transform -1 0 4508 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_1_
timestamp 1649977179
transform -1 0 4508 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_2_
timestamp 1649977179
transform 1 0 4508 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_0_
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_1_
timestamp 1649977179
transform 1 0 4140 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_2_
timestamp 1649977179
transform -1 0 4692 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_3_
timestamp 1649977179
transform -1 0 3588 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_7.mux_l2_in_3__142
timestamp 1649977179
transform 1 0 3864 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l3_in_0_
timestamp 1649977179
transform -1 0 4416 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l3_in_1_
timestamp 1649977179
transform -1 0 4876 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l4_in_0_
timestamp 1649977179
transform -1 0 6164 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 6900 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_0_
timestamp 1649977179
transform -1 0 7820 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_1_
timestamp 1649977179
transform -1 0 7544 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_2_
timestamp 1649977179
transform -1 0 7084 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_0_
timestamp 1649977179
transform 1 0 7544 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_1_
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_2_
timestamp 1649977179
transform -1 0 6256 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_8.mux_l2_in_3__143
timestamp 1649977179
transform -1 0 6992 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_3_
timestamp 1649977179
transform 1 0 7084 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l3_in_0_
timestamp 1649977179
transform -1 0 6164 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l3_in_1_
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l4_in_0_
timestamp 1649977179
transform -1 0 6992 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 8096 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l1_in_0_
timestamp 1649977179
transform 1 0 13156 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_0_
timestamp 1649977179
transform -1 0 13156 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_1_
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_2_
timestamp 1649977179
transform -1 0 14168 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_3_
timestamp 1649977179
transform -1 0 13340 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_9.mux_l2_in_3__144
timestamp 1649977179
transform 1 0 12972 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l3_in_0_
timestamp 1649977179
transform 1 0 12972 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l3_in_1_
timestamp 1649977179
transform 1 0 13984 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l4_in_0_
timestamp 1649977179
transform 1 0 12144 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 11132 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l1_in_0_
timestamp 1649977179
transform 1 0 16560 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_0_
timestamp 1649977179
transform -1 0 15732 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_1_
timestamp 1649977179
transform -1 0 16284 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_2_
timestamp 1649977179
transform 1 0 16652 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_3_
timestamp 1649977179
transform 1 0 17572 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_10.mux_l2_in_3__147
timestamp 1649977179
transform -1 0 16192 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l3_in_0_
timestamp 1649977179
transform 1 0 15732 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l3_in_1_
timestamp 1649977179
transform 1 0 15548 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l4_in_0_
timestamp 1649977179
transform 1 0 14720 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_0_
timestamp 1649977179
transform 1 0 9844 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_1_
timestamp 1649977179
transform 1 0 8740 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_2_
timestamp 1649977179
transform 1 0 12236 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_0_
timestamp 1649977179
transform -1 0 9292 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_1_
timestamp 1649977179
transform 1 0 10304 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_2_
timestamp 1649977179
transform 1 0 11408 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_3_
timestamp 1649977179
transform 1 0 10764 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_11.mux_l2_in_3__148
timestamp 1649977179
transform 1 0 12328 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l3_in_0_
timestamp 1649977179
transform -1 0 10120 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l3_in_1_
timestamp 1649977179
transform -1 0 11408 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l4_in_0_
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 11776 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_0_
timestamp 1649977179
transform 1 0 14812 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_1_
timestamp 1649977179
transform 1 0 13984 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_2_
timestamp 1649977179
transform 1 0 16652 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_0_
timestamp 1649977179
transform -1 0 13984 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_1_
timestamp 1649977179
transform -1 0 14904 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_2_
timestamp 1649977179
transform 1 0 17204 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_12.mux_l2_in_3__149
timestamp 1649977179
transform 1 0 13340 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_3_
timestamp 1649977179
transform -1 0 13524 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l3_in_0_
timestamp 1649977179
transform 1 0 14352 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l3_in_1_
timestamp 1649977179
transform 1 0 13524 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l4_in_0_
timestamp 1649977179
transform 1 0 13064 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 12512 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l1_in_0_
timestamp 1649977179
transform -1 0 17296 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_0_
timestamp 1649977179
transform 1 0 17480 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_1_
timestamp 1649977179
transform 1 0 17480 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_2_
timestamp 1649977179
transform 1 0 15824 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_3_
timestamp 1649977179
transform 1 0 15824 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_13.mux_l2_in_3__150
timestamp 1649977179
transform 1 0 16284 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l3_in_0_
timestamp 1649977179
transform -1 0 15824 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l3_in_1_
timestamp 1649977179
transform -1 0 15824 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l4_in_0_
timestamp 1649977179
transform 1 0 15640 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 14260 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l1_in_0_
timestamp 1649977179
transform -1 0 17940 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_0_
timestamp 1649977179
transform 1 0 17480 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_1_
timestamp 1649977179
transform 1 0 17480 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_2_
timestamp 1649977179
transform 1 0 17296 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_14.mux_l2_in_3__151
timestamp 1649977179
transform 1 0 18308 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_3_
timestamp 1649977179
transform -1 0 17480 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l3_in_0_
timestamp 1649977179
transform 1 0 15180 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l3_in_1_
timestamp 1649977179
transform 1 0 16652 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l4_in_0_
timestamp 1649977179
transform -1 0 14996 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 14812 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_0_
timestamp 1649977179
transform 1 0 11776 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_1_
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_2_
timestamp 1649977179
transform -1 0 13156 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_0_
timestamp 1649977179
transform -1 0 11316 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_1_
timestamp 1649977179
transform 1 0 12604 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_2_
timestamp 1649977179
transform 1 0 11684 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_15.mux_l2_in_3__152
timestamp 1649977179
transform -1 0 12604 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_3_
timestamp 1649977179
transform 1 0 12512 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l3_in_0_
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l3_in_1_
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l4_in_0_
timestamp 1649977179
transform -1 0 11500 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 12052 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output51 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 3496 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output52
timestamp 1649977179
transform 1 0 17020 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp 1649977179
transform -1 0 6716 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp 1649977179
transform -1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp 1649977179
transform 1 0 12052 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp 1649977179
transform 1 0 12880 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp 1649977179
transform -1 0 14444 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp 1649977179
transform -1 0 14904 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp 1649977179
transform 1 0 15364 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp 1649977179
transform 1 0 3772 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 1649977179
transform -1 0 4968 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp 1649977179
transform 1 0 5428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1649977179
transform -1 0 6716 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1649977179
transform -1 0 7452 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1649977179
transform 1 0 7912 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 1649977179
transform 1 0 9568 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 1649977179
transform -1 0 10764 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1649977179
transform -1 0 2484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1649977179
transform -1 0 2852 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 1649977179
transform -1 0 2852 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1649977179
transform -1 0 2116 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1649977179
transform -1 0 2484 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1649977179
transform -1 0 1748 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1649977179
transform -1 0 3036 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1649977179
transform -1 0 2116 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1649977179
transform -1 0 1748 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1649977179
transform -1 0 1748 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1649977179
transform -1 0 2668 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1649977179
transform -1 0 1748 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1649977179
transform -1 0 2484 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1649977179
transform -1 0 2852 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1649977179
transform -1 0 2116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1649977179
transform -1 0 1748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1649977179
transform -1 0 2116 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1649977179
transform -1 0 1748 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1649977179
transform 1 0 1748 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1649977179
transform -1 0 2484 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1649977179
transform -1 0 1748 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1649977179
transform 1 0 17848 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1649977179
transform 1 0 18216 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1649977179
transform 1 0 17848 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1649977179
transform 1 0 18216 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1649977179
transform 1 0 14168 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1649977179
transform 1 0 16192 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1649977179
transform -1 0 16560 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1649977179
transform -1 0 17112 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1649977179
transform 1 0 18216 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp 1649977179
transform 1 0 18216 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1649977179
transform -1 0 17204 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp 1649977179
transform 1 0 17480 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp 1649977179
transform 1 0 18216 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output104
timestamp 1649977179
transform 1 0 16744 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output105
timestamp 1649977179
transform 1 0 17112 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output106
timestamp 1649977179
transform 1 0 17848 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output107
timestamp 1649977179
transform 1 0 17480 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output108
timestamp 1649977179
transform 1 0 18216 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output109
timestamp 1649977179
transform 1 0 17848 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output110
timestamp 1649977179
transform 1 0 17480 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output111
timestamp 1649977179
transform 1 0 10396 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output112
timestamp 1649977179
transform 1 0 17848 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output113
timestamp 1649977179
transform 1 0 17112 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output114
timestamp 1649977179
transform -1 0 4416 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output115
timestamp 1649977179
transform 1 0 16744 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output116
timestamp 1649977179
transform -1 0 3588 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  output117
timestamp 1649977179
transform 1 0 18308 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output118
timestamp 1649977179
transform 1 0 18216 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output119
timestamp 1649977179
transform 1 0 17480 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output120
timestamp 1649977179
transform 1 0 17480 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output121
timestamp 1649977179
transform 1 0 4140 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output122
timestamp 1649977179
transform 1 0 17112 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output123
timestamp 1649977179
transform -1 0 4140 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 17204 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_W_FTB01 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 14352 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  prog_clk_1_N_FTB01
timestamp 1649977179
transform -1 0 15732 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  prog_clk_1_S_FTB01
timestamp 1649977179
transform -1 0 16008 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  prog_clk_2_E_FTB01
timestamp 1649977179
transform -1 0 16008 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  prog_clk_2_W_FTB01
timestamp 1649977179
transform -1 0 3404 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  prog_clk_3_E_FTB01
timestamp 1649977179
transform -1 0 11224 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  prog_clk_3_W_FTB01
timestamp 1649977179
transform 1 0 4784 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater124
timestamp 1649977179
transform 1 0 10212 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  repeater125
timestamp 1649977179
transform -1 0 6624 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater126
timestamp 1649977179
transform 1 0 6532 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater127
timestamp 1649977179
transform 1 0 14812 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  repeater128
timestamp 1649977179
transform -1 0 10764 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater129
timestamp 1649977179
transform 1 0 16652 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  repeater130
timestamp 1649977179
transform -1 0 10580 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater131
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  repeater132
timestamp 1649977179
transform 1 0 11132 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater133
timestamp 1649977179
transform 1 0 13708 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater134
timestamp 1649977179
transform -1 0 10856 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  repeater135
timestamp 1649977179
transform 1 0 3220 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater136
timestamp 1649977179
transform 1 0 9936 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  repeater137
timestamp 1649977179
transform -1 0 6808 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater138
timestamp 1649977179
transform 1 0 10856 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  repeater139
timestamp 1649977179
transform -1 0 3680 0 -1 9792
box -38 -48 314 592
<< labels >>
flabel metal3 s 0 12656 800 12776 0 FreeSans 480 0 0 0 REGIN_FEEDTHROUGH
port 0 nsew signal input
flabel metal3 s 0 12384 800 12504 0 FreeSans 480 0 0 0 REGOUT_FEEDTHROUGH
port 1 nsew signal tristate
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 SC_IN_BOT
port 2 nsew signal input
flabel metal2 s 2042 16400 2098 17200 0 FreeSans 224 90 0 0 SC_IN_TOP
port 3 nsew signal input
flabel metal2 s 16946 0 17002 800 0 FreeSans 224 90 0 0 SC_OUT_BOT
port 4 nsew signal tristate
flabel metal2 s 5998 16400 6054 17200 0 FreeSans 224 90 0 0 SC_OUT_TOP
port 5 nsew signal tristate
flabel metal4 s 5392 2128 5712 14736 0 FreeSans 1920 90 0 0 VGND
port 6 nsew ground bidirectional
flabel metal4 s 9840 2128 10160 14736 0 FreeSans 1920 90 0 0 VGND
port 6 nsew ground bidirectional
flabel metal4 s 14288 2128 14608 14736 0 FreeSans 1920 90 0 0 VGND
port 6 nsew ground bidirectional
flabel metal4 s 3168 2128 3488 14736 0 FreeSans 1920 90 0 0 VPWR
port 7 nsew power bidirectional
flabel metal4 s 7616 2128 7936 14736 0 FreeSans 1920 90 0 0 VPWR
port 7 nsew power bidirectional
flabel metal4 s 12064 2128 12384 14736 0 FreeSans 1920 90 0 0 VPWR
port 7 nsew power bidirectional
flabel metal4 s 16512 2128 16832 14736 0 FreeSans 1920 90 0 0 VPWR
port 7 nsew power bidirectional
flabel metal2 s 2870 0 2926 800 0 FreeSans 224 90 0 0 bottom_grid_pin_0_
port 8 nsew signal tristate
flabel metal2 s 11150 0 11206 800 0 FreeSans 224 90 0 0 bottom_grid_pin_10_
port 9 nsew signal tristate
flabel metal2 s 11978 0 12034 800 0 FreeSans 224 90 0 0 bottom_grid_pin_11_
port 10 nsew signal tristate
flabel metal2 s 12806 0 12862 800 0 FreeSans 224 90 0 0 bottom_grid_pin_12_
port 11 nsew signal tristate
flabel metal2 s 13634 0 13690 800 0 FreeSans 224 90 0 0 bottom_grid_pin_13_
port 12 nsew signal tristate
flabel metal2 s 14462 0 14518 800 0 FreeSans 224 90 0 0 bottom_grid_pin_14_
port 13 nsew signal tristate
flabel metal2 s 15290 0 15346 800 0 FreeSans 224 90 0 0 bottom_grid_pin_15_
port 14 nsew signal tristate
flabel metal2 s 3698 0 3754 800 0 FreeSans 224 90 0 0 bottom_grid_pin_1_
port 15 nsew signal tristate
flabel metal2 s 4526 0 4582 800 0 FreeSans 224 90 0 0 bottom_grid_pin_2_
port 16 nsew signal tristate
flabel metal2 s 5354 0 5410 800 0 FreeSans 224 90 0 0 bottom_grid_pin_3_
port 17 nsew signal tristate
flabel metal2 s 6182 0 6238 800 0 FreeSans 224 90 0 0 bottom_grid_pin_4_
port 18 nsew signal tristate
flabel metal2 s 7010 0 7066 800 0 FreeSans 224 90 0 0 bottom_grid_pin_5_
port 19 nsew signal tristate
flabel metal2 s 7838 0 7894 800 0 FreeSans 224 90 0 0 bottom_grid_pin_6_
port 20 nsew signal tristate
flabel metal2 s 8666 0 8722 800 0 FreeSans 224 90 0 0 bottom_grid_pin_7_
port 21 nsew signal tristate
flabel metal2 s 9494 0 9550 800 0 FreeSans 224 90 0 0 bottom_grid_pin_8_
port 22 nsew signal tristate
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 bottom_grid_pin_9_
port 23 nsew signal tristate
flabel metal2 s 1214 0 1270 800 0 FreeSans 224 90 0 0 ccff_head
port 24 nsew signal input
flabel metal2 s 2042 0 2098 800 0 FreeSans 224 90 0 0 ccff_tail
port 25 nsew signal tristate
flabel metal3 s 0 6944 800 7064 0 FreeSans 480 0 0 0 chanx_left_in[0]
port 26 nsew signal input
flabel metal3 s 0 9664 800 9784 0 FreeSans 480 0 0 0 chanx_left_in[10]
port 27 nsew signal input
flabel metal3 s 0 9936 800 10056 0 FreeSans 480 0 0 0 chanx_left_in[11]
port 28 nsew signal input
flabel metal3 s 0 10208 800 10328 0 FreeSans 480 0 0 0 chanx_left_in[12]
port 29 nsew signal input
flabel metal3 s 0 10480 800 10600 0 FreeSans 480 0 0 0 chanx_left_in[13]
port 30 nsew signal input
flabel metal3 s 0 10752 800 10872 0 FreeSans 480 0 0 0 chanx_left_in[14]
port 31 nsew signal input
flabel metal3 s 0 11024 800 11144 0 FreeSans 480 0 0 0 chanx_left_in[15]
port 32 nsew signal input
flabel metal3 s 0 11296 800 11416 0 FreeSans 480 0 0 0 chanx_left_in[16]
port 33 nsew signal input
flabel metal3 s 0 11568 800 11688 0 FreeSans 480 0 0 0 chanx_left_in[17]
port 34 nsew signal input
flabel metal3 s 0 11840 800 11960 0 FreeSans 480 0 0 0 chanx_left_in[18]
port 35 nsew signal input
flabel metal3 s 0 12112 800 12232 0 FreeSans 480 0 0 0 chanx_left_in[19]
port 36 nsew signal input
flabel metal3 s 0 7216 800 7336 0 FreeSans 480 0 0 0 chanx_left_in[1]
port 37 nsew signal input
flabel metal3 s 0 7488 800 7608 0 FreeSans 480 0 0 0 chanx_left_in[2]
port 38 nsew signal input
flabel metal3 s 0 7760 800 7880 0 FreeSans 480 0 0 0 chanx_left_in[3]
port 39 nsew signal input
flabel metal3 s 0 8032 800 8152 0 FreeSans 480 0 0 0 chanx_left_in[4]
port 40 nsew signal input
flabel metal3 s 0 8304 800 8424 0 FreeSans 480 0 0 0 chanx_left_in[5]
port 41 nsew signal input
flabel metal3 s 0 8576 800 8696 0 FreeSans 480 0 0 0 chanx_left_in[6]
port 42 nsew signal input
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 chanx_left_in[7]
port 43 nsew signal input
flabel metal3 s 0 9120 800 9240 0 FreeSans 480 0 0 0 chanx_left_in[8]
port 44 nsew signal input
flabel metal3 s 0 9392 800 9512 0 FreeSans 480 0 0 0 chanx_left_in[9]
port 45 nsew signal input
flabel metal3 s 0 1504 800 1624 0 FreeSans 480 0 0 0 chanx_left_out[0]
port 46 nsew signal tristate
flabel metal3 s 0 4224 800 4344 0 FreeSans 480 0 0 0 chanx_left_out[10]
port 47 nsew signal tristate
flabel metal3 s 0 4496 800 4616 0 FreeSans 480 0 0 0 chanx_left_out[11]
port 48 nsew signal tristate
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 chanx_left_out[12]
port 49 nsew signal tristate
flabel metal3 s 0 5040 800 5160 0 FreeSans 480 0 0 0 chanx_left_out[13]
port 50 nsew signal tristate
flabel metal3 s 0 5312 800 5432 0 FreeSans 480 0 0 0 chanx_left_out[14]
port 51 nsew signal tristate
flabel metal3 s 0 5584 800 5704 0 FreeSans 480 0 0 0 chanx_left_out[15]
port 52 nsew signal tristate
flabel metal3 s 0 5856 800 5976 0 FreeSans 480 0 0 0 chanx_left_out[16]
port 53 nsew signal tristate
flabel metal3 s 0 6128 800 6248 0 FreeSans 480 0 0 0 chanx_left_out[17]
port 54 nsew signal tristate
flabel metal3 s 0 6400 800 6520 0 FreeSans 480 0 0 0 chanx_left_out[18]
port 55 nsew signal tristate
flabel metal3 s 0 6672 800 6792 0 FreeSans 480 0 0 0 chanx_left_out[19]
port 56 nsew signal tristate
flabel metal3 s 0 1776 800 1896 0 FreeSans 480 0 0 0 chanx_left_out[1]
port 57 nsew signal tristate
flabel metal3 s 0 2048 800 2168 0 FreeSans 480 0 0 0 chanx_left_out[2]
port 58 nsew signal tristate
flabel metal3 s 0 2320 800 2440 0 FreeSans 480 0 0 0 chanx_left_out[3]
port 59 nsew signal tristate
flabel metal3 s 0 2592 800 2712 0 FreeSans 480 0 0 0 chanx_left_out[4]
port 60 nsew signal tristate
flabel metal3 s 0 2864 800 2984 0 FreeSans 480 0 0 0 chanx_left_out[5]
port 61 nsew signal tristate
flabel metal3 s 0 3136 800 3256 0 FreeSans 480 0 0 0 chanx_left_out[6]
port 62 nsew signal tristate
flabel metal3 s 0 3408 800 3528 0 FreeSans 480 0 0 0 chanx_left_out[7]
port 63 nsew signal tristate
flabel metal3 s 0 3680 800 3800 0 FreeSans 480 0 0 0 chanx_left_out[8]
port 64 nsew signal tristate
flabel metal3 s 0 3952 800 4072 0 FreeSans 480 0 0 0 chanx_left_out[9]
port 65 nsew signal tristate
flabel metal3 s 19200 9256 20000 9376 0 FreeSans 480 0 0 0 chanx_right_in[0]
port 66 nsew signal input
flabel metal3 s 19200 11976 20000 12096 0 FreeSans 480 0 0 0 chanx_right_in[10]
port 67 nsew signal input
flabel metal3 s 19200 12248 20000 12368 0 FreeSans 480 0 0 0 chanx_right_in[11]
port 68 nsew signal input
flabel metal3 s 19200 12520 20000 12640 0 FreeSans 480 0 0 0 chanx_right_in[12]
port 69 nsew signal input
flabel metal3 s 19200 12792 20000 12912 0 FreeSans 480 0 0 0 chanx_right_in[13]
port 70 nsew signal input
flabel metal3 s 19200 13064 20000 13184 0 FreeSans 480 0 0 0 chanx_right_in[14]
port 71 nsew signal input
flabel metal3 s 19200 13336 20000 13456 0 FreeSans 480 0 0 0 chanx_right_in[15]
port 72 nsew signal input
flabel metal3 s 19200 13608 20000 13728 0 FreeSans 480 0 0 0 chanx_right_in[16]
port 73 nsew signal input
flabel metal3 s 19200 13880 20000 14000 0 FreeSans 480 0 0 0 chanx_right_in[17]
port 74 nsew signal input
flabel metal3 s 19200 14152 20000 14272 0 FreeSans 480 0 0 0 chanx_right_in[18]
port 75 nsew signal input
flabel metal3 s 19200 14424 20000 14544 0 FreeSans 480 0 0 0 chanx_right_in[19]
port 76 nsew signal input
flabel metal3 s 19200 9528 20000 9648 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 77 nsew signal input
flabel metal3 s 19200 9800 20000 9920 0 FreeSans 480 0 0 0 chanx_right_in[2]
port 78 nsew signal input
flabel metal3 s 19200 10072 20000 10192 0 FreeSans 480 0 0 0 chanx_right_in[3]
port 79 nsew signal input
flabel metal3 s 19200 10344 20000 10464 0 FreeSans 480 0 0 0 chanx_right_in[4]
port 80 nsew signal input
flabel metal3 s 19200 10616 20000 10736 0 FreeSans 480 0 0 0 chanx_right_in[5]
port 81 nsew signal input
flabel metal3 s 19200 10888 20000 11008 0 FreeSans 480 0 0 0 chanx_right_in[6]
port 82 nsew signal input
flabel metal3 s 19200 11160 20000 11280 0 FreeSans 480 0 0 0 chanx_right_in[7]
port 83 nsew signal input
flabel metal3 s 19200 11432 20000 11552 0 FreeSans 480 0 0 0 chanx_right_in[8]
port 84 nsew signal input
flabel metal3 s 19200 11704 20000 11824 0 FreeSans 480 0 0 0 chanx_right_in[9]
port 85 nsew signal input
flabel metal3 s 19200 3816 20000 3936 0 FreeSans 480 0 0 0 chanx_right_out[0]
port 86 nsew signal tristate
flabel metal3 s 19200 6536 20000 6656 0 FreeSans 480 0 0 0 chanx_right_out[10]
port 87 nsew signal tristate
flabel metal3 s 19200 6808 20000 6928 0 FreeSans 480 0 0 0 chanx_right_out[11]
port 88 nsew signal tristate
flabel metal3 s 19200 7080 20000 7200 0 FreeSans 480 0 0 0 chanx_right_out[12]
port 89 nsew signal tristate
flabel metal3 s 19200 7352 20000 7472 0 FreeSans 480 0 0 0 chanx_right_out[13]
port 90 nsew signal tristate
flabel metal3 s 19200 7624 20000 7744 0 FreeSans 480 0 0 0 chanx_right_out[14]
port 91 nsew signal tristate
flabel metal3 s 19200 7896 20000 8016 0 FreeSans 480 0 0 0 chanx_right_out[15]
port 92 nsew signal tristate
flabel metal3 s 19200 8168 20000 8288 0 FreeSans 480 0 0 0 chanx_right_out[16]
port 93 nsew signal tristate
flabel metal3 s 19200 8440 20000 8560 0 FreeSans 480 0 0 0 chanx_right_out[17]
port 94 nsew signal tristate
flabel metal3 s 19200 8712 20000 8832 0 FreeSans 480 0 0 0 chanx_right_out[18]
port 95 nsew signal tristate
flabel metal3 s 19200 8984 20000 9104 0 FreeSans 480 0 0 0 chanx_right_out[19]
port 96 nsew signal tristate
flabel metal3 s 19200 4088 20000 4208 0 FreeSans 480 0 0 0 chanx_right_out[1]
port 97 nsew signal tristate
flabel metal3 s 19200 4360 20000 4480 0 FreeSans 480 0 0 0 chanx_right_out[2]
port 98 nsew signal tristate
flabel metal3 s 19200 4632 20000 4752 0 FreeSans 480 0 0 0 chanx_right_out[3]
port 99 nsew signal tristate
flabel metal3 s 19200 4904 20000 5024 0 FreeSans 480 0 0 0 chanx_right_out[4]
port 100 nsew signal tristate
flabel metal3 s 19200 5176 20000 5296 0 FreeSans 480 0 0 0 chanx_right_out[5]
port 101 nsew signal tristate
flabel metal3 s 19200 5448 20000 5568 0 FreeSans 480 0 0 0 chanx_right_out[6]
port 102 nsew signal tristate
flabel metal3 s 19200 5720 20000 5840 0 FreeSans 480 0 0 0 chanx_right_out[7]
port 103 nsew signal tristate
flabel metal3 s 19200 5992 20000 6112 0 FreeSans 480 0 0 0 chanx_right_out[8]
port 104 nsew signal tristate
flabel metal3 s 19200 6264 20000 6384 0 FreeSans 480 0 0 0 chanx_right_out[9]
port 105 nsew signal tristate
flabel metal2 s 9954 16400 10010 17200 0 FreeSans 224 90 0 0 clk_1_N_out
port 106 nsew signal tristate
flabel metal2 s 17774 0 17830 800 0 FreeSans 224 90 0 0 clk_1_S_out
port 107 nsew signal tristate
flabel metal3 s 0 15376 800 15496 0 FreeSans 480 0 0 0 clk_1_W_in
port 108 nsew signal input
flabel metal3 s 19200 3544 20000 3664 0 FreeSans 480 0 0 0 clk_2_E_out
port 109 nsew signal tristate
flabel metal3 s 0 15104 800 15224 0 FreeSans 480 0 0 0 clk_2_W_in
port 110 nsew signal input
flabel metal3 s 0 13744 800 13864 0 FreeSans 480 0 0 0 clk_2_W_out
port 111 nsew signal tristate
flabel metal3 s 19200 3272 20000 3392 0 FreeSans 480 0 0 0 clk_3_E_out
port 112 nsew signal tristate
flabel metal3 s 0 14832 800 14952 0 FreeSans 480 0 0 0 clk_3_W_in
port 113 nsew signal input
flabel metal3 s 0 13472 800 13592 0 FreeSans 480 0 0 0 clk_3_W_out
port 114 nsew signal tristate
flabel metal2 s 13910 16400 13966 17200 0 FreeSans 224 90 0 0 prog_clk_0_N_in
port 115 nsew signal input
flabel metal2 s 17866 16400 17922 17200 0 FreeSans 224 90 0 0 prog_clk_0_W_out
port 116 nsew signal tristate
flabel metal3 s 19200 3000 20000 3120 0 FreeSans 480 0 0 0 prog_clk_1_N_out
port 117 nsew signal tristate
flabel metal2 s 18602 0 18658 800 0 FreeSans 224 90 0 0 prog_clk_1_S_out
port 118 nsew signal tristate
flabel metal3 s 0 14560 800 14680 0 FreeSans 480 0 0 0 prog_clk_1_W_in
port 119 nsew signal input
flabel metal3 s 19200 2728 20000 2848 0 FreeSans 480 0 0 0 prog_clk_2_E_out
port 120 nsew signal tristate
flabel metal3 s 0 14288 800 14408 0 FreeSans 480 0 0 0 prog_clk_2_W_in
port 121 nsew signal input
flabel metal3 s 0 13200 800 13320 0 FreeSans 480 0 0 0 prog_clk_2_W_out
port 122 nsew signal tristate
flabel metal3 s 19200 2456 20000 2576 0 FreeSans 480 0 0 0 prog_clk_3_E_out
port 123 nsew signal tristate
flabel metal3 s 0 14016 800 14136 0 FreeSans 480 0 0 0 prog_clk_3_W_in
port 124 nsew signal input
flabel metal3 s 0 12928 800 13048 0 FreeSans 480 0 0 0 prog_clk_3_W_out
port 125 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 20000 17200
<< end >>
