magic
tech sky130A
magscale 1 2
timestamp 1656242772
<< obsli1 >>
rect 1104 2159 21896 20689
<< obsm1 >>
rect 198 2128 22802 20800
<< metal2 >>
rect 202 22200 258 23000
rect 662 22200 718 23000
rect 1122 22200 1178 23000
rect 1582 22200 1638 23000
rect 2042 22200 2098 23000
rect 2502 22200 2558 23000
rect 2962 22200 3018 23000
rect 3422 22200 3478 23000
rect 3882 22200 3938 23000
rect 4342 22200 4398 23000
rect 4802 22200 4858 23000
rect 5262 22200 5318 23000
rect 5722 22200 5778 23000
rect 6182 22200 6238 23000
rect 6642 22200 6698 23000
rect 7102 22200 7158 23000
rect 7562 22200 7618 23000
rect 8022 22200 8078 23000
rect 8482 22200 8538 23000
rect 8942 22200 8998 23000
rect 9402 22200 9458 23000
rect 9862 22200 9918 23000
rect 10322 22200 10378 23000
rect 10782 22200 10838 23000
rect 11242 22200 11298 23000
rect 11702 22200 11758 23000
rect 12162 22200 12218 23000
rect 12622 22200 12678 23000
rect 13082 22200 13138 23000
rect 13542 22200 13598 23000
rect 14002 22200 14058 23000
rect 14462 22200 14518 23000
rect 14922 22200 14978 23000
rect 15382 22200 15438 23000
rect 15842 22200 15898 23000
rect 16302 22200 16358 23000
rect 16762 22200 16818 23000
rect 17222 22200 17278 23000
rect 17682 22200 17738 23000
rect 18142 22200 18198 23000
rect 18602 22200 18658 23000
rect 19062 22200 19118 23000
rect 19522 22200 19578 23000
rect 19982 22200 20038 23000
rect 20442 22200 20498 23000
rect 20902 22200 20958 23000
rect 21362 22200 21418 23000
rect 21822 22200 21878 23000
rect 22282 22200 22338 23000
rect 22742 22200 22798 23000
rect 11426 0 11482 800
<< obsm2 >>
rect 314 22144 606 22250
rect 774 22144 1066 22250
rect 1234 22144 1526 22250
rect 1694 22144 1986 22250
rect 2154 22144 2446 22250
rect 2614 22144 2906 22250
rect 3074 22144 3366 22250
rect 3534 22144 3826 22250
rect 3994 22144 4286 22250
rect 4454 22144 4746 22250
rect 4914 22144 5206 22250
rect 5374 22144 5666 22250
rect 5834 22144 6126 22250
rect 6294 22144 6586 22250
rect 6754 22144 7046 22250
rect 7214 22144 7506 22250
rect 7674 22144 7966 22250
rect 8134 22144 8426 22250
rect 8594 22144 8886 22250
rect 9054 22144 9346 22250
rect 9514 22144 9806 22250
rect 9974 22144 10266 22250
rect 10434 22144 10726 22250
rect 10894 22144 11186 22250
rect 11354 22144 11646 22250
rect 11814 22144 12106 22250
rect 12274 22144 12566 22250
rect 12734 22144 13026 22250
rect 13194 22144 13486 22250
rect 13654 22144 13946 22250
rect 14114 22144 14406 22250
rect 14574 22144 14866 22250
rect 15034 22144 15326 22250
rect 15494 22144 15786 22250
rect 15954 22144 16246 22250
rect 16414 22144 16706 22250
rect 16874 22144 17166 22250
rect 17334 22144 17626 22250
rect 17794 22144 18086 22250
rect 18254 22144 18546 22250
rect 18714 22144 19006 22250
rect 19174 22144 19466 22250
rect 19634 22144 19926 22250
rect 20094 22144 20386 22250
rect 20554 22144 20846 22250
rect 21014 22144 21306 22250
rect 21474 22144 21766 22250
rect 21934 22144 22226 22250
rect 22394 22144 22686 22250
rect 204 856 22796 22144
rect 204 734 11370 856
rect 11538 734 22796 856
<< metal3 >>
rect 0 21224 800 21344
rect 0 20816 800 20936
rect 0 20408 800 20528
rect 0 20000 800 20120
rect 0 19592 800 19712
rect 0 19184 800 19304
rect 0 18776 800 18896
rect 0 18368 800 18488
rect 0 17960 800 18080
rect 0 17552 800 17672
rect 0 17144 800 17264
rect 0 16736 800 16856
rect 0 16328 800 16448
rect 0 15920 800 16040
rect 0 15512 800 15632
rect 0 15104 800 15224
rect 0 14696 800 14816
rect 0 14288 800 14408
rect 0 13880 800 14000
rect 0 13472 800 13592
rect 0 13064 800 13184
rect 0 12656 800 12776
rect 0 12248 800 12368
rect 0 11840 800 11960
rect 0 11432 800 11552
rect 22200 11432 23000 11552
rect 0 11024 800 11144
rect 0 10616 800 10736
rect 0 10208 800 10328
rect 0 9800 800 9920
rect 0 9392 800 9512
rect 0 8984 800 9104
rect 0 8576 800 8696
rect 0 8168 800 8288
rect 0 7760 800 7880
rect 0 7352 800 7472
rect 0 6944 800 7064
rect 0 6536 800 6656
rect 0 6128 800 6248
rect 0 5720 800 5840
rect 0 5312 800 5432
rect 0 4904 800 5024
rect 0 4496 800 4616
rect 0 4088 800 4208
rect 0 3680 800 3800
rect 0 3272 800 3392
rect 0 2864 800 2984
rect 0 2456 800 2576
rect 0 2048 800 2168
rect 0 1640 800 1760
<< obsm3 >>
rect 880 21144 22200 21317
rect 800 21016 22200 21144
rect 880 20736 22200 21016
rect 800 20608 22200 20736
rect 880 20328 22200 20608
rect 800 20200 22200 20328
rect 880 19920 22200 20200
rect 800 19792 22200 19920
rect 880 19512 22200 19792
rect 800 19384 22200 19512
rect 880 19104 22200 19384
rect 800 18976 22200 19104
rect 880 18696 22200 18976
rect 800 18568 22200 18696
rect 880 18288 22200 18568
rect 800 18160 22200 18288
rect 880 17880 22200 18160
rect 800 17752 22200 17880
rect 880 17472 22200 17752
rect 800 17344 22200 17472
rect 880 17064 22200 17344
rect 800 16936 22200 17064
rect 880 16656 22200 16936
rect 800 16528 22200 16656
rect 880 16248 22200 16528
rect 800 16120 22200 16248
rect 880 15840 22200 16120
rect 800 15712 22200 15840
rect 880 15432 22200 15712
rect 800 15304 22200 15432
rect 880 15024 22200 15304
rect 800 14896 22200 15024
rect 880 14616 22200 14896
rect 800 14488 22200 14616
rect 880 14208 22200 14488
rect 800 14080 22200 14208
rect 880 13800 22200 14080
rect 800 13672 22200 13800
rect 880 13392 22200 13672
rect 800 13264 22200 13392
rect 880 12984 22200 13264
rect 800 12856 22200 12984
rect 880 12576 22200 12856
rect 800 12448 22200 12576
rect 880 12168 22200 12448
rect 800 12040 22200 12168
rect 880 11760 22200 12040
rect 800 11632 22200 11760
rect 880 11352 22120 11632
rect 800 11224 22200 11352
rect 880 10944 22200 11224
rect 800 10816 22200 10944
rect 880 10536 22200 10816
rect 800 10408 22200 10536
rect 880 10128 22200 10408
rect 800 10000 22200 10128
rect 880 9720 22200 10000
rect 800 9592 22200 9720
rect 880 9312 22200 9592
rect 800 9184 22200 9312
rect 880 8904 22200 9184
rect 800 8776 22200 8904
rect 880 8496 22200 8776
rect 800 8368 22200 8496
rect 880 8088 22200 8368
rect 800 7960 22200 8088
rect 880 7680 22200 7960
rect 800 7552 22200 7680
rect 880 7272 22200 7552
rect 800 7144 22200 7272
rect 880 6864 22200 7144
rect 800 6736 22200 6864
rect 880 6456 22200 6736
rect 800 6328 22200 6456
rect 880 6048 22200 6328
rect 800 5920 22200 6048
rect 880 5640 22200 5920
rect 800 5512 22200 5640
rect 880 5232 22200 5512
rect 800 5104 22200 5232
rect 880 4824 22200 5104
rect 800 4696 22200 4824
rect 880 4416 22200 4696
rect 800 4288 22200 4416
rect 880 4008 22200 4288
rect 800 3880 22200 4008
rect 880 3600 22200 3880
rect 800 3472 22200 3600
rect 880 3192 22200 3472
rect 800 3064 22200 3192
rect 880 2784 22200 3064
rect 800 2656 22200 2784
rect 880 2376 22200 2656
rect 800 2248 22200 2376
rect 880 1968 22200 2248
rect 800 1840 22200 1968
rect 880 1667 22200 1840
<< metal4 >>
rect 3543 2128 3863 20720
rect 6142 2128 6462 20720
rect 8741 2128 9061 20720
rect 11340 2128 11660 20720
rect 13939 2128 14259 20720
rect 16538 2128 16858 20720
rect 19137 2128 19457 20720
rect 21736 2128 22056 20720
<< obsm4 >>
rect 2083 6699 3463 19549
rect 3943 6699 6062 19549
rect 6542 6699 8661 19549
rect 9141 6699 11260 19549
rect 11740 6699 13189 19549
<< labels >>
rlabel metal4 s 6142 2128 6462 20720 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 11340 2128 11660 20720 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 16538 2128 16858 20720 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 21736 2128 22056 20720 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 3543 2128 3863 20720 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 8741 2128 9061 20720 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 13939 2128 14259 20720 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 19137 2128 19457 20720 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 22200 11432 23000 11552 6 ccff_head
port 3 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 ccff_tail
port 4 nsew signal output
rlabel metal3 s 0 5312 800 5432 6 chanx_left_in[0]
port 5 nsew signal input
rlabel metal3 s 0 9392 800 9512 6 chanx_left_in[10]
port 6 nsew signal input
rlabel metal3 s 0 9800 800 9920 6 chanx_left_in[11]
port 7 nsew signal input
rlabel metal3 s 0 10208 800 10328 6 chanx_left_in[12]
port 8 nsew signal input
rlabel metal3 s 0 10616 800 10736 6 chanx_left_in[13]
port 9 nsew signal input
rlabel metal3 s 0 11024 800 11144 6 chanx_left_in[14]
port 10 nsew signal input
rlabel metal3 s 0 11432 800 11552 6 chanx_left_in[15]
port 11 nsew signal input
rlabel metal3 s 0 11840 800 11960 6 chanx_left_in[16]
port 12 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 chanx_left_in[17]
port 13 nsew signal input
rlabel metal3 s 0 12656 800 12776 6 chanx_left_in[18]
port 14 nsew signal input
rlabel metal3 s 0 13064 800 13184 6 chanx_left_in[19]
port 15 nsew signal input
rlabel metal3 s 0 5720 800 5840 6 chanx_left_in[1]
port 16 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 chanx_left_in[2]
port 17 nsew signal input
rlabel metal3 s 0 6536 800 6656 6 chanx_left_in[3]
port 18 nsew signal input
rlabel metal3 s 0 6944 800 7064 6 chanx_left_in[4]
port 19 nsew signal input
rlabel metal3 s 0 7352 800 7472 6 chanx_left_in[5]
port 20 nsew signal input
rlabel metal3 s 0 7760 800 7880 6 chanx_left_in[6]
port 21 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 chanx_left_in[7]
port 22 nsew signal input
rlabel metal3 s 0 8576 800 8696 6 chanx_left_in[8]
port 23 nsew signal input
rlabel metal3 s 0 8984 800 9104 6 chanx_left_in[9]
port 24 nsew signal input
rlabel metal3 s 0 13472 800 13592 6 chanx_left_out[0]
port 25 nsew signal output
rlabel metal3 s 0 17552 800 17672 6 chanx_left_out[10]
port 26 nsew signal output
rlabel metal3 s 0 17960 800 18080 6 chanx_left_out[11]
port 27 nsew signal output
rlabel metal3 s 0 18368 800 18488 6 chanx_left_out[12]
port 28 nsew signal output
rlabel metal3 s 0 18776 800 18896 6 chanx_left_out[13]
port 29 nsew signal output
rlabel metal3 s 0 19184 800 19304 6 chanx_left_out[14]
port 30 nsew signal output
rlabel metal3 s 0 19592 800 19712 6 chanx_left_out[15]
port 31 nsew signal output
rlabel metal3 s 0 20000 800 20120 6 chanx_left_out[16]
port 32 nsew signal output
rlabel metal3 s 0 20408 800 20528 6 chanx_left_out[17]
port 33 nsew signal output
rlabel metal3 s 0 20816 800 20936 6 chanx_left_out[18]
port 34 nsew signal output
rlabel metal3 s 0 21224 800 21344 6 chanx_left_out[19]
port 35 nsew signal output
rlabel metal3 s 0 13880 800 14000 6 chanx_left_out[1]
port 36 nsew signal output
rlabel metal3 s 0 14288 800 14408 6 chanx_left_out[2]
port 37 nsew signal output
rlabel metal3 s 0 14696 800 14816 6 chanx_left_out[3]
port 38 nsew signal output
rlabel metal3 s 0 15104 800 15224 6 chanx_left_out[4]
port 39 nsew signal output
rlabel metal3 s 0 15512 800 15632 6 chanx_left_out[5]
port 40 nsew signal output
rlabel metal3 s 0 15920 800 16040 6 chanx_left_out[6]
port 41 nsew signal output
rlabel metal3 s 0 16328 800 16448 6 chanx_left_out[7]
port 42 nsew signal output
rlabel metal3 s 0 16736 800 16856 6 chanx_left_out[8]
port 43 nsew signal output
rlabel metal3 s 0 17144 800 17264 6 chanx_left_out[9]
port 44 nsew signal output
rlabel metal2 s 3882 22200 3938 23000 6 chany_top_in[0]
port 45 nsew signal input
rlabel metal2 s 8482 22200 8538 23000 6 chany_top_in[10]
port 46 nsew signal input
rlabel metal2 s 8942 22200 8998 23000 6 chany_top_in[11]
port 47 nsew signal input
rlabel metal2 s 9402 22200 9458 23000 6 chany_top_in[12]
port 48 nsew signal input
rlabel metal2 s 9862 22200 9918 23000 6 chany_top_in[13]
port 49 nsew signal input
rlabel metal2 s 10322 22200 10378 23000 6 chany_top_in[14]
port 50 nsew signal input
rlabel metal2 s 10782 22200 10838 23000 6 chany_top_in[15]
port 51 nsew signal input
rlabel metal2 s 11242 22200 11298 23000 6 chany_top_in[16]
port 52 nsew signal input
rlabel metal2 s 11702 22200 11758 23000 6 chany_top_in[17]
port 53 nsew signal input
rlabel metal2 s 12162 22200 12218 23000 6 chany_top_in[18]
port 54 nsew signal input
rlabel metal2 s 12622 22200 12678 23000 6 chany_top_in[19]
port 55 nsew signal input
rlabel metal2 s 4342 22200 4398 23000 6 chany_top_in[1]
port 56 nsew signal input
rlabel metal2 s 4802 22200 4858 23000 6 chany_top_in[2]
port 57 nsew signal input
rlabel metal2 s 5262 22200 5318 23000 6 chany_top_in[3]
port 58 nsew signal input
rlabel metal2 s 5722 22200 5778 23000 6 chany_top_in[4]
port 59 nsew signal input
rlabel metal2 s 6182 22200 6238 23000 6 chany_top_in[5]
port 60 nsew signal input
rlabel metal2 s 6642 22200 6698 23000 6 chany_top_in[6]
port 61 nsew signal input
rlabel metal2 s 7102 22200 7158 23000 6 chany_top_in[7]
port 62 nsew signal input
rlabel metal2 s 7562 22200 7618 23000 6 chany_top_in[8]
port 63 nsew signal input
rlabel metal2 s 8022 22200 8078 23000 6 chany_top_in[9]
port 64 nsew signal input
rlabel metal2 s 13082 22200 13138 23000 6 chany_top_out[0]
port 65 nsew signal output
rlabel metal2 s 17682 22200 17738 23000 6 chany_top_out[10]
port 66 nsew signal output
rlabel metal2 s 18142 22200 18198 23000 6 chany_top_out[11]
port 67 nsew signal output
rlabel metal2 s 18602 22200 18658 23000 6 chany_top_out[12]
port 68 nsew signal output
rlabel metal2 s 19062 22200 19118 23000 6 chany_top_out[13]
port 69 nsew signal output
rlabel metal2 s 19522 22200 19578 23000 6 chany_top_out[14]
port 70 nsew signal output
rlabel metal2 s 19982 22200 20038 23000 6 chany_top_out[15]
port 71 nsew signal output
rlabel metal2 s 20442 22200 20498 23000 6 chany_top_out[16]
port 72 nsew signal output
rlabel metal2 s 20902 22200 20958 23000 6 chany_top_out[17]
port 73 nsew signal output
rlabel metal2 s 21362 22200 21418 23000 6 chany_top_out[18]
port 74 nsew signal output
rlabel metal2 s 21822 22200 21878 23000 6 chany_top_out[19]
port 75 nsew signal output
rlabel metal2 s 13542 22200 13598 23000 6 chany_top_out[1]
port 76 nsew signal output
rlabel metal2 s 14002 22200 14058 23000 6 chany_top_out[2]
port 77 nsew signal output
rlabel metal2 s 14462 22200 14518 23000 6 chany_top_out[3]
port 78 nsew signal output
rlabel metal2 s 14922 22200 14978 23000 6 chany_top_out[4]
port 79 nsew signal output
rlabel metal2 s 15382 22200 15438 23000 6 chany_top_out[5]
port 80 nsew signal output
rlabel metal2 s 15842 22200 15898 23000 6 chany_top_out[6]
port 81 nsew signal output
rlabel metal2 s 16302 22200 16358 23000 6 chany_top_out[7]
port 82 nsew signal output
rlabel metal2 s 16762 22200 16818 23000 6 chany_top_out[8]
port 83 nsew signal output
rlabel metal2 s 17222 22200 17278 23000 6 chany_top_out[9]
port 84 nsew signal output
rlabel metal3 s 0 3680 800 3800 6 left_bottom_grid_pin_11_
port 85 nsew signal input
rlabel metal3 s 0 4088 800 4208 6 left_bottom_grid_pin_13_
port 86 nsew signal input
rlabel metal3 s 0 4496 800 4616 6 left_bottom_grid_pin_15_
port 87 nsew signal input
rlabel metal3 s 0 4904 800 5024 6 left_bottom_grid_pin_17_
port 88 nsew signal input
rlabel metal3 s 0 1640 800 1760 6 left_bottom_grid_pin_1_
port 89 nsew signal input
rlabel metal3 s 0 2048 800 2168 6 left_bottom_grid_pin_3_
port 90 nsew signal input
rlabel metal3 s 0 2456 800 2576 6 left_bottom_grid_pin_5_
port 91 nsew signal input
rlabel metal3 s 0 2864 800 2984 6 left_bottom_grid_pin_7_
port 92 nsew signal input
rlabel metal3 s 0 3272 800 3392 6 left_bottom_grid_pin_9_
port 93 nsew signal input
rlabel metal2 s 22282 22200 22338 23000 6 prog_clk_0_N_in
port 94 nsew signal input
rlabel metal2 s 202 22200 258 23000 6 top_left_grid_pin_42_
port 95 nsew signal input
rlabel metal2 s 662 22200 718 23000 6 top_left_grid_pin_43_
port 96 nsew signal input
rlabel metal2 s 1122 22200 1178 23000 6 top_left_grid_pin_44_
port 97 nsew signal input
rlabel metal2 s 1582 22200 1638 23000 6 top_left_grid_pin_45_
port 98 nsew signal input
rlabel metal2 s 2042 22200 2098 23000 6 top_left_grid_pin_46_
port 99 nsew signal input
rlabel metal2 s 2502 22200 2558 23000 6 top_left_grid_pin_47_
port 100 nsew signal input
rlabel metal2 s 2962 22200 3018 23000 6 top_left_grid_pin_48_
port 101 nsew signal input
rlabel metal2 s 3422 22200 3478 23000 6 top_left_grid_pin_49_
port 102 nsew signal input
rlabel metal2 s 22742 22200 22798 23000 6 top_right_grid_pin_1_
port 103 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 23000 23000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1259728
string GDS_FILE /home/marwan/clear_signoff_final/openlane/sb_2__0_/runs/sb_2__0_/results/signoff/sb_2__0_.magic.gds
string GDS_START 75876
<< end >>

